module tt_um_a1k0n_vgadonut (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire clknet_leaf_0_clk;
 wire net299;
 wire hsync;
 wire \vgadonut.bayer_j[0] ;
 wire \vgadonut.bayer_j[1] ;
 wire \vgadonut.donut.cA[0] ;
 wire \vgadonut.donut.cA[10] ;
 wire \vgadonut.donut.cA[11] ;
 wire \vgadonut.donut.cA[12] ;
 wire \vgadonut.donut.cA[13] ;
 wire \vgadonut.donut.cA[14] ;
 wire \vgadonut.donut.cA[15] ;
 wire \vgadonut.donut.cA[1] ;
 wire \vgadonut.donut.cA[2] ;
 wire \vgadonut.donut.cA[3] ;
 wire \vgadonut.donut.cA[4] ;
 wire \vgadonut.donut.cA[5] ;
 wire \vgadonut.donut.cA[6] ;
 wire \vgadonut.donut.cA[7] ;
 wire \vgadonut.donut.cA[8] ;
 wire \vgadonut.donut.cA[9] ;
 wire \vgadonut.donut.cAcB[0] ;
 wire \vgadonut.donut.cAcB[10] ;
 wire \vgadonut.donut.cAcB[11] ;
 wire \vgadonut.donut.cAcB[12] ;
 wire \vgadonut.donut.cAcB[13] ;
 wire \vgadonut.donut.cAcB[14] ;
 wire \vgadonut.donut.cAcB[15] ;
 wire \vgadonut.donut.cAcB[1] ;
 wire \vgadonut.donut.cAcB[2] ;
 wire \vgadonut.donut.cAcB[3] ;
 wire \vgadonut.donut.cAcB[4] ;
 wire \vgadonut.donut.cAcB[5] ;
 wire \vgadonut.donut.cAcB[6] ;
 wire \vgadonut.donut.cAcB[7] ;
 wire \vgadonut.donut.cAcB[8] ;
 wire \vgadonut.donut.cAcB[9] ;
 wire \vgadonut.donut.cAsB[0] ;
 wire \vgadonut.donut.cAsB[10] ;
 wire \vgadonut.donut.cAsB[11] ;
 wire \vgadonut.donut.cAsB[12] ;
 wire \vgadonut.donut.cAsB[13] ;
 wire \vgadonut.donut.cAsB[14] ;
 wire \vgadonut.donut.cAsB[15] ;
 wire \vgadonut.donut.cAsB[1] ;
 wire \vgadonut.donut.cAsB[2] ;
 wire \vgadonut.donut.cAsB[3] ;
 wire \vgadonut.donut.cAsB[4] ;
 wire \vgadonut.donut.cAsB[5] ;
 wire \vgadonut.donut.cAsB[6] ;
 wire \vgadonut.donut.cAsB[7] ;
 wire \vgadonut.donut.cAsB[8] ;
 wire \vgadonut.donut.cAsB[9] ;
 wire \vgadonut.donut.cB[0] ;
 wire \vgadonut.donut.cB[10] ;
 wire \vgadonut.donut.cB[11] ;
 wire \vgadonut.donut.cB[12] ;
 wire \vgadonut.donut.cB[13] ;
 wire \vgadonut.donut.cB[14] ;
 wire \vgadonut.donut.cB[15] ;
 wire \vgadonut.donut.cB[1] ;
 wire \vgadonut.donut.cB[2] ;
 wire \vgadonut.donut.cB[3] ;
 wire \vgadonut.donut.cB[4] ;
 wire \vgadonut.donut.cB[5] ;
 wire \vgadonut.donut.cB[6] ;
 wire \vgadonut.donut.cB[7] ;
 wire \vgadonut.donut.cB[8] ;
 wire \vgadonut.donut.cB[9] ;
 wire \vgadonut.donut.donut_luma[0] ;
 wire \vgadonut.donut.donut_luma[1] ;
 wire \vgadonut.donut.donut_luma[2] ;
 wire \vgadonut.donut.donut_luma[3] ;
 wire \vgadonut.donut.donut_luma[4] ;
 wire \vgadonut.donut.donut_luma[5] ;
 wire \vgadonut.donut.donut_visible ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[0] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[10] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[11] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[12] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[13] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[1] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[2] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[3] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[4] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[5] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[6] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[7] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[8] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[9] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[0] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[10] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[11] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[12] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[13] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[14] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[15] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[1] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[2] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[3] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[4] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[5] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[6] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[7] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[8] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[9] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[0] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[10] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[11] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[12] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[13] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[14] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[15] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[1] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[2] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[3] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[4] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[5] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[6] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[7] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[8] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[9] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[10] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[11] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[12] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[13] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[8] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[9] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[0] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[10] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[11] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[12] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[13] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[14] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[15] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[1] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[2] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[3] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[4] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[5] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[6] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[7] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[8] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[9] ;
 wire \vgadonut.donut.donuthit.hit ;
 wire \vgadonut.donut.donuthit.light[10] ;
 wire \vgadonut.donut.donuthit.light[11] ;
 wire \vgadonut.donut.donuthit.light[12] ;
 wire \vgadonut.donut.donuthit.light[13] ;
 wire \vgadonut.donut.donuthit.light[8] ;
 wire \vgadonut.donut.donuthit.light[9] ;
 wire \vgadonut.donut.donuthit.rx[10] ;
 wire \vgadonut.donut.donuthit.rx[11] ;
 wire \vgadonut.donut.donuthit.rx[12] ;
 wire \vgadonut.donut.donuthit.rx[13] ;
 wire \vgadonut.donut.donuthit.rx[14] ;
 wire \vgadonut.donut.donuthit.rx[15] ;
 wire \vgadonut.donut.donuthit.rx[5] ;
 wire \vgadonut.donut.donuthit.rx[6] ;
 wire \vgadonut.donut.donuthit.rx[7] ;
 wire \vgadonut.donut.donuthit.rx[8] ;
 wire \vgadonut.donut.donuthit.rx[9] ;
 wire \vgadonut.donut.donuthit.rxin[0] ;
 wire \vgadonut.donut.donuthit.rxin[10] ;
 wire \vgadonut.donut.donuthit.rxin[11] ;
 wire \vgadonut.donut.donuthit.rxin[12] ;
 wire \vgadonut.donut.donuthit.rxin[13] ;
 wire \vgadonut.donut.donuthit.rxin[14] ;
 wire \vgadonut.donut.donuthit.rxin[15] ;
 wire \vgadonut.donut.donuthit.rxin[1] ;
 wire \vgadonut.donut.donuthit.rxin[2] ;
 wire \vgadonut.donut.donuthit.rxin[3] ;
 wire \vgadonut.donut.donuthit.rxin[4] ;
 wire \vgadonut.donut.donuthit.rxin[5] ;
 wire \vgadonut.donut.donuthit.rxin[6] ;
 wire \vgadonut.donut.donuthit.rxin[7] ;
 wire \vgadonut.donut.donuthit.rxin[8] ;
 wire \vgadonut.donut.donuthit.rxin[9] ;
 wire \vgadonut.donut.donuthit.ry[10] ;
 wire \vgadonut.donut.donuthit.ry[11] ;
 wire \vgadonut.donut.donuthit.ry[12] ;
 wire \vgadonut.donut.donuthit.ry[13] ;
 wire \vgadonut.donut.donuthit.ry[14] ;
 wire \vgadonut.donut.donuthit.ry[15] ;
 wire \vgadonut.donut.donuthit.ry[5] ;
 wire \vgadonut.donut.donuthit.ry[6] ;
 wire \vgadonut.donut.donuthit.ry[7] ;
 wire \vgadonut.donut.donuthit.ry[8] ;
 wire \vgadonut.donut.donuthit.ry[9] ;
 wire \vgadonut.donut.donuthit.ryin[0] ;
 wire \vgadonut.donut.donuthit.ryin[10] ;
 wire \vgadonut.donut.donuthit.ryin[11] ;
 wire \vgadonut.donut.donuthit.ryin[12] ;
 wire \vgadonut.donut.donuthit.ryin[13] ;
 wire \vgadonut.donut.donuthit.ryin[14] ;
 wire \vgadonut.donut.donuthit.ryin[15] ;
 wire \vgadonut.donut.donuthit.ryin[1] ;
 wire \vgadonut.donut.donuthit.ryin[2] ;
 wire \vgadonut.donut.donuthit.ryin[3] ;
 wire \vgadonut.donut.donuthit.ryin[4] ;
 wire \vgadonut.donut.donuthit.ryin[5] ;
 wire \vgadonut.donut.donuthit.ryin[6] ;
 wire \vgadonut.donut.donuthit.ryin[7] ;
 wire \vgadonut.donut.donuthit.ryin[8] ;
 wire \vgadonut.donut.donuthit.ryin[9] ;
 wire \vgadonut.donut.donuthit.rz[10] ;
 wire \vgadonut.donut.donuthit.rz[11] ;
 wire \vgadonut.donut.donuthit.rz[12] ;
 wire \vgadonut.donut.donuthit.rz[13] ;
 wire \vgadonut.donut.donuthit.rz[14] ;
 wire \vgadonut.donut.donuthit.rz[15] ;
 wire \vgadonut.donut.donuthit.rz[5] ;
 wire \vgadonut.donut.donuthit.rz[6] ;
 wire \vgadonut.donut.donuthit.rz[7] ;
 wire \vgadonut.donut.donuthit.rz[8] ;
 wire \vgadonut.donut.donuthit.rz[9] ;
 wire \vgadonut.donut.donuthit.rzin[0] ;
 wire \vgadonut.donut.donuthit.rzin[10] ;
 wire \vgadonut.donut.donuthit.rzin[11] ;
 wire \vgadonut.donut.donuthit.rzin[12] ;
 wire \vgadonut.donut.donuthit.rzin[13] ;
 wire \vgadonut.donut.donuthit.rzin[14] ;
 wire \vgadonut.donut.donuthit.rzin[15] ;
 wire \vgadonut.donut.donuthit.rzin[1] ;
 wire \vgadonut.donut.donuthit.rzin[2] ;
 wire \vgadonut.donut.donuthit.rzin[3] ;
 wire \vgadonut.donut.donuthit.rzin[4] ;
 wire \vgadonut.donut.donuthit.rzin[5] ;
 wire \vgadonut.donut.donuthit.rzin[6] ;
 wire \vgadonut.donut.donuthit.rzin[7] ;
 wire \vgadonut.donut.donuthit.rzin[8] ;
 wire \vgadonut.donut.donuthit.rzin[9] ;
 wire \vgadonut.donut.donuthit.t[0] ;
 wire \vgadonut.donut.donuthit.t[10] ;
 wire \vgadonut.donut.donuthit.t[11] ;
 wire \vgadonut.donut.donuthit.t[12] ;
 wire \vgadonut.donut.donuthit.t[13] ;
 wire \vgadonut.donut.donuthit.t[14] ;
 wire \vgadonut.donut.donuthit.t[15] ;
 wire \vgadonut.donut.donuthit.t[1] ;
 wire \vgadonut.donut.donuthit.t[2] ;
 wire \vgadonut.donut.donuthit.t[3] ;
 wire \vgadonut.donut.donuthit.t[4] ;
 wire \vgadonut.donut.donuthit.t[5] ;
 wire \vgadonut.donut.donuthit.t[6] ;
 wire \vgadonut.donut.donuthit.t[7] ;
 wire \vgadonut.donut.donuthit.t[8] ;
 wire \vgadonut.donut.donuthit.t[9] ;
 wire \vgadonut.donut.frame ;
 wire \vgadonut.donut.h_count[0] ;
 wire \vgadonut.donut.h_count[10] ;
 wire \vgadonut.donut.h_count[1] ;
 wire \vgadonut.donut.h_count[2] ;
 wire \vgadonut.donut.h_count[3] ;
 wire \vgadonut.donut.h_count[4] ;
 wire \vgadonut.donut.h_count[5] ;
 wire \vgadonut.donut.h_count[6] ;
 wire \vgadonut.donut.h_count[7] ;
 wire \vgadonut.donut.h_count[8] ;
 wire \vgadonut.donut.h_count[9] ;
 wire \vgadonut.donut.rx6[0] ;
 wire \vgadonut.donut.rx6[1] ;
 wire \vgadonut.donut.rx6[2] ;
 wire \vgadonut.donut.rx6[3] ;
 wire \vgadonut.donut.rx6[4] ;
 wire \vgadonut.donut.rx6[5] ;
 wire \vgadonut.donut.ry6[0] ;
 wire \vgadonut.donut.ry6[1] ;
 wire \vgadonut.donut.ry6[2] ;
 wire \vgadonut.donut.ry6[3] ;
 wire \vgadonut.donut.ry6[4] ;
 wire \vgadonut.donut.ry6[5] ;
 wire \vgadonut.donut.rz6[0] ;
 wire \vgadonut.donut.rz6[1] ;
 wire \vgadonut.donut.rz6[2] ;
 wire \vgadonut.donut.rz6[3] ;
 wire \vgadonut.donut.rz6[4] ;
 wire \vgadonut.donut.rz6[5] ;
 wire \vgadonut.donut.sA[0] ;
 wire \vgadonut.donut.sA[10] ;
 wire \vgadonut.donut.sA[11] ;
 wire \vgadonut.donut.sA[12] ;
 wire \vgadonut.donut.sA[13] ;
 wire \vgadonut.donut.sA[14] ;
 wire \vgadonut.donut.sA[15] ;
 wire \vgadonut.donut.sA[1] ;
 wire \vgadonut.donut.sA[2] ;
 wire \vgadonut.donut.sA[3] ;
 wire \vgadonut.donut.sA[4] ;
 wire \vgadonut.donut.sA[5] ;
 wire \vgadonut.donut.sA[6] ;
 wire \vgadonut.donut.sA[7] ;
 wire \vgadonut.donut.sA[8] ;
 wire \vgadonut.donut.sA[9] ;
 wire \vgadonut.donut.sAcB[0] ;
 wire \vgadonut.donut.sAcB[10] ;
 wire \vgadonut.donut.sAcB[11] ;
 wire \vgadonut.donut.sAcB[12] ;
 wire \vgadonut.donut.sAcB[13] ;
 wire \vgadonut.donut.sAcB[14] ;
 wire \vgadonut.donut.sAcB[15] ;
 wire \vgadonut.donut.sAcB[1] ;
 wire \vgadonut.donut.sAcB[2] ;
 wire \vgadonut.donut.sAcB[3] ;
 wire \vgadonut.donut.sAcB[4] ;
 wire \vgadonut.donut.sAcB[5] ;
 wire \vgadonut.donut.sAcB[6] ;
 wire \vgadonut.donut.sAcB[7] ;
 wire \vgadonut.donut.sAcB[8] ;
 wire \vgadonut.donut.sAcB[9] ;
 wire \vgadonut.donut.sAsB[0] ;
 wire \vgadonut.donut.sAsB[10] ;
 wire \vgadonut.donut.sAsB[11] ;
 wire \vgadonut.donut.sAsB[12] ;
 wire \vgadonut.donut.sAsB[13] ;
 wire \vgadonut.donut.sAsB[14] ;
 wire \vgadonut.donut.sAsB[15] ;
 wire \vgadonut.donut.sAsB[1] ;
 wire \vgadonut.donut.sAsB[2] ;
 wire \vgadonut.donut.sAsB[3] ;
 wire \vgadonut.donut.sAsB[4] ;
 wire \vgadonut.donut.sAsB[5] ;
 wire \vgadonut.donut.sAsB[6] ;
 wire \vgadonut.donut.sAsB[7] ;
 wire \vgadonut.donut.sAsB[8] ;
 wire \vgadonut.donut.sAsB[9] ;
 wire \vgadonut.donut.sB[0] ;
 wire \vgadonut.donut.sB[1] ;
 wire \vgadonut.donut.v_count[2] ;
 wire \vgadonut.donut.v_count[3] ;
 wire \vgadonut.donut.v_count[4] ;
 wire \vgadonut.donut.v_count[5] ;
 wire \vgadonut.donut.v_count[6] ;
 wire \vgadonut.donut.v_count[7] ;
 wire \vgadonut.donut.v_count[8] ;
 wire \vgadonut.donut.v_count[9] ;
 wire \vgadonut.donut.ycA[0] ;
 wire \vgadonut.donut.ycA[10] ;
 wire \vgadonut.donut.ycA[11] ;
 wire \vgadonut.donut.ycA[12] ;
 wire \vgadonut.donut.ycA[13] ;
 wire \vgadonut.donut.ycA[14] ;
 wire \vgadonut.donut.ycA[15] ;
 wire \vgadonut.donut.ycA[16] ;
 wire \vgadonut.donut.ycA[17] ;
 wire \vgadonut.donut.ycA[18] ;
 wire \vgadonut.donut.ycA[19] ;
 wire \vgadonut.donut.ycA[1] ;
 wire \vgadonut.donut.ycA[20] ;
 wire \vgadonut.donut.ycA[21] ;
 wire \vgadonut.donut.ycA[2] ;
 wire \vgadonut.donut.ycA[3] ;
 wire \vgadonut.donut.ycA[4] ;
 wire \vgadonut.donut.ycA[5] ;
 wire \vgadonut.donut.ycA[6] ;
 wire \vgadonut.donut.ycA[7] ;
 wire \vgadonut.donut.ycA[8] ;
 wire \vgadonut.donut.ycA[9] ;
 wire \vgadonut.donut.ysA[0] ;
 wire \vgadonut.donut.ysA[10] ;
 wire \vgadonut.donut.ysA[11] ;
 wire \vgadonut.donut.ysA[12] ;
 wire \vgadonut.donut.ysA[13] ;
 wire \vgadonut.donut.ysA[14] ;
 wire \vgadonut.donut.ysA[15] ;
 wire \vgadonut.donut.ysA[16] ;
 wire \vgadonut.donut.ysA[17] ;
 wire \vgadonut.donut.ysA[18] ;
 wire \vgadonut.donut.ysA[19] ;
 wire \vgadonut.donut.ysA[1] ;
 wire \vgadonut.donut.ysA[20] ;
 wire \vgadonut.donut.ysA[21] ;
 wire \vgadonut.donut.ysA[2] ;
 wire \vgadonut.donut.ysA[3] ;
 wire \vgadonut.donut.ysA[4] ;
 wire \vgadonut.donut.ysA[5] ;
 wire \vgadonut.donut.ysA[6] ;
 wire \vgadonut.donut.ysA[7] ;
 wire \vgadonut.donut.ysA[8] ;
 wire \vgadonut.donut.ysA[9] ;
 wire \vgadonut.frame[1] ;
 wire \vgadonut.frame[2] ;
 wire \vgadonut.frame[3] ;
 wire \vgadonut.frame[4] ;
 wire \vgadonut.frame[5] ;
 wire \vgadonut.frame[6] ;
 wire \vgadonut.frame[7] ;
 wire \vgadonut.vsync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _10709_ (.A(\vgadonut.donut.h_count[6] ),
    .X(_09637_));
 sg13g2_buf_2 _10710_ (.A(\vgadonut.donut.h_count[9] ),
    .X(_09645_));
 sg13g2_buf_1 _10711_ (.A(\vgadonut.donut.h_count[8] ),
    .X(_09654_));
 sg13g2_inv_1 _10712_ (.Y(_09663_),
    .A(\vgadonut.donut.h_count[7] ));
 sg13g2_inv_1 _10713_ (.Y(_09672_),
    .A(\vgadonut.donut.h_count[10] ));
 sg13g2_nor4_1 _10714_ (.A(_09645_),
    .B(_09654_),
    .C(_09663_),
    .D(_09672_),
    .Y(_09683_));
 sg13g2_buf_1 _10715_ (.A(\vgadonut.donut.h_count[5] ),
    .X(_09694_));
 sg13g2_inv_1 _10716_ (.Y(_09705_),
    .A(_09694_));
 sg13g2_buf_2 _10717_ (.A(\vgadonut.donut.h_count[3] ),
    .X(_09716_));
 sg13g2_buf_1 _10718_ (.A(\vgadonut.donut.h_count[4] ),
    .X(_09726_));
 sg13g2_nand2_1 _10719_ (.Y(_09737_),
    .A(_09716_),
    .B(_09726_));
 sg13g2_inv_1 _10720_ (.Y(_09748_),
    .A(_09683_));
 sg13g2_nor4_1 _10721_ (.A(_09705_),
    .B(net255),
    .C(_09737_),
    .D(_09748_),
    .Y(_09759_));
 sg13g2_buf_1 _10722_ (.A(\vgadonut.donut.h_count[2] ),
    .X(_09769_));
 sg13g2_inv_1 _10723_ (.Y(_09780_),
    .A(_09645_));
 sg13g2_a21oi_1 _10724_ (.A1(_09780_),
    .A2(_00172_),
    .Y(_09790_),
    .B1(_09672_));
 sg13g2_a221oi_1 _10725_ (.B2(net254),
    .C1(_09790_),
    .B1(_09759_),
    .A1(net255),
    .Y(_09800_),
    .A2(_09683_));
 sg13g2_buf_2 _10726_ (.A(\vgadonut.donut.frame ),
    .X(_09811_));
 sg13g2_xnor2_1 _10727_ (.Y(_09821_),
    .A(_09811_),
    .B(_00170_));
 sg13g2_buf_1 _10728_ (.A(\vgadonut.bayer_j[0] ),
    .X(_09832_));
 sg13g2_nand3_1 _10729_ (.B(net254),
    .C(_09832_),
    .A(_09821_),
    .Y(_09842_));
 sg13g2_inv_1 _10730_ (.Y(_09853_),
    .A(net254));
 sg13g2_inv_1 _10731_ (.Y(_09863_),
    .A(_09832_));
 sg13g2_nand3b_1 _10732_ (.B(_09853_),
    .C(_09863_),
    .Y(_09874_),
    .A_N(_09821_));
 sg13g2_buf_2 _10733_ (.A(\vgadonut.donut.h_count[0] ),
    .X(_09884_));
 sg13g2_buf_2 _10734_ (.A(\vgadonut.bayer_j[1] ),
    .X(_09894_));
 sg13g2_buf_1 _10735_ (.A(\vgadonut.donut.h_count[1] ),
    .X(_09905_));
 sg13g2_xnor2_1 _10736_ (.Y(_09915_),
    .A(_09905_),
    .B(_09811_));
 sg13g2_buf_1 _10737_ (.A(_09915_),
    .X(_09925_));
 sg13g2_xnor2_1 _10738_ (.Y(_09935_),
    .A(_09894_),
    .B(_09925_));
 sg13g2_inv_1 _10739_ (.Y(_09946_),
    .A(_09935_));
 sg13g2_nand2b_1 _10740_ (.Y(_09954_),
    .B(_09946_),
    .A_N(_09884_));
 sg13g2_a21oi_1 _10741_ (.A1(_09842_),
    .A2(_09874_),
    .Y(_09962_),
    .B1(_09954_));
 sg13g2_nand2_1 _10742_ (.Y(_09971_),
    .A(_09800_),
    .B(_09962_));
 sg13g2_buf_2 _10743_ (.A(_09971_),
    .X(_09979_));
 sg13g2_inv_1 _10744_ (.Y(_09988_),
    .A(_09979_));
 sg13g2_buf_2 _10745_ (.A(_09988_),
    .X(_09996_));
 sg13g2_inv_1 _10746_ (.Y(_10004_),
    .A(net275));
 sg13g2_buf_1 _10747_ (.A(_00169_),
    .X(_10011_));
 sg13g2_inv_1 _10748_ (.Y(_10020_),
    .A(_09654_));
 sg13g2_nor3_1 _10749_ (.A(_09645_),
    .B(_10011_),
    .C(_10020_),
    .Y(_10029_));
 sg13g2_nor2b_1 _10750_ (.A(_09716_),
    .B_N(_10029_),
    .Y(_10040_));
 sg13g2_nand2_1 _10751_ (.Y(_10051_),
    .A(_09694_),
    .B(net255));
 sg13g2_nor3_1 _10752_ (.A(_09726_),
    .B(_09663_),
    .C(_10051_),
    .Y(_10062_));
 sg13g2_inv_1 _10753_ (.Y(_10073_),
    .A(_09905_));
 sg13g2_nor3_1 _10754_ (.A(_09884_),
    .B(_10073_),
    .C(_09853_),
    .Y(_10084_));
 sg13g2_nand3_1 _10755_ (.B(_10062_),
    .C(_10084_),
    .A(_10040_),
    .Y(_10095_));
 sg13g2_buf_2 _10756_ (.A(_10095_),
    .X(_10106_));
 sg13g2_inv_2 _10757_ (.Y(_10117_),
    .A(_10106_));
 sg13g2_nor2_1 _10758_ (.A(_10004_),
    .B(_10117_),
    .Y(_10128_));
 sg13g2_nand2_1 _10759_ (.Y(_10139_),
    .A(_09996_),
    .B(_10128_));
 sg13g2_buf_1 _10760_ (.A(_10139_),
    .X(_10150_));
 sg13g2_buf_1 _10761_ (.A(_10150_),
    .X(_10161_));
 sg13g2_nor2_1 _10762_ (.A(_00046_),
    .B(net106),
    .Y(_10172_));
 sg13g2_nand2b_1 _10763_ (.Y(_10183_),
    .B(net106),
    .A_N(\vgadonut.donut.donut_luma[5] ));
 sg13g2_nand2b_1 _10764_ (.Y(_10192_),
    .B(_10183_),
    .A_N(_10172_));
 sg13g2_buf_1 _10765_ (.A(_10192_),
    .X(_10196_));
 sg13g2_inv_1 _10766_ (.Y(_10203_),
    .A(_10196_));
 sg13g2_buf_1 _10767_ (.A(_10203_),
    .X(_00014_));
 sg13g2_nor2_1 _10768_ (.A(\vgadonut.donut.donuthit.light[12] ),
    .B(net106),
    .Y(_10217_));
 sg13g2_nand2b_1 _10769_ (.Y(_10228_),
    .B(net106),
    .A_N(\vgadonut.donut.donut_luma[4] ));
 sg13g2_nand2b_1 _10770_ (.Y(_10239_),
    .B(_10228_),
    .A_N(_10217_));
 sg13g2_buf_2 _10771_ (.A(_10239_),
    .X(_10250_));
 sg13g2_inv_2 _10772_ (.Y(_10261_),
    .A(_10250_));
 sg13g2_buf_1 _10773_ (.A(_10261_),
    .X(_00173_));
 sg13g2_nor2_1 _10774_ (.A(\vgadonut.donut.donuthit.light[9] ),
    .B(_10150_),
    .Y(_10282_));
 sg13g2_nand2b_1 _10775_ (.Y(_10293_),
    .B(_10150_),
    .A_N(\vgadonut.donut.donut_luma[1] ));
 sg13g2_nand2b_1 _10776_ (.Y(_10304_),
    .B(_10293_),
    .A_N(_10282_));
 sg13g2_buf_2 _10777_ (.A(_10304_),
    .X(_10315_));
 sg13g2_inv_1 _10778_ (.Y(_10324_),
    .A(_10315_));
 sg13g2_buf_1 _10779_ (.A(_10324_),
    .X(_00177_));
 sg13g2_nor2_1 _10780_ (.A(\vgadonut.donut.donuthit.light[8] ),
    .B(_10150_),
    .Y(_10345_));
 sg13g2_nand2b_1 _10781_ (.Y(_10356_),
    .B(_10150_),
    .A_N(\vgadonut.donut.donut_luma[0] ));
 sg13g2_nand2b_1 _10782_ (.Y(_10367_),
    .B(_10356_),
    .A_N(_10345_));
 sg13g2_buf_2 _10783_ (.A(_10367_),
    .X(_10377_));
 sg13g2_inv_2 _10784_ (.Y(_00178_),
    .A(_10377_));
 sg13g2_nor2_1 _10785_ (.A(\vgadonut.donut.donuthit.light[10] ),
    .B(net106),
    .Y(_10397_));
 sg13g2_nand2b_1 _10786_ (.Y(_10408_),
    .B(net106),
    .A_N(\vgadonut.donut.donut_luma[2] ));
 sg13g2_nand2b_1 _10787_ (.Y(_10419_),
    .B(_10408_),
    .A_N(_10397_));
 sg13g2_buf_2 _10788_ (.A(_10419_),
    .X(_00543_));
 sg13g2_inv_1 _10789_ (.Y(_00179_),
    .A(_00543_));
 sg13g2_nor2_1 _10790_ (.A(\vgadonut.donut.donuthit.light[11] ),
    .B(_10161_),
    .Y(_00562_));
 sg13g2_nand2b_1 _10791_ (.Y(_00573_),
    .B(_10161_),
    .A_N(\vgadonut.donut.donut_luma[3] ));
 sg13g2_nand2b_1 _10792_ (.Y(_00584_),
    .B(_00573_),
    .A_N(_00562_));
 sg13g2_buf_1 _10793_ (.A(_00584_),
    .X(_00595_));
 sg13g2_inv_1 _10794_ (.Y(_00606_),
    .A(_00595_));
 sg13g2_buf_1 _10795_ (.A(_00606_),
    .X(_00617_));
 sg13g2_buf_1 _10796_ (.A(net79),
    .X(_00180_));
 sg13g2_nor2_2 _10797_ (.A(_10377_),
    .B(net88),
    .Y(_00638_));
 sg13g2_nor2_1 _10798_ (.A(_10377_),
    .B(_00543_),
    .Y(_00649_));
 sg13g2_nor2_1 _10799_ (.A(_00178_),
    .B(net87),
    .Y(_00660_));
 sg13g2_nor2_1 _10800_ (.A(_00649_),
    .B(_00660_),
    .Y(_00671_));
 sg13g2_inv_1 _10801_ (.Y(_00682_),
    .A(_00671_));
 sg13g2_o21ai_1 _10802_ (.B1(net78),
    .Y(_00693_),
    .A1(_00638_),
    .A2(_00682_));
 sg13g2_nor2_1 _10803_ (.A(_10196_),
    .B(_10261_),
    .Y(_00704_));
 sg13g2_inv_1 _10804_ (.Y(_00715_),
    .A(_00704_));
 sg13g2_nor2_2 _10805_ (.A(_10315_),
    .B(_00178_),
    .Y(_00726_));
 sg13g2_nor3_1 _10806_ (.A(net78),
    .B(_00649_),
    .C(_00726_),
    .Y(_00737_));
 sg13g2_nor2_1 _10807_ (.A(_00715_),
    .B(_00737_),
    .Y(_00748_));
 sg13g2_nor2_2 _10808_ (.A(net88),
    .B(net87),
    .Y(_00759_));
 sg13g2_nor2_1 _10809_ (.A(_00595_),
    .B(_00759_),
    .Y(_00770_));
 sg13g2_inv_1 _10810_ (.Y(_00781_),
    .A(_00770_));
 sg13g2_nor2_1 _10811_ (.A(_00178_),
    .B(_00781_),
    .Y(_00792_));
 sg13g2_buf_1 _10812_ (.A(_10196_),
    .X(_00803_));
 sg13g2_o21ai_1 _10813_ (.B1(net86),
    .Y(_00814_),
    .A1(_10377_),
    .A2(_00770_));
 sg13g2_nand2_1 _10814_ (.Y(_00825_),
    .A(net80),
    .B(net86));
 sg13g2_o21ai_1 _10815_ (.B1(_00825_),
    .Y(_00836_),
    .A1(_00792_),
    .A2(_00814_));
 sg13g2_nor2_1 _10816_ (.A(_10315_),
    .B(net87),
    .Y(_00847_));
 sg13g2_buf_1 _10817_ (.A(_00595_),
    .X(_00858_));
 sg13g2_o21ai_1 _10818_ (.B1(_00858_),
    .Y(_00869_),
    .A1(_00847_),
    .A2(_00682_));
 sg13g2_nor2_1 _10819_ (.A(_00595_),
    .B(_00847_),
    .Y(_00880_));
 sg13g2_nand2_1 _10820_ (.Y(_00891_),
    .A(_00671_),
    .B(_00880_));
 sg13g2_buf_1 _10821_ (.A(_10250_),
    .X(_00902_));
 sg13g2_a21o_1 _10822_ (.A2(_00891_),
    .A1(_00869_),
    .B1(net84),
    .X(_00913_));
 sg13g2_a22oi_1 _10823_ (.Y(_00009_),
    .B1(_00836_),
    .B2(_00913_),
    .A2(_00748_),
    .A1(_00693_));
 sg13g2_nand2_1 _10824_ (.Y(_00934_),
    .A(net87),
    .B(_00858_));
 sg13g2_nand2_1 _10825_ (.Y(_00945_),
    .A(_00934_),
    .B(net88));
 sg13g2_nor2_1 _10826_ (.A(_00715_),
    .B(_00682_),
    .Y(_00956_));
 sg13g2_nor2_1 _10827_ (.A(_00543_),
    .B(net88),
    .Y(_00967_));
 sg13g2_nor2_1 _10828_ (.A(_00649_),
    .B(_00967_),
    .Y(_00978_));
 sg13g2_nor2_1 _10829_ (.A(_00638_),
    .B(_00978_),
    .Y(_00989_));
 sg13g2_inv_1 _10830_ (.Y(_01000_),
    .A(_00989_));
 sg13g2_nor2_1 _10831_ (.A(net87),
    .B(_00726_),
    .Y(_01011_));
 sg13g2_inv_1 _10832_ (.Y(_01022_),
    .A(_01011_));
 sg13g2_a21oi_1 _10833_ (.A1(_01000_),
    .A2(_01022_),
    .Y(_01033_),
    .B1(net85));
 sg13g2_nor2_1 _10834_ (.A(net88),
    .B(_00606_),
    .Y(_01044_));
 sg13g2_inv_1 _10835_ (.Y(_01055_),
    .A(_01044_));
 sg13g2_nand3b_1 _10836_ (.B(net84),
    .C(_01055_),
    .Y(_01066_),
    .A_N(_01033_));
 sg13g2_nor2_1 _10837_ (.A(_10250_),
    .B(_00606_),
    .Y(_01077_));
 sg13g2_inv_1 _10838_ (.Y(_01088_),
    .A(_01077_));
 sg13g2_nor2_1 _10839_ (.A(_10315_),
    .B(_00543_),
    .Y(_01099_));
 sg13g2_buf_1 _10840_ (.A(_01099_),
    .X(_01110_));
 sg13g2_inv_1 _10841_ (.Y(_01121_),
    .A(_01110_));
 sg13g2_o21ai_1 _10842_ (.B1(_01121_),
    .Y(_01132_),
    .A1(_00638_),
    .A2(_01022_));
 sg13g2_o21ai_1 _10843_ (.B1(net86),
    .Y(_01143_),
    .A1(_01088_),
    .A2(_01132_));
 sg13g2_a21oi_1 _10844_ (.A1(net80),
    .A2(_01033_),
    .Y(_01154_),
    .B1(_01143_));
 sg13g2_a22oi_1 _10845_ (.Y(_00010_),
    .B1(_01066_),
    .B2(_01154_),
    .A2(_00956_),
    .A1(_00945_));
 sg13g2_nor2_1 _10846_ (.A(_00638_),
    .B(_01022_),
    .Y(_01175_));
 sg13g2_nand2_1 _10847_ (.Y(_01186_),
    .A(_01175_),
    .B(net78));
 sg13g2_nor2_1 _10848_ (.A(_00177_),
    .B(_00178_),
    .Y(_01197_));
 sg13g2_nor2_1 _10849_ (.A(net79),
    .B(_00967_),
    .Y(_01208_));
 sg13g2_nand2b_1 _10850_ (.Y(_01219_),
    .B(_01208_),
    .A_N(_01197_));
 sg13g2_a21oi_1 _10851_ (.A1(_01110_),
    .A2(_00180_),
    .Y(_01230_),
    .B1(_00173_));
 sg13g2_nand3_1 _10852_ (.B(_01219_),
    .C(_01230_),
    .A(_01186_),
    .Y(_01241_));
 sg13g2_nor2_1 _10853_ (.A(_00543_),
    .B(_01197_),
    .Y(_01252_));
 sg13g2_o21ai_1 _10854_ (.B1(_10261_),
    .Y(_01263_),
    .A1(_00759_),
    .A2(_01252_));
 sg13g2_nor2_1 _10855_ (.A(_10315_),
    .B(_10377_),
    .Y(_01274_));
 sg13g2_a21oi_1 _10856_ (.A1(_01274_),
    .A2(_00543_),
    .Y(_01285_),
    .B1(_00967_));
 sg13g2_nor2_1 _10857_ (.A(net79),
    .B(_01285_),
    .Y(_01296_));
 sg13g2_a21oi_1 _10858_ (.A1(_01263_),
    .A2(_01088_),
    .Y(_01307_),
    .B1(_01296_));
 sg13g2_a21oi_1 _10859_ (.A1(_00682_),
    .A2(net88),
    .Y(_01318_),
    .B1(_00759_));
 sg13g2_nand2_1 _10860_ (.Y(_01329_),
    .A(_00934_),
    .B(_10250_));
 sg13g2_a21oi_1 _10861_ (.A1(_01318_),
    .A2(net78),
    .Y(_01340_),
    .B1(_01329_));
 sg13g2_nor3_1 _10862_ (.A(_10203_),
    .B(_01307_),
    .C(_01340_),
    .Y(_01351_));
 sg13g2_a21o_1 _10863_ (.A2(_01241_),
    .A1(_00014_),
    .B1(_01351_),
    .X(_00011_));
 sg13g2_nor2_1 _10864_ (.A(_10377_),
    .B(_01121_),
    .Y(_01372_));
 sg13g2_inv_1 _10865_ (.Y(_01383_),
    .A(_01372_));
 sg13g2_nor2_1 _10866_ (.A(net85),
    .B(_10261_),
    .Y(_01394_));
 sg13g2_inv_1 _10867_ (.Y(_01405_),
    .A(_00649_));
 sg13g2_nand3_1 _10868_ (.B(_01121_),
    .C(net79),
    .A(_01405_),
    .Y(_01416_));
 sg13g2_nand2_1 _10869_ (.Y(_01427_),
    .A(_01110_),
    .B(net85));
 sg13g2_nand2_1 _10870_ (.Y(_01438_),
    .A(_01416_),
    .B(_01427_));
 sg13g2_a22oi_1 _10871_ (.Y(_01449_),
    .B1(net80),
    .B2(_01438_),
    .A2(_01394_),
    .A1(_01383_));
 sg13g2_a21oi_1 _10872_ (.A1(_01197_),
    .A2(net78),
    .Y(_01460_),
    .B1(net87));
 sg13g2_a21o_1 _10873_ (.A2(_00902_),
    .A1(_01460_),
    .B1(_00803_),
    .X(_01471_));
 sg13g2_o21ai_1 _10874_ (.B1(_01471_),
    .Y(_00012_),
    .A1(net81),
    .A2(_01449_));
 sg13g2_a21oi_1 _10875_ (.A1(_01372_),
    .A2(net78),
    .Y(_01492_),
    .B1(net80));
 sg13g2_nand2_1 _10876_ (.Y(_01503_),
    .A(_01252_),
    .B(net79));
 sg13g2_o21ai_1 _10877_ (.B1(net86),
    .Y(_01514_),
    .A1(_10250_),
    .A2(_01503_));
 sg13g2_buf_1 _10878_ (.A(_01514_),
    .X(_00228_));
 sg13g2_nor3_1 _10879_ (.A(net88),
    .B(_00178_),
    .C(net87),
    .Y(_01535_));
 sg13g2_o21ai_1 _10880_ (.B1(_00902_),
    .Y(_01546_),
    .A1(net85),
    .A2(_01535_));
 sg13g2_nand2_1 _10881_ (.Y(_01557_),
    .A(_01546_),
    .B(net81));
 sg13g2_o21ai_1 _10882_ (.B1(_01557_),
    .Y(_00013_),
    .A1(_01492_),
    .A2(_00228_));
 sg13g2_a21oi_1 _10883_ (.A1(_00726_),
    .A2(net78),
    .Y(_01578_),
    .B1(net84));
 sg13g2_a22oi_1 _10884_ (.Y(_01589_),
    .B1(_01578_),
    .B2(_01318_),
    .A2(_00179_),
    .A1(net84));
 sg13g2_nor2_1 _10885_ (.A(_10315_),
    .B(net78),
    .Y(_01600_));
 sg13g2_nor2_1 _10886_ (.A(net79),
    .B(_00671_),
    .Y(_01611_));
 sg13g2_inv_1 _10887_ (.Y(_01622_),
    .A(_01611_));
 sg13g2_o21ai_1 _10888_ (.B1(_01622_),
    .Y(_01633_),
    .A1(_00660_),
    .A2(_01600_));
 sg13g2_nand2_1 _10889_ (.Y(_01644_),
    .A(_10203_),
    .B(_10261_));
 sg13g2_a21oi_1 _10890_ (.A1(_00660_),
    .A2(_01044_),
    .Y(_01655_),
    .B1(_01644_));
 sg13g2_a21oi_1 _10891_ (.A1(_01633_),
    .A2(_00704_),
    .Y(_01666_),
    .B1(_01655_));
 sg13g2_o21ai_1 _10892_ (.B1(_01666_),
    .Y(_00000_),
    .A1(net81),
    .A2(_01589_));
 sg13g2_a21oi_1 _10893_ (.A1(_01405_),
    .A2(_00880_),
    .Y(_01687_),
    .B1(_01296_));
 sg13g2_nor3_1 _10894_ (.A(_10250_),
    .B(_00726_),
    .C(_01622_),
    .Y(_01698_));
 sg13g2_a21o_1 _10895_ (.A2(net84),
    .A1(_01687_),
    .B1(_01698_),
    .X(_01709_));
 sg13g2_nand2_1 _10896_ (.Y(_01720_),
    .A(_01110_),
    .B(net79));
 sg13g2_nand2_1 _10897_ (.Y(_01731_),
    .A(_01720_),
    .B(_10261_));
 sg13g2_a21oi_1 _10898_ (.A1(_01383_),
    .A2(net85),
    .Y(_01742_),
    .B1(_01731_));
 sg13g2_nor3_1 _10899_ (.A(net81),
    .B(_01394_),
    .C(_01742_),
    .Y(_01753_));
 sg13g2_a21oi_1 _10900_ (.A1(_01709_),
    .A2(net81),
    .Y(_00001_),
    .B1(_01753_));
 sg13g2_nand2_1 _10901_ (.Y(_01774_),
    .A(_01000_),
    .B(_00880_));
 sg13g2_nand3_1 _10902_ (.B(net84),
    .C(_01427_),
    .A(_01774_),
    .Y(_01785_));
 sg13g2_nand3_1 _10903_ (.B(_01121_),
    .C(_01077_),
    .A(_01022_),
    .Y(_01796_));
 sg13g2_nand3_1 _10904_ (.B(net81),
    .C(_01796_),
    .A(_01785_),
    .Y(_01806_));
 sg13g2_o21ai_1 _10905_ (.B1(_01806_),
    .Y(_00002_),
    .A1(net81),
    .A2(_01731_));
 sg13g2_a22oi_1 _10906_ (.Y(_01827_),
    .B1(_01077_),
    .B2(_01000_),
    .A2(_01394_),
    .A1(_01383_));
 sg13g2_o21ai_1 _10907_ (.B1(net81),
    .Y(_01838_),
    .A1(_00759_),
    .A2(_01827_));
 sg13g2_o21ai_1 _10908_ (.B1(_01838_),
    .Y(_00003_),
    .A1(_00825_),
    .A2(_01720_));
 sg13g2_a221oi_1 _10909_ (.B2(_01208_),
    .C1(_00715_),
    .B1(_00671_),
    .A1(_00770_),
    .Y(_01856_),
    .A2(_01405_));
 sg13g2_nand3b_1 _10910_ (.B(_01022_),
    .C(net85),
    .Y(_01857_),
    .A_N(_00638_));
 sg13g2_nand3b_1 _10911_ (.B(_00978_),
    .C(net79),
    .Y(_01858_),
    .A_N(_00660_));
 sg13g2_nand3_1 _10912_ (.B(_01858_),
    .C(net84),
    .A(_01857_),
    .Y(_01859_));
 sg13g2_nand3_1 _10913_ (.B(net80),
    .C(_00891_),
    .A(_01622_),
    .Y(_01860_));
 sg13g2_nand3_1 _10914_ (.B(net86),
    .C(_01860_),
    .A(_01859_),
    .Y(_01861_));
 sg13g2_a21oi_1 _10915_ (.A1(_00759_),
    .A2(net85),
    .Y(_01862_),
    .B1(_10250_));
 sg13g2_nand2_1 _10916_ (.Y(_01863_),
    .A(_01862_),
    .B(_10203_));
 sg13g2_nand3b_1 _10917_ (.B(_01861_),
    .C(_01863_),
    .Y(_00004_),
    .A_N(_01856_));
 sg13g2_nor3_1 _10918_ (.A(_00178_),
    .B(_01110_),
    .C(_01044_),
    .Y(_01864_));
 sg13g2_a21oi_1 _10919_ (.A1(_01720_),
    .A2(_01055_),
    .Y(_01865_),
    .B1(_10377_));
 sg13g2_nor3_1 _10920_ (.A(_00715_),
    .B(_01864_),
    .C(_01865_),
    .Y(_01866_));
 sg13g2_o21ai_1 _10921_ (.B1(net88),
    .Y(_01867_),
    .A1(_00543_),
    .A2(_00178_));
 sg13g2_inv_1 _10922_ (.Y(_01868_),
    .A(_01274_));
 sg13g2_nand2_1 _10923_ (.Y(_01869_),
    .A(_01868_),
    .B(_00543_));
 sg13g2_nor2_2 _10924_ (.A(_00606_),
    .B(_01252_),
    .Y(_01870_));
 sg13g2_a22oi_1 _10925_ (.Y(_01871_),
    .B1(_01869_),
    .B2(_01870_),
    .A2(_01867_),
    .A1(_00617_));
 sg13g2_o21ai_1 _10926_ (.B1(net85),
    .Y(_01872_),
    .A1(_00967_),
    .A2(_01175_));
 sg13g2_nand3_1 _10927_ (.B(_10261_),
    .C(_01774_),
    .A(_01872_),
    .Y(_01873_));
 sg13g2_o21ai_1 _10928_ (.B1(_01873_),
    .Y(_01874_),
    .A1(net80),
    .A2(_01871_));
 sg13g2_nand2_1 _10929_ (.Y(_01875_),
    .A(_01874_),
    .B(net86));
 sg13g2_nand3b_1 _10930_ (.B(_01875_),
    .C(_01863_),
    .Y(_00005_),
    .A_N(_01866_));
 sg13g2_nor2_1 _10931_ (.A(_01110_),
    .B(_00781_),
    .Y(_01876_));
 sg13g2_nor3_1 _10932_ (.A(_01870_),
    .B(_00792_),
    .C(_01876_),
    .Y(_01877_));
 sg13g2_nor2_1 _10933_ (.A(_00617_),
    .B(_01869_),
    .Y(_01878_));
 sg13g2_nor2_1 _10934_ (.A(_10250_),
    .B(_01878_),
    .Y(_01879_));
 sg13g2_a21oi_1 _10935_ (.A1(_01879_),
    .A2(_01416_),
    .Y(_01880_),
    .B1(_10203_));
 sg13g2_o21ai_1 _10936_ (.B1(_01880_),
    .Y(_01881_),
    .A1(net80),
    .A2(_01877_));
 sg13g2_inv_1 _10937_ (.Y(_01882_),
    .A(_01870_));
 sg13g2_nand2b_1 _10938_ (.Y(_01883_),
    .B(_00880_),
    .A_N(_00726_));
 sg13g2_o21ai_1 _10939_ (.B1(_01883_),
    .Y(_01884_),
    .A1(_01535_),
    .A2(_01882_));
 sg13g2_a21oi_1 _10940_ (.A1(_01884_),
    .A2(_00704_),
    .Y(_01885_),
    .B1(_01655_));
 sg13g2_nand2_1 _10941_ (.Y(_00006_),
    .A(_01881_),
    .B(_01885_));
 sg13g2_nor2_1 _10942_ (.A(_01870_),
    .B(_01876_),
    .Y(_01886_));
 sg13g2_inv_1 _10943_ (.Y(_01887_),
    .A(_00228_));
 sg13g2_inv_1 _10944_ (.Y(_01888_),
    .A(_01879_));
 sg13g2_o21ai_1 _10945_ (.B1(_01888_),
    .Y(_01889_),
    .A1(net80),
    .A2(_00770_));
 sg13g2_a22oi_1 _10946_ (.Y(_00007_),
    .B1(_01887_),
    .B2(_01889_),
    .A2(_01886_),
    .A1(_00704_));
 sg13g2_a22oi_1 _10947_ (.Y(_00008_),
    .B1(_00803_),
    .B2(_01888_),
    .A2(_01882_),
    .A1(_01230_));
 sg13g2_buf_2 _10948_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[8] ),
    .X(_01890_));
 sg13g2_buf_2 _10949_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[8] ),
    .X(_01891_));
 sg13g2_xor2_1 _10950_ (.B(_01891_),
    .A(_01890_),
    .X(_01892_));
 sg13g2_buf_2 _10951_ (.A(_01892_),
    .X(_01893_));
 sg13g2_buf_8 _10952_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[7] ),
    .X(_01894_));
 sg13g2_buf_2 _10953_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[7] ),
    .X(_01895_));
 sg13g2_nand2_1 _10954_ (.Y(_01896_),
    .A(_01894_),
    .B(_01895_));
 sg13g2_inv_1 _10955_ (.Y(_01897_),
    .A(_01896_));
 sg13g2_nand2_1 _10956_ (.Y(_01898_),
    .A(_01893_),
    .B(_01897_));
 sg13g2_nand2_1 _10957_ (.Y(_01899_),
    .A(_01890_),
    .B(_01891_));
 sg13g2_nand2_1 _10958_ (.Y(_01900_),
    .A(_01898_),
    .B(_01899_));
 sg13g2_buf_8 _10959_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[9] ),
    .X(_01901_));
 sg13g2_buf_8 _10960_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[9] ),
    .X(_01902_));
 sg13g2_xnor2_1 _10961_ (.Y(_01903_),
    .A(_01901_),
    .B(_01902_));
 sg13g2_inv_2 _10962_ (.Y(_01904_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[10] ));
 sg13g2_inv_4 _10963_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[10] ),
    .Y(_01905_));
 sg13g2_nand2_1 _10964_ (.Y(_01906_),
    .A(_01904_),
    .B(_01905_));
 sg13g2_nand2_1 _10965_ (.Y(_01907_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[10] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[10] ));
 sg13g2_nand2_1 _10966_ (.Y(_01908_),
    .A(_01906_),
    .B(_01907_));
 sg13g2_buf_2 _10967_ (.A(_01908_),
    .X(_01909_));
 sg13g2_nor2_1 _10968_ (.A(_01903_),
    .B(_01909_),
    .Y(_01910_));
 sg13g2_nand2_1 _10969_ (.Y(_01911_),
    .A(_01900_),
    .B(_01910_));
 sg13g2_nand2_1 _10970_ (.Y(_01912_),
    .A(_01901_),
    .B(_01902_));
 sg13g2_inv_1 _10971_ (.Y(_01913_),
    .A(_01906_));
 sg13g2_a21oi_1 _10972_ (.A1(_01912_),
    .A2(_01907_),
    .Y(_01914_),
    .B1(_01913_));
 sg13g2_inv_1 _10973_ (.Y(_01915_),
    .A(_01914_));
 sg13g2_nand2_1 _10974_ (.Y(_01916_),
    .A(_01911_),
    .B(_01915_));
 sg13g2_buf_8 _10975_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[12] ),
    .X(_01917_));
 sg13g2_buf_2 _10976_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[12] ),
    .X(_01918_));
 sg13g2_xor2_1 _10977_ (.B(_01918_),
    .A(_01917_),
    .X(_01919_));
 sg13g2_buf_8 _10978_ (.A(_01919_),
    .X(_01920_));
 sg13g2_buf_8 _10979_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[11] ),
    .X(_01921_));
 sg13g2_buf_2 _10980_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[11] ),
    .X(_01922_));
 sg13g2_xor2_1 _10981_ (.B(_01922_),
    .A(_01921_),
    .X(_01923_));
 sg13g2_buf_8 _10982_ (.A(_01923_),
    .X(_01924_));
 sg13g2_nand2_1 _10983_ (.Y(_01925_),
    .A(_01920_),
    .B(_01924_));
 sg13g2_inv_1 _10984_ (.Y(_01926_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[13] ));
 sg13g2_nor2_1 _10985_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[13] ),
    .B(_01926_),
    .Y(_01927_));
 sg13g2_inv_1 _10986_ (.Y(_01928_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[13] ));
 sg13g2_nor2_1 _10987_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[13] ),
    .B(_01928_),
    .Y(_01929_));
 sg13g2_nor2_2 _10988_ (.A(_01927_),
    .B(_01929_),
    .Y(_01930_));
 sg13g2_inv_4 _10989_ (.A(_01930_),
    .Y(_01931_));
 sg13g2_nor2_1 _10990_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[14] ),
    .B(\vgadonut.donut.donuthit.cordicxy.yin[14] ),
    .Y(_01932_));
 sg13g2_nand2_1 _10991_ (.Y(_01933_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[14] ),
    .B(\vgadonut.donut.donuthit.cordicxy.yin[14] ));
 sg13g2_inv_1 _10992_ (.Y(_01934_),
    .A(_01933_));
 sg13g2_nor2_1 _10993_ (.A(_01932_),
    .B(_01934_),
    .Y(_01935_));
 sg13g2_buf_2 _10994_ (.A(_01935_),
    .X(_01936_));
 sg13g2_nand2_1 _10995_ (.Y(_01937_),
    .A(_01931_),
    .B(_01936_));
 sg13g2_nor2_1 _10996_ (.A(_01925_),
    .B(_01937_),
    .Y(_01938_));
 sg13g2_nand2_1 _10997_ (.Y(_01939_),
    .A(_01921_),
    .B(_01922_));
 sg13g2_inv_1 _10998_ (.Y(_01940_),
    .A(_01939_));
 sg13g2_nand2_1 _10999_ (.Y(_01941_),
    .A(_01917_),
    .B(_01918_));
 sg13g2_inv_1 _11000_ (.Y(_01942_),
    .A(_01941_));
 sg13g2_a21oi_1 _11001_ (.A1(_01920_),
    .A2(_01940_),
    .Y(_01943_),
    .B1(_01942_));
 sg13g2_nand2_1 _11002_ (.Y(_01944_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[13] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[13] ));
 sg13g2_inv_1 _11003_ (.Y(_01945_),
    .A(_01944_));
 sg13g2_a21oi_1 _11004_ (.A1(_01936_),
    .A2(_01945_),
    .Y(_01946_),
    .B1(_01934_));
 sg13g2_o21ai_1 _11005_ (.B1(_01946_),
    .Y(_01947_),
    .A1(_01937_),
    .A2(_01943_));
 sg13g2_a21oi_1 _11006_ (.A1(_01916_),
    .A2(_01938_),
    .Y(_01948_),
    .B1(_01947_));
 sg13g2_buf_8 _11007_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[1] ),
    .X(_01949_));
 sg13g2_buf_8 _11008_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[1] ),
    .X(_01950_));
 sg13g2_nor2_1 _11009_ (.A(_01949_),
    .B(_01950_),
    .Y(_01951_));
 sg13g2_nand2_1 _11010_ (.Y(_01952_),
    .A(_01949_),
    .B(_01950_));
 sg13g2_inv_1 _11011_ (.Y(_01953_),
    .A(_01952_));
 sg13g2_nor2_1 _11012_ (.A(_01951_),
    .B(_01953_),
    .Y(_01954_));
 sg13g2_buf_8 _11013_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[2] ),
    .X(_01955_));
 sg13g2_buf_8 _11014_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[2] ),
    .X(_01956_));
 sg13g2_xor2_1 _11015_ (.B(net253),
    .A(_01955_),
    .X(_01957_));
 sg13g2_buf_2 _11016_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[0] ),
    .X(_01958_));
 sg13g2_buf_2 _11017_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[0] ),
    .X(_01959_));
 sg13g2_nand2_1 _11018_ (.Y(_01960_),
    .A(_01958_),
    .B(_01959_));
 sg13g2_inv_1 _11019_ (.Y(_01961_),
    .A(_01960_));
 sg13g2_nand3_1 _11020_ (.B(_01957_),
    .C(_01961_),
    .A(_01954_),
    .Y(_01962_));
 sg13g2_nor2_1 _11021_ (.A(_01955_),
    .B(net253),
    .Y(_01963_));
 sg13g2_nand2_1 _11022_ (.Y(_01964_),
    .A(_01955_),
    .B(net253));
 sg13g2_o21ai_1 _11023_ (.B1(_01964_),
    .Y(_01965_),
    .A1(_01952_),
    .A2(_01963_));
 sg13g2_inv_1 _11024_ (.Y(_01966_),
    .A(_01965_));
 sg13g2_nand2_1 _11025_ (.Y(_01967_),
    .A(_01962_),
    .B(_01966_));
 sg13g2_buf_8 _11026_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[4] ),
    .X(_01968_));
 sg13g2_buf_8 _11027_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[4] ),
    .X(_01969_));
 sg13g2_xnor2_1 _11028_ (.Y(_01970_),
    .A(_01968_),
    .B(_01969_));
 sg13g2_buf_2 _11029_ (.A(_01970_),
    .X(_01971_));
 sg13g2_inv_2 _11030_ (.Y(_01972_),
    .A(_01971_));
 sg13g2_buf_2 _11031_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[3] ),
    .X(_01973_));
 sg13g2_inv_2 _11032_ (.Y(_01974_),
    .A(_01973_));
 sg13g2_buf_2 _11033_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[3] ),
    .X(_01975_));
 sg13g2_nand2_1 _11034_ (.Y(_01976_),
    .A(_01974_),
    .B(_01975_));
 sg13g2_inv_2 _11035_ (.Y(_01977_),
    .A(_01975_));
 sg13g2_nand2_1 _11036_ (.Y(_01978_),
    .A(_01977_),
    .B(_01973_));
 sg13g2_nand2_1 _11037_ (.Y(_01979_),
    .A(_01976_),
    .B(_01978_));
 sg13g2_nand2_1 _11038_ (.Y(_01980_),
    .A(_01972_),
    .B(_01979_));
 sg13g2_buf_8 _11039_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[5] ),
    .X(_01981_));
 sg13g2_buf_8 _11040_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[5] ),
    .X(_01982_));
 sg13g2_xnor2_1 _11041_ (.Y(_01983_),
    .A(_01981_),
    .B(_01982_));
 sg13g2_buf_2 _11042_ (.A(_01983_),
    .X(_01984_));
 sg13g2_inv_4 _11043_ (.A(_01984_),
    .Y(_01985_));
 sg13g2_buf_8 _11044_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[6] ),
    .X(_01986_));
 sg13g2_buf_8 _11045_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[6] ),
    .X(_01987_));
 sg13g2_nor2_1 _11046_ (.A(_01986_),
    .B(_01987_),
    .Y(_01988_));
 sg13g2_nand2_1 _11047_ (.Y(_01989_),
    .A(_01986_),
    .B(_01987_));
 sg13g2_inv_1 _11048_ (.Y(_01990_),
    .A(_01989_));
 sg13g2_nor2_1 _11049_ (.A(_01988_),
    .B(_01990_),
    .Y(_01991_));
 sg13g2_nand2_1 _11050_ (.Y(_01992_),
    .A(_01985_),
    .B(_01991_));
 sg13g2_nor2_1 _11051_ (.A(_01980_),
    .B(_01992_),
    .Y(_01993_));
 sg13g2_nand2_1 _11052_ (.Y(_01994_),
    .A(_01967_),
    .B(_01993_));
 sg13g2_inv_4 _11053_ (.A(_01987_),
    .Y(_01995_));
 sg13g2_nor2_1 _11054_ (.A(_01986_),
    .B(_01995_),
    .Y(_01996_));
 sg13g2_nand2_1 _11055_ (.Y(_01997_),
    .A(_01995_),
    .B(_01986_));
 sg13g2_inv_2 _11056_ (.Y(_01998_),
    .A(_01997_));
 sg13g2_nor2_2 _11057_ (.A(_01996_),
    .B(_01998_),
    .Y(_01999_));
 sg13g2_nor2_1 _11058_ (.A(_01984_),
    .B(_01999_),
    .Y(_02000_));
 sg13g2_nand2_1 _11059_ (.Y(_02001_),
    .A(_01975_),
    .B(_01973_));
 sg13g2_nor2_1 _11060_ (.A(_01968_),
    .B(_01969_),
    .Y(_02002_));
 sg13g2_nand2_1 _11061_ (.Y(_02003_),
    .A(_01968_),
    .B(_01969_));
 sg13g2_o21ai_1 _11062_ (.B1(_02003_),
    .Y(_02004_),
    .A1(_02001_),
    .A2(_02002_));
 sg13g2_nand2_1 _11063_ (.Y(_02005_),
    .A(_01981_),
    .B(_01982_));
 sg13g2_a21oi_1 _11064_ (.A1(_02005_),
    .A2(_01989_),
    .Y(_02006_),
    .B1(_01988_));
 sg13g2_a21oi_1 _11065_ (.A1(_02000_),
    .A2(_02004_),
    .Y(_02007_),
    .B1(_02006_));
 sg13g2_nand2_1 _11066_ (.Y(_02008_),
    .A(_01994_),
    .B(_02007_));
 sg13g2_xnor2_1 _11067_ (.Y(_02009_),
    .A(_01894_),
    .B(_01895_));
 sg13g2_buf_4 _11068_ (.X(_02010_),
    .A(_02009_));
 sg13g2_inv_1 _11069_ (.Y(_02011_),
    .A(_01891_));
 sg13g2_nor2_1 _11070_ (.A(_01890_),
    .B(_02011_),
    .Y(_02012_));
 sg13g2_inv_2 _11071_ (.Y(_02013_),
    .A(_01890_));
 sg13g2_nor2_1 _11072_ (.A(_01891_),
    .B(_02013_),
    .Y(_02014_));
 sg13g2_nor2_1 _11073_ (.A(_02012_),
    .B(_02014_),
    .Y(_02015_));
 sg13g2_nor2_1 _11074_ (.A(_02010_),
    .B(_02015_),
    .Y(_02016_));
 sg13g2_nand2_1 _11075_ (.Y(_02017_),
    .A(_02016_),
    .B(_01910_));
 sg13g2_nor3_1 _11076_ (.A(_01925_),
    .B(_01937_),
    .C(_02017_),
    .Y(_02018_));
 sg13g2_nand2_1 _11077_ (.Y(_02019_),
    .A(_02008_),
    .B(_02018_));
 sg13g2_buf_2 _11078_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[15] ),
    .X(_02020_));
 sg13g2_xnor2_1 _11079_ (.Y(_02021_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[15] ),
    .B(_02020_));
 sg13g2_buf_1 _11080_ (.A(_02021_),
    .X(_02022_));
 sg13g2_inv_1 _11081_ (.Y(_02023_),
    .A(net187));
 sg13g2_nand3_1 _11082_ (.B(_02019_),
    .C(_02023_),
    .A(_01948_),
    .Y(_02024_));
 sg13g2_buf_1 _11083_ (.A(_02024_),
    .X(_02025_));
 sg13g2_xnor2_1 _11084_ (.Y(_02026_),
    .A(_01949_),
    .B(_01950_));
 sg13g2_xnor2_1 _11085_ (.Y(_02027_),
    .A(_01955_),
    .B(net253));
 sg13g2_buf_1 _11086_ (.A(_02027_),
    .X(_02028_));
 sg13g2_inv_2 _11087_ (.Y(_02029_),
    .A(_01958_));
 sg13g2_nand2_1 _11088_ (.Y(_02030_),
    .A(_02029_),
    .B(_01959_));
 sg13g2_nand3_1 _11089_ (.B(_02028_),
    .C(_02030_),
    .A(_02026_),
    .Y(_02031_));
 sg13g2_inv_2 _11090_ (.Y(_02032_),
    .A(_01949_));
 sg13g2_nor2_1 _11091_ (.A(_01950_),
    .B(_02032_),
    .Y(_02033_));
 sg13g2_inv_2 _11092_ (.Y(_02034_),
    .A(_01955_));
 sg13g2_nand2_1 _11093_ (.Y(_02035_),
    .A(_02034_),
    .B(net253));
 sg13g2_nor2_1 _11094_ (.A(net253),
    .B(_02034_),
    .Y(_02036_));
 sg13g2_a21oi_1 _11095_ (.A1(_02033_),
    .A2(_02035_),
    .Y(_02037_),
    .B1(_02036_));
 sg13g2_nand2_1 _11096_ (.Y(_02038_),
    .A(_02031_),
    .B(_02037_));
 sg13g2_xnor2_1 _11097_ (.Y(_02039_),
    .A(_01975_),
    .B(_01973_));
 sg13g2_buf_2 _11098_ (.A(_02039_),
    .X(_02040_));
 sg13g2_nand2_1 _11099_ (.Y(_02041_),
    .A(_01971_),
    .B(_02040_));
 sg13g2_nand2_1 _11100_ (.Y(_02042_),
    .A(_01999_),
    .B(_01984_));
 sg13g2_nor2_1 _11101_ (.A(_02041_),
    .B(_02042_),
    .Y(_02043_));
 sg13g2_nand2_1 _11102_ (.Y(_02044_),
    .A(_02038_),
    .B(_02043_));
 sg13g2_nor2_1 _11103_ (.A(_01991_),
    .B(_01985_),
    .Y(_02045_));
 sg13g2_inv_1 _11104_ (.Y(_02046_),
    .A(_01969_));
 sg13g2_nand2_1 _11105_ (.Y(_02047_),
    .A(_02046_),
    .B(_01968_));
 sg13g2_inv_1 _11106_ (.Y(_02048_),
    .A(_01968_));
 sg13g2_nand2_1 _11107_ (.Y(_02049_),
    .A(_02048_),
    .B(_01969_));
 sg13g2_inv_1 _11108_ (.Y(_02050_),
    .A(_02049_));
 sg13g2_a21oi_1 _11109_ (.A1(_02047_),
    .A2(_01976_),
    .Y(_02051_),
    .B1(_02050_));
 sg13g2_inv_1 _11110_ (.Y(_02052_),
    .A(_01982_));
 sg13g2_nand2_1 _11111_ (.Y(_02053_),
    .A(_02052_),
    .B(_01981_));
 sg13g2_a21oi_1 _11112_ (.A1(_01997_),
    .A2(_02053_),
    .Y(_02054_),
    .B1(_01996_));
 sg13g2_a21oi_1 _11113_ (.A1(_02045_),
    .A2(_02051_),
    .Y(_02055_),
    .B1(_02054_));
 sg13g2_nand2_1 _11114_ (.Y(_02056_),
    .A(_02044_),
    .B(_02055_));
 sg13g2_xor2_1 _11115_ (.B(_01902_),
    .A(_01901_),
    .X(_02057_));
 sg13g2_inv_4 _11116_ (.A(_01909_),
    .Y(_02058_));
 sg13g2_nor2_1 _11117_ (.A(_02057_),
    .B(_02058_),
    .Y(_02059_));
 sg13g2_inv_8 _11118_ (.Y(_02060_),
    .A(_02010_));
 sg13g2_nor2_1 _11119_ (.A(_01893_),
    .B(_02060_),
    .Y(_02061_));
 sg13g2_nand2_1 _11120_ (.Y(_02062_),
    .A(_02059_),
    .B(_02061_));
 sg13g2_inv_2 _11121_ (.Y(_02063_),
    .A(_01936_));
 sg13g2_nand2_1 _11122_ (.Y(_02064_),
    .A(_02063_),
    .B(_01930_));
 sg13g2_nor2_1 _11123_ (.A(_01920_),
    .B(_01924_),
    .Y(_02065_));
 sg13g2_nor2b_1 _11124_ (.A(_02064_),
    .B_N(_02065_),
    .Y(_02066_));
 sg13g2_nor2b_1 _11125_ (.A(_02062_),
    .B_N(_02066_),
    .Y(_02067_));
 sg13g2_nand2_1 _11126_ (.Y(_02068_),
    .A(_02056_),
    .B(_02067_));
 sg13g2_inv_1 _11127_ (.Y(_02069_),
    .A(_02014_));
 sg13g2_inv_1 _11128_ (.Y(_02070_),
    .A(_01895_));
 sg13g2_nand2_1 _11129_ (.Y(_02071_),
    .A(_02070_),
    .B(_01894_));
 sg13g2_a21oi_1 _11130_ (.A1(_02069_),
    .A2(_02071_),
    .Y(_02072_),
    .B1(_02012_));
 sg13g2_nand2_1 _11131_ (.Y(_02073_),
    .A(_02059_),
    .B(_02072_));
 sg13g2_inv_1 _11132_ (.Y(_02074_),
    .A(_01901_));
 sg13g2_nor2_1 _11133_ (.A(_01902_),
    .B(_02074_),
    .Y(_02075_));
 sg13g2_nand2_1 _11134_ (.Y(_02076_),
    .A(_01905_),
    .B(\vgadonut.donut.donuthit.cordicxy.yin[10] ));
 sg13g2_inv_1 _11135_ (.Y(_02077_),
    .A(_02076_));
 sg13g2_a21oi_1 _11136_ (.A1(_01909_),
    .A2(_02075_),
    .Y(_02078_),
    .B1(_02077_));
 sg13g2_nand2_1 _11137_ (.Y(_02079_),
    .A(_02073_),
    .B(_02078_));
 sg13g2_inv_1 _11138_ (.Y(_02080_),
    .A(_02064_));
 sg13g2_inv_1 _11139_ (.Y(_02081_),
    .A(_01918_));
 sg13g2_nand2_1 _11140_ (.Y(_02082_),
    .A(_02081_),
    .B(_01917_));
 sg13g2_inv_1 _11141_ (.Y(_02083_),
    .A(_01922_));
 sg13g2_nand2_1 _11142_ (.Y(_02084_),
    .A(_02083_),
    .B(_01921_));
 sg13g2_nor2_1 _11143_ (.A(_01917_),
    .B(_02081_),
    .Y(_02085_));
 sg13g2_a21oi_1 _11144_ (.A1(_02082_),
    .A2(_02084_),
    .Y(_02086_),
    .B1(_02085_));
 sg13g2_nand2_1 _11145_ (.Y(_02087_),
    .A(_02080_),
    .B(_02086_));
 sg13g2_nor2b_1 _11146_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[14] ),
    .B_N(\vgadonut.donut.donuthit.cordicxy.yin[14] ),
    .Y(_02088_));
 sg13g2_a21oi_1 _11147_ (.A1(_02063_),
    .A2(_01927_),
    .Y(_02089_),
    .B1(_02088_));
 sg13g2_nand2_1 _11148_ (.Y(_02090_),
    .A(_02087_),
    .B(_02089_));
 sg13g2_a21oi_1 _11149_ (.A1(_02079_),
    .A2(_02066_),
    .Y(_02091_),
    .B1(_02090_));
 sg13g2_nand3_1 _11150_ (.B(net187),
    .C(_02091_),
    .A(_02068_),
    .Y(_02092_));
 sg13g2_buf_8 _11151_ (.A(_02092_),
    .X(_02093_));
 sg13g2_nand2_1 _11152_ (.Y(_02094_),
    .A(_02025_),
    .B(_02093_));
 sg13g2_buf_8 _11153_ (.A(_02094_),
    .X(_02095_));
 sg13g2_buf_8 _11154_ (.A(_02020_),
    .X(_02096_));
 sg13g2_nand2_1 _11155_ (.Y(_02097_),
    .A(_02095_),
    .B(net214));
 sg13g2_inv_4 _11156_ (.A(_02020_),
    .Y(_02098_));
 sg13g2_nand3_1 _11157_ (.B(_02098_),
    .C(_02093_),
    .A(_02025_),
    .Y(_02099_));
 sg13g2_nand2_1 _11158_ (.Y(_02100_),
    .A(_02097_),
    .B(_02099_));
 sg13g2_buf_8 _11159_ (.A(_02100_),
    .X(_02101_));
 sg13g2_nor2_1 _11160_ (.A(_01903_),
    .B(_02015_),
    .Y(_02102_));
 sg13g2_nor2_1 _11161_ (.A(_01894_),
    .B(_01895_),
    .Y(_02103_));
 sg13g2_a21oi_1 _11162_ (.A1(_01989_),
    .A2(_01896_),
    .Y(_02104_),
    .B1(_02103_));
 sg13g2_nand2_1 _11163_ (.Y(_02105_),
    .A(_02102_),
    .B(_02104_));
 sg13g2_nand2_1 _11164_ (.Y(_02106_),
    .A(_01912_),
    .B(_01899_));
 sg13g2_o21ai_1 _11165_ (.B1(_02106_),
    .Y(_02107_),
    .A1(_01901_),
    .A2(_01902_));
 sg13g2_nand2_1 _11166_ (.Y(_02108_),
    .A(_02105_),
    .B(_02107_));
 sg13g2_nor2_1 _11167_ (.A(_01975_),
    .B(_01973_),
    .Y(_02109_));
 sg13g2_o21ai_1 _11168_ (.B1(_02001_),
    .Y(_02110_),
    .A1(_01964_),
    .A2(_02109_));
 sg13g2_nor2_1 _11169_ (.A(_01984_),
    .B(_01971_),
    .Y(_02111_));
 sg13g2_nor2_1 _11170_ (.A(_01981_),
    .B(_01982_),
    .Y(_02112_));
 sg13g2_a21oi_1 _11171_ (.A1(_02005_),
    .A2(_02003_),
    .Y(_02113_),
    .B1(_02112_));
 sg13g2_a21oi_1 _11172_ (.A1(_02110_),
    .A2(_02111_),
    .Y(_02114_),
    .B1(_02113_));
 sg13g2_o21ai_1 _11173_ (.B1(_01952_),
    .Y(_02115_),
    .A1(_01960_),
    .A2(_01951_));
 sg13g2_buf_1 _11174_ (.A(_02115_),
    .X(_02116_));
 sg13g2_nor2_1 _11175_ (.A(_02028_),
    .B(_02040_),
    .Y(_02117_));
 sg13g2_nand3_1 _11176_ (.B(_02116_),
    .C(_02117_),
    .A(_02111_),
    .Y(_02118_));
 sg13g2_nand2_1 _11177_ (.Y(_02119_),
    .A(_02114_),
    .B(_02118_));
 sg13g2_inv_1 _11178_ (.Y(_02120_),
    .A(_02102_));
 sg13g2_nor2_1 _11179_ (.A(_02010_),
    .B(_01999_),
    .Y(_02121_));
 sg13g2_inv_1 _11180_ (.Y(_02122_),
    .A(_02121_));
 sg13g2_nor2_1 _11181_ (.A(_02120_),
    .B(_02122_),
    .Y(_02123_));
 sg13g2_nand2_1 _11182_ (.Y(_02124_),
    .A(_02119_),
    .B(_02123_));
 sg13g2_nand2b_1 _11183_ (.Y(_02125_),
    .B(_02124_),
    .A_N(_02108_));
 sg13g2_xnor2_1 _11184_ (.Y(_02126_),
    .A(_01909_),
    .B(_02125_));
 sg13g2_buf_1 _11185_ (.A(net187),
    .X(_02127_));
 sg13g2_buf_1 _11186_ (.A(net179),
    .X(_02128_));
 sg13g2_nand2_1 _11187_ (.Y(_02129_),
    .A(_02126_),
    .B(net176));
 sg13g2_nor2_1 _11188_ (.A(_01981_),
    .B(_02052_),
    .Y(_02130_));
 sg13g2_a21oi_1 _11189_ (.A1(_02053_),
    .A2(_02047_),
    .Y(_02131_),
    .B1(_02130_));
 sg13g2_nand2_1 _11190_ (.Y(_02132_),
    .A(_01971_),
    .B(_01984_));
 sg13g2_inv_1 _11191_ (.Y(_02133_),
    .A(_01976_));
 sg13g2_a21oi_1 _11192_ (.A1(_02036_),
    .A2(_01978_),
    .Y(_02134_),
    .B1(_02133_));
 sg13g2_nor2_1 _11193_ (.A(_02132_),
    .B(_02134_),
    .Y(_02135_));
 sg13g2_nor2_1 _11194_ (.A(_02131_),
    .B(_02135_),
    .Y(_02136_));
 sg13g2_nand2_1 _11195_ (.Y(_02137_),
    .A(_02028_),
    .B(_02040_));
 sg13g2_nor2_1 _11196_ (.A(_02132_),
    .B(_02137_),
    .Y(_02138_));
 sg13g2_nand2_1 _11197_ (.Y(_02139_),
    .A(_02032_),
    .B(_01950_));
 sg13g2_a21oi_1 _11198_ (.A1(_02139_),
    .A2(_02030_),
    .Y(_02140_),
    .B1(_02033_));
 sg13g2_inv_1 _11199_ (.Y(_02141_),
    .A(_02140_));
 sg13g2_nand2_1 _11200_ (.Y(_02142_),
    .A(_02138_),
    .B(_02141_));
 sg13g2_nand2_1 _11201_ (.Y(_02143_),
    .A(_02136_),
    .B(_02142_));
 sg13g2_nor2_1 _11202_ (.A(_01893_),
    .B(_02057_),
    .Y(_02144_));
 sg13g2_inv_1 _11203_ (.Y(_02145_),
    .A(_02144_));
 sg13g2_nor2_1 _11204_ (.A(_01991_),
    .B(_02060_),
    .Y(_02146_));
 sg13g2_inv_1 _11205_ (.Y(_02147_),
    .A(_02146_));
 sg13g2_nor2_1 _11206_ (.A(_02145_),
    .B(_02147_),
    .Y(_02148_));
 sg13g2_nand2_1 _11207_ (.Y(_02149_),
    .A(_02143_),
    .B(_02148_));
 sg13g2_nor2_1 _11208_ (.A(_01894_),
    .B(_02070_),
    .Y(_02150_));
 sg13g2_a21oi_1 _11209_ (.A1(_01997_),
    .A2(_02071_),
    .Y(_02151_),
    .B1(_02150_));
 sg13g2_nor2_1 _11210_ (.A(_02014_),
    .B(_02075_),
    .Y(_02152_));
 sg13g2_a21oi_1 _11211_ (.A1(_02074_),
    .A2(_01902_),
    .Y(_02153_),
    .B1(_02152_));
 sg13g2_a21oi_1 _11212_ (.A1(_02144_),
    .A2(_02151_),
    .Y(_02154_),
    .B1(_02153_));
 sg13g2_nand2_1 _11213_ (.Y(_02155_),
    .A(_02149_),
    .B(_02154_));
 sg13g2_xnor2_1 _11214_ (.Y(_02156_),
    .A(_02058_),
    .B(_02155_));
 sg13g2_buf_1 _11215_ (.A(_02023_),
    .X(_02157_));
 sg13g2_nand2_1 _11216_ (.Y(_02158_),
    .A(_02156_),
    .B(net175));
 sg13g2_nand2_1 _11217_ (.Y(_02159_),
    .A(_02129_),
    .B(_02158_));
 sg13g2_nand2_1 _11218_ (.Y(_02160_),
    .A(_02101_),
    .B(_02159_));
 sg13g2_nand2_1 _11219_ (.Y(_02161_),
    .A(_01948_),
    .B(_02019_));
 sg13g2_nand2_1 _11220_ (.Y(_02162_),
    .A(_02161_),
    .B(_02023_));
 sg13g2_nand2_1 _11221_ (.Y(_02163_),
    .A(_02068_),
    .B(_02091_));
 sg13g2_nand2_1 _11222_ (.Y(_02164_),
    .A(_02163_),
    .B(net187));
 sg13g2_nand3_1 _11223_ (.B(_02164_),
    .C(_02098_),
    .A(_02162_),
    .Y(_02165_));
 sg13g2_nand3_1 _11224_ (.B(_02020_),
    .C(_02093_),
    .A(_02025_),
    .Y(_02166_));
 sg13g2_nand2_1 _11225_ (.Y(_02167_),
    .A(_02165_),
    .B(_02166_));
 sg13g2_buf_2 _11226_ (.A(_02167_),
    .X(_02168_));
 sg13g2_xnor2_1 _11227_ (.Y(_02169_),
    .A(_02058_),
    .B(_02125_));
 sg13g2_nand2_1 _11228_ (.Y(_02170_),
    .A(_02169_),
    .B(net176));
 sg13g2_xnor2_1 _11229_ (.Y(_02171_),
    .A(_01909_),
    .B(_02155_));
 sg13g2_buf_1 _11230_ (.A(net175),
    .X(_02172_));
 sg13g2_nand2_1 _11231_ (.Y(_02173_),
    .A(_02171_),
    .B(net173));
 sg13g2_nand2_1 _11232_ (.Y(_02174_),
    .A(_02170_),
    .B(_02173_));
 sg13g2_nand2_1 _11233_ (.Y(_02175_),
    .A(_02168_),
    .B(_02174_));
 sg13g2_nand2_1 _11234_ (.Y(_02176_),
    .A(_02160_),
    .B(_02175_));
 sg13g2_buf_1 _11235_ (.A(net179),
    .X(_02177_));
 sg13g2_nand2_1 _11236_ (.Y(_02178_),
    .A(_02016_),
    .B(_02006_));
 sg13g2_nand2b_1 _11237_ (.Y(_02179_),
    .B(_02178_),
    .A_N(_01900_));
 sg13g2_nor2_1 _11238_ (.A(_01971_),
    .B(_02040_),
    .Y(_02180_));
 sg13g2_a21oi_1 _11239_ (.A1(_01965_),
    .A2(_02180_),
    .Y(_02181_),
    .B1(_02004_));
 sg13g2_nor2b_1 _11240_ (.A(_01992_),
    .B_N(_02016_),
    .Y(_02182_));
 sg13g2_nor2b_1 _11241_ (.A(_02181_),
    .B_N(_02182_),
    .Y(_02183_));
 sg13g2_nor2_1 _11242_ (.A(_02179_),
    .B(_02183_),
    .Y(_02184_));
 sg13g2_nand2_1 _11243_ (.Y(_02185_),
    .A(_01954_),
    .B(_01957_));
 sg13g2_nor2_1 _11244_ (.A(_02185_),
    .B(_01980_),
    .Y(_02186_));
 sg13g2_nand3_1 _11245_ (.B(_01961_),
    .C(_02186_),
    .A(_02182_),
    .Y(_02187_));
 sg13g2_nand2_1 _11246_ (.Y(_02188_),
    .A(_02184_),
    .B(_02187_));
 sg13g2_nand2_1 _11247_ (.Y(_02189_),
    .A(_02188_),
    .B(_02057_));
 sg13g2_nand3_1 _11248_ (.B(_01903_),
    .C(_02187_),
    .A(_02184_),
    .Y(_02190_));
 sg13g2_nand2_1 _11249_ (.Y(_02191_),
    .A(_02189_),
    .B(_02190_));
 sg13g2_nand2b_1 _11250_ (.Y(_02192_),
    .B(_02038_),
    .A_N(_02041_));
 sg13g2_inv_1 _11251_ (.Y(_02193_),
    .A(_02051_));
 sg13g2_nand2_1 _11252_ (.Y(_02194_),
    .A(_02192_),
    .B(_02193_));
 sg13g2_nand2_1 _11253_ (.Y(_02195_),
    .A(_02045_),
    .B(_02061_));
 sg13g2_inv_1 _11254_ (.Y(_02196_),
    .A(_02195_));
 sg13g2_nand2_1 _11255_ (.Y(_02197_),
    .A(_02194_),
    .B(_02196_));
 sg13g2_a21oi_1 _11256_ (.A1(_02061_),
    .A2(_02054_),
    .Y(_02198_),
    .B1(_02072_));
 sg13g2_nand2_1 _11257_ (.Y(_02199_),
    .A(_02197_),
    .B(_02198_));
 sg13g2_nand2_1 _11258_ (.Y(_02200_),
    .A(_02199_),
    .B(_01903_));
 sg13g2_nand3_1 _11259_ (.B(_02057_),
    .C(_02198_),
    .A(_02197_),
    .Y(_02201_));
 sg13g2_buf_1 _11260_ (.A(_02201_),
    .X(_02202_));
 sg13g2_nand3_1 _11261_ (.B(_02202_),
    .C(net176),
    .A(_02200_),
    .Y(_02203_));
 sg13g2_o21ai_1 _11262_ (.B1(_02203_),
    .Y(_02204_),
    .A1(net174),
    .A2(_02191_));
 sg13g2_buf_1 _11263_ (.A(_02204_),
    .X(_02205_));
 sg13g2_inv_1 _11264_ (.Y(_02206_),
    .A(_02205_));
 sg13g2_nand2_1 _11265_ (.Y(_02207_),
    .A(_02176_),
    .B(_02206_));
 sg13g2_nand3_1 _11266_ (.B(_02175_),
    .C(_02205_),
    .A(_02160_),
    .Y(_02208_));
 sg13g2_buf_1 _11267_ (.A(_02208_),
    .X(_02209_));
 sg13g2_nand2_2 _11268_ (.Y(_02210_),
    .A(_02207_),
    .B(_02209_));
 sg13g2_inv_1 _11269_ (.Y(_02211_),
    .A(_02062_));
 sg13g2_nand2_1 _11270_ (.Y(_02212_),
    .A(_02056_),
    .B(_02211_));
 sg13g2_inv_1 _11271_ (.Y(_02213_),
    .A(_02079_));
 sg13g2_nand2_1 _11272_ (.Y(_02214_),
    .A(_02212_),
    .B(_02213_));
 sg13g2_xnor2_1 _11273_ (.Y(_02215_),
    .A(_01921_),
    .B(_01922_));
 sg13g2_nand2_1 _11274_ (.Y(_02216_),
    .A(_02214_),
    .B(_02215_));
 sg13g2_nand3_1 _11275_ (.B(_01924_),
    .C(_02213_),
    .A(_02212_),
    .Y(_02217_));
 sg13g2_nand2_1 _11276_ (.Y(_02218_),
    .A(_02216_),
    .B(_02217_));
 sg13g2_nand2_1 _11277_ (.Y(_02219_),
    .A(_02218_),
    .B(net173));
 sg13g2_inv_1 _11278_ (.Y(_02220_),
    .A(_02017_));
 sg13g2_nand2_1 _11279_ (.Y(_02221_),
    .A(_02008_),
    .B(_02220_));
 sg13g2_inv_1 _11280_ (.Y(_02222_),
    .A(_01916_));
 sg13g2_nand2_1 _11281_ (.Y(_02223_),
    .A(_02221_),
    .B(_02222_));
 sg13g2_nand2_1 _11282_ (.Y(_02224_),
    .A(_02223_),
    .B(_02215_));
 sg13g2_nand3_1 _11283_ (.B(_01924_),
    .C(_02222_),
    .A(_02221_),
    .Y(_02225_));
 sg13g2_nand3_1 _11284_ (.B(_02225_),
    .C(net176),
    .A(_02224_),
    .Y(_02226_));
 sg13g2_nand2_1 _11285_ (.Y(_02227_),
    .A(_02219_),
    .B(_02226_));
 sg13g2_nand2_1 _11286_ (.Y(_02228_),
    .A(_02168_),
    .B(_02227_));
 sg13g2_nand2_1 _11287_ (.Y(_02229_),
    .A(_02223_),
    .B(_01924_));
 sg13g2_nand3_1 _11288_ (.B(_02215_),
    .C(_02222_),
    .A(_02221_),
    .Y(_02230_));
 sg13g2_nand3_1 _11289_ (.B(_02230_),
    .C(net179),
    .A(_02229_),
    .Y(_02231_));
 sg13g2_nand3_1 _11290_ (.B(_02217_),
    .C(net175),
    .A(_02216_),
    .Y(_02232_));
 sg13g2_nand2_1 _11291_ (.Y(_02233_),
    .A(_02231_),
    .B(_02232_));
 sg13g2_nand2_1 _11292_ (.Y(_02234_),
    .A(_02101_),
    .B(_02233_));
 sg13g2_nand2_1 _11293_ (.Y(_02235_),
    .A(_02228_),
    .B(_02234_));
 sg13g2_buf_1 _11294_ (.A(net175),
    .X(_02236_));
 sg13g2_buf_1 _11295_ (.A(net172),
    .X(_02237_));
 sg13g2_nor2_1 _11296_ (.A(net172),
    .B(_02156_),
    .Y(_02238_));
 sg13g2_a21oi_2 _11297_ (.B1(_02238_),
    .Y(_02239_),
    .A2(_02169_),
    .A1(_02237_));
 sg13g2_inv_1 _11298_ (.Y(_02240_),
    .A(_02239_));
 sg13g2_nand2_1 _11299_ (.Y(_02241_),
    .A(_02235_),
    .B(_02240_));
 sg13g2_nand3_1 _11300_ (.B(_02234_),
    .C(_02239_),
    .A(_02228_),
    .Y(_02242_));
 sg13g2_nand2_2 _11301_ (.Y(_02243_),
    .A(_02241_),
    .B(_02242_));
 sg13g2_nor2_1 _11302_ (.A(_02210_),
    .B(_02243_),
    .Y(_02244_));
 sg13g2_nand2_1 _11303_ (.Y(_02245_),
    .A(_02056_),
    .B(_02010_));
 sg13g2_nand3_1 _11304_ (.B(_02060_),
    .C(_02055_),
    .A(_02044_),
    .Y(_02246_));
 sg13g2_nand2_1 _11305_ (.Y(_02247_),
    .A(_02245_),
    .B(_02246_));
 sg13g2_inv_1 _11306_ (.Y(_02248_),
    .A(_02247_));
 sg13g2_nand2_1 _11307_ (.Y(_02249_),
    .A(_02008_),
    .B(_02010_));
 sg13g2_nand3_1 _11308_ (.B(_02007_),
    .C(_02060_),
    .A(_01994_),
    .Y(_02250_));
 sg13g2_a21oi_1 _11309_ (.A1(_02249_),
    .A2(_02250_),
    .Y(_02251_),
    .B1(net176));
 sg13g2_a21o_1 _11310_ (.A2(_02248_),
    .A1(net174),
    .B1(_02251_),
    .X(_02252_));
 sg13g2_buf_1 _11311_ (.A(_02252_),
    .X(_02253_));
 sg13g2_inv_1 _11312_ (.Y(_02254_),
    .A(_02253_));
 sg13g2_o21ai_1 _11313_ (.B1(_02134_),
    .Y(_02255_),
    .A1(_02137_),
    .A2(_02140_));
 sg13g2_nor2_1 _11314_ (.A(_02132_),
    .B(_02147_),
    .Y(_02256_));
 sg13g2_nand2_1 _11315_ (.Y(_02257_),
    .A(_02146_),
    .B(_02131_));
 sg13g2_nand2b_1 _11316_ (.Y(_02258_),
    .B(_02257_),
    .A_N(_02151_));
 sg13g2_a21oi_1 _11317_ (.A1(_02255_),
    .A2(_02256_),
    .Y(_02259_),
    .B1(_02258_));
 sg13g2_xnor2_1 _11318_ (.Y(_02260_),
    .A(_01893_),
    .B(_02259_));
 sg13g2_nand2_1 _11319_ (.Y(_02261_),
    .A(_02116_),
    .B(_02117_));
 sg13g2_inv_1 _11320_ (.Y(_02262_),
    .A(_02110_));
 sg13g2_nand2_1 _11321_ (.Y(_02263_),
    .A(_02261_),
    .B(_02262_));
 sg13g2_nor2b_1 _11322_ (.A(_02122_),
    .B_N(_02111_),
    .Y(_02264_));
 sg13g2_nand2_1 _11323_ (.Y(_02265_),
    .A(_02263_),
    .B(_02264_));
 sg13g2_a21oi_1 _11324_ (.A1(_02121_),
    .A2(_02113_),
    .Y(_02266_),
    .B1(_02104_));
 sg13g2_nand2_1 _11325_ (.Y(_02267_),
    .A(_02265_),
    .B(_02266_));
 sg13g2_nor2_1 _11326_ (.A(_01893_),
    .B(_02267_),
    .Y(_02268_));
 sg13g2_inv_1 _11327_ (.Y(_02269_),
    .A(_02268_));
 sg13g2_nand2_1 _11328_ (.Y(_02270_),
    .A(_02267_),
    .B(_01893_));
 sg13g2_nand3_1 _11329_ (.B(net179),
    .C(_02270_),
    .A(_02269_),
    .Y(_02271_));
 sg13g2_o21ai_1 _11330_ (.B1(_02271_),
    .Y(_02272_),
    .A1(net179),
    .A2(_02260_));
 sg13g2_buf_1 _11331_ (.A(_02272_),
    .X(_02273_));
 sg13g2_nand2_1 _11332_ (.Y(_02274_),
    .A(_02101_),
    .B(_02273_));
 sg13g2_inv_1 _11333_ (.Y(_02275_),
    .A(_02273_));
 sg13g2_nand2_1 _11334_ (.Y(_02276_),
    .A(_02168_),
    .B(_02275_));
 sg13g2_nand2_1 _11335_ (.Y(_02277_),
    .A(_02274_),
    .B(_02276_));
 sg13g2_nor2_1 _11336_ (.A(_02254_),
    .B(_02277_),
    .Y(_02278_));
 sg13g2_nand2_1 _11337_ (.Y(_02279_),
    .A(_02200_),
    .B(_02202_));
 sg13g2_nand2_1 _11338_ (.Y(_02280_),
    .A(_02279_),
    .B(net173));
 sg13g2_nand2_1 _11339_ (.Y(_02281_),
    .A(_02191_),
    .B(net174));
 sg13g2_nand2_1 _11340_ (.Y(_02282_),
    .A(_02280_),
    .B(_02281_));
 sg13g2_nand2_1 _11341_ (.Y(_02283_),
    .A(_02101_),
    .B(_02282_));
 sg13g2_nand3_1 _11342_ (.B(_02202_),
    .C(net175),
    .A(_02200_),
    .Y(_02284_));
 sg13g2_nand3_1 _11343_ (.B(_02190_),
    .C(net179),
    .A(_02189_),
    .Y(_02285_));
 sg13g2_nand2_1 _11344_ (.Y(_02286_),
    .A(_02284_),
    .B(_02285_));
 sg13g2_nand2_1 _11345_ (.Y(_02287_),
    .A(_02168_),
    .B(_02286_));
 sg13g2_nand3_1 _11346_ (.B(net173),
    .C(_02270_),
    .A(_02269_),
    .Y(_02288_));
 sg13g2_o21ai_1 _11347_ (.B1(_02288_),
    .Y(_02289_),
    .A1(net173),
    .A2(_02260_));
 sg13g2_buf_1 _11348_ (.A(_02289_),
    .X(_02290_));
 sg13g2_inv_1 _11349_ (.Y(_02291_),
    .A(_02290_));
 sg13g2_nand3_1 _11350_ (.B(_02287_),
    .C(_02291_),
    .A(_02283_),
    .Y(_02292_));
 sg13g2_nand2_1 _11351_ (.Y(_02293_),
    .A(_02278_),
    .B(_02292_));
 sg13g2_nand2_1 _11352_ (.Y(_02294_),
    .A(_02283_),
    .B(_02287_));
 sg13g2_nand2_1 _11353_ (.Y(_02295_),
    .A(_02294_),
    .B(_02290_));
 sg13g2_nand2_1 _11354_ (.Y(_02296_),
    .A(_02293_),
    .B(_02295_));
 sg13g2_nand2_1 _11355_ (.Y(_02297_),
    .A(_02244_),
    .B(_02296_));
 sg13g2_inv_1 _11356_ (.Y(_02298_),
    .A(_02209_));
 sg13g2_inv_1 _11357_ (.Y(_02299_),
    .A(_02242_));
 sg13g2_a21oi_1 _11358_ (.A1(_02298_),
    .A2(_02241_),
    .Y(_02300_),
    .B1(_02299_));
 sg13g2_nand2_1 _11359_ (.Y(_02301_),
    .A(_02297_),
    .B(_02300_));
 sg13g2_nor2_1 _11360_ (.A(_01924_),
    .B(_02058_),
    .Y(_02302_));
 sg13g2_nor2b_1 _11361_ (.A(_02145_),
    .B_N(_02302_),
    .Y(_02303_));
 sg13g2_o21ai_1 _11362_ (.B1(_02084_),
    .Y(_02304_),
    .A1(_02076_),
    .A2(_01924_));
 sg13g2_nand2_1 _11363_ (.Y(_02305_),
    .A(_02153_),
    .B(_02302_));
 sg13g2_nand2b_1 _11364_ (.Y(_02306_),
    .B(_02305_),
    .A_N(_02304_));
 sg13g2_a21oi_1 _11365_ (.A1(_02303_),
    .A2(_02258_),
    .Y(_02307_),
    .B1(_02306_));
 sg13g2_nand3_1 _11366_ (.B(_02303_),
    .C(_02256_),
    .A(_02255_),
    .Y(_02308_));
 sg13g2_nand2_1 _11367_ (.Y(_02309_),
    .A(_02307_),
    .B(_02308_));
 sg13g2_inv_1 _11368_ (.Y(_02310_),
    .A(_01920_));
 sg13g2_nand2_1 _11369_ (.Y(_02311_),
    .A(_02309_),
    .B(_02310_));
 sg13g2_nand3_1 _11370_ (.B(_01920_),
    .C(_02308_),
    .A(_02307_),
    .Y(_02312_));
 sg13g2_nand3_1 _11371_ (.B(_02312_),
    .C(net174),
    .A(_02311_),
    .Y(_02313_));
 sg13g2_nand2_1 _11372_ (.Y(_02314_),
    .A(_02058_),
    .B(_01924_));
 sg13g2_o21ai_1 _11373_ (.B1(_01939_),
    .Y(_02315_),
    .A1(_01907_),
    .A2(_02215_));
 sg13g2_inv_1 _11374_ (.Y(_02316_),
    .A(_02315_));
 sg13g2_o21ai_1 _11375_ (.B1(_02316_),
    .Y(_02317_),
    .A1(_02314_),
    .A2(_02107_));
 sg13g2_nor2_1 _11376_ (.A(_02314_),
    .B(_02120_),
    .Y(_02318_));
 sg13g2_nor2b_1 _11377_ (.A(_02266_),
    .B_N(_02318_),
    .Y(_02319_));
 sg13g2_nor2_1 _11378_ (.A(_02317_),
    .B(_02319_),
    .Y(_02320_));
 sg13g2_nand3_1 _11379_ (.B(_02318_),
    .C(_02264_),
    .A(_02263_),
    .Y(_02321_));
 sg13g2_nand2_1 _11380_ (.Y(_02322_),
    .A(_02320_),
    .B(_02321_));
 sg13g2_nand2_1 _11381_ (.Y(_02323_),
    .A(_02322_),
    .B(_01920_));
 sg13g2_nand3_1 _11382_ (.B(_02310_),
    .C(_02321_),
    .A(_02320_),
    .Y(_02324_));
 sg13g2_nand3_1 _11383_ (.B(_02324_),
    .C(net172),
    .A(_02323_),
    .Y(_02325_));
 sg13g2_nand2_1 _11384_ (.Y(_02326_),
    .A(_02313_),
    .B(_02325_));
 sg13g2_inv_1 _11385_ (.Y(_02327_),
    .A(_02326_));
 sg13g2_buf_8 _11386_ (.A(_02168_),
    .X(_02328_));
 sg13g2_nand2_1 _11387_ (.Y(_02329_),
    .A(_02186_),
    .B(_01961_));
 sg13g2_nand2_1 _11388_ (.Y(_02330_),
    .A(_02181_),
    .B(_02329_));
 sg13g2_nor2b_1 _11389_ (.A(_01925_),
    .B_N(_01910_),
    .Y(_02331_));
 sg13g2_nand3_1 _11390_ (.B(_02331_),
    .C(_02182_),
    .A(_02330_),
    .Y(_02332_));
 sg13g2_o21ai_1 _11391_ (.B1(_01943_),
    .Y(_02333_),
    .A1(_01925_),
    .A2(_01915_));
 sg13g2_a21oi_1 _11392_ (.A1(_02179_),
    .A2(_02331_),
    .Y(_02334_),
    .B1(_02333_));
 sg13g2_nand2_1 _11393_ (.Y(_02335_),
    .A(_02332_),
    .B(_02334_));
 sg13g2_nand2_1 _11394_ (.Y(_02336_),
    .A(_02335_),
    .B(_01931_));
 sg13g2_nand3_1 _11395_ (.B(_01930_),
    .C(_02334_),
    .A(_02332_),
    .Y(_02337_));
 sg13g2_nand3_1 _11396_ (.B(_02337_),
    .C(net174),
    .A(_02336_),
    .Y(_02338_));
 sg13g2_nand2_1 _11397_ (.Y(_02339_),
    .A(_02059_),
    .B(_02065_));
 sg13g2_nor2_1 _11398_ (.A(_02339_),
    .B(_02198_),
    .Y(_02340_));
 sg13g2_nor2b_1 _11399_ (.A(_02078_),
    .B_N(_02065_),
    .Y(_02341_));
 sg13g2_nor2_1 _11400_ (.A(_02086_),
    .B(_02341_),
    .Y(_02342_));
 sg13g2_nor2b_1 _11401_ (.A(_02340_),
    .B_N(_02342_),
    .Y(_02343_));
 sg13g2_nor2_1 _11402_ (.A(_02195_),
    .B(_02339_),
    .Y(_02344_));
 sg13g2_nand2_1 _11403_ (.Y(_02345_),
    .A(_02194_),
    .B(_02344_));
 sg13g2_nand2_1 _11404_ (.Y(_02346_),
    .A(_02343_),
    .B(_02345_));
 sg13g2_nand2_1 _11405_ (.Y(_02347_),
    .A(_02346_),
    .B(_01930_));
 sg13g2_nand3_1 _11406_ (.B(_02345_),
    .C(_01931_),
    .A(_02343_),
    .Y(_02348_));
 sg13g2_nand3_1 _11407_ (.B(_02348_),
    .C(_02236_),
    .A(_02347_),
    .Y(_02349_));
 sg13g2_nand2_2 _11408_ (.Y(_02350_),
    .A(_02338_),
    .B(_02349_));
 sg13g2_xnor2_1 _11409_ (.Y(_02351_),
    .A(net102),
    .B(_02350_));
 sg13g2_xnor2_1 _11410_ (.Y(_02352_),
    .A(_02327_),
    .B(_02351_));
 sg13g2_nand3_1 _11411_ (.B(_02230_),
    .C(net172),
    .A(_02229_),
    .Y(_02353_));
 sg13g2_o21ai_1 _11412_ (.B1(_02353_),
    .Y(_02354_),
    .A1(net172),
    .A2(_02218_));
 sg13g2_buf_1 _11413_ (.A(_02354_),
    .X(_02355_));
 sg13g2_nand3_1 _11414_ (.B(_02312_),
    .C(net173),
    .A(_02311_),
    .Y(_02356_));
 sg13g2_nand3_1 _11415_ (.B(_02324_),
    .C(net176),
    .A(_02323_),
    .Y(_02357_));
 sg13g2_nand2_1 _11416_ (.Y(_02358_),
    .A(_02356_),
    .B(_02357_));
 sg13g2_xnor2_1 _11417_ (.Y(_02359_),
    .A(_02358_),
    .B(_02101_));
 sg13g2_xnor2_1 _11418_ (.Y(_02360_),
    .A(_02355_),
    .B(_02359_));
 sg13g2_nand2_1 _11419_ (.Y(_02361_),
    .A(_02352_),
    .B(_02360_));
 sg13g2_nor2_1 _11420_ (.A(_01920_),
    .B(_01931_),
    .Y(_02362_));
 sg13g2_nand2_1 _11421_ (.Y(_02363_),
    .A(_02362_),
    .B(_02302_));
 sg13g2_nand3b_1 _11422_ (.B(_02143_),
    .C(_02148_),
    .Y(_02364_),
    .A_N(_02363_));
 sg13g2_nand2_1 _11423_ (.Y(_02365_),
    .A(_02304_),
    .B(_02362_));
 sg13g2_nor2_1 _11424_ (.A(_02082_),
    .B(_01929_),
    .Y(_02366_));
 sg13g2_nor2_1 _11425_ (.A(_01927_),
    .B(_02366_),
    .Y(_02367_));
 sg13g2_nand2_1 _11426_ (.Y(_02368_),
    .A(_02365_),
    .B(_02367_));
 sg13g2_nor2_1 _11427_ (.A(_02363_),
    .B(_02154_),
    .Y(_02369_));
 sg13g2_nor2_1 _11428_ (.A(_02368_),
    .B(_02369_),
    .Y(_02370_));
 sg13g2_nand2_1 _11429_ (.Y(_02371_),
    .A(_02364_),
    .B(_02370_));
 sg13g2_nand2_1 _11430_ (.Y(_02372_),
    .A(_02371_),
    .B(_02063_));
 sg13g2_nand3_1 _11431_ (.B(_02370_),
    .C(_01936_),
    .A(_02364_),
    .Y(_02373_));
 sg13g2_buf_1 _11432_ (.A(net176),
    .X(_02374_));
 sg13g2_nand3_1 _11433_ (.B(_02373_),
    .C(_02374_),
    .A(_02372_),
    .Y(_02375_));
 sg13g2_nor2_1 _11434_ (.A(_01930_),
    .B(_02310_),
    .Y(_02376_));
 sg13g2_nor2b_1 _11435_ (.A(_02314_),
    .B_N(_02376_),
    .Y(_02377_));
 sg13g2_nand3_1 _11436_ (.B(_02377_),
    .C(_02123_),
    .A(_02119_),
    .Y(_02378_));
 sg13g2_nand2_1 _11437_ (.Y(_02379_),
    .A(_02315_),
    .B(_02376_));
 sg13g2_a21oi_1 _11438_ (.A1(_01931_),
    .A2(_01942_),
    .Y(_02380_),
    .B1(_01945_));
 sg13g2_nand2_1 _11439_ (.Y(_02381_),
    .A(_02379_),
    .B(_02380_));
 sg13g2_a21oi_1 _11440_ (.A1(_02108_),
    .A2(_02377_),
    .Y(_02382_),
    .B1(_02381_));
 sg13g2_nand2_1 _11441_ (.Y(_02383_),
    .A(_02378_),
    .B(_02382_));
 sg13g2_nand2_1 _11442_ (.Y(_02384_),
    .A(_02383_),
    .B(_01936_));
 sg13g2_nand3_1 _11443_ (.B(_02382_),
    .C(_02063_),
    .A(_02378_),
    .Y(_02385_));
 sg13g2_nand3_1 _11444_ (.B(_02385_),
    .C(_02237_),
    .A(_02384_),
    .Y(_02386_));
 sg13g2_nand2_1 _11445_ (.Y(_02387_),
    .A(_02375_),
    .B(_02386_));
 sg13g2_mux2_1 _11446_ (.A0(_02163_),
    .A1(_02161_),
    .S(_02127_),
    .X(_02388_));
 sg13g2_buf_1 _11447_ (.A(_02388_),
    .X(_02389_));
 sg13g2_nand2b_1 _11448_ (.Y(_02390_),
    .B(net102),
    .A_N(_02389_));
 sg13g2_buf_8 _11449_ (.A(_02101_),
    .X(_02391_));
 sg13g2_nand2_1 _11450_ (.Y(_02392_),
    .A(net83),
    .B(_02389_));
 sg13g2_nand2_1 _11451_ (.Y(_02393_),
    .A(_02390_),
    .B(_02392_));
 sg13g2_nand2b_1 _11452_ (.Y(_02394_),
    .B(_02393_),
    .A_N(_02387_));
 sg13g2_nand3_1 _11453_ (.B(_02392_),
    .C(_02387_),
    .A(_02390_),
    .Y(_02395_));
 sg13g2_nand2_2 _11454_ (.Y(_02396_),
    .A(_02394_),
    .B(_02395_));
 sg13g2_nand3_1 _11455_ (.B(_02373_),
    .C(net172),
    .A(_02372_),
    .Y(_02397_));
 sg13g2_nand3_1 _11456_ (.B(_02385_),
    .C(net174),
    .A(_02384_),
    .Y(_02398_));
 sg13g2_nand2_2 _11457_ (.Y(_02399_),
    .A(_02397_),
    .B(_02398_));
 sg13g2_xnor2_1 _11458_ (.Y(_02400_),
    .A(net102),
    .B(_02399_));
 sg13g2_nand3_1 _11459_ (.B(_02337_),
    .C(_02236_),
    .A(_02336_),
    .Y(_02401_));
 sg13g2_nand3_1 _11460_ (.B(_02348_),
    .C(net174),
    .A(_02347_),
    .Y(_02402_));
 sg13g2_nand2_1 _11461_ (.Y(_02403_),
    .A(_02401_),
    .B(_02402_));
 sg13g2_nand2_1 _11462_ (.Y(_02404_),
    .A(_02400_),
    .B(_02403_));
 sg13g2_xnor2_1 _11463_ (.Y(_02405_),
    .A(net83),
    .B(_02399_));
 sg13g2_inv_1 _11464_ (.Y(_02406_),
    .A(_02403_));
 sg13g2_nand2_1 _11465_ (.Y(_02407_),
    .A(_02405_),
    .B(_02406_));
 sg13g2_nand2_2 _11466_ (.Y(_02408_),
    .A(_02404_),
    .B(_02407_));
 sg13g2_inv_1 _11467_ (.Y(_02409_),
    .A(_02408_));
 sg13g2_nand2b_1 _11468_ (.Y(_02410_),
    .B(_02409_),
    .A_N(_02396_));
 sg13g2_nor2_1 _11469_ (.A(_02361_),
    .B(_02410_),
    .Y(_02411_));
 sg13g2_nor2_1 _11470_ (.A(_02396_),
    .B(_02408_),
    .Y(_02412_));
 sg13g2_xnor2_1 _11471_ (.Y(_02413_),
    .A(net83),
    .B(_02350_));
 sg13g2_nand2_1 _11472_ (.Y(_02414_),
    .A(_02413_),
    .B(_02327_));
 sg13g2_inv_1 _11473_ (.Y(_02415_),
    .A(_02355_));
 sg13g2_nor2_1 _11474_ (.A(_02415_),
    .B(_02359_),
    .Y(_02416_));
 sg13g2_nand2_1 _11475_ (.Y(_02417_),
    .A(_02414_),
    .B(_02416_));
 sg13g2_nand2_1 _11476_ (.Y(_02418_),
    .A(_02351_),
    .B(_02326_));
 sg13g2_nand2_1 _11477_ (.Y(_02419_),
    .A(_02417_),
    .B(_02418_));
 sg13g2_nand2_1 _11478_ (.Y(_02420_),
    .A(_02412_),
    .B(_02419_));
 sg13g2_inv_1 _11479_ (.Y(_02421_),
    .A(_02404_));
 sg13g2_inv_1 _11480_ (.Y(_02422_),
    .A(_02395_));
 sg13g2_a21oi_1 _11481_ (.A1(_02421_),
    .A2(_02394_),
    .Y(_02423_),
    .B1(_02422_));
 sg13g2_nand2_1 _11482_ (.Y(_02424_),
    .A(_02420_),
    .B(_02423_));
 sg13g2_a21oi_1 _11483_ (.A1(_02301_),
    .A2(_02411_),
    .Y(_02425_),
    .B1(_02424_));
 sg13g2_xnor2_1 _11484_ (.Y(_02426_),
    .A(_01999_),
    .B(_02119_));
 sg13g2_nand2_1 _11485_ (.Y(_02427_),
    .A(_02426_),
    .B(net187));
 sg13g2_nand2_1 _11486_ (.Y(_02428_),
    .A(_02143_),
    .B(_01991_));
 sg13g2_nand3_1 _11487_ (.B(_02142_),
    .C(_01999_),
    .A(_02136_),
    .Y(_02429_));
 sg13g2_nand2_1 _11488_ (.Y(_02430_),
    .A(_02428_),
    .B(_02429_));
 sg13g2_nand2_1 _11489_ (.Y(_02431_),
    .A(_02430_),
    .B(_02023_));
 sg13g2_nand2_1 _11490_ (.Y(_02432_),
    .A(_02427_),
    .B(_02431_));
 sg13g2_nand2_1 _11491_ (.Y(_02433_),
    .A(_02432_),
    .B(net214));
 sg13g2_nand3_1 _11492_ (.B(_02431_),
    .C(_02098_),
    .A(_02427_),
    .Y(_02434_));
 sg13g2_nand2_1 _11493_ (.Y(_02435_),
    .A(_02433_),
    .B(_02434_));
 sg13g2_buf_8 _11494_ (.A(_02095_),
    .X(_02436_));
 sg13g2_nand2_1 _11495_ (.Y(_02437_),
    .A(_02435_),
    .B(net103));
 sg13g2_inv_4 _11496_ (.A(_02095_),
    .Y(_02438_));
 sg13g2_nand3_1 _11497_ (.B(_02438_),
    .C(_02434_),
    .A(_02433_),
    .Y(_02439_));
 sg13g2_nand2_1 _11498_ (.Y(_02440_),
    .A(_02437_),
    .B(_02439_));
 sg13g2_nand2_1 _11499_ (.Y(_02441_),
    .A(_02194_),
    .B(_01984_));
 sg13g2_nand3_1 _11500_ (.B(_01985_),
    .C(_02193_),
    .A(_02192_),
    .Y(_02442_));
 sg13g2_and2_1 _11501_ (.A(_02441_),
    .B(_02442_),
    .X(_02443_));
 sg13g2_nand2_1 _11502_ (.Y(_02444_),
    .A(_02330_),
    .B(_01984_));
 sg13g2_nand3_1 _11503_ (.B(_02329_),
    .C(_01985_),
    .A(_02181_),
    .Y(_02445_));
 sg13g2_a21oi_1 _11504_ (.A1(_02444_),
    .A2(_02445_),
    .Y(_02446_),
    .B1(net176));
 sg13g2_a21o_1 _11505_ (.A2(net174),
    .A1(_02443_),
    .B1(_02446_),
    .X(_02447_));
 sg13g2_buf_1 _11506_ (.A(_02447_),
    .X(_02448_));
 sg13g2_inv_1 _11507_ (.Y(_02449_),
    .A(_02448_));
 sg13g2_nand2_1 _11508_ (.Y(_02450_),
    .A(_02440_),
    .B(_02449_));
 sg13g2_nand3_1 _11509_ (.B(_02439_),
    .C(_02448_),
    .A(_02437_),
    .Y(_02451_));
 sg13g2_buf_1 _11510_ (.A(_02451_),
    .X(_02452_));
 sg13g2_nand2_1 _11511_ (.Y(_02453_),
    .A(_02450_),
    .B(_02452_));
 sg13g2_nand2_1 _11512_ (.Y(_02454_),
    .A(_02008_),
    .B(_02060_));
 sg13g2_nand3_1 _11513_ (.B(_02007_),
    .C(_02010_),
    .A(_01994_),
    .Y(_02455_));
 sg13g2_nand3_1 _11514_ (.B(_02455_),
    .C(_02022_),
    .A(_02454_),
    .Y(_02456_));
 sg13g2_buf_1 _11515_ (.A(_02456_),
    .X(_02457_));
 sg13g2_nand3_1 _11516_ (.B(_02246_),
    .C(net175),
    .A(_02245_),
    .Y(_02458_));
 sg13g2_buf_1 _11517_ (.A(_02458_),
    .X(_02459_));
 sg13g2_nand2_1 _11518_ (.Y(_02460_),
    .A(_02457_),
    .B(_02459_));
 sg13g2_buf_8 _11519_ (.A(_02098_),
    .X(_02461_));
 sg13g2_nand2_1 _11520_ (.Y(_02462_),
    .A(_02460_),
    .B(net186));
 sg13g2_nand3_1 _11521_ (.B(_02459_),
    .C(net214),
    .A(_02457_),
    .Y(_02463_));
 sg13g2_nand3_1 _11522_ (.B(_02463_),
    .C(_02095_),
    .A(_02462_),
    .Y(_02464_));
 sg13g2_nand3_1 _11523_ (.B(_02459_),
    .C(net186),
    .A(_02457_),
    .Y(_02465_));
 sg13g2_nand3_1 _11524_ (.B(_02250_),
    .C(_02128_),
    .A(_02249_),
    .Y(_02466_));
 sg13g2_nand2_1 _11525_ (.Y(_02467_),
    .A(_02056_),
    .B(_02060_));
 sg13g2_nand3_1 _11526_ (.B(_02010_),
    .C(_02055_),
    .A(_02044_),
    .Y(_02468_));
 sg13g2_nand3_1 _11527_ (.B(_02468_),
    .C(net175),
    .A(_02467_),
    .Y(_02469_));
 sg13g2_nand3_1 _11528_ (.B(_02469_),
    .C(_02096_),
    .A(_02466_),
    .Y(_02470_));
 sg13g2_buf_8 _11529_ (.A(_02438_),
    .X(_02471_));
 sg13g2_nand3_1 _11530_ (.B(_02470_),
    .C(_02471_),
    .A(_02465_),
    .Y(_02472_));
 sg13g2_nand2_1 _11531_ (.Y(_02473_),
    .A(_02464_),
    .B(_02472_));
 sg13g2_inv_1 _11532_ (.Y(_02474_),
    .A(_02430_));
 sg13g2_nand2_1 _11533_ (.Y(_02475_),
    .A(_02426_),
    .B(net173));
 sg13g2_o21ai_1 _11534_ (.B1(_02475_),
    .Y(_02476_),
    .A1(net173),
    .A2(_02474_));
 sg13g2_buf_1 _11535_ (.A(_02476_),
    .X(_02477_));
 sg13g2_inv_1 _11536_ (.Y(_02478_),
    .A(_02477_));
 sg13g2_nand2_1 _11537_ (.Y(_02479_),
    .A(_02473_),
    .B(_02478_));
 sg13g2_nand3_1 _11538_ (.B(_02472_),
    .C(_02477_),
    .A(_02464_),
    .Y(_02480_));
 sg13g2_buf_1 _11539_ (.A(_02480_),
    .X(_02481_));
 sg13g2_nand2_1 _11540_ (.Y(_02482_),
    .A(_02479_),
    .B(_02481_));
 sg13g2_nor2_1 _11541_ (.A(_02453_),
    .B(_02482_),
    .Y(_02483_));
 sg13g2_nand3_1 _11542_ (.B(_02442_),
    .C(net175),
    .A(_02441_),
    .Y(_02484_));
 sg13g2_buf_1 _11543_ (.A(_02484_),
    .X(_02485_));
 sg13g2_nand2_1 _11544_ (.Y(_02486_),
    .A(_02444_),
    .B(_02445_));
 sg13g2_nand2_1 _11545_ (.Y(_02487_),
    .A(_02486_),
    .B(net179));
 sg13g2_nand2_1 _11546_ (.Y(_02488_),
    .A(_02485_),
    .B(_02487_));
 sg13g2_nand2_1 _11547_ (.Y(_02489_),
    .A(_02488_),
    .B(net186));
 sg13g2_nand3_1 _11548_ (.B(_02487_),
    .C(net214),
    .A(_02485_),
    .Y(_02490_));
 sg13g2_nand3_1 _11549_ (.B(_02490_),
    .C(net101),
    .A(_02489_),
    .Y(_02491_));
 sg13g2_nand2_1 _11550_ (.Y(_02492_),
    .A(_02488_),
    .B(net214));
 sg13g2_nand3_1 _11551_ (.B(_02487_),
    .C(net186),
    .A(_02485_),
    .Y(_02493_));
 sg13g2_nand3_1 _11552_ (.B(_02493_),
    .C(net103),
    .A(_02492_),
    .Y(_02494_));
 sg13g2_nand2_1 _11553_ (.Y(_02495_),
    .A(_02491_),
    .B(_02494_));
 sg13g2_xnor2_1 _11554_ (.Y(_02496_),
    .A(_01972_),
    .B(_02255_));
 sg13g2_inv_1 _11555_ (.Y(_02497_),
    .A(_02496_));
 sg13g2_nand2_1 _11556_ (.Y(_02498_),
    .A(_02263_),
    .B(_01972_));
 sg13g2_nand3_1 _11557_ (.B(_02262_),
    .C(_01971_),
    .A(_02261_),
    .Y(_02499_));
 sg13g2_nand3_1 _11558_ (.B(_02499_),
    .C(_02172_),
    .A(_02498_),
    .Y(_02500_));
 sg13g2_o21ai_1 _11559_ (.B1(_02500_),
    .Y(_02501_),
    .A1(net172),
    .A2(_02497_));
 sg13g2_nand2_1 _11560_ (.Y(_02502_),
    .A(_02495_),
    .B(_02501_));
 sg13g2_nand2_1 _11561_ (.Y(_02503_),
    .A(_02496_),
    .B(_02157_));
 sg13g2_nand3_1 _11562_ (.B(_02499_),
    .C(_02127_),
    .A(_02498_),
    .Y(_02504_));
 sg13g2_nand2_1 _11563_ (.Y(_02505_),
    .A(_02503_),
    .B(_02504_));
 sg13g2_xnor2_1 _11564_ (.Y(_02506_),
    .A(net186),
    .B(_02505_));
 sg13g2_xnor2_1 _11565_ (.Y(_02507_),
    .A(net103),
    .B(_02506_));
 sg13g2_nand2_1 _11566_ (.Y(_02508_),
    .A(_02038_),
    .B(_02040_));
 sg13g2_nand3_1 _11567_ (.B(_01979_),
    .C(_02037_),
    .A(_02031_),
    .Y(_02509_));
 sg13g2_and2_1 _11568_ (.A(_02508_),
    .B(_02509_),
    .X(_02510_));
 sg13g2_xnor2_1 _11569_ (.Y(_02511_),
    .A(_02040_),
    .B(_01967_));
 sg13g2_nor2b_1 _11570_ (.A(_02128_),
    .B_N(_02511_),
    .Y(_02512_));
 sg13g2_a21o_1 _11571_ (.A2(_02510_),
    .A1(_02177_),
    .B1(_02512_),
    .X(_02513_));
 sg13g2_buf_1 _11572_ (.A(_02513_),
    .X(_02514_));
 sg13g2_nand2_1 _11573_ (.Y(_02515_),
    .A(_02507_),
    .B(_02514_));
 sg13g2_buf_1 _11574_ (.A(_02515_),
    .X(_02516_));
 sg13g2_inv_1 _11575_ (.Y(_02517_),
    .A(_02501_));
 sg13g2_nand3_1 _11576_ (.B(_02494_),
    .C(_02517_),
    .A(_02491_),
    .Y(_02518_));
 sg13g2_inv_1 _11577_ (.Y(_02519_),
    .A(_02518_));
 sg13g2_a21oi_1 _11578_ (.A1(_02502_),
    .A2(_02516_),
    .Y(_02520_),
    .B1(_02519_));
 sg13g2_nand2b_1 _11579_ (.Y(_02521_),
    .B(_02479_),
    .A_N(_02452_));
 sg13g2_nand2_1 _11580_ (.Y(_02522_),
    .A(_02521_),
    .B(_02481_));
 sg13g2_a21oi_1 _11581_ (.A1(_02483_),
    .A2(_02520_),
    .Y(_02523_),
    .B1(_02522_));
 sg13g2_xnor2_1 _11582_ (.Y(_02524_),
    .A(net101),
    .B(_02506_));
 sg13g2_nand2b_1 _11583_ (.Y(_02525_),
    .B(_02524_),
    .A_N(_02514_));
 sg13g2_buf_1 _11584_ (.A(_02525_),
    .X(_02526_));
 sg13g2_nand2_1 _11585_ (.Y(_02527_),
    .A(_02526_),
    .B(_02516_));
 sg13g2_nand2_2 _11586_ (.Y(_02528_),
    .A(_02502_),
    .B(_02518_));
 sg13g2_nor2_1 _11587_ (.A(_02527_),
    .B(_02528_),
    .Y(_02529_));
 sg13g2_xnor2_1 _11588_ (.Y(_02530_),
    .A(_02028_),
    .B(_02116_));
 sg13g2_nand2_1 _11589_ (.Y(_02531_),
    .A(_02530_),
    .B(net187));
 sg13g2_nand2_1 _11590_ (.Y(_02532_),
    .A(_02141_),
    .B(_02028_));
 sg13g2_nand2_1 _11591_ (.Y(_02533_),
    .A(_02140_),
    .B(_01957_));
 sg13g2_nand3_1 _11592_ (.B(_02023_),
    .C(_02533_),
    .A(_02532_),
    .Y(_02534_));
 sg13g2_nand2_1 _11593_ (.Y(_02535_),
    .A(_02531_),
    .B(_02534_));
 sg13g2_xnor2_1 _11594_ (.Y(_02536_),
    .A(_02098_),
    .B(_02535_));
 sg13g2_inv_1 _11595_ (.Y(_02537_),
    .A(_02536_));
 sg13g2_nand2_1 _11596_ (.Y(_02538_),
    .A(net103),
    .B(_02537_));
 sg13g2_nand3_1 _11597_ (.B(_02536_),
    .C(_02093_),
    .A(_02025_),
    .Y(_02539_));
 sg13g2_xor2_1 _11598_ (.B(_02026_),
    .A(_02030_),
    .X(_02540_));
 sg13g2_xnor2_1 _11599_ (.Y(_02541_),
    .A(_01960_),
    .B(_02026_));
 sg13g2_nor2_1 _11600_ (.A(_02177_),
    .B(_02541_),
    .Y(_02542_));
 sg13g2_a21o_1 _11601_ (.A2(_02540_),
    .A1(_02374_),
    .B1(_02542_),
    .X(_02543_));
 sg13g2_nand3_1 _11602_ (.B(_02539_),
    .C(_02543_),
    .A(_02538_),
    .Y(_02544_));
 sg13g2_nor2_1 _11603_ (.A(net187),
    .B(_02540_),
    .Y(_02545_));
 sg13g2_a21oi_1 _11604_ (.A1(net179),
    .A2(_02541_),
    .Y(_02546_),
    .B1(_02545_));
 sg13g2_xnor2_1 _11605_ (.Y(_02547_),
    .A(_02461_),
    .B(_02546_));
 sg13g2_inv_1 _11606_ (.Y(_02548_),
    .A(_02547_));
 sg13g2_nand2_1 _11607_ (.Y(_02549_),
    .A(net103),
    .B(_02548_));
 sg13g2_nand3_1 _11608_ (.B(_02093_),
    .C(_02547_),
    .A(_02025_),
    .Y(_02550_));
 sg13g2_xor2_1 _11609_ (.B(_01959_),
    .A(_01958_),
    .X(_02551_));
 sg13g2_nand3_1 _11610_ (.B(_02550_),
    .C(_02551_),
    .A(_02549_),
    .Y(_02552_));
 sg13g2_nand2_1 _11611_ (.Y(_02553_),
    .A(_02544_),
    .B(_02552_));
 sg13g2_nand2_1 _11612_ (.Y(_02554_),
    .A(_02511_),
    .B(net187));
 sg13g2_nand3_1 _11613_ (.B(_02509_),
    .C(_02157_),
    .A(_02508_),
    .Y(_02555_));
 sg13g2_nand2_1 _11614_ (.Y(_02556_),
    .A(_02554_),
    .B(_02555_));
 sg13g2_xnor2_1 _11615_ (.Y(_02557_),
    .A(_02096_),
    .B(_02556_));
 sg13g2_inv_1 _11616_ (.Y(_02558_),
    .A(_02557_));
 sg13g2_nand2_1 _11617_ (.Y(_02559_),
    .A(_02558_),
    .B(net103));
 sg13g2_nand2_1 _11618_ (.Y(_02560_),
    .A(_02557_),
    .B(net101));
 sg13g2_nand2_1 _11619_ (.Y(_02561_),
    .A(_02532_),
    .B(_02533_));
 sg13g2_nand2_1 _11620_ (.Y(_02562_),
    .A(_02530_),
    .B(_02172_));
 sg13g2_o21ai_1 _11621_ (.B1(_02562_),
    .Y(_02563_),
    .A1(net172),
    .A2(_02561_));
 sg13g2_inv_1 _11622_ (.Y(_02564_),
    .A(_02563_));
 sg13g2_nand3_1 _11623_ (.B(_02560_),
    .C(_02564_),
    .A(_02559_),
    .Y(_02565_));
 sg13g2_nand2_1 _11624_ (.Y(_02566_),
    .A(_02538_),
    .B(_02539_));
 sg13g2_inv_1 _11625_ (.Y(_02567_),
    .A(_02543_));
 sg13g2_nand2_1 _11626_ (.Y(_02568_),
    .A(_02566_),
    .B(_02567_));
 sg13g2_nand3_1 _11627_ (.B(_02565_),
    .C(_02568_),
    .A(_02553_),
    .Y(_02569_));
 sg13g2_nand2_1 _11628_ (.Y(_02570_),
    .A(_02559_),
    .B(_02560_));
 sg13g2_nand2_1 _11629_ (.Y(_02571_),
    .A(_02570_),
    .B(_02563_));
 sg13g2_nand2_1 _11630_ (.Y(_02572_),
    .A(_02569_),
    .B(_02571_));
 sg13g2_nand3_1 _11631_ (.B(_02529_),
    .C(_02572_),
    .A(_02483_),
    .Y(_02573_));
 sg13g2_nand2_2 _11632_ (.Y(_02574_),
    .A(_02523_),
    .B(_02573_));
 sg13g2_nand2_1 _11633_ (.Y(_02575_),
    .A(_02277_),
    .B(_02254_));
 sg13g2_nand3_1 _11634_ (.B(_02276_),
    .C(_02253_),
    .A(_02274_),
    .Y(_02576_));
 sg13g2_nand2_1 _11635_ (.Y(_02577_),
    .A(_02575_),
    .B(_02576_));
 sg13g2_nand2_2 _11636_ (.Y(_02578_),
    .A(_02295_),
    .B(_02292_));
 sg13g2_nor2_1 _11637_ (.A(_02577_),
    .B(_02578_),
    .Y(_02579_));
 sg13g2_nand2_1 _11638_ (.Y(_02580_),
    .A(_02579_),
    .B(_02244_));
 sg13g2_xnor2_1 _11639_ (.Y(_02581_),
    .A(_02415_),
    .B(_02359_));
 sg13g2_nand2_1 _11640_ (.Y(_02582_),
    .A(_02414_),
    .B(_02418_));
 sg13g2_nor2_1 _11641_ (.A(_02581_),
    .B(_02582_),
    .Y(_02583_));
 sg13g2_nand2_1 _11642_ (.Y(_02584_),
    .A(_02583_),
    .B(_02412_));
 sg13g2_nor2_1 _11643_ (.A(_02580_),
    .B(_02584_),
    .Y(_02585_));
 sg13g2_nand2_1 _11644_ (.Y(_02586_),
    .A(_02574_),
    .B(_02585_));
 sg13g2_nand2_1 _11645_ (.Y(_02587_),
    .A(_02425_),
    .B(_02586_));
 sg13g2_xnor2_1 _11646_ (.Y(_02588_),
    .A(net186),
    .B(_02389_));
 sg13g2_nand2_1 _11647_ (.Y(_02589_),
    .A(_02587_),
    .B(_02588_));
 sg13g2_inv_1 _11648_ (.Y(_02590_),
    .A(_02588_));
 sg13g2_nand3_1 _11649_ (.B(_02590_),
    .C(_02586_),
    .A(_02425_),
    .Y(_02591_));
 sg13g2_buf_8 _11650_ (.A(_02591_),
    .X(_02592_));
 sg13g2_nand2_1 _11651_ (.Y(_02593_),
    .A(_02589_),
    .B(_02592_));
 sg13g2_buf_1 _11652_ (.A(_02593_),
    .X(_02594_));
 sg13g2_xnor2_1 _11653_ (.Y(_02595_),
    .A(_02527_),
    .B(_02572_));
 sg13g2_inv_1 _11654_ (.Y(_02596_),
    .A(_02595_));
 sg13g2_nand2_1 _11655_ (.Y(_02597_),
    .A(net73),
    .B(_02596_));
 sg13g2_nand3_1 _11656_ (.B(_02592_),
    .C(_02595_),
    .A(_02589_),
    .Y(_02598_));
 sg13g2_nand3_1 _11657_ (.B(_02598_),
    .C(_02548_),
    .A(_02597_),
    .Y(_02599_));
 sg13g2_buf_1 _11658_ (.A(_02599_),
    .X(_02600_));
 sg13g2_xnor2_1 _11659_ (.Y(_02601_),
    .A(_02564_),
    .B(_02436_));
 sg13g2_a21oi_1 _11660_ (.A1(_02597_),
    .A2(_02598_),
    .Y(_02602_),
    .B1(_02548_));
 sg13g2_a21oi_1 _11661_ (.A1(_02600_),
    .A2(_02601_),
    .Y(_02603_),
    .B1(_02602_));
 sg13g2_inv_1 _11662_ (.Y(_02604_),
    .A(_02603_));
 sg13g2_nand2_1 _11663_ (.Y(_02605_),
    .A(_02572_),
    .B(_02526_));
 sg13g2_nand2_1 _11664_ (.Y(_02606_),
    .A(_02605_),
    .B(_02516_));
 sg13g2_xnor2_1 _11665_ (.Y(_02607_),
    .A(_02528_),
    .B(_02606_));
 sg13g2_inv_1 _11666_ (.Y(_02608_),
    .A(_02607_));
 sg13g2_nand2_1 _11667_ (.Y(_02609_),
    .A(net73),
    .B(_02608_));
 sg13g2_nand3_1 _11668_ (.B(_02592_),
    .C(_02607_),
    .A(_02589_),
    .Y(_02610_));
 sg13g2_buf_1 _11669_ (.A(_02610_),
    .X(_02611_));
 sg13g2_nand2_1 _11670_ (.Y(_02612_),
    .A(_02609_),
    .B(_02611_));
 sg13g2_nand2_1 _11671_ (.Y(_02613_),
    .A(_02612_),
    .B(_02536_));
 sg13g2_nand3_1 _11672_ (.B(_02611_),
    .C(_02537_),
    .A(_02609_),
    .Y(_02614_));
 sg13g2_buf_1 _11673_ (.A(_02614_),
    .X(_02615_));
 sg13g2_xnor2_1 _11674_ (.Y(_02616_),
    .A(net101),
    .B(_02514_));
 sg13g2_nand3_1 _11675_ (.B(_02615_),
    .C(_02616_),
    .A(_02613_),
    .Y(_02617_));
 sg13g2_buf_1 _11676_ (.A(_02617_),
    .X(_02618_));
 sg13g2_nand2_1 _11677_ (.Y(_02619_),
    .A(_02613_),
    .B(_02615_));
 sg13g2_inv_1 _11678_ (.Y(_02620_),
    .A(_02616_));
 sg13g2_nand2_1 _11679_ (.Y(_02621_),
    .A(_02619_),
    .B(_02620_));
 sg13g2_nand3_1 _11680_ (.B(_02618_),
    .C(_02621_),
    .A(_02604_),
    .Y(_02622_));
 sg13g2_buf_1 _11681_ (.A(_02622_),
    .X(_02623_));
 sg13g2_nand2_1 _11682_ (.Y(_02624_),
    .A(_02621_),
    .B(_02618_));
 sg13g2_nand2_1 _11683_ (.Y(_02625_),
    .A(_02624_),
    .B(_02603_));
 sg13g2_nand2_1 _11684_ (.Y(_02626_),
    .A(_02623_),
    .B(_02625_));
 sg13g2_buf_8 _11685_ (.A(net73),
    .X(_02627_));
 sg13g2_nand2_1 _11686_ (.Y(_02628_),
    .A(net71),
    .B(_02595_));
 sg13g2_nand2_1 _11687_ (.Y(_02629_),
    .A(_02587_),
    .B(_02590_));
 sg13g2_nand3_1 _11688_ (.B(_02588_),
    .C(_02586_),
    .A(_02425_),
    .Y(_02630_));
 sg13g2_nand2_1 _11689_ (.Y(_02631_),
    .A(_02629_),
    .B(_02630_));
 sg13g2_buf_8 _11690_ (.A(_02631_),
    .X(_02632_));
 sg13g2_nand2_1 _11691_ (.Y(_02633_),
    .A(net72),
    .B(_02596_));
 sg13g2_nand3_1 _11692_ (.B(_02633_),
    .C(_02547_),
    .A(_02628_),
    .Y(_02634_));
 sg13g2_nand2_1 _11693_ (.Y(_02635_),
    .A(_02634_),
    .B(_02600_));
 sg13g2_inv_1 _11694_ (.Y(_02636_),
    .A(_02601_));
 sg13g2_nand2_1 _11695_ (.Y(_02637_),
    .A(_02635_),
    .B(_02636_));
 sg13g2_nand3_1 _11696_ (.B(_02600_),
    .C(_02601_),
    .A(_02634_),
    .Y(_02638_));
 sg13g2_xnor2_1 _11697_ (.Y(_02639_),
    .A(_02461_),
    .B(_02551_));
 sg13g2_xnor2_1 _11698_ (.Y(_02640_),
    .A(_02567_),
    .B(_02436_));
 sg13g2_nor2_1 _11699_ (.A(_02639_),
    .B(_02640_),
    .Y(_02641_));
 sg13g2_nand2_1 _11700_ (.Y(_02642_),
    .A(_02571_),
    .B(_02565_));
 sg13g2_nand2_1 _11701_ (.Y(_02643_),
    .A(_02553_),
    .B(_02568_));
 sg13g2_xnor2_1 _11702_ (.Y(_02644_),
    .A(_02642_),
    .B(_02643_));
 sg13g2_buf_1 _11703_ (.A(net72),
    .X(_02645_));
 sg13g2_xnor2_1 _11704_ (.Y(_02646_),
    .A(_02644_),
    .B(_02645_));
 sg13g2_nand2_1 _11705_ (.Y(_02647_),
    .A(_02640_),
    .B(_02639_));
 sg13g2_o21ai_1 _11706_ (.B1(_02647_),
    .Y(_02648_),
    .A1(_02641_),
    .A2(_02646_));
 sg13g2_buf_1 _11707_ (.A(_02648_),
    .X(_02649_));
 sg13g2_nand3_1 _11708_ (.B(_02638_),
    .C(_02649_),
    .A(_02637_),
    .Y(_02650_));
 sg13g2_nand2_1 _11709_ (.Y(_02651_),
    .A(_02626_),
    .B(_02650_));
 sg13g2_nand2_1 _11710_ (.Y(_02652_),
    .A(_02637_),
    .B(_02638_));
 sg13g2_nor2b_1 _11711_ (.A(_02652_),
    .B_N(_02649_),
    .Y(_02653_));
 sg13g2_nand3_1 _11712_ (.B(_02653_),
    .C(_02625_),
    .A(_02623_),
    .Y(_02654_));
 sg13g2_nand2_1 _11713_ (.Y(_02655_),
    .A(_02651_),
    .B(_02654_));
 sg13g2_nor2_1 _11714_ (.A(_02603_),
    .B(_02624_),
    .Y(_02656_));
 sg13g2_a21oi_1 _11715_ (.A1(_02609_),
    .A2(_02611_),
    .Y(_02657_),
    .B1(_02537_));
 sg13g2_a21oi_2 _11716_ (.B1(_02657_),
    .Y(_02658_),
    .A2(_02616_),
    .A1(_02615_));
 sg13g2_xnor2_1 _11717_ (.Y(_02659_),
    .A(_02517_),
    .B(net103));
 sg13g2_inv_1 _11718_ (.Y(_02660_),
    .A(_02528_));
 sg13g2_nand4_1 _11719_ (.B(_02660_),
    .C(_02516_),
    .A(_02572_),
    .Y(_02661_),
    .D(_02526_));
 sg13g2_nand2b_1 _11720_ (.Y(_02662_),
    .B(_02661_),
    .A_N(_02520_));
 sg13g2_xnor2_1 _11721_ (.Y(_02663_),
    .A(_02453_),
    .B(_02662_));
 sg13g2_nand2b_1 _11722_ (.Y(_02664_),
    .B(net73),
    .A_N(_02663_));
 sg13g2_nand3_1 _11723_ (.B(_02592_),
    .C(_02663_),
    .A(_02589_),
    .Y(_02665_));
 sg13g2_buf_1 _11724_ (.A(_02665_),
    .X(_02666_));
 sg13g2_nand2_1 _11725_ (.Y(_02667_),
    .A(_02664_),
    .B(_02666_));
 sg13g2_nand2_1 _11726_ (.Y(_02668_),
    .A(_02667_),
    .B(_02558_));
 sg13g2_nand3_1 _11727_ (.B(_02666_),
    .C(_02557_),
    .A(_02664_),
    .Y(_02669_));
 sg13g2_buf_1 _11728_ (.A(_02669_),
    .X(_02670_));
 sg13g2_nand2_1 _11729_ (.Y(_02671_),
    .A(_02668_),
    .B(_02670_));
 sg13g2_nand2b_1 _11730_ (.Y(_02672_),
    .B(_02671_),
    .A_N(_02659_));
 sg13g2_nand3_1 _11731_ (.B(_02670_),
    .C(_02659_),
    .A(_02668_),
    .Y(_02673_));
 sg13g2_buf_1 _11732_ (.A(_02673_),
    .X(_02674_));
 sg13g2_nand2_1 _11733_ (.Y(_02675_),
    .A(_02672_),
    .B(_02674_));
 sg13g2_nor2_1 _11734_ (.A(_02658_),
    .B(_02675_),
    .Y(_02676_));
 sg13g2_nor2_1 _11735_ (.A(_02656_),
    .B(_02676_),
    .Y(_02677_));
 sg13g2_nand2_1 _11736_ (.Y(_02678_),
    .A(_02654_),
    .B(_02677_));
 sg13g2_nand2_1 _11737_ (.Y(_02679_),
    .A(_02675_),
    .B(_02658_));
 sg13g2_nand2_1 _11738_ (.Y(_02680_),
    .A(_02678_),
    .B(_02679_));
 sg13g2_a21oi_1 _11739_ (.A1(_02664_),
    .A2(_02666_),
    .Y(_02681_),
    .B1(_02557_));
 sg13g2_a21oi_1 _11740_ (.A1(_02670_),
    .A2(_02659_),
    .Y(_02682_),
    .B1(_02681_));
 sg13g2_inv_1 _11741_ (.Y(_02683_),
    .A(_02682_));
 sg13g2_inv_1 _11742_ (.Y(_02684_),
    .A(_02450_));
 sg13g2_a21oi_1 _11743_ (.A1(_02502_),
    .A2(_02452_),
    .Y(_02685_),
    .B1(_02684_));
 sg13g2_inv_1 _11744_ (.Y(_02686_),
    .A(_02526_));
 sg13g2_o21ai_1 _11745_ (.B1(_02516_),
    .Y(_02687_),
    .A1(_02571_),
    .A2(_02686_));
 sg13g2_nor2_1 _11746_ (.A(_02453_),
    .B(_02528_),
    .Y(_02688_));
 sg13g2_nand2_1 _11747_ (.Y(_02689_),
    .A(_02687_),
    .B(_02688_));
 sg13g2_nand2b_1 _11748_ (.Y(_02690_),
    .B(_02689_),
    .A_N(_02685_));
 sg13g2_inv_1 _11749_ (.Y(_02691_),
    .A(_02688_));
 sg13g2_nor2_1 _11750_ (.A(_02642_),
    .B(_02527_),
    .Y(_02692_));
 sg13g2_nor2b_1 _11751_ (.A(_02691_),
    .B_N(_02692_),
    .Y(_02693_));
 sg13g2_inv_1 _11752_ (.Y(_02694_),
    .A(_02643_));
 sg13g2_nand2_1 _11753_ (.Y(_02695_),
    .A(_02693_),
    .B(_02694_));
 sg13g2_nand2b_1 _11754_ (.Y(_02696_),
    .B(_02695_),
    .A_N(_02690_));
 sg13g2_xnor2_1 _11755_ (.Y(_02697_),
    .A(_02482_),
    .B(_02696_));
 sg13g2_nand2_1 _11756_ (.Y(_02698_),
    .A(net72),
    .B(_02697_));
 sg13g2_inv_1 _11757_ (.Y(_02699_),
    .A(_02697_));
 sg13g2_nand2_1 _11758_ (.Y(_02700_),
    .A(_02594_),
    .B(_02699_));
 sg13g2_nand2_1 _11759_ (.Y(_02701_),
    .A(_02698_),
    .B(_02700_));
 sg13g2_nand2_1 _11760_ (.Y(_02702_),
    .A(_02701_),
    .B(_02506_));
 sg13g2_inv_1 _11761_ (.Y(_02703_),
    .A(_02506_));
 sg13g2_nand3_1 _11762_ (.B(_02700_),
    .C(_02703_),
    .A(_02698_),
    .Y(_02704_));
 sg13g2_buf_1 _11763_ (.A(_02704_),
    .X(_02705_));
 sg13g2_nand2_1 _11764_ (.Y(_02706_),
    .A(_02702_),
    .B(_02705_));
 sg13g2_xnor2_1 _11765_ (.Y(_02707_),
    .A(_02471_),
    .B(_02448_));
 sg13g2_inv_1 _11766_ (.Y(_02708_),
    .A(_02707_));
 sg13g2_nand2_1 _11767_ (.Y(_02709_),
    .A(_02706_),
    .B(_02708_));
 sg13g2_nand3_1 _11768_ (.B(_02705_),
    .C(_02707_),
    .A(_02702_),
    .Y(_02710_));
 sg13g2_nand2_1 _11769_ (.Y(_02711_),
    .A(_02709_),
    .B(_02710_));
 sg13g2_xnor2_1 _11770_ (.Y(_02712_),
    .A(_02683_),
    .B(_02711_));
 sg13g2_nand2_1 _11771_ (.Y(_02713_),
    .A(_02680_),
    .B(_02712_));
 sg13g2_nand2_1 _11772_ (.Y(_02714_),
    .A(_02711_),
    .B(_02682_));
 sg13g2_nand3_1 _11773_ (.B(_02709_),
    .C(_02710_),
    .A(_02683_),
    .Y(_02715_));
 sg13g2_buf_1 _11774_ (.A(_02715_),
    .X(_02716_));
 sg13g2_nand2_1 _11775_ (.Y(_02717_),
    .A(_02714_),
    .B(_02716_));
 sg13g2_nand3_1 _11776_ (.B(_02717_),
    .C(_02679_),
    .A(_02678_),
    .Y(_02718_));
 sg13g2_nand2_1 _11777_ (.Y(_02719_),
    .A(_02713_),
    .B(_02718_));
 sg13g2_nand2b_1 _11778_ (.Y(_02720_),
    .B(_02719_),
    .A_N(_02655_));
 sg13g2_buf_1 _11779_ (.A(_02720_),
    .X(_02721_));
 sg13g2_nand3_1 _11780_ (.B(_02718_),
    .C(_02655_),
    .A(_02713_),
    .Y(_02722_));
 sg13g2_xor2_1 _11781_ (.B(_02652_),
    .A(_02649_),
    .X(_02723_));
 sg13g2_inv_1 _11782_ (.Y(_02724_),
    .A(_02658_));
 sg13g2_nand2_1 _11783_ (.Y(_02725_),
    .A(_02675_),
    .B(_02724_));
 sg13g2_nand3_1 _11784_ (.B(_02658_),
    .C(_02674_),
    .A(_02672_),
    .Y(_02726_));
 sg13g2_nand2_1 _11785_ (.Y(_02727_),
    .A(_02725_),
    .B(_02726_));
 sg13g2_a21oi_1 _11786_ (.A1(_02621_),
    .A2(_02618_),
    .Y(_02728_),
    .B1(_02604_));
 sg13g2_o21ai_1 _11787_ (.B1(_02623_),
    .Y(_02729_),
    .A1(_02650_),
    .A2(_02728_));
 sg13g2_buf_1 _11788_ (.A(_02729_),
    .X(_02730_));
 sg13g2_xnor2_1 _11789_ (.Y(_02731_),
    .A(_02727_),
    .B(_02730_));
 sg13g2_nor2_1 _11790_ (.A(_02723_),
    .B(_02731_),
    .Y(_02732_));
 sg13g2_nand3_1 _11791_ (.B(_02722_),
    .C(_02732_),
    .A(_02721_),
    .Y(_02733_));
 sg13g2_buf_1 _11792_ (.A(_02733_),
    .X(_02734_));
 sg13g2_inv_1 _11793_ (.Y(_02735_),
    .A(_02702_));
 sg13g2_a21oi_2 _11794_ (.B1(_02735_),
    .Y(_02736_),
    .A2(_02707_),
    .A1(_02705_));
 sg13g2_xor2_1 _11795_ (.B(_02477_),
    .A(net103),
    .X(_02737_));
 sg13g2_inv_1 _11796_ (.Y(_02738_),
    .A(_02577_));
 sg13g2_xnor2_1 _11797_ (.Y(_02739_),
    .A(_02738_),
    .B(_02574_));
 sg13g2_nand2_1 _11798_ (.Y(_02740_),
    .A(net71),
    .B(_02739_));
 sg13g2_inv_1 _11799_ (.Y(_02741_),
    .A(_02739_));
 sg13g2_nand2_1 _11800_ (.Y(_02742_),
    .A(_02632_),
    .B(_02741_));
 sg13g2_nand2_1 _11801_ (.Y(_02743_),
    .A(_02740_),
    .B(_02742_));
 sg13g2_nand2_1 _11802_ (.Y(_02744_),
    .A(_02489_),
    .B(_02490_));
 sg13g2_nand2_1 _11803_ (.Y(_02745_),
    .A(_02743_),
    .B(_02744_));
 sg13g2_inv_1 _11804_ (.Y(_02746_),
    .A(_02744_));
 sg13g2_nand3_1 _11805_ (.B(_02742_),
    .C(_02746_),
    .A(_02740_),
    .Y(_02747_));
 sg13g2_buf_1 _11806_ (.A(_02747_),
    .X(_02748_));
 sg13g2_nand2_1 _11807_ (.Y(_02749_),
    .A(_02745_),
    .B(_02748_));
 sg13g2_nand2b_1 _11808_ (.Y(_02750_),
    .B(_02749_),
    .A_N(_02737_));
 sg13g2_nand3_1 _11809_ (.B(_02748_),
    .C(_02737_),
    .A(_02745_),
    .Y(_02751_));
 sg13g2_buf_1 _11810_ (.A(_02751_),
    .X(_02752_));
 sg13g2_nand2_1 _11811_ (.Y(_02753_),
    .A(_02750_),
    .B(_02752_));
 sg13g2_xnor2_1 _11812_ (.Y(_02754_),
    .A(_02736_),
    .B(_02753_));
 sg13g2_nand2_1 _11813_ (.Y(_02755_),
    .A(_02714_),
    .B(_02676_));
 sg13g2_nand2_1 _11814_ (.Y(_02756_),
    .A(_02755_),
    .B(_02716_));
 sg13g2_nand3_1 _11815_ (.B(_02672_),
    .C(_02674_),
    .A(_02724_),
    .Y(_02757_));
 sg13g2_nand2_1 _11816_ (.Y(_02758_),
    .A(_02757_),
    .B(_02679_));
 sg13g2_nor2_1 _11817_ (.A(_02758_),
    .B(_02717_),
    .Y(_02759_));
 sg13g2_nand2_1 _11818_ (.Y(_02760_),
    .A(_02730_),
    .B(_02759_));
 sg13g2_nand2b_1 _11819_ (.Y(_02761_),
    .B(_02760_),
    .A_N(_02756_));
 sg13g2_buf_1 _11820_ (.A(_02761_),
    .X(_02762_));
 sg13g2_xnor2_1 _11821_ (.Y(_02763_),
    .A(_02754_),
    .B(_02762_));
 sg13g2_nand2b_1 _11822_ (.Y(_02764_),
    .B(_02763_),
    .A_N(_02731_));
 sg13g2_buf_1 _11823_ (.A(_02764_),
    .X(_02765_));
 sg13g2_inv_1 _11824_ (.Y(_02766_),
    .A(_02736_));
 sg13g2_xnor2_1 _11825_ (.Y(_02767_),
    .A(_02766_),
    .B(_02753_));
 sg13g2_xnor2_1 _11826_ (.Y(_02768_),
    .A(_02767_),
    .B(_02762_));
 sg13g2_nand2_1 _11827_ (.Y(_02769_),
    .A(_02768_),
    .B(_02731_));
 sg13g2_nand2_1 _11828_ (.Y(_02770_),
    .A(_02765_),
    .B(_02769_));
 sg13g2_a21oi_2 _11829_ (.B1(_02770_),
    .Y(_02771_),
    .A2(_02721_),
    .A1(_02734_));
 sg13g2_nand3_1 _11830_ (.B(_02750_),
    .C(_02752_),
    .A(_02766_),
    .Y(_02772_));
 sg13g2_a21oi_1 _11831_ (.A1(_02750_),
    .A2(_02752_),
    .Y(_02773_),
    .B1(_02766_));
 sg13g2_a21oi_1 _11832_ (.A1(_02772_),
    .A2(_02716_),
    .Y(_02774_),
    .B1(_02773_));
 sg13g2_a21oi_1 _11833_ (.A1(_02656_),
    .A2(_02679_),
    .Y(_02775_),
    .B1(_02676_));
 sg13g2_nand2_1 _11834_ (.Y(_02776_),
    .A(_02767_),
    .B(_02712_));
 sg13g2_nor2_1 _11835_ (.A(_02775_),
    .B(_02776_),
    .Y(_02777_));
 sg13g2_nor2_1 _11836_ (.A(_02774_),
    .B(_02777_),
    .Y(_02778_));
 sg13g2_nor2_1 _11837_ (.A(_02717_),
    .B(_02754_),
    .Y(_02779_));
 sg13g2_nor2_1 _11838_ (.A(_02626_),
    .B(_02758_),
    .Y(_02780_));
 sg13g2_nand3_1 _11839_ (.B(_02780_),
    .C(_02653_),
    .A(_02779_),
    .Y(_02781_));
 sg13g2_nand2_2 _11840_ (.Y(_02782_),
    .A(_02778_),
    .B(_02781_));
 sg13g2_inv_1 _11841_ (.Y(_02783_),
    .A(_02745_));
 sg13g2_a21oi_2 _11842_ (.B1(_02783_),
    .Y(_02784_),
    .A2(_02737_),
    .A1(_02748_));
 sg13g2_buf_1 _11843_ (.A(net101),
    .X(_02785_));
 sg13g2_xnor2_1 _11844_ (.Y(_02786_),
    .A(net94),
    .B(_02253_));
 sg13g2_nor2_1 _11845_ (.A(_02482_),
    .B(_02577_),
    .Y(_02787_));
 sg13g2_inv_1 _11846_ (.Y(_02788_),
    .A(_02787_));
 sg13g2_nor2_1 _11847_ (.A(_02691_),
    .B(_02788_),
    .Y(_02789_));
 sg13g2_inv_1 _11848_ (.Y(_02790_),
    .A(_02575_));
 sg13g2_a21oi_1 _11849_ (.A1(_02576_),
    .A2(_02481_),
    .Y(_02791_),
    .B1(_02790_));
 sg13g2_nand2_1 _11850_ (.Y(_02792_),
    .A(_02787_),
    .B(_02685_));
 sg13g2_nand2b_1 _11851_ (.Y(_02793_),
    .B(_02792_),
    .A_N(_02791_));
 sg13g2_a21o_1 _11852_ (.A2(_02789_),
    .A1(_02606_),
    .B1(_02793_),
    .X(_02794_));
 sg13g2_xor2_1 _11853_ (.B(_02794_),
    .A(_02578_),
    .X(_02795_));
 sg13g2_nand2_1 _11854_ (.Y(_02796_),
    .A(net71),
    .B(_02795_));
 sg13g2_xnor2_1 _11855_ (.Y(_02797_),
    .A(_02578_),
    .B(_02794_));
 sg13g2_nand2_1 _11856_ (.Y(_02798_),
    .A(net72),
    .B(_02797_));
 sg13g2_nand2_1 _11857_ (.Y(_02799_),
    .A(_02796_),
    .B(_02798_));
 sg13g2_nand2b_1 _11858_ (.Y(_02800_),
    .B(_02799_),
    .A_N(_02435_));
 sg13g2_nand3_1 _11859_ (.B(_02798_),
    .C(_02435_),
    .A(_02796_),
    .Y(_02801_));
 sg13g2_buf_1 _11860_ (.A(_02801_),
    .X(_02802_));
 sg13g2_nand2_1 _11861_ (.Y(_02803_),
    .A(_02800_),
    .B(_02802_));
 sg13g2_nand2b_1 _11862_ (.Y(_02804_),
    .B(_02803_),
    .A_N(_02786_));
 sg13g2_nand3_1 _11863_ (.B(_02802_),
    .C(_02786_),
    .A(_02800_),
    .Y(_02805_));
 sg13g2_nand2_2 _11864_ (.Y(_02806_),
    .A(_02804_),
    .B(_02805_));
 sg13g2_xnor2_1 _11865_ (.Y(_02807_),
    .A(_02784_),
    .B(_02806_));
 sg13g2_nand2_1 _11866_ (.Y(_02808_),
    .A(_02782_),
    .B(_02807_));
 sg13g2_xor2_1 _11867_ (.B(_02806_),
    .A(_02784_),
    .X(_02809_));
 sg13g2_nand3_1 _11868_ (.B(_02781_),
    .C(_02809_),
    .A(_02778_),
    .Y(_02810_));
 sg13g2_nand2_1 _11869_ (.Y(_02811_),
    .A(_02808_),
    .B(_02810_));
 sg13g2_inv_1 _11870_ (.Y(_02812_),
    .A(_02719_));
 sg13g2_nand2_1 _11871_ (.Y(_02813_),
    .A(_02811_),
    .B(_02812_));
 sg13g2_nand3_1 _11872_ (.B(_02810_),
    .C(_02719_),
    .A(_02808_),
    .Y(_02814_));
 sg13g2_buf_1 _11873_ (.A(_02814_),
    .X(_02815_));
 sg13g2_nand3_1 _11874_ (.B(_02815_),
    .C(_02765_),
    .A(_02813_),
    .Y(_02816_));
 sg13g2_a21oi_1 _11875_ (.A1(_02813_),
    .A2(_02815_),
    .Y(_02817_),
    .B1(_02765_));
 sg13g2_a21oi_1 _11876_ (.A1(_02771_),
    .A2(_02816_),
    .Y(_02818_),
    .B1(_02817_));
 sg13g2_inv_1 _11877_ (.Y(_02819_),
    .A(_02818_));
 sg13g2_nand2_1 _11878_ (.Y(_02820_),
    .A(_02811_),
    .B(_02719_));
 sg13g2_inv_1 _11879_ (.Y(_02821_),
    .A(_02820_));
 sg13g2_inv_1 _11880_ (.Y(_02822_),
    .A(_02800_));
 sg13g2_a21oi_2 _11881_ (.B1(_02822_),
    .Y(_02823_),
    .A2(_02786_),
    .A1(_02802_));
 sg13g2_xnor2_1 _11882_ (.Y(_02824_),
    .A(net101),
    .B(_02290_));
 sg13g2_a21oi_1 _11883_ (.A1(_02574_),
    .A2(_02579_),
    .Y(_02825_),
    .B1(_02296_));
 sg13g2_xnor2_1 _11884_ (.Y(_02826_),
    .A(_02210_),
    .B(_02825_));
 sg13g2_nand2_1 _11885_ (.Y(_02827_),
    .A(net73),
    .B(_02826_));
 sg13g2_inv_1 _11886_ (.Y(_02828_),
    .A(_02210_));
 sg13g2_xnor2_1 _11887_ (.Y(_02829_),
    .A(_02828_),
    .B(_02825_));
 sg13g2_nand2_1 _11888_ (.Y(_02830_),
    .A(_02632_),
    .B(_02829_));
 sg13g2_nand2_1 _11889_ (.Y(_02831_),
    .A(_02827_),
    .B(_02830_));
 sg13g2_nand2_1 _11890_ (.Y(_02832_),
    .A(_02462_),
    .B(_02463_));
 sg13g2_nand2_1 _11891_ (.Y(_02833_),
    .A(_02831_),
    .B(_02832_));
 sg13g2_inv_1 _11892_ (.Y(_02834_),
    .A(_02832_));
 sg13g2_nand3_1 _11893_ (.B(_02830_),
    .C(_02834_),
    .A(_02827_),
    .Y(_02835_));
 sg13g2_buf_1 _11894_ (.A(_02835_),
    .X(_02836_));
 sg13g2_nand2_1 _11895_ (.Y(_02837_),
    .A(_02833_),
    .B(_02836_));
 sg13g2_nand2b_1 _11896_ (.Y(_02838_),
    .B(_02837_),
    .A_N(_02824_));
 sg13g2_nand3_1 _11897_ (.B(_02836_),
    .C(_02824_),
    .A(_02833_),
    .Y(_02839_));
 sg13g2_nand2_1 _11898_ (.Y(_02840_),
    .A(_02838_),
    .B(_02839_));
 sg13g2_xnor2_1 _11899_ (.Y(_02841_),
    .A(_02823_),
    .B(_02840_));
 sg13g2_inv_2 _11900_ (.Y(_02842_),
    .A(_02841_));
 sg13g2_nor2_1 _11901_ (.A(_02754_),
    .B(_02807_),
    .Y(_02843_));
 sg13g2_nor2_1 _11902_ (.A(_02784_),
    .B(_02806_),
    .Y(_02844_));
 sg13g2_nor2_1 _11903_ (.A(_02736_),
    .B(_02753_),
    .Y(_02845_));
 sg13g2_nand2_1 _11904_ (.Y(_02846_),
    .A(_02806_),
    .B(_02784_));
 sg13g2_nand2_1 _11905_ (.Y(_02847_),
    .A(_02845_),
    .B(_02846_));
 sg13g2_nand2b_1 _11906_ (.Y(_02848_),
    .B(_02847_),
    .A_N(_02844_));
 sg13g2_a21oi_1 _11907_ (.A1(_02843_),
    .A2(_02756_),
    .Y(_02849_),
    .B1(_02848_));
 sg13g2_nand3_1 _11908_ (.B(_02730_),
    .C(_02759_),
    .A(_02843_),
    .Y(_02850_));
 sg13g2_nand2_1 _11909_ (.Y(_02851_),
    .A(_02849_),
    .B(_02850_));
 sg13g2_xnor2_1 _11910_ (.Y(_02852_),
    .A(_02842_),
    .B(_02851_));
 sg13g2_nand2_1 _11911_ (.Y(_02853_),
    .A(_02852_),
    .B(_02768_));
 sg13g2_nand2_1 _11912_ (.Y(_02854_),
    .A(_02851_),
    .B(_02842_));
 sg13g2_nand3_1 _11913_ (.B(_02850_),
    .C(_02841_),
    .A(_02849_),
    .Y(_02855_));
 sg13g2_nand3_1 _11914_ (.B(_02854_),
    .C(_02855_),
    .A(_02763_),
    .Y(_02856_));
 sg13g2_buf_1 _11915_ (.A(_02856_),
    .X(_02857_));
 sg13g2_nand3_1 _11916_ (.B(_02853_),
    .C(_02857_),
    .A(_02821_),
    .Y(_02858_));
 sg13g2_nand2_1 _11917_ (.Y(_02859_),
    .A(_02853_),
    .B(_02857_));
 sg13g2_nand2_1 _11918_ (.Y(_02860_),
    .A(_02859_),
    .B(_02820_));
 sg13g2_nand2_1 _11919_ (.Y(_02861_),
    .A(_02858_),
    .B(_02860_));
 sg13g2_nor2_1 _11920_ (.A(_02656_),
    .B(_02728_),
    .Y(_02862_));
 sg13g2_nand3_1 _11921_ (.B(_02727_),
    .C(_02653_),
    .A(_02862_),
    .Y(_02863_));
 sg13g2_nand2_1 _11922_ (.Y(_02864_),
    .A(_02863_),
    .B(_02775_));
 sg13g2_nand2_1 _11923_ (.Y(_02865_),
    .A(_02842_),
    .B(_02809_));
 sg13g2_nor2_1 _11924_ (.A(_02776_),
    .B(_02865_),
    .Y(_02866_));
 sg13g2_nand2_1 _11925_ (.Y(_02867_),
    .A(_02864_),
    .B(_02866_));
 sg13g2_nor2_1 _11926_ (.A(_02807_),
    .B(_02841_),
    .Y(_02868_));
 sg13g2_nor2_1 _11927_ (.A(_02823_),
    .B(_02840_),
    .Y(_02869_));
 sg13g2_nor2_1 _11928_ (.A(_02844_),
    .B(_02869_),
    .Y(_02870_));
 sg13g2_nand2_1 _11929_ (.Y(_02871_),
    .A(_02840_),
    .B(_02823_));
 sg13g2_nor2b_1 _11930_ (.A(_02870_),
    .B_N(_02871_),
    .Y(_02872_));
 sg13g2_a21oi_1 _11931_ (.A1(_02868_),
    .A2(_02774_),
    .Y(_02873_),
    .B1(_02872_));
 sg13g2_nand2_1 _11932_ (.Y(_02874_),
    .A(_02867_),
    .B(_02873_));
 sg13g2_inv_1 _11933_ (.Y(_02875_),
    .A(_02833_));
 sg13g2_a21oi_2 _11934_ (.B1(_02875_),
    .Y(_02876_),
    .A2(_02824_),
    .A1(_02836_));
 sg13g2_xnor2_1 _11935_ (.Y(_02877_),
    .A(net101),
    .B(_02205_));
 sg13g2_xnor2_1 _11936_ (.Y(_02878_),
    .A(net214),
    .B(_02273_));
 sg13g2_nor2_1 _11937_ (.A(_02210_),
    .B(_02578_),
    .Y(_02879_));
 sg13g2_inv_1 _11938_ (.Y(_02880_),
    .A(_02879_));
 sg13g2_nor2_1 _11939_ (.A(_02788_),
    .B(_02880_),
    .Y(_02881_));
 sg13g2_inv_1 _11940_ (.Y(_02882_),
    .A(_02207_));
 sg13g2_a21oi_1 _11941_ (.A1(_02295_),
    .A2(_02209_),
    .Y(_02883_),
    .B1(_02882_));
 sg13g2_nand2_1 _11942_ (.Y(_02884_),
    .A(_02879_),
    .B(_02791_));
 sg13g2_nand2b_1 _11943_ (.Y(_02885_),
    .B(_02884_),
    .A_N(_02883_));
 sg13g2_a21oi_1 _11944_ (.A1(_02690_),
    .A2(_02881_),
    .Y(_02886_),
    .B1(_02885_));
 sg13g2_nand3_1 _11945_ (.B(_02694_),
    .C(_02693_),
    .A(_02881_),
    .Y(_02887_));
 sg13g2_nand2_1 _11946_ (.Y(_02888_),
    .A(_02886_),
    .B(_02887_));
 sg13g2_xnor2_1 _11947_ (.Y(_02889_),
    .A(_02243_),
    .B(_02888_));
 sg13g2_nand2_1 _11948_ (.Y(_02890_),
    .A(_02889_),
    .B(net72));
 sg13g2_xor2_1 _11949_ (.B(_02888_),
    .A(_02243_),
    .X(_02891_));
 sg13g2_nand2_1 _11950_ (.Y(_02892_),
    .A(_02891_),
    .B(net73));
 sg13g2_nand2_1 _11951_ (.Y(_02893_),
    .A(_02890_),
    .B(_02892_));
 sg13g2_nand2b_1 _11952_ (.Y(_02894_),
    .B(_02893_),
    .A_N(_02878_));
 sg13g2_nand3_1 _11953_ (.B(_02892_),
    .C(_02878_),
    .A(_02890_),
    .Y(_02895_));
 sg13g2_buf_1 _11954_ (.A(_02895_),
    .X(_02896_));
 sg13g2_nand2_1 _11955_ (.Y(_02897_),
    .A(_02894_),
    .B(_02896_));
 sg13g2_nand2b_1 _11956_ (.Y(_02898_),
    .B(_02897_),
    .A_N(_02877_));
 sg13g2_nand3_1 _11957_ (.B(_02896_),
    .C(_02877_),
    .A(_02894_),
    .Y(_02899_));
 sg13g2_nand2_1 _11958_ (.Y(_02900_),
    .A(_02898_),
    .B(_02899_));
 sg13g2_xnor2_1 _11959_ (.Y(_02901_),
    .A(_02876_),
    .B(_02900_));
 sg13g2_buf_2 _11960_ (.A(_02901_),
    .X(_02902_));
 sg13g2_nand2_1 _11961_ (.Y(_02903_),
    .A(_02874_),
    .B(_02902_));
 sg13g2_inv_1 _11962_ (.Y(_02904_),
    .A(_02902_));
 sg13g2_nand3_1 _11963_ (.B(_02904_),
    .C(_02873_),
    .A(_02867_),
    .Y(_02905_));
 sg13g2_nand2_1 _11964_ (.Y(_02906_),
    .A(_02903_),
    .B(_02905_));
 sg13g2_nand2_1 _11965_ (.Y(_02907_),
    .A(_02906_),
    .B(_02811_));
 sg13g2_nand2_1 _11966_ (.Y(_02908_),
    .A(_02874_),
    .B(_02904_));
 sg13g2_nand3_1 _11967_ (.B(_02902_),
    .C(_02873_),
    .A(_02867_),
    .Y(_02909_));
 sg13g2_nand2_1 _11968_ (.Y(_02910_),
    .A(_02908_),
    .B(_02909_));
 sg13g2_xnor2_1 _11969_ (.Y(_02911_),
    .A(_02809_),
    .B(_02782_));
 sg13g2_nand2_1 _11970_ (.Y(_02912_),
    .A(_02910_),
    .B(_02911_));
 sg13g2_nand3b_1 _11971_ (.B(_02907_),
    .C(_02912_),
    .Y(_02913_),
    .A_N(_02857_));
 sg13g2_buf_1 _11972_ (.A(_02913_),
    .X(_02914_));
 sg13g2_nand2_1 _11973_ (.Y(_02915_),
    .A(_02906_),
    .B(_02911_));
 sg13g2_nand2_1 _11974_ (.Y(_02916_),
    .A(_02910_),
    .B(_02811_));
 sg13g2_nand3_1 _11975_ (.B(_02916_),
    .C(_02857_),
    .A(_02915_),
    .Y(_02917_));
 sg13g2_nand2_1 _11976_ (.Y(_02918_),
    .A(_02914_),
    .B(_02917_));
 sg13g2_nor2_1 _11977_ (.A(_02861_),
    .B(_02918_),
    .Y(_02919_));
 sg13g2_nand2_1 _11978_ (.Y(_02920_),
    .A(_02819_),
    .B(_02919_));
 sg13g2_inv_1 _11979_ (.Y(_02921_),
    .A(_02858_));
 sg13g2_inv_1 _11980_ (.Y(_02922_),
    .A(_02914_));
 sg13g2_a21oi_1 _11981_ (.A1(_02921_),
    .A2(_02917_),
    .Y(_02923_),
    .B1(_02922_));
 sg13g2_nand2_1 _11982_ (.Y(_02924_),
    .A(_02920_),
    .B(_02923_));
 sg13g2_inv_1 _11983_ (.Y(_02925_),
    .A(_02907_));
 sg13g2_inv_1 _11984_ (.Y(_02926_),
    .A(_02894_));
 sg13g2_a21oi_2 _11985_ (.B1(_02926_),
    .Y(_02927_),
    .A2(_02877_),
    .A1(_02896_));
 sg13g2_xnor2_1 _11986_ (.Y(_02928_),
    .A(net94),
    .B(_02239_));
 sg13g2_xnor2_1 _11987_ (.Y(_02929_),
    .A(net186),
    .B(_02286_));
 sg13g2_nand2b_1 _11988_ (.Y(_02930_),
    .B(_02574_),
    .A_N(_02580_));
 sg13g2_nand2b_1 _11989_ (.Y(_02931_),
    .B(_02930_),
    .A_N(_02301_));
 sg13g2_xnor2_1 _11990_ (.Y(_02932_),
    .A(_02581_),
    .B(_02931_));
 sg13g2_xnor2_1 _11991_ (.Y(_02933_),
    .A(net71),
    .B(_02932_));
 sg13g2_xnor2_1 _11992_ (.Y(_02934_),
    .A(_02929_),
    .B(_02933_));
 sg13g2_xnor2_1 _11993_ (.Y(_02935_),
    .A(_02928_),
    .B(_02934_));
 sg13g2_xnor2_1 _11994_ (.Y(_02936_),
    .A(_02927_),
    .B(_02935_));
 sg13g2_nor2_1 _11995_ (.A(_02876_),
    .B(_02900_),
    .Y(_02937_));
 sg13g2_nor2_1 _11996_ (.A(_02869_),
    .B(_02937_),
    .Y(_02938_));
 sg13g2_nand2_1 _11997_ (.Y(_02939_),
    .A(_02900_),
    .B(_02876_));
 sg13g2_nor2b_1 _11998_ (.A(_02938_),
    .B_N(_02939_),
    .Y(_02940_));
 sg13g2_nor2_1 _11999_ (.A(_02841_),
    .B(_02902_),
    .Y(_02941_));
 sg13g2_nand2_1 _12000_ (.Y(_02942_),
    .A(_02941_),
    .B(_02848_));
 sg13g2_nand2b_1 _12001_ (.Y(_02943_),
    .B(_02942_),
    .A_N(_02940_));
 sg13g2_inv_1 _12002_ (.Y(_02944_),
    .A(_02941_));
 sg13g2_nor2b_1 _12003_ (.A(_02944_),
    .B_N(_02843_),
    .Y(_02945_));
 sg13g2_nand2_1 _12004_ (.Y(_02946_),
    .A(_02762_),
    .B(_02945_));
 sg13g2_nand2b_1 _12005_ (.Y(_02947_),
    .B(_02946_),
    .A_N(_02943_));
 sg13g2_xnor2_1 _12006_ (.Y(_02948_),
    .A(_02936_),
    .B(_02947_));
 sg13g2_xnor2_1 _12007_ (.Y(_02949_),
    .A(_02852_),
    .B(_02948_));
 sg13g2_nor2_1 _12008_ (.A(_02925_),
    .B(_02949_),
    .Y(_02950_));
 sg13g2_nand2_1 _12009_ (.Y(_02951_),
    .A(_02949_),
    .B(_02925_));
 sg13g2_nand2b_1 _12010_ (.Y(_02952_),
    .B(_02951_),
    .A_N(_02950_));
 sg13g2_nand2_1 _12011_ (.Y(_02953_),
    .A(_02924_),
    .B(_02952_));
 sg13g2_nor2b_1 _12012_ (.A(_02950_),
    .B_N(_02951_),
    .Y(_02954_));
 sg13g2_nand3_1 _12013_ (.B(_02954_),
    .C(_02923_),
    .A(_02920_),
    .Y(_02955_));
 sg13g2_nand2_1 _12014_ (.Y(_02956_),
    .A(_02953_),
    .B(_02955_));
 sg13g2_buf_1 _12015_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[6] ),
    .X(_02957_));
 sg13g2_nand2_1 _12016_ (.Y(_02958_),
    .A(_02956_),
    .B(_02957_));
 sg13g2_inv_1 _12017_ (.Y(_02959_),
    .A(_02957_));
 sg13g2_nand3_1 _12018_ (.B(_02955_),
    .C(_02959_),
    .A(_02953_),
    .Y(_02960_));
 sg13g2_buf_1 _12019_ (.A(_02960_),
    .X(_02961_));
 sg13g2_nand2_1 _12020_ (.Y(_02962_),
    .A(_02958_),
    .B(_02961_));
 sg13g2_buf_2 _12021_ (.A(_02962_),
    .X(_02963_));
 sg13g2_buf_1 _12022_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[5] ),
    .X(_02964_));
 sg13g2_inv_1 _12023_ (.Y(_02965_),
    .A(_02918_));
 sg13g2_xnor2_1 _12024_ (.Y(_02966_),
    .A(_02821_),
    .B(_02859_));
 sg13g2_nand2_1 _12025_ (.Y(_02967_),
    .A(_02813_),
    .B(_02815_));
 sg13g2_xnor2_1 _12026_ (.Y(_02968_),
    .A(_02765_),
    .B(_02967_));
 sg13g2_nand3_1 _12027_ (.B(_02968_),
    .C(_02771_),
    .A(_02966_),
    .Y(_02969_));
 sg13g2_a21oi_1 _12028_ (.A1(_02860_),
    .A2(_02817_),
    .Y(_02970_),
    .B1(_02921_));
 sg13g2_nand2_1 _12029_ (.Y(_02971_),
    .A(_02969_),
    .B(_02970_));
 sg13g2_xnor2_1 _12030_ (.Y(_02972_),
    .A(_02965_),
    .B(_02971_));
 sg13g2_nor2_1 _12031_ (.A(_02964_),
    .B(_02972_),
    .Y(_02973_));
 sg13g2_nand2_1 _12032_ (.Y(_02974_),
    .A(_02963_),
    .B(_02973_));
 sg13g2_nand2_1 _12033_ (.Y(_02975_),
    .A(_02956_),
    .B(_02959_));
 sg13g2_nand2_1 _12034_ (.Y(_02976_),
    .A(_02974_),
    .B(_02975_));
 sg13g2_inv_1 _12035_ (.Y(_02977_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[4] ));
 sg13g2_xnor2_1 _12036_ (.Y(_02978_),
    .A(_02861_),
    .B(_02818_));
 sg13g2_xnor2_1 _12037_ (.Y(_02979_),
    .A(_02977_),
    .B(_02978_));
 sg13g2_buf_2 _12038_ (.A(_02979_),
    .X(_02980_));
 sg13g2_inv_1 _12039_ (.Y(_02981_),
    .A(_02968_));
 sg13g2_nand2b_1 _12040_ (.Y(_02982_),
    .B(_02981_),
    .A_N(_02771_));
 sg13g2_buf_1 _12041_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[3] ),
    .X(_02983_));
 sg13g2_inv_1 _12042_ (.Y(_02984_),
    .A(_02983_));
 sg13g2_nand2_1 _12043_ (.Y(_02985_),
    .A(_02968_),
    .B(_02771_));
 sg13g2_nand3_1 _12044_ (.B(_02984_),
    .C(_02985_),
    .A(_02982_),
    .Y(_02986_));
 sg13g2_inv_1 _12045_ (.Y(_02987_),
    .A(_02986_));
 sg13g2_nor2_1 _12046_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[4] ),
    .B(_02978_),
    .Y(_02988_));
 sg13g2_a21oi_1 _12047_ (.A1(_02980_),
    .A2(_02987_),
    .Y(_02989_),
    .B1(_02988_));
 sg13g2_xnor2_1 _12048_ (.Y(_02990_),
    .A(_00160_),
    .B(_02972_));
 sg13g2_nand2_1 _12049_ (.Y(_02991_),
    .A(_02963_),
    .B(_02990_));
 sg13g2_nor2_1 _12050_ (.A(_02989_),
    .B(_02991_),
    .Y(_02992_));
 sg13g2_nor2_1 _12051_ (.A(_02976_),
    .B(_02992_),
    .Y(_02993_));
 sg13g2_buf_2 _12052_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[2] ),
    .X(_02994_));
 sg13g2_xnor2_1 _12053_ (.Y(_02995_),
    .A(_02721_),
    .B(_02770_));
 sg13g2_nand2_1 _12054_ (.Y(_02996_),
    .A(_02995_),
    .B(_02734_));
 sg13g2_nor2_1 _12055_ (.A(_02770_),
    .B(_02734_),
    .Y(_02997_));
 sg13g2_inv_1 _12056_ (.Y(_02998_),
    .A(_02997_));
 sg13g2_nand2_1 _12057_ (.Y(_02999_),
    .A(_02996_),
    .B(_02998_));
 sg13g2_buf_1 _12058_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[1] ),
    .X(_03000_));
 sg13g2_inv_1 _12059_ (.Y(_03001_),
    .A(_03000_));
 sg13g2_a21oi_1 _12060_ (.A1(_02721_),
    .A2(_02722_),
    .Y(_03002_),
    .B1(_02732_));
 sg13g2_nand2b_1 _12061_ (.Y(_03003_),
    .B(_02734_),
    .A_N(_03002_));
 sg13g2_nor2_1 _12062_ (.A(_03001_),
    .B(_03003_),
    .Y(_03004_));
 sg13g2_nand2_1 _12063_ (.Y(_03005_),
    .A(_03003_),
    .B(_03001_));
 sg13g2_nand2b_1 _12064_ (.Y(_03006_),
    .B(_03005_),
    .A_N(_03004_));
 sg13g2_xnor2_1 _12065_ (.Y(_03007_),
    .A(_02723_),
    .B(_02731_));
 sg13g2_inv_1 _12066_ (.Y(_03008_),
    .A(_00163_));
 sg13g2_nand2_1 _12067_ (.Y(_03009_),
    .A(_03007_),
    .B(_03008_));
 sg13g2_nor2_1 _12068_ (.A(_03000_),
    .B(_03003_),
    .Y(_03010_));
 sg13g2_a21oi_1 _12069_ (.A1(_03006_),
    .A2(_03009_),
    .Y(_03011_),
    .B1(_03010_));
 sg13g2_xnor2_1 _12070_ (.Y(_03012_),
    .A(_00162_),
    .B(_02999_));
 sg13g2_nand2b_1 _12071_ (.Y(_03013_),
    .B(_03012_),
    .A_N(_03011_));
 sg13g2_o21ai_1 _12072_ (.B1(_03013_),
    .Y(_03014_),
    .A1(_02994_),
    .A2(_02999_));
 sg13g2_nand2_1 _12073_ (.Y(_03015_),
    .A(_02982_),
    .B(_02985_));
 sg13g2_xor2_1 _12074_ (.B(_03015_),
    .A(_00161_),
    .X(_03016_));
 sg13g2_inv_2 _12075_ (.Y(_03017_),
    .A(_02980_));
 sg13g2_nor2_1 _12076_ (.A(_03016_),
    .B(_03017_),
    .Y(_03018_));
 sg13g2_nand4_1 _12077_ (.B(_02990_),
    .C(_03014_),
    .A(_02963_),
    .Y(_03019_),
    .D(_03018_));
 sg13g2_nand2_1 _12078_ (.Y(_03020_),
    .A(_02993_),
    .B(_03019_));
 sg13g2_xor2_1 _12079_ (.B(_02935_),
    .A(_02927_),
    .X(_03021_));
 sg13g2_nand2_1 _12080_ (.Y(_03022_),
    .A(_03021_),
    .B(_02904_));
 sg13g2_nor2_1 _12081_ (.A(_02865_),
    .B(_03022_),
    .Y(_03023_));
 sg13g2_nand2_1 _12082_ (.Y(_03024_),
    .A(_02782_),
    .B(_03023_));
 sg13g2_nor2_1 _12083_ (.A(_02902_),
    .B(_02936_),
    .Y(_03025_));
 sg13g2_nor2_1 _12084_ (.A(_02927_),
    .B(_02935_),
    .Y(_03026_));
 sg13g2_nand2_1 _12085_ (.Y(_03027_),
    .A(_02935_),
    .B(_02927_));
 sg13g2_nand2_1 _12086_ (.Y(_03028_),
    .A(_03027_),
    .B(_02937_));
 sg13g2_nand2b_1 _12087_ (.Y(_03029_),
    .B(_03028_),
    .A_N(_03026_));
 sg13g2_a21oi_2 _12088_ (.B1(_03029_),
    .Y(_03030_),
    .A2(_02872_),
    .A1(_03025_));
 sg13g2_nand2_1 _12089_ (.Y(_03031_),
    .A(_03024_),
    .B(_03030_));
 sg13g2_inv_1 _12090_ (.Y(_03032_),
    .A(_02929_));
 sg13g2_nand2_1 _12091_ (.Y(_03033_),
    .A(_02933_),
    .B(_03032_));
 sg13g2_nor2_1 _12092_ (.A(_03032_),
    .B(_02933_),
    .Y(_03034_));
 sg13g2_a21oi_2 _12093_ (.B1(_03034_),
    .Y(_03035_),
    .A2(_02928_),
    .A1(_03033_));
 sg13g2_xnor2_1 _12094_ (.Y(_03036_),
    .A(net101),
    .B(_02355_));
 sg13g2_buf_1 _12095_ (.A(net214),
    .X(_03037_));
 sg13g2_xnor2_1 _12096_ (.Y(_03038_),
    .A(_03037_),
    .B(_02159_));
 sg13g2_nor2_1 _12097_ (.A(_02243_),
    .B(_02581_),
    .Y(_03039_));
 sg13g2_inv_1 _12098_ (.Y(_03040_),
    .A(_03039_));
 sg13g2_nor2_1 _12099_ (.A(_02880_),
    .B(_03040_),
    .Y(_03041_));
 sg13g2_nand2_1 _12100_ (.Y(_03042_),
    .A(_03039_),
    .B(_02883_));
 sg13g2_nand2_1 _12101_ (.Y(_03043_),
    .A(_02359_),
    .B(_02415_));
 sg13g2_a21oi_1 _12102_ (.A1(_02299_),
    .A2(_03043_),
    .Y(_03044_),
    .B1(_02416_));
 sg13g2_nand2_1 _12103_ (.Y(_03045_),
    .A(_03042_),
    .B(_03044_));
 sg13g2_a21oi_1 _12104_ (.A1(_02793_),
    .A2(_03041_),
    .Y(_03046_),
    .B1(_03045_));
 sg13g2_nand3_1 _12105_ (.B(_02606_),
    .C(_02789_),
    .A(_03041_),
    .Y(_03047_));
 sg13g2_nand2_1 _12106_ (.Y(_03048_),
    .A(_03046_),
    .B(_03047_));
 sg13g2_xnor2_1 _12107_ (.Y(_03049_),
    .A(_02582_),
    .B(_03048_));
 sg13g2_inv_1 _12108_ (.Y(_03050_),
    .A(_03049_));
 sg13g2_nand2_1 _12109_ (.Y(_03051_),
    .A(_03050_),
    .B(net73));
 sg13g2_nand2_1 _12110_ (.Y(_03052_),
    .A(_03049_),
    .B(net72));
 sg13g2_nand2_1 _12111_ (.Y(_03053_),
    .A(_03051_),
    .B(_03052_));
 sg13g2_nand2b_1 _12112_ (.Y(_03054_),
    .B(_03053_),
    .A_N(_03038_));
 sg13g2_nand3_1 _12113_ (.B(_03052_),
    .C(_03038_),
    .A(_03051_),
    .Y(_03055_));
 sg13g2_buf_1 _12114_ (.A(_03055_),
    .X(_03056_));
 sg13g2_nand2_1 _12115_ (.Y(_03057_),
    .A(_03054_),
    .B(_03056_));
 sg13g2_nand2b_1 _12116_ (.Y(_03058_),
    .B(_03057_),
    .A_N(_03036_));
 sg13g2_nand3_1 _12117_ (.B(_03056_),
    .C(_03036_),
    .A(_03054_),
    .Y(_03059_));
 sg13g2_nand2_1 _12118_ (.Y(_03060_),
    .A(_03058_),
    .B(_03059_));
 sg13g2_xnor2_1 _12119_ (.Y(_03061_),
    .A(_03035_),
    .B(_03060_));
 sg13g2_buf_1 _12120_ (.A(_03061_),
    .X(_03062_));
 sg13g2_inv_1 _12121_ (.Y(_03063_),
    .A(_03062_));
 sg13g2_nand2_1 _12122_ (.Y(_03064_),
    .A(_03031_),
    .B(_03063_));
 sg13g2_nand3_1 _12123_ (.B(_03062_),
    .C(_03030_),
    .A(_03024_),
    .Y(_03065_));
 sg13g2_nand2_1 _12124_ (.Y(_03066_),
    .A(_03064_),
    .B(_03065_));
 sg13g2_nand2_1 _12125_ (.Y(_03067_),
    .A(_03066_),
    .B(_02906_));
 sg13g2_nand2_1 _12126_ (.Y(_03068_),
    .A(_03031_),
    .B(_03062_));
 sg13g2_nand3_1 _12127_ (.B(_03063_),
    .C(_03030_),
    .A(_03024_),
    .Y(_03069_));
 sg13g2_nand2_1 _12128_ (.Y(_03070_),
    .A(_03068_),
    .B(_03069_));
 sg13g2_nand2_1 _12129_ (.Y(_03071_),
    .A(_03070_),
    .B(_02910_));
 sg13g2_nand2_1 _12130_ (.Y(_03072_),
    .A(_03067_),
    .B(_03071_));
 sg13g2_inv_1 _12131_ (.Y(_03073_),
    .A(_02948_));
 sg13g2_nor2_1 _12132_ (.A(_02852_),
    .B(_03073_),
    .Y(_03074_));
 sg13g2_nand2_1 _12133_ (.Y(_03075_),
    .A(_03072_),
    .B(_03074_));
 sg13g2_inv_1 _12134_ (.Y(_03076_),
    .A(_03074_));
 sg13g2_nand3_1 _12135_ (.B(_03067_),
    .C(_03071_),
    .A(_03076_),
    .Y(_03077_));
 sg13g2_nand2_1 _12136_ (.Y(_03078_),
    .A(_03075_),
    .B(_03077_));
 sg13g2_nor2_1 _12137_ (.A(_03078_),
    .B(_02952_),
    .Y(_03079_));
 sg13g2_nand2_1 _12138_ (.Y(_03080_),
    .A(_02924_),
    .B(_03079_));
 sg13g2_nand2_1 _12139_ (.Y(_03081_),
    .A(_03075_),
    .B(_02951_));
 sg13g2_nand2_1 _12140_ (.Y(_03082_),
    .A(_03081_),
    .B(_03077_));
 sg13g2_nand2_1 _12141_ (.Y(_03083_),
    .A(_03080_),
    .B(_03082_));
 sg13g2_inv_1 _12142_ (.Y(_03084_),
    .A(_03054_));
 sg13g2_a21oi_2 _12143_ (.B1(_03084_),
    .Y(_03085_),
    .A2(_03036_),
    .A1(_03056_));
 sg13g2_xnor2_1 _12144_ (.Y(_03086_),
    .A(net94),
    .B(_02326_));
 sg13g2_nand2_1 _12145_ (.Y(_03087_),
    .A(_02579_),
    .B(_02522_));
 sg13g2_nand2b_1 _12146_ (.Y(_03088_),
    .B(_03087_),
    .A_N(_02296_));
 sg13g2_nand2_1 _12147_ (.Y(_03089_),
    .A(_02583_),
    .B(_02244_));
 sg13g2_inv_1 _12148_ (.Y(_03090_),
    .A(_03089_));
 sg13g2_inv_1 _12149_ (.Y(_03091_),
    .A(_02419_));
 sg13g2_o21ai_1 _12150_ (.B1(_03091_),
    .Y(_03092_),
    .A1(_02300_),
    .A2(_02361_));
 sg13g2_a21oi_1 _12151_ (.A1(_03088_),
    .A2(_03090_),
    .Y(_03093_),
    .B1(_03092_));
 sg13g2_nand2_1 _12152_ (.Y(_03094_),
    .A(_02579_),
    .B(_02483_));
 sg13g2_nor2_1 _12153_ (.A(_03094_),
    .B(_03089_),
    .Y(_03095_));
 sg13g2_nand2_1 _12154_ (.Y(_03096_),
    .A(_02662_),
    .B(_03095_));
 sg13g2_nand2_1 _12155_ (.Y(_03097_),
    .A(_03093_),
    .B(_03096_));
 sg13g2_xnor2_1 _12156_ (.Y(_03098_),
    .A(_02408_),
    .B(_03097_));
 sg13g2_nand2_1 _12157_ (.Y(_03099_),
    .A(_03098_),
    .B(net72));
 sg13g2_nand2_1 _12158_ (.Y(_03100_),
    .A(_03097_),
    .B(_02409_));
 sg13g2_nand3_1 _12159_ (.B(_03096_),
    .C(_02408_),
    .A(_03093_),
    .Y(_03101_));
 sg13g2_nand2_1 _12160_ (.Y(_03102_),
    .A(_03100_),
    .B(_03101_));
 sg13g2_nand2_1 _12161_ (.Y(_03103_),
    .A(_03102_),
    .B(net73));
 sg13g2_nand2_1 _12162_ (.Y(_03104_),
    .A(_03099_),
    .B(_03103_));
 sg13g2_xnor2_1 _12163_ (.Y(_03105_),
    .A(net214),
    .B(_02233_));
 sg13g2_inv_1 _12164_ (.Y(_03106_),
    .A(_03105_));
 sg13g2_nand2_1 _12165_ (.Y(_03107_),
    .A(_03104_),
    .B(_03106_));
 sg13g2_nand3_1 _12166_ (.B(_03103_),
    .C(_03105_),
    .A(_03099_),
    .Y(_03108_));
 sg13g2_buf_1 _12167_ (.A(_03108_),
    .X(_03109_));
 sg13g2_nand2_1 _12168_ (.Y(_03110_),
    .A(_03107_),
    .B(_03109_));
 sg13g2_nand2b_1 _12169_ (.Y(_03111_),
    .B(_03110_),
    .A_N(_03086_));
 sg13g2_nand3_1 _12170_ (.B(_03109_),
    .C(_03086_),
    .A(_03107_),
    .Y(_03112_));
 sg13g2_nand2_1 _12171_ (.Y(_03113_),
    .A(_03111_),
    .B(_03112_));
 sg13g2_xnor2_1 _12172_ (.Y(_03114_),
    .A(_03085_),
    .B(_03113_));
 sg13g2_buf_2 _12173_ (.A(_03114_),
    .X(_03115_));
 sg13g2_nand2_1 _12174_ (.Y(_03116_),
    .A(_03063_),
    .B(_03021_));
 sg13g2_nor2_1 _12175_ (.A(_02944_),
    .B(_03116_),
    .Y(_03117_));
 sg13g2_nand2_1 _12176_ (.Y(_03118_),
    .A(_02851_),
    .B(_03117_));
 sg13g2_nor2_1 _12177_ (.A(_03062_),
    .B(_02936_),
    .Y(_03119_));
 sg13g2_nor2_1 _12178_ (.A(_03035_),
    .B(_03060_),
    .Y(_03120_));
 sg13g2_nor2_1 _12179_ (.A(_03120_),
    .B(_03026_),
    .Y(_03121_));
 sg13g2_nand2_1 _12180_ (.Y(_03122_),
    .A(_03060_),
    .B(_03035_));
 sg13g2_nor2b_1 _12181_ (.A(_03121_),
    .B_N(_03122_),
    .Y(_03123_));
 sg13g2_a21oi_1 _12182_ (.A1(_03119_),
    .A2(_02940_),
    .Y(_03124_),
    .B1(_03123_));
 sg13g2_nand2_1 _12183_ (.Y(_03125_),
    .A(_03118_),
    .B(_03124_));
 sg13g2_xnor2_1 _12184_ (.Y(_03126_),
    .A(_03115_),
    .B(_03125_));
 sg13g2_nand2_1 _12185_ (.Y(_03127_),
    .A(_03126_),
    .B(_02948_));
 sg13g2_buf_2 _12186_ (.A(_03127_),
    .X(_03128_));
 sg13g2_nand2b_1 _12187_ (.Y(_03129_),
    .B(_03125_),
    .A_N(_03115_));
 sg13g2_nand3_1 _12188_ (.B(_03115_),
    .C(_03124_),
    .A(_03118_),
    .Y(_03130_));
 sg13g2_nand2_1 _12189_ (.Y(_03131_),
    .A(_03129_),
    .B(_03130_));
 sg13g2_nand2_1 _12190_ (.Y(_03132_),
    .A(_03131_),
    .B(_03073_));
 sg13g2_nand2_1 _12191_ (.Y(_03133_),
    .A(_03128_),
    .B(_03132_));
 sg13g2_nand2_1 _12192_ (.Y(_03134_),
    .A(_03070_),
    .B(_02906_));
 sg13g2_nand2_1 _12193_ (.Y(_03135_),
    .A(_03133_),
    .B(_03134_));
 sg13g2_nor2_1 _12194_ (.A(_02910_),
    .B(_03066_),
    .Y(_03136_));
 sg13g2_nand3_1 _12195_ (.B(_03132_),
    .C(_03136_),
    .A(_03128_),
    .Y(_03137_));
 sg13g2_buf_1 _12196_ (.A(_03137_),
    .X(_03138_));
 sg13g2_nand2_1 _12197_ (.Y(_03139_),
    .A(_03135_),
    .B(_03138_));
 sg13g2_nand2_1 _12198_ (.Y(_03140_),
    .A(_03083_),
    .B(_03139_));
 sg13g2_nand2_1 _12199_ (.Y(_03141_),
    .A(_03133_),
    .B(_03136_));
 sg13g2_nand3_1 _12200_ (.B(_03132_),
    .C(_03134_),
    .A(_03128_),
    .Y(_03142_));
 sg13g2_nand2_1 _12201_ (.Y(_03143_),
    .A(_03141_),
    .B(_03142_));
 sg13g2_nand3_1 _12202_ (.B(_03143_),
    .C(_03082_),
    .A(_03080_),
    .Y(_03144_));
 sg13g2_nand2_1 _12203_ (.Y(_03145_),
    .A(_03140_),
    .B(_03144_));
 sg13g2_inv_1 _12204_ (.Y(_03146_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[8] ));
 sg13g2_nand2_1 _12205_ (.Y(_03147_),
    .A(_03145_),
    .B(_03146_));
 sg13g2_nand3_1 _12206_ (.B(_03144_),
    .C(\vgadonut.donut.donuthit.cordicxz.xin[8] ),
    .A(_03140_),
    .Y(_03148_));
 sg13g2_nand2_1 _12207_ (.Y(_03149_),
    .A(_03147_),
    .B(_03148_));
 sg13g2_buf_2 _12208_ (.A(_03149_),
    .X(_03150_));
 sg13g2_a21oi_1 _12209_ (.A1(_02951_),
    .A2(_02914_),
    .Y(_03151_),
    .B1(_02950_));
 sg13g2_nor2_1 _12210_ (.A(_02918_),
    .B(_02952_),
    .Y(_03152_));
 sg13g2_nand2_1 _12211_ (.Y(_03153_),
    .A(_03152_),
    .B(_02971_));
 sg13g2_nand2b_1 _12212_ (.Y(_03154_),
    .B(_03153_),
    .A_N(_03151_));
 sg13g2_xor2_1 _12213_ (.B(_03154_),
    .A(_03078_),
    .X(_03155_));
 sg13g2_xor2_1 _12214_ (.B(_03155_),
    .A(_00159_),
    .X(_03156_));
 sg13g2_nor2_1 _12215_ (.A(_03150_),
    .B(_03156_),
    .Y(_03157_));
 sg13g2_nand2_1 _12216_ (.Y(_03158_),
    .A(_03020_),
    .B(_03157_));
 sg13g2_nand2_1 _12217_ (.Y(_03159_),
    .A(_02868_),
    .B(_02774_));
 sg13g2_nand2b_1 _12218_ (.Y(_03160_),
    .B(_03159_),
    .A_N(_02872_));
 sg13g2_nor2_1 _12219_ (.A(_03115_),
    .B(_03062_),
    .Y(_03161_));
 sg13g2_inv_1 _12220_ (.Y(_03162_),
    .A(_03161_));
 sg13g2_nor2_1 _12221_ (.A(_03022_),
    .B(_03162_),
    .Y(_03163_));
 sg13g2_nand2_1 _12222_ (.Y(_03164_),
    .A(_03161_),
    .B(_03029_));
 sg13g2_nor2_1 _12223_ (.A(_03085_),
    .B(_03113_),
    .Y(_03165_));
 sg13g2_nand2_1 _12224_ (.Y(_03166_),
    .A(_03113_),
    .B(_03085_));
 sg13g2_o21ai_1 _12225_ (.B1(_03166_),
    .Y(_03167_),
    .A1(_03165_),
    .A2(_03120_));
 sg13g2_nand2_1 _12226_ (.Y(_03168_),
    .A(_03164_),
    .B(_03167_));
 sg13g2_a21oi_1 _12227_ (.A1(_03160_),
    .A2(_03163_),
    .Y(_03169_),
    .B1(_03168_));
 sg13g2_nand3_1 _12228_ (.B(_02864_),
    .C(_02866_),
    .A(_03163_),
    .Y(_03170_));
 sg13g2_buf_1 _12229_ (.A(_03170_),
    .X(_03171_));
 sg13g2_nand2_1 _12230_ (.Y(_03172_),
    .A(_03169_),
    .B(_03171_));
 sg13g2_inv_1 _12231_ (.Y(_03173_),
    .A(_03107_));
 sg13g2_a21oi_1 _12232_ (.A1(_03109_),
    .A2(_03086_),
    .Y(_03174_),
    .B1(_03173_));
 sg13g2_inv_1 _12233_ (.Y(_03175_),
    .A(_03174_));
 sg13g2_xnor2_1 _12234_ (.Y(_03176_),
    .A(net94),
    .B(_02403_));
 sg13g2_xnor2_1 _12235_ (.Y(_03177_),
    .A(_03037_),
    .B(_02358_));
 sg13g2_nor2_1 _12236_ (.A(_02582_),
    .B(_02408_),
    .Y(_03178_));
 sg13g2_nand2_1 _12237_ (.Y(_03179_),
    .A(_03178_),
    .B(_03039_));
 sg13g2_inv_1 _12238_ (.Y(_03180_),
    .A(_03179_));
 sg13g2_nand2b_1 _12239_ (.Y(_03181_),
    .B(_03178_),
    .A_N(_03044_));
 sg13g2_inv_1 _12240_ (.Y(_03182_),
    .A(_02418_));
 sg13g2_a21oi_1 _12241_ (.A1(_03182_),
    .A2(_02407_),
    .Y(_03183_),
    .B1(_02421_));
 sg13g2_nand2_1 _12242_ (.Y(_03184_),
    .A(_03181_),
    .B(_03183_));
 sg13g2_a21oi_1 _12243_ (.A1(_03180_),
    .A2(_02885_),
    .Y(_03185_),
    .B1(_03184_));
 sg13g2_nor2b_1 _12244_ (.A(_03179_),
    .B_N(_02881_),
    .Y(_03186_));
 sg13g2_nand2_1 _12245_ (.Y(_03187_),
    .A(_02696_),
    .B(_03186_));
 sg13g2_nand2_1 _12246_ (.Y(_03188_),
    .A(_03185_),
    .B(_03187_));
 sg13g2_xor2_1 _12247_ (.B(_03188_),
    .A(_02396_),
    .X(_03189_));
 sg13g2_nand2_1 _12248_ (.Y(_03190_),
    .A(_03189_),
    .B(net71));
 sg13g2_xnor2_1 _12249_ (.Y(_03191_),
    .A(_02396_),
    .B(_03188_));
 sg13g2_nand2_1 _12250_ (.Y(_03192_),
    .A(_03191_),
    .B(net72));
 sg13g2_nand2_1 _12251_ (.Y(_03193_),
    .A(_03190_),
    .B(_03192_));
 sg13g2_nand2b_1 _12252_ (.Y(_03194_),
    .B(_03193_),
    .A_N(_03177_));
 sg13g2_nand3_1 _12253_ (.B(_03192_),
    .C(_03177_),
    .A(_03190_),
    .Y(_03195_));
 sg13g2_buf_1 _12254_ (.A(_03195_),
    .X(_03196_));
 sg13g2_nand2_1 _12255_ (.Y(_03197_),
    .A(_03194_),
    .B(_03196_));
 sg13g2_nand2b_1 _12256_ (.Y(_03198_),
    .B(_03197_),
    .A_N(_03176_));
 sg13g2_nand3_1 _12257_ (.B(_03196_),
    .C(_03176_),
    .A(_03194_),
    .Y(_03199_));
 sg13g2_nand2_1 _12258_ (.Y(_03200_),
    .A(_03198_),
    .B(_03199_));
 sg13g2_xnor2_1 _12259_ (.Y(_03201_),
    .A(_03175_),
    .B(_03200_));
 sg13g2_nand2_1 _12260_ (.Y(_03202_),
    .A(_03172_),
    .B(_03201_));
 sg13g2_nand3_1 _12261_ (.B(_03175_),
    .C(_03199_),
    .A(_03198_),
    .Y(_03203_));
 sg13g2_nand2_1 _12262_ (.Y(_03204_),
    .A(_03200_),
    .B(_03174_));
 sg13g2_nand2_1 _12263_ (.Y(_03205_),
    .A(_03203_),
    .B(_03204_));
 sg13g2_nand3_1 _12264_ (.B(_03205_),
    .C(_03171_),
    .A(_03169_),
    .Y(_03206_));
 sg13g2_nand2_1 _12265_ (.Y(_03207_),
    .A(_03202_),
    .B(_03206_));
 sg13g2_nand2_1 _12266_ (.Y(_03208_),
    .A(_03207_),
    .B(_03066_));
 sg13g2_buf_2 _12267_ (.A(_03208_),
    .X(_03209_));
 sg13g2_nand2_1 _12268_ (.Y(_03210_),
    .A(_03172_),
    .B(_03205_));
 sg13g2_nand3_1 _12269_ (.B(_03201_),
    .C(_03171_),
    .A(_03169_),
    .Y(_03211_));
 sg13g2_nand2_1 _12270_ (.Y(_03212_),
    .A(_03210_),
    .B(_03211_));
 sg13g2_nand2_1 _12271_ (.Y(_03213_),
    .A(_03212_),
    .B(_03070_));
 sg13g2_nand2_1 _12272_ (.Y(_03214_),
    .A(_03209_),
    .B(_03213_));
 sg13g2_inv_1 _12273_ (.Y(_03215_),
    .A(_03128_));
 sg13g2_nand2_1 _12274_ (.Y(_03216_),
    .A(_03214_),
    .B(_03215_));
 sg13g2_nand3_1 _12275_ (.B(_03209_),
    .C(_03213_),
    .A(_03128_),
    .Y(_03217_));
 sg13g2_nand2_1 _12276_ (.Y(_03218_),
    .A(_03216_),
    .B(_03217_));
 sg13g2_nor2_1 _12277_ (.A(_03139_),
    .B(_03218_),
    .Y(_03219_));
 sg13g2_nand3_1 _12278_ (.B(_03219_),
    .C(_03079_),
    .A(_02924_),
    .Y(_03220_));
 sg13g2_xnor2_1 _12279_ (.Y(_03221_),
    .A(_03128_),
    .B(_03214_));
 sg13g2_nand2_1 _12280_ (.Y(_03222_),
    .A(_03221_),
    .B(_03143_));
 sg13g2_nor2_1 _12281_ (.A(_03082_),
    .B(_03222_),
    .Y(_03223_));
 sg13g2_nand2_1 _12282_ (.Y(_03224_),
    .A(_03216_),
    .B(_03138_));
 sg13g2_nand2_1 _12283_ (.Y(_03225_),
    .A(_03224_),
    .B(_03217_));
 sg13g2_nor2b_1 _12284_ (.A(_03223_),
    .B_N(_03225_),
    .Y(_03226_));
 sg13g2_nand2_1 _12285_ (.Y(_03227_),
    .A(_03220_),
    .B(_03226_));
 sg13g2_buf_1 _12286_ (.A(net186),
    .X(_03228_));
 sg13g2_xnor2_1 _12287_ (.Y(_03229_),
    .A(net178),
    .B(_02350_));
 sg13g2_xnor2_1 _12288_ (.Y(_03230_),
    .A(net94),
    .B(_02387_));
 sg13g2_xnor2_1 _12289_ (.Y(_03231_),
    .A(_03229_),
    .B(_03230_));
 sg13g2_inv_1 _12290_ (.Y(_03232_),
    .A(_03194_));
 sg13g2_a21oi_1 _12291_ (.A1(_03196_),
    .A2(_03176_),
    .Y(_03233_),
    .B1(_03232_));
 sg13g2_nor2_1 _12292_ (.A(_03231_),
    .B(_03233_),
    .Y(_03234_));
 sg13g2_nand2_1 _12293_ (.Y(_03235_),
    .A(_03233_),
    .B(_03231_));
 sg13g2_nor2b_1 _12294_ (.A(_03234_),
    .B_N(_03235_),
    .Y(_03236_));
 sg13g2_buf_2 _12295_ (.A(_03236_),
    .X(_03237_));
 sg13g2_nor2_1 _12296_ (.A(_03115_),
    .B(_03205_),
    .Y(_03238_));
 sg13g2_inv_1 _12297_ (.Y(_03239_),
    .A(_03238_));
 sg13g2_nor2_1 _12298_ (.A(_03116_),
    .B(_03239_),
    .Y(_03240_));
 sg13g2_nand2_1 _12299_ (.Y(_03241_),
    .A(_03238_),
    .B(_03123_));
 sg13g2_inv_1 _12300_ (.Y(_03242_),
    .A(_03203_));
 sg13g2_o21ai_1 _12301_ (.B1(_03204_),
    .Y(_03243_),
    .A1(_03165_),
    .A2(_03242_));
 sg13g2_nand2_1 _12302_ (.Y(_03244_),
    .A(_03241_),
    .B(_03243_));
 sg13g2_a21oi_1 _12303_ (.A1(_02943_),
    .A2(_03240_),
    .Y(_03245_),
    .B1(_03244_));
 sg13g2_nand3_1 _12304_ (.B(_02762_),
    .C(_02945_),
    .A(_03240_),
    .Y(_03246_));
 sg13g2_nand2_1 _12305_ (.Y(_03247_),
    .A(_03245_),
    .B(_03246_));
 sg13g2_xnor2_1 _12306_ (.Y(_03248_),
    .A(_03237_),
    .B(_03247_));
 sg13g2_nand2_1 _12307_ (.Y(_03249_),
    .A(_03248_),
    .B(_03131_));
 sg13g2_inv_1 _12308_ (.Y(_03250_),
    .A(_03237_));
 sg13g2_xnor2_1 _12309_ (.Y(_03251_),
    .A(_03250_),
    .B(_03247_));
 sg13g2_nand2_1 _12310_ (.Y(_03252_),
    .A(_03251_),
    .B(_03126_));
 sg13g2_nand2_1 _12311_ (.Y(_03253_),
    .A(_03249_),
    .B(_03252_));
 sg13g2_xor2_1 _12312_ (.B(_03253_),
    .A(_03209_),
    .X(_03254_));
 sg13g2_nand2_1 _12313_ (.Y(_03255_),
    .A(_03227_),
    .B(_03254_));
 sg13g2_xnor2_1 _12314_ (.Y(_03256_),
    .A(_03209_),
    .B(_03253_));
 sg13g2_nand3_1 _12315_ (.B(_03226_),
    .C(_03256_),
    .A(_03220_),
    .Y(_03257_));
 sg13g2_inv_1 _12316_ (.Y(_03258_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[10] ));
 sg13g2_nand3_1 _12317_ (.B(_03257_),
    .C(_03258_),
    .A(_03255_),
    .Y(_03259_));
 sg13g2_buf_1 _12318_ (.A(_03259_),
    .X(_03260_));
 sg13g2_nor2_1 _12319_ (.A(_03078_),
    .B(_03139_),
    .Y(_03261_));
 sg13g2_nand2_1 _12320_ (.Y(_03262_),
    .A(_03138_),
    .B(_03075_));
 sg13g2_nand2_1 _12321_ (.Y(_03263_),
    .A(_03262_),
    .B(_03135_));
 sg13g2_inv_1 _12322_ (.Y(_03264_),
    .A(_03263_));
 sg13g2_a21oi_1 _12323_ (.A1(_03261_),
    .A2(_03151_),
    .Y(_03265_),
    .B1(_03264_));
 sg13g2_nand3_1 _12324_ (.B(_03152_),
    .C(_02971_),
    .A(_03261_),
    .Y(_03266_));
 sg13g2_nand2_1 _12325_ (.Y(_03267_),
    .A(_03265_),
    .B(_03266_));
 sg13g2_nand2_1 _12326_ (.Y(_03268_),
    .A(_03267_),
    .B(_03221_));
 sg13g2_nand3_1 _12327_ (.B(_03266_),
    .C(_03218_),
    .A(_03265_),
    .Y(_03269_));
 sg13g2_inv_1 _12328_ (.Y(_03270_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[9] ));
 sg13g2_nand3_1 _12329_ (.B(_03269_),
    .C(_03270_),
    .A(_03268_),
    .Y(_03271_));
 sg13g2_nand2_1 _12330_ (.Y(_03272_),
    .A(_03260_),
    .B(_03271_));
 sg13g2_nand2_1 _12331_ (.Y(_03273_),
    .A(_03255_),
    .B(_03257_));
 sg13g2_nand2_1 _12332_ (.Y(_03274_),
    .A(_03273_),
    .B(\vgadonut.donut.donuthit.cordicxz.xin[10] ));
 sg13g2_buf_2 _12333_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[7] ),
    .X(_03275_));
 sg13g2_nor2_1 _12334_ (.A(_03275_),
    .B(_03155_),
    .Y(_03276_));
 sg13g2_nand2_1 _12335_ (.Y(_03277_),
    .A(_03276_),
    .B(_03148_));
 sg13g2_nand2_1 _12336_ (.Y(_03278_),
    .A(_03277_),
    .B(_03147_));
 sg13g2_a21oi_1 _12337_ (.A1(_03272_),
    .A2(_03274_),
    .Y(_03279_),
    .B1(_03278_));
 sg13g2_nand2_1 _12338_ (.Y(_03280_),
    .A(_03268_),
    .B(_03269_));
 sg13g2_nand3_1 _12339_ (.B(\vgadonut.donut.donuthit.cordicxz.xin[9] ),
    .C(_03280_),
    .A(_03260_),
    .Y(_03281_));
 sg13g2_nand2_1 _12340_ (.Y(_03282_),
    .A(_03281_),
    .B(_03274_));
 sg13g2_a21oi_1 _12341_ (.A1(_03158_),
    .A2(_03279_),
    .Y(_03283_),
    .B1(_03282_));
 sg13g2_nand2_1 _12342_ (.Y(_03284_),
    .A(_03201_),
    .B(_03237_));
 sg13g2_a21oi_1 _12343_ (.A1(_03242_),
    .A2(_03235_),
    .Y(_03285_),
    .B1(_03234_));
 sg13g2_o21ai_1 _12344_ (.B1(_03285_),
    .Y(_03286_),
    .A1(_03167_),
    .A2(_03284_));
 sg13g2_nand3_1 _12345_ (.B(_03237_),
    .C(_03201_),
    .A(_03161_),
    .Y(_03287_));
 sg13g2_nor2_1 _12346_ (.A(_03287_),
    .B(_03030_),
    .Y(_03288_));
 sg13g2_nor2_1 _12347_ (.A(_03286_),
    .B(_03288_),
    .Y(_03289_));
 sg13g2_nor2b_1 _12348_ (.A(_03287_),
    .B_N(_03023_),
    .Y(_03290_));
 sg13g2_nand2_1 _12349_ (.Y(_03291_),
    .A(_03290_),
    .B(_02782_));
 sg13g2_nand2_1 _12350_ (.Y(_03292_),
    .A(_03289_),
    .B(_03291_));
 sg13g2_xnor2_1 _12351_ (.Y(_03293_),
    .A(net178),
    .B(_02399_));
 sg13g2_nand2_1 _12352_ (.Y(_03294_),
    .A(_03230_),
    .B(_03229_));
 sg13g2_xnor2_1 _12353_ (.Y(_03295_),
    .A(_03293_),
    .B(_03294_));
 sg13g2_inv_1 _12354_ (.Y(_03296_),
    .A(_03295_));
 sg13g2_nand2_1 _12355_ (.Y(_03297_),
    .A(_03292_),
    .B(_03296_));
 sg13g2_nand3_1 _12356_ (.B(_03295_),
    .C(_03291_),
    .A(_03289_),
    .Y(_03298_));
 sg13g2_nand2_1 _12357_ (.Y(_03299_),
    .A(_03297_),
    .B(_03298_));
 sg13g2_buf_8 _12358_ (.A(_03299_),
    .X(_03300_));
 sg13g2_inv_4 _12359_ (.A(_03300_),
    .Y(_03301_));
 sg13g2_nand2_2 _12360_ (.Y(_03302_),
    .A(_03301_),
    .B(_03207_));
 sg13g2_inv_1 _12361_ (.Y(_03303_),
    .A(_03249_));
 sg13g2_nand2_1 _12362_ (.Y(_03304_),
    .A(_03300_),
    .B(_03212_));
 sg13g2_nand3_1 _12363_ (.B(_03303_),
    .C(_03304_),
    .A(_03302_),
    .Y(_03305_));
 sg13g2_nand2_1 _12364_ (.Y(_03306_),
    .A(_03301_),
    .B(_03212_));
 sg13g2_nand2_1 _12365_ (.Y(_03307_),
    .A(_03300_),
    .B(_03207_));
 sg13g2_nand3_1 _12366_ (.B(_03307_),
    .C(_03249_),
    .A(_03306_),
    .Y(_03308_));
 sg13g2_buf_1 _12367_ (.A(_03308_),
    .X(_03309_));
 sg13g2_nand2_2 _12368_ (.Y(_03310_),
    .A(_03305_),
    .B(_03309_));
 sg13g2_nand2_1 _12369_ (.Y(_03311_),
    .A(_03237_),
    .B(_03295_));
 sg13g2_nor2b_1 _12370_ (.A(_03294_),
    .B_N(_03293_),
    .Y(_03312_));
 sg13g2_a21oi_1 _12371_ (.A1(_03234_),
    .A2(_03295_),
    .Y(_03313_),
    .B1(_03312_));
 sg13g2_o21ai_1 _12372_ (.B1(_03313_),
    .Y(_03314_),
    .A1(_03311_),
    .A2(_03243_));
 sg13g2_nor2_1 _12373_ (.A(_03311_),
    .B(_03239_),
    .Y(_03315_));
 sg13g2_nor2b_1 _12374_ (.A(_03124_),
    .B_N(_03315_),
    .Y(_03316_));
 sg13g2_nor2_1 _12375_ (.A(_03314_),
    .B(_03316_),
    .Y(_03317_));
 sg13g2_nand3_1 _12376_ (.B(_03315_),
    .C(_03117_),
    .A(_02851_),
    .Y(_03318_));
 sg13g2_nand2_1 _12377_ (.Y(_03319_),
    .A(_03317_),
    .B(_03318_));
 sg13g2_xnor2_1 _12378_ (.Y(_03320_),
    .A(_02588_),
    .B(_03319_));
 sg13g2_xnor2_1 _12379_ (.Y(_03321_),
    .A(_03248_),
    .B(_03320_));
 sg13g2_xnor2_1 _12380_ (.Y(_03322_),
    .A(_03302_),
    .B(_03321_));
 sg13g2_buf_2 _12381_ (.A(_03322_),
    .X(_03323_));
 sg13g2_nand2_1 _12382_ (.Y(_03324_),
    .A(_03254_),
    .B(_03221_));
 sg13g2_nor3_1 _12383_ (.A(_03310_),
    .B(_03323_),
    .C(_03324_),
    .Y(_03325_));
 sg13g2_nand2_1 _12384_ (.Y(_03326_),
    .A(_03267_),
    .B(_03325_));
 sg13g2_nand2_1 _12385_ (.Y(_03327_),
    .A(_03253_),
    .B(_03209_));
 sg13g2_o21ai_1 _12386_ (.B1(_03327_),
    .Y(_03328_),
    .A1(_03216_),
    .A2(_03256_));
 sg13g2_nor2_1 _12387_ (.A(_03310_),
    .B(_03323_),
    .Y(_03329_));
 sg13g2_nand2_1 _12388_ (.Y(_03330_),
    .A(_03321_),
    .B(_03302_));
 sg13g2_nor2_1 _12389_ (.A(_03302_),
    .B(_03321_),
    .Y(_03331_));
 sg13g2_a21oi_1 _12390_ (.A1(_03330_),
    .A2(_03309_),
    .Y(_03332_),
    .B1(_03331_));
 sg13g2_a21oi_1 _12391_ (.A1(_03328_),
    .A2(_03329_),
    .Y(_03333_),
    .B1(_03332_));
 sg13g2_nand2_1 _12392_ (.Y(_03334_),
    .A(_03326_),
    .B(_03333_));
 sg13g2_nor2b_1 _12393_ (.A(_03300_),
    .B_N(_03320_),
    .Y(_03335_));
 sg13g2_nand2_1 _12394_ (.Y(_03336_),
    .A(_03335_),
    .B(_03251_));
 sg13g2_nand3_1 _12395_ (.B(_03300_),
    .C(_03248_),
    .A(_03320_),
    .Y(_03337_));
 sg13g2_nand2b_1 _12396_ (.Y(_03338_),
    .B(_03300_),
    .A_N(_03320_));
 sg13g2_nand3_1 _12397_ (.B(_03337_),
    .C(_03338_),
    .A(_03336_),
    .Y(_03339_));
 sg13g2_buf_1 _12398_ (.A(_03339_),
    .X(_03340_));
 sg13g2_nand2_1 _12399_ (.Y(_03341_),
    .A(_03334_),
    .B(_03340_));
 sg13g2_inv_1 _12400_ (.Y(_03342_),
    .A(_03340_));
 sg13g2_nand3_1 _12401_ (.B(_03333_),
    .C(_03342_),
    .A(_03326_),
    .Y(_03343_));
 sg13g2_buf_1 _12402_ (.A(_03343_),
    .X(_03344_));
 sg13g2_nand2_1 _12403_ (.Y(_03345_),
    .A(_03341_),
    .B(_03344_));
 sg13g2_buf_2 _12404_ (.A(_00166_),
    .X(_03346_));
 sg13g2_nand2_1 _12405_ (.Y(_03347_),
    .A(_03345_),
    .B(_03346_));
 sg13g2_inv_1 _12406_ (.Y(_03348_),
    .A(_03346_));
 sg13g2_nand3_1 _12407_ (.B(_03344_),
    .C(_03348_),
    .A(_03341_),
    .Y(_03349_));
 sg13g2_nand2_2 _12408_ (.Y(_03350_),
    .A(_03347_),
    .B(_03349_));
 sg13g2_inv_2 _12409_ (.Y(_03351_),
    .A(_03310_));
 sg13g2_nand2_1 _12410_ (.Y(_03352_),
    .A(_03351_),
    .B(_03254_));
 sg13g2_nor3_1 _12411_ (.A(_03323_),
    .B(_03340_),
    .C(_03352_),
    .Y(_03353_));
 sg13g2_nand2_1 _12412_ (.Y(_03354_),
    .A(_03227_),
    .B(_03353_));
 sg13g2_o21ai_1 _12413_ (.B1(_03309_),
    .Y(_03355_),
    .A1(_03327_),
    .A2(_03310_));
 sg13g2_nor2_1 _12414_ (.A(_03323_),
    .B(_03340_),
    .Y(_03356_));
 sg13g2_inv_1 _12415_ (.Y(_03357_),
    .A(_03337_));
 sg13g2_nand2_1 _12416_ (.Y(_03358_),
    .A(_03336_),
    .B(_03338_));
 sg13g2_inv_1 _12417_ (.Y(_03359_),
    .A(_03358_));
 sg13g2_o21ai_1 _12418_ (.B1(_03359_),
    .Y(_03360_),
    .A1(_03330_),
    .A2(_03357_));
 sg13g2_a21oi_1 _12419_ (.A1(_03355_),
    .A2(_03356_),
    .Y(_03361_),
    .B1(_03360_));
 sg13g2_nand2_1 _12420_ (.Y(_03362_),
    .A(_03354_),
    .B(_03361_));
 sg13g2_inv_1 _12421_ (.Y(_03363_),
    .A(_03335_));
 sg13g2_nand2_1 _12422_ (.Y(_03364_),
    .A(_03362_),
    .B(_03363_));
 sg13g2_nand3_1 _12423_ (.B(_03335_),
    .C(_03361_),
    .A(_03354_),
    .Y(_03365_));
 sg13g2_nand2_1 _12424_ (.Y(_03366_),
    .A(_03364_),
    .B(_03365_));
 sg13g2_inv_1 _12425_ (.Y(_03367_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[14] ));
 sg13g2_nand2_1 _12426_ (.Y(_03368_),
    .A(_03366_),
    .B(_03367_));
 sg13g2_nand3_1 _12427_ (.B(_03365_),
    .C(\vgadonut.donut.donuthit.cordicxz.xin[14] ),
    .A(_03364_),
    .Y(_03369_));
 sg13g2_nand2_1 _12428_ (.Y(_03370_),
    .A(_03368_),
    .B(_03369_));
 sg13g2_nor2_1 _12429_ (.A(_03222_),
    .B(_03352_),
    .Y(_03371_));
 sg13g2_nand2_1 _12430_ (.Y(_03372_),
    .A(_03083_),
    .B(_03371_));
 sg13g2_nor2_1 _12431_ (.A(_03225_),
    .B(_03352_),
    .Y(_03373_));
 sg13g2_nor2_1 _12432_ (.A(_03355_),
    .B(_03373_),
    .Y(_03374_));
 sg13g2_nand2_1 _12433_ (.Y(_03375_),
    .A(_03372_),
    .B(_03374_));
 sg13g2_nand2_1 _12434_ (.Y(_03376_),
    .A(_03375_),
    .B(_03323_));
 sg13g2_inv_1 _12435_ (.Y(_03377_),
    .A(_03323_));
 sg13g2_nand3_1 _12436_ (.B(_03374_),
    .C(_03377_),
    .A(_03372_),
    .Y(_03378_));
 sg13g2_buf_1 _12437_ (.A(_03378_),
    .X(_03379_));
 sg13g2_nand2_1 _12438_ (.Y(_03380_),
    .A(_03376_),
    .B(_03379_));
 sg13g2_inv_1 _12439_ (.Y(_03381_),
    .A(_00167_));
 sg13g2_nand2_1 _12440_ (.Y(_03382_),
    .A(_03380_),
    .B(_03381_));
 sg13g2_nand3_1 _12441_ (.B(_03379_),
    .C(_00167_),
    .A(_03376_),
    .Y(_03383_));
 sg13g2_nand2_1 _12442_ (.Y(_03384_),
    .A(_03382_),
    .B(_03383_));
 sg13g2_nor2b_1 _12443_ (.A(_03324_),
    .B_N(_03261_),
    .Y(_03385_));
 sg13g2_nand2_1 _12444_ (.Y(_03386_),
    .A(_03154_),
    .B(_03385_));
 sg13g2_nor2_1 _12445_ (.A(_03263_),
    .B(_03324_),
    .Y(_03387_));
 sg13g2_nor2_1 _12446_ (.A(_03387_),
    .B(_03328_),
    .Y(_03388_));
 sg13g2_nand2_1 _12447_ (.Y(_03389_),
    .A(_03386_),
    .B(_03388_));
 sg13g2_nand2_1 _12448_ (.Y(_03390_),
    .A(_03389_),
    .B(_03351_));
 sg13g2_nand3_1 _12449_ (.B(_03388_),
    .C(_03310_),
    .A(_03386_),
    .Y(_03391_));
 sg13g2_nand2_1 _12450_ (.Y(_03392_),
    .A(_03390_),
    .B(_03391_));
 sg13g2_xnor2_1 _12451_ (.Y(_03393_),
    .A(_00158_),
    .B(_03392_));
 sg13g2_nand2_1 _12452_ (.Y(_03394_),
    .A(_03384_),
    .B(_03393_));
 sg13g2_nor3_1 _12453_ (.A(_03350_),
    .B(_03370_),
    .C(_03394_),
    .Y(_03395_));
 sg13g2_nand2_1 _12454_ (.Y(_03396_),
    .A(_03283_),
    .B(_03395_));
 sg13g2_nor2_1 _12455_ (.A(_03350_),
    .B(_03370_),
    .Y(_03397_));
 sg13g2_buf_1 _12456_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[12] ),
    .X(_03398_));
 sg13g2_nand3_1 _12457_ (.B(_03379_),
    .C(_03398_),
    .A(_03376_),
    .Y(_03399_));
 sg13g2_nor2_1 _12458_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[11] ),
    .B(_03392_),
    .Y(_03400_));
 sg13g2_nand2_1 _12459_ (.Y(_03401_),
    .A(_03399_),
    .B(_03400_));
 sg13g2_inv_1 _12460_ (.Y(_03402_),
    .A(_03398_));
 sg13g2_nand2_1 _12461_ (.Y(_03403_),
    .A(_03380_),
    .B(_03402_));
 sg13g2_nand2_1 _12462_ (.Y(_03404_),
    .A(_03401_),
    .B(_03403_));
 sg13g2_inv_1 _12463_ (.Y(_03405_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[13] ));
 sg13g2_nand2_1 _12464_ (.Y(_03406_),
    .A(_03345_),
    .B(_03405_));
 sg13g2_inv_1 _12465_ (.Y(_03407_),
    .A(_03369_));
 sg13g2_a21oi_1 _12466_ (.A1(_03368_),
    .A2(_03406_),
    .Y(_03408_),
    .B1(_03407_));
 sg13g2_a21oi_1 _12467_ (.A1(_03397_),
    .A2(_03404_),
    .Y(_03409_),
    .B1(_03408_));
 sg13g2_nand2_1 _12468_ (.Y(_03410_),
    .A(_03396_),
    .B(_03409_));
 sg13g2_nor3_1 _12469_ (.A(_03300_),
    .B(_03251_),
    .C(_03332_),
    .Y(_03411_));
 sg13g2_o21ai_1 _12470_ (.B1(_03411_),
    .Y(_03412_),
    .A1(_03323_),
    .A2(_03390_));
 sg13g2_nand2_1 _12471_ (.Y(_03413_),
    .A(_03412_),
    .B(_03320_));
 sg13g2_buf_2 _12472_ (.A(_03413_),
    .X(_03414_));
 sg13g2_xnor2_1 _12473_ (.Y(_03415_),
    .A(_00165_),
    .B(_03414_));
 sg13g2_inv_1 _12474_ (.Y(_03416_),
    .A(_03415_));
 sg13g2_nand2_1 _12475_ (.Y(_03417_),
    .A(_03410_),
    .B(_03416_));
 sg13g2_nand3_1 _12476_ (.B(_03409_),
    .C(_03415_),
    .A(_03396_),
    .Y(_03418_));
 sg13g2_inv_1 _12477_ (.Y(_03419_),
    .A(_03414_));
 sg13g2_nand2_1 _12478_ (.Y(_03420_),
    .A(_03419_),
    .B(\vgadonut.donut.donuthit.cordicxz.xin[15] ));
 sg13g2_nand2b_1 _12479_ (.Y(_03421_),
    .B(_03414_),
    .A_N(\vgadonut.donut.donuthit.cordicxz.xin[15] ));
 sg13g2_nand2_1 _12480_ (.Y(_03422_),
    .A(_03420_),
    .B(_03421_));
 sg13g2_buf_8 _12481_ (.A(_03422_),
    .X(_03423_));
 sg13g2_inv_2 _12482_ (.Y(_03424_),
    .A(_03423_));
 sg13g2_nand3_1 _12483_ (.B(_03418_),
    .C(_03424_),
    .A(_03417_),
    .Y(_03425_));
 sg13g2_buf_1 _12484_ (.A(_03425_),
    .X(_03426_));
 sg13g2_inv_1 _12485_ (.Y(_03427_),
    .A(_03150_));
 sg13g2_nor2_1 _12486_ (.A(_02977_),
    .B(_02978_),
    .Y(_03428_));
 sg13g2_nor2_1 _12487_ (.A(_02984_),
    .B(_03015_),
    .Y(_03429_));
 sg13g2_nor2b_1 _12488_ (.A(_03007_),
    .B_N(\vgadonut.donut.donuthit.cordicxz.xin[0] ),
    .Y(_03430_));
 sg13g2_a21oi_1 _12489_ (.A1(_03005_),
    .A2(_03430_),
    .Y(_03431_),
    .B1(_03004_));
 sg13g2_a21oi_1 _12490_ (.A1(_02996_),
    .A2(_02998_),
    .Y(_03432_),
    .B1(_02994_));
 sg13g2_nand3_1 _12491_ (.B(_02994_),
    .C(_02998_),
    .A(_02996_),
    .Y(_03433_));
 sg13g2_o21ai_1 _12492_ (.B1(_03433_),
    .Y(_03434_),
    .A1(_03431_),
    .A2(_03432_));
 sg13g2_nand2_1 _12493_ (.Y(_03435_),
    .A(_03015_),
    .B(_02983_));
 sg13g2_nand2_1 _12494_ (.Y(_03436_),
    .A(_03435_),
    .B(_02986_));
 sg13g2_nand2_1 _12495_ (.Y(_03437_),
    .A(_03434_),
    .B(_03436_));
 sg13g2_nand2b_1 _12496_ (.Y(_03438_),
    .B(_03437_),
    .A_N(_03429_));
 sg13g2_nand2_1 _12497_ (.Y(_03439_),
    .A(_03438_),
    .B(_03017_));
 sg13g2_nand2b_1 _12498_ (.Y(_03440_),
    .B(_03439_),
    .A_N(_03428_));
 sg13g2_inv_1 _12499_ (.Y(_03441_),
    .A(_02964_));
 sg13g2_nor2_1 _12500_ (.A(_03441_),
    .B(_02972_),
    .Y(_03442_));
 sg13g2_nand2_1 _12501_ (.Y(_03443_),
    .A(_02972_),
    .B(_03441_));
 sg13g2_nor2b_1 _12502_ (.A(_03442_),
    .B_N(_03443_),
    .Y(_03444_));
 sg13g2_nand2_1 _12503_ (.Y(_03445_),
    .A(_03440_),
    .B(_03444_));
 sg13g2_inv_1 _12504_ (.Y(_03446_),
    .A(_02958_));
 sg13g2_nor2_1 _12505_ (.A(_03442_),
    .B(_03446_),
    .Y(_03447_));
 sg13g2_nand2_1 _12506_ (.Y(_03448_),
    .A(_03445_),
    .B(_03447_));
 sg13g2_inv_1 _12507_ (.Y(_03449_),
    .A(_03275_));
 sg13g2_nor2_1 _12508_ (.A(_03449_),
    .B(_03155_),
    .Y(_03450_));
 sg13g2_inv_1 _12509_ (.Y(_03451_),
    .A(_03155_));
 sg13g2_nor2_1 _12510_ (.A(_03275_),
    .B(_03451_),
    .Y(_03452_));
 sg13g2_nor2_1 _12511_ (.A(_03450_),
    .B(_03452_),
    .Y(_03453_));
 sg13g2_nand3_1 _12512_ (.B(_02961_),
    .C(_03453_),
    .A(_03448_),
    .Y(_03454_));
 sg13g2_nor2_1 _12513_ (.A(_03427_),
    .B(_03454_),
    .Y(_03455_));
 sg13g2_inv_1 _12514_ (.Y(_03456_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[11] ));
 sg13g2_nor2_1 _12515_ (.A(_03456_),
    .B(_03392_),
    .Y(_03457_));
 sg13g2_inv_1 _12516_ (.Y(_03458_),
    .A(_03457_));
 sg13g2_nand2_1 _12517_ (.Y(_03459_),
    .A(_03392_),
    .B(_03456_));
 sg13g2_nand2_1 _12518_ (.Y(_03460_),
    .A(_03458_),
    .B(_03459_));
 sg13g2_nand2_1 _12519_ (.Y(_03461_),
    .A(_03403_),
    .B(_03399_));
 sg13g2_buf_2 _12520_ (.A(_03461_),
    .X(_03462_));
 sg13g2_nor2b_1 _12521_ (.A(_03460_),
    .B_N(_03462_),
    .Y(_03463_));
 sg13g2_nor2_1 _12522_ (.A(_03270_),
    .B(_03280_),
    .Y(_03464_));
 sg13g2_nand2_1 _12523_ (.Y(_03465_),
    .A(_03280_),
    .B(_03270_));
 sg13g2_nand2b_1 _12524_ (.Y(_03466_),
    .B(_03465_),
    .A_N(_03464_));
 sg13g2_buf_1 _12525_ (.A(_03466_),
    .X(_03467_));
 sg13g2_nand2_1 _12526_ (.Y(_03468_),
    .A(_03274_),
    .B(_03260_));
 sg13g2_buf_8 _12527_ (.A(_03468_),
    .X(_03469_));
 sg13g2_nor2b_1 _12528_ (.A(_03467_),
    .B_N(_03469_),
    .Y(_03470_));
 sg13g2_nand3_1 _12529_ (.B(_03463_),
    .C(_03470_),
    .A(_03455_),
    .Y(_03471_));
 sg13g2_a22oi_1 _12530_ (.Y(_03472_),
    .B1(_03457_),
    .B2(_03462_),
    .A2(_03380_),
    .A1(_03381_));
 sg13g2_nand2_1 _12531_ (.Y(_03473_),
    .A(_03471_),
    .B(_03472_));
 sg13g2_nand2_1 _12532_ (.Y(_03474_),
    .A(_03345_),
    .B(\vgadonut.donut.donuthit.cordicxz.xin[13] ));
 sg13g2_nand3_1 _12533_ (.B(_03344_),
    .C(_03405_),
    .A(_03341_),
    .Y(_03475_));
 sg13g2_nand2_1 _12534_ (.Y(_03476_),
    .A(_03474_),
    .B(_03475_));
 sg13g2_inv_2 _12535_ (.Y(_03477_),
    .A(_00168_));
 sg13g2_xnor2_1 _12536_ (.Y(_03478_),
    .A(_03477_),
    .B(_03366_));
 sg13g2_nor2_1 _12537_ (.A(_03476_),
    .B(_03478_),
    .Y(_03479_));
 sg13g2_nand2_1 _12538_ (.Y(_03480_),
    .A(_03473_),
    .B(_03479_));
 sg13g2_nand2_1 _12539_ (.Y(_03481_),
    .A(_03479_),
    .B(_03463_));
 sg13g2_inv_1 _12540_ (.Y(_03482_),
    .A(_03145_));
 sg13g2_nor2_1 _12541_ (.A(_03146_),
    .B(_03482_),
    .Y(_03483_));
 sg13g2_a21oi_1 _12542_ (.A1(_03150_),
    .A2(_03450_),
    .Y(_03484_),
    .B1(_03483_));
 sg13g2_inv_1 _12543_ (.Y(_03485_),
    .A(_03484_));
 sg13g2_nand2_1 _12544_ (.Y(_03486_),
    .A(_03470_),
    .B(_03485_));
 sg13g2_nor2_1 _12545_ (.A(_00164_),
    .B(_03273_),
    .Y(_03487_));
 sg13g2_a21oi_1 _12546_ (.A1(_03469_),
    .A2(_03464_),
    .Y(_03488_),
    .B1(_03487_));
 sg13g2_nand2_1 _12547_ (.Y(_03489_),
    .A(_03486_),
    .B(_03488_));
 sg13g2_nor2b_1 _12548_ (.A(_03481_),
    .B_N(_03489_),
    .Y(_03490_));
 sg13g2_inv_1 _12549_ (.Y(_03491_),
    .A(_03366_));
 sg13g2_a21oi_1 _12550_ (.A1(_03491_),
    .A2(_00168_),
    .Y(_03492_),
    .B1(_03474_));
 sg13g2_a21oi_1 _12551_ (.A1(_03477_),
    .A2(_03366_),
    .Y(_03493_),
    .B1(_03492_));
 sg13g2_nor2b_1 _12552_ (.A(_03490_),
    .B_N(_03493_),
    .Y(_03494_));
 sg13g2_nand3_1 _12553_ (.B(_03423_),
    .C(_03494_),
    .A(_03480_),
    .Y(_03495_));
 sg13g2_buf_8 _12554_ (.A(_03495_),
    .X(_03496_));
 sg13g2_nand2_1 _12555_ (.Y(_03497_),
    .A(_03426_),
    .B(_03496_));
 sg13g2_buf_8 _12556_ (.A(_03497_),
    .X(_03498_));
 sg13g2_buf_8 _12557_ (.A(_03498_),
    .X(_03499_));
 sg13g2_nand2_1 _12558_ (.Y(_03500_),
    .A(_03448_),
    .B(_02961_));
 sg13g2_inv_1 _12559_ (.Y(_03501_),
    .A(_03450_));
 sg13g2_a21oi_1 _12560_ (.A1(_03500_),
    .A2(_03501_),
    .Y(_03502_),
    .B1(_03452_));
 sg13g2_inv_1 _12561_ (.Y(_03503_),
    .A(_03467_));
 sg13g2_nand3_1 _12562_ (.B(_03150_),
    .C(_03503_),
    .A(_03502_),
    .Y(_03504_));
 sg13g2_o21ai_1 _12563_ (.B1(_03465_),
    .Y(_03505_),
    .A1(_03483_),
    .A2(_03464_));
 sg13g2_nand2_1 _12564_ (.Y(_03506_),
    .A(_03504_),
    .B(_03505_));
 sg13g2_xnor2_1 _12565_ (.Y(_03507_),
    .A(_03469_),
    .B(_03506_));
 sg13g2_buf_8 _12566_ (.A(_03423_),
    .X(_03508_));
 sg13g2_buf_2 _12567_ (.A(_03508_),
    .X(_03509_));
 sg13g2_buf_8 _12568_ (.A(_03509_),
    .X(_03510_));
 sg13g2_nand2b_1 _12569_ (.Y(_03511_),
    .B(_03158_),
    .A_N(_03278_));
 sg13g2_nand2_1 _12570_ (.Y(_03512_),
    .A(_03511_),
    .B(_03467_));
 sg13g2_nand2_1 _12571_ (.Y(_03513_),
    .A(_03512_),
    .B(_03271_));
 sg13g2_xnor2_1 _12572_ (.Y(_03514_),
    .A(_03469_),
    .B(_03513_));
 sg13g2_nor2_1 _12573_ (.A(_03509_),
    .B(_03514_),
    .Y(_03515_));
 sg13g2_a21oi_1 _12574_ (.A1(_03507_),
    .A2(net47),
    .Y(_03516_),
    .B1(_03515_));
 sg13g2_xor2_1 _12575_ (.B(_03516_),
    .A(net40),
    .X(_03517_));
 sg13g2_buf_1 _12576_ (.A(_03419_),
    .X(_03518_));
 sg13g2_nor2_1 _12577_ (.A(_03485_),
    .B(_03455_),
    .Y(_03519_));
 sg13g2_xnor2_1 _12578_ (.Y(_03520_),
    .A(_03503_),
    .B(_03519_));
 sg13g2_xnor2_1 _12579_ (.Y(_03521_),
    .A(_03503_),
    .B(_03511_));
 sg13g2_nand2b_1 _12580_ (.Y(_03522_),
    .B(net49),
    .A_N(_03521_));
 sg13g2_o21ai_1 _12581_ (.B1(_03522_),
    .Y(_03523_),
    .A1(_03510_),
    .A2(_03520_));
 sg13g2_xnor2_1 _12582_ (.Y(_03524_),
    .A(net52),
    .B(_03523_));
 sg13g2_nand2b_1 _12583_ (.Y(_03525_),
    .B(_03524_),
    .A_N(_03517_));
 sg13g2_nand2b_1 _12584_ (.Y(_03526_),
    .B(_03517_),
    .A_N(_03524_));
 sg13g2_nand2_2 _12585_ (.Y(_03527_),
    .A(_03525_),
    .B(_03526_));
 sg13g2_xnor2_1 _12586_ (.Y(_03528_),
    .A(_03009_),
    .B(_03006_));
 sg13g2_xor2_1 _12587_ (.B(_03006_),
    .A(_03430_),
    .X(_03529_));
 sg13g2_nor2b_1 _12588_ (.A(net50),
    .B_N(_03529_),
    .Y(_03530_));
 sg13g2_a21oi_1 _12589_ (.A1(net50),
    .A2(_03528_),
    .Y(_03531_),
    .B1(_03530_));
 sg13g2_xnor2_1 _12590_ (.Y(_03532_),
    .A(_03414_),
    .B(_03531_));
 sg13g2_inv_1 _12591_ (.Y(_03533_),
    .A(_03433_));
 sg13g2_nor2_1 _12592_ (.A(_03432_),
    .B(_03533_),
    .Y(_03534_));
 sg13g2_xor2_1 _12593_ (.B(_03534_),
    .A(_03431_),
    .X(_03535_));
 sg13g2_xor2_1 _12594_ (.B(_03011_),
    .A(_03012_),
    .X(_03536_));
 sg13g2_nor2b_1 _12595_ (.A(_03423_),
    .B_N(_03536_),
    .Y(_03537_));
 sg13g2_a21oi_1 _12596_ (.A1(_03423_),
    .A2(_03535_),
    .Y(_03538_),
    .B1(_03537_));
 sg13g2_inv_1 _12597_ (.Y(_03539_),
    .A(_03538_));
 sg13g2_nand2_1 _12598_ (.Y(_03540_),
    .A(_03498_),
    .B(_03539_));
 sg13g2_nand3_1 _12599_ (.B(_03496_),
    .C(_03538_),
    .A(_03426_),
    .Y(_03541_));
 sg13g2_nand2_1 _12600_ (.Y(_03542_),
    .A(_03540_),
    .B(_03541_));
 sg13g2_nand2b_1 _12601_ (.Y(_03543_),
    .B(_03542_),
    .A_N(_03532_));
 sg13g2_buf_1 _12602_ (.A(_03543_),
    .X(_03544_));
 sg13g2_nor2b_1 _12603_ (.A(_03423_),
    .B_N(_03528_),
    .Y(_03545_));
 sg13g2_a21oi_1 _12604_ (.A1(_03508_),
    .A2(_03529_),
    .Y(_03546_),
    .B1(_03545_));
 sg13g2_inv_1 _12605_ (.Y(_03547_),
    .A(_03546_));
 sg13g2_nand3_1 _12606_ (.B(_03496_),
    .C(_03547_),
    .A(_03426_),
    .Y(_03548_));
 sg13g2_xnor2_1 _12607_ (.Y(_03549_),
    .A(_00163_),
    .B(_03007_));
 sg13g2_xnor2_1 _12608_ (.Y(_03550_),
    .A(_03549_),
    .B(_03414_));
 sg13g2_nand2_1 _12609_ (.Y(_03551_),
    .A(_03548_),
    .B(_03550_));
 sg13g2_nand2_1 _12610_ (.Y(_03552_),
    .A(net40),
    .B(_03546_));
 sg13g2_nor2b_1 _12611_ (.A(_03551_),
    .B_N(_03552_),
    .Y(_03553_));
 sg13g2_nand3_1 _12612_ (.B(_03541_),
    .C(_03532_),
    .A(_03540_),
    .Y(_03554_));
 sg13g2_nand3_1 _12613_ (.B(_03553_),
    .C(_03554_),
    .A(_03544_),
    .Y(_03555_));
 sg13g2_nor2b_1 _12614_ (.A(_03423_),
    .B_N(_03535_),
    .Y(_03556_));
 sg13g2_a21oi_1 _12615_ (.A1(net50),
    .A2(_03536_),
    .Y(_03557_),
    .B1(_03556_));
 sg13g2_xnor2_1 _12616_ (.Y(_03558_),
    .A(_03414_),
    .B(_03557_));
 sg13g2_xnor2_1 _12617_ (.Y(_03559_),
    .A(_03436_),
    .B(_03434_));
 sg13g2_inv_1 _12618_ (.Y(_03560_),
    .A(_03016_));
 sg13g2_xnor2_1 _12619_ (.Y(_03561_),
    .A(_03560_),
    .B(_03014_));
 sg13g2_nor2b_1 _12620_ (.A(_03423_),
    .B_N(_03561_),
    .Y(_03562_));
 sg13g2_a21oi_1 _12621_ (.A1(net50),
    .A2(_03559_),
    .Y(_03563_),
    .B1(_03562_));
 sg13g2_inv_1 _12622_ (.Y(_03564_),
    .A(_03563_));
 sg13g2_nand2_1 _12623_ (.Y(_03565_),
    .A(_03498_),
    .B(_03564_));
 sg13g2_nand3_1 _12624_ (.B(_03496_),
    .C(_03563_),
    .A(_03426_),
    .Y(_03566_));
 sg13g2_nand2_1 _12625_ (.Y(_03567_),
    .A(_03565_),
    .B(_03566_));
 sg13g2_nand2b_1 _12626_ (.Y(_03568_),
    .B(_03567_),
    .A_N(_03558_));
 sg13g2_and2_1 _12627_ (.A(_03544_),
    .B(_03568_),
    .X(_03569_));
 sg13g2_nand2_1 _12628_ (.Y(_03570_),
    .A(_03555_),
    .B(_03569_));
 sg13g2_nand3_1 _12629_ (.B(_03566_),
    .C(_03558_),
    .A(_03565_),
    .Y(_03571_));
 sg13g2_buf_1 _12630_ (.A(_03571_),
    .X(_03572_));
 sg13g2_buf_1 _12631_ (.A(_03414_),
    .X(_03573_));
 sg13g2_nor2b_1 _12632_ (.A(net50),
    .B_N(_03559_),
    .Y(_03574_));
 sg13g2_a21oi_1 _12633_ (.A1(net50),
    .A2(_03561_),
    .Y(_03575_),
    .B1(_03574_));
 sg13g2_xnor2_1 _12634_ (.Y(_03576_),
    .A(net53),
    .B(_03575_));
 sg13g2_a21o_1 _12635_ (.A2(_03560_),
    .A1(_03014_),
    .B1(_02987_),
    .X(_03577_));
 sg13g2_xnor2_1 _12636_ (.Y(_03578_),
    .A(_02980_),
    .B(_03577_));
 sg13g2_xnor2_1 _12637_ (.Y(_03579_),
    .A(_02980_),
    .B(_03438_));
 sg13g2_nor2_1 _12638_ (.A(_03579_),
    .B(_03424_),
    .Y(_03580_));
 sg13g2_a21oi_1 _12639_ (.A1(_03424_),
    .A2(_03578_),
    .Y(_03581_),
    .B1(_03580_));
 sg13g2_inv_1 _12640_ (.Y(_03582_),
    .A(_03581_));
 sg13g2_nand2_1 _12641_ (.Y(_03583_),
    .A(_03498_),
    .B(_03582_));
 sg13g2_nand3_1 _12642_ (.B(_03496_),
    .C(_03581_),
    .A(_03426_),
    .Y(_03584_));
 sg13g2_nand2_1 _12643_ (.Y(_03585_),
    .A(_03583_),
    .B(_03584_));
 sg13g2_nand2b_1 _12644_ (.Y(_03586_),
    .B(_03585_),
    .A_N(_03576_));
 sg13g2_nand3_1 _12645_ (.B(_03584_),
    .C(_03576_),
    .A(_03583_),
    .Y(_03587_));
 sg13g2_nand2_1 _12646_ (.Y(_03588_),
    .A(_03586_),
    .B(_03587_));
 sg13g2_nor2_1 _12647_ (.A(_03579_),
    .B(net50),
    .Y(_03589_));
 sg13g2_a21oi_1 _12648_ (.A1(net50),
    .A2(_03578_),
    .Y(_03590_),
    .B1(_03589_));
 sg13g2_xnor2_1 _12649_ (.Y(_03591_),
    .A(net52),
    .B(_03590_));
 sg13g2_xnor2_1 _12650_ (.Y(_03592_),
    .A(_03444_),
    .B(_03440_));
 sg13g2_a21o_1 _12651_ (.A2(_02980_),
    .A1(_03577_),
    .B1(_02988_),
    .X(_03593_));
 sg13g2_xnor2_1 _12652_ (.Y(_03594_),
    .A(_02990_),
    .B(_03593_));
 sg13g2_mux2_1 _12653_ (.A0(_03592_),
    .A1(_03594_),
    .S(_03424_),
    .X(_03595_));
 sg13g2_xor2_1 _12654_ (.B(_03498_),
    .A(_03595_),
    .X(_03596_));
 sg13g2_nand2b_1 _12655_ (.Y(_03597_),
    .B(_03596_),
    .A_N(_03591_));
 sg13g2_xnor2_1 _12656_ (.Y(_03598_),
    .A(_03595_),
    .B(net40));
 sg13g2_nand2_1 _12657_ (.Y(_03599_),
    .A(_03598_),
    .B(_03591_));
 sg13g2_nand2_1 _12658_ (.Y(_03600_),
    .A(_03597_),
    .B(_03599_));
 sg13g2_nor2_1 _12659_ (.A(_03588_),
    .B(_03600_),
    .Y(_03601_));
 sg13g2_nand3_1 _12660_ (.B(_03572_),
    .C(_03601_),
    .A(_03570_),
    .Y(_03602_));
 sg13g2_buf_1 _12661_ (.A(_03602_),
    .X(_03603_));
 sg13g2_inv_1 _12662_ (.Y(_03604_),
    .A(_03586_));
 sg13g2_nor2b_1 _12663_ (.A(_03596_),
    .B_N(_03591_),
    .Y(_03605_));
 sg13g2_a21oi_1 _12664_ (.A1(_03604_),
    .A2(_03597_),
    .Y(_03606_),
    .B1(_03605_));
 sg13g2_nand2_1 _12665_ (.Y(_03607_),
    .A(_03603_),
    .B(_03606_));
 sg13g2_nor2b_1 _12666_ (.A(net49),
    .B_N(_03592_),
    .Y(_03608_));
 sg13g2_a21oi_1 _12667_ (.A1(_03594_),
    .A2(net49),
    .Y(_03609_),
    .B1(_03608_));
 sg13g2_xnor2_1 _12668_ (.Y(_03610_),
    .A(net53),
    .B(_03609_));
 sg13g2_a21oi_1 _12669_ (.A1(_03593_),
    .A2(_02990_),
    .Y(_03611_),
    .B1(_02973_));
 sg13g2_xor2_1 _12670_ (.B(_03611_),
    .A(_02963_),
    .X(_03612_));
 sg13g2_buf_8 _12671_ (.A(_03424_),
    .X(_03613_));
 sg13g2_a21o_1 _12672_ (.A2(_03443_),
    .A1(_03440_),
    .B1(_03442_),
    .X(_03614_));
 sg13g2_xnor2_1 _12673_ (.Y(_03615_),
    .A(_02963_),
    .B(_03614_));
 sg13g2_nor2_1 _12674_ (.A(_03615_),
    .B(_03424_),
    .Y(_03616_));
 sg13g2_a21oi_1 _12675_ (.A1(_03612_),
    .A2(_03613_),
    .Y(_03617_),
    .B1(_03616_));
 sg13g2_xnor2_1 _12676_ (.Y(_03618_),
    .A(_03617_),
    .B(net40));
 sg13g2_nor2_1 _12677_ (.A(_03610_),
    .B(_03618_),
    .Y(_03619_));
 sg13g2_nand2_1 _12678_ (.Y(_03620_),
    .A(_03618_),
    .B(_03610_));
 sg13g2_nor2b_1 _12679_ (.A(_03619_),
    .B_N(_03620_),
    .Y(_03621_));
 sg13g2_inv_2 _12680_ (.Y(_03622_),
    .A(_03621_));
 sg13g2_nor2_1 _12681_ (.A(_03615_),
    .B(net49),
    .Y(_03623_));
 sg13g2_a21oi_1 _12682_ (.A1(_03612_),
    .A2(net49),
    .Y(_03624_),
    .B1(_03623_));
 sg13g2_xnor2_1 _12683_ (.Y(_03625_),
    .A(net53),
    .B(_03624_));
 sg13g2_xnor2_1 _12684_ (.Y(_03626_),
    .A(_03156_),
    .B(_03020_));
 sg13g2_inv_1 _12685_ (.Y(_03627_),
    .A(_03453_));
 sg13g2_nand2_1 _12686_ (.Y(_03628_),
    .A(_03500_),
    .B(_03627_));
 sg13g2_nand2_1 _12687_ (.Y(_03629_),
    .A(_03628_),
    .B(_03454_));
 sg13g2_nand2_1 _12688_ (.Y(_03630_),
    .A(net49),
    .B(_03629_));
 sg13g2_o21ai_1 _12689_ (.B1(_03630_),
    .Y(_03631_),
    .A1(net49),
    .A2(_03626_));
 sg13g2_xor2_1 _12690_ (.B(net40),
    .A(_03631_),
    .X(_03632_));
 sg13g2_nor2_1 _12691_ (.A(_03625_),
    .B(_03632_),
    .Y(_03633_));
 sg13g2_nand2_1 _12692_ (.Y(_03634_),
    .A(_03632_),
    .B(_03625_));
 sg13g2_nor2b_1 _12693_ (.A(_03633_),
    .B_N(_03634_),
    .Y(_03635_));
 sg13g2_inv_1 _12694_ (.Y(_03636_),
    .A(_03635_));
 sg13g2_nor2_1 _12695_ (.A(_03622_),
    .B(_03636_),
    .Y(_03637_));
 sg13g2_nand2_1 _12696_ (.Y(_03638_),
    .A(_03607_),
    .B(_03637_));
 sg13g2_a21o_1 _12697_ (.A2(_03619_),
    .A1(_03634_),
    .B1(_03633_),
    .X(_03639_));
 sg13g2_buf_1 _12698_ (.A(_03639_),
    .X(_03640_));
 sg13g2_nand2b_1 _12699_ (.Y(_03641_),
    .B(net48),
    .A_N(_03521_));
 sg13g2_o21ai_1 _12700_ (.B1(_03641_),
    .Y(_03642_),
    .A1(net48),
    .A2(_03520_));
 sg13g2_xnor2_1 _12701_ (.Y(_03643_),
    .A(_03642_),
    .B(net40));
 sg13g2_xnor2_1 _12702_ (.Y(_03644_),
    .A(_03150_),
    .B(_03502_));
 sg13g2_inv_1 _12703_ (.Y(_03645_),
    .A(_03156_));
 sg13g2_a21oi_1 _12704_ (.A1(_03020_),
    .A2(_03645_),
    .Y(_03646_),
    .B1(_03276_));
 sg13g2_xnor2_1 _12705_ (.Y(_03647_),
    .A(_03150_),
    .B(_03646_));
 sg13g2_mux2_1 _12706_ (.A0(_03644_),
    .A1(_03647_),
    .S(net49),
    .X(_03648_));
 sg13g2_xnor2_1 _12707_ (.Y(_03649_),
    .A(net52),
    .B(_03648_));
 sg13g2_nand2b_1 _12708_ (.Y(_03650_),
    .B(_03649_),
    .A_N(_03643_));
 sg13g2_nor2_1 _12709_ (.A(_03626_),
    .B(net48),
    .Y(_03651_));
 sg13g2_a21oi_1 _12710_ (.A1(net48),
    .A2(_03629_),
    .Y(_03652_),
    .B1(_03651_));
 sg13g2_xnor2_1 _12711_ (.Y(_03653_),
    .A(_03573_),
    .B(_03652_));
 sg13g2_mux2_1 _12712_ (.A0(_03644_),
    .A1(_03647_),
    .S(net48),
    .X(_03654_));
 sg13g2_xnor2_1 _12713_ (.Y(_03655_),
    .A(_03654_),
    .B(net40));
 sg13g2_nand2b_1 _12714_ (.Y(_03656_),
    .B(_03655_),
    .A_N(_03653_));
 sg13g2_inv_1 _12715_ (.Y(_03657_),
    .A(_03656_));
 sg13g2_nand2b_1 _12716_ (.Y(_03658_),
    .B(_03643_),
    .A_N(_03649_));
 sg13g2_inv_2 _12717_ (.Y(_03659_),
    .A(_03658_));
 sg13g2_a21oi_1 _12718_ (.A1(_03650_),
    .A2(_03657_),
    .Y(_03660_),
    .B1(_03659_));
 sg13g2_inv_1 _12719_ (.Y(_03661_),
    .A(_03660_));
 sg13g2_nor2_1 _12720_ (.A(_03640_),
    .B(_03661_),
    .Y(_03662_));
 sg13g2_nand2_1 _12721_ (.Y(_03663_),
    .A(_03638_),
    .B(_03662_));
 sg13g2_nor2b_1 _12722_ (.A(_03659_),
    .B_N(_03650_),
    .Y(_03664_));
 sg13g2_xnor2_1 _12723_ (.Y(_03665_),
    .A(_03653_),
    .B(_03655_));
 sg13g2_nand2_1 _12724_ (.Y(_03666_),
    .A(_03664_),
    .B(_03665_));
 sg13g2_nand2_1 _12725_ (.Y(_03667_),
    .A(_03666_),
    .B(_03660_));
 sg13g2_nand2_1 _12726_ (.Y(_03668_),
    .A(_03663_),
    .B(_03667_));
 sg13g2_xnor2_1 _12727_ (.Y(_03669_),
    .A(_03527_),
    .B(_03668_));
 sg13g2_nor2b_1 _12728_ (.A(_03640_),
    .B_N(_03606_),
    .Y(_03670_));
 sg13g2_nand2_1 _12729_ (.Y(_03671_),
    .A(_03603_),
    .B(_03670_));
 sg13g2_or2_1 _12730_ (.X(_03672_),
    .B(_03637_),
    .A(_03640_));
 sg13g2_buf_1 _12731_ (.A(_03672_),
    .X(_03673_));
 sg13g2_inv_4 _12732_ (.A(_03499_),
    .Y(_03674_));
 sg13g2_buf_8 _12733_ (.A(_03674_),
    .X(_03675_));
 sg13g2_a21o_1 _12734_ (.A2(_03470_),
    .A1(_03455_),
    .B1(_03489_),
    .X(_03676_));
 sg13g2_xnor2_1 _12735_ (.Y(_03677_),
    .A(_03460_),
    .B(_03676_));
 sg13g2_xnor2_1 _12736_ (.Y(_03678_),
    .A(_03393_),
    .B(_03283_));
 sg13g2_nor2_1 _12737_ (.A(_03510_),
    .B(_03678_),
    .Y(_03679_));
 sg13g2_a21oi_1 _12738_ (.A1(_03677_),
    .A2(net47),
    .Y(_03680_),
    .B1(_03679_));
 sg13g2_xnor2_1 _12739_ (.Y(_03681_),
    .A(net38),
    .B(_03680_));
 sg13g2_nor2_1 _12740_ (.A(net48),
    .B(_03514_),
    .Y(_03682_));
 sg13g2_a21oi_1 _12741_ (.A1(_03507_),
    .A2(_03613_),
    .Y(_03683_),
    .B1(_03682_));
 sg13g2_xnor2_1 _12742_ (.Y(_03684_),
    .A(net52),
    .B(_03683_));
 sg13g2_nand2b_1 _12743_ (.Y(_03685_),
    .B(_03684_),
    .A_N(_03681_));
 sg13g2_inv_2 _12744_ (.Y(_03686_),
    .A(_03685_));
 sg13g2_nand2b_1 _12745_ (.Y(_03687_),
    .B(_03681_),
    .A_N(_03684_));
 sg13g2_nor2b_1 _12746_ (.A(_03686_),
    .B_N(_03687_),
    .Y(_03688_));
 sg13g2_inv_2 _12747_ (.Y(_03689_),
    .A(_03527_));
 sg13g2_nand2_1 _12748_ (.Y(_03690_),
    .A(_03688_),
    .B(_03689_));
 sg13g2_nor2_1 _12749_ (.A(_03666_),
    .B(_03690_),
    .Y(_03691_));
 sg13g2_nand3_1 _12750_ (.B(_03673_),
    .C(_03691_),
    .A(_03671_),
    .Y(_03692_));
 sg13g2_inv_1 _12751_ (.Y(_03693_),
    .A(_03690_));
 sg13g2_inv_1 _12752_ (.Y(_03694_),
    .A(_03526_));
 sg13g2_a21oi_1 _12753_ (.A1(_03687_),
    .A2(_03694_),
    .Y(_03695_),
    .B1(_03686_));
 sg13g2_inv_1 _12754_ (.Y(_03696_),
    .A(_03695_));
 sg13g2_a21oi_1 _12755_ (.A1(_03693_),
    .A2(_03661_),
    .Y(_03697_),
    .B1(_03696_));
 sg13g2_nand2_1 _12756_ (.Y(_03698_),
    .A(_03692_),
    .B(_03697_));
 sg13g2_nand2_1 _12757_ (.Y(_03699_),
    .A(_03678_),
    .B(net47));
 sg13g2_o21ai_1 _12758_ (.B1(_03699_),
    .Y(_03700_),
    .A1(net47),
    .A2(_03677_));
 sg13g2_xnor2_1 _12759_ (.Y(_03701_),
    .A(_03518_),
    .B(_03700_));
 sg13g2_inv_1 _12760_ (.Y(_03702_),
    .A(_03701_));
 sg13g2_buf_1 _12761_ (.A(net48),
    .X(_03703_));
 sg13g2_nand3_1 _12762_ (.B(_03458_),
    .C(_03459_),
    .A(_03469_),
    .Y(_03704_));
 sg13g2_nor3_1 _12763_ (.A(_03427_),
    .B(_03467_),
    .C(_03704_),
    .Y(_03705_));
 sg13g2_a21oi_1 _12764_ (.A1(_03443_),
    .A2(_03428_),
    .Y(_03706_),
    .B1(_03442_));
 sg13g2_nor2_1 _12765_ (.A(_02963_),
    .B(_03627_),
    .Y(_03707_));
 sg13g2_inv_1 _12766_ (.Y(_03708_),
    .A(_03707_));
 sg13g2_a21oi_1 _12767_ (.A1(_03453_),
    .A2(_03446_),
    .Y(_03709_),
    .B1(_03450_));
 sg13g2_o21ai_1 _12768_ (.B1(_03709_),
    .Y(_03710_),
    .A1(_03706_),
    .A2(_03708_));
 sg13g2_o21ai_1 _12769_ (.B1(_03459_),
    .Y(_03711_),
    .A1(_03487_),
    .A2(_03457_));
 sg13g2_o21ai_1 _12770_ (.B1(_03711_),
    .Y(_03712_),
    .A1(_03505_),
    .A2(_03704_));
 sg13g2_a21oi_1 _12771_ (.A1(_03705_),
    .A2(_03710_),
    .Y(_03713_),
    .B1(_03712_));
 sg13g2_nand2_1 _12772_ (.Y(_03714_),
    .A(_03444_),
    .B(_03017_));
 sg13g2_nor2_1 _12773_ (.A(_03714_),
    .B(_03708_),
    .Y(_03715_));
 sg13g2_nand3_1 _12774_ (.B(_03438_),
    .C(_03715_),
    .A(_03705_),
    .Y(_03716_));
 sg13g2_nand2_1 _12775_ (.Y(_03717_),
    .A(_03713_),
    .B(_03716_));
 sg13g2_xnor2_1 _12776_ (.Y(_03718_),
    .A(_03462_),
    .B(_03717_));
 sg13g2_inv_1 _12777_ (.Y(_03719_),
    .A(_03718_));
 sg13g2_nor2b_1 _12778_ (.A(_03469_),
    .B_N(_03393_),
    .Y(_03720_));
 sg13g2_inv_1 _12779_ (.Y(_03721_),
    .A(_03260_));
 sg13g2_a21o_1 _12780_ (.A2(_03721_),
    .A1(_03393_),
    .B1(_03400_),
    .X(_03722_));
 sg13g2_a21oi_1 _12781_ (.A1(_03513_),
    .A2(_03720_),
    .Y(_03723_),
    .B1(_03722_));
 sg13g2_xnor2_1 _12782_ (.Y(_03724_),
    .A(_03462_),
    .B(_03723_));
 sg13g2_nand2_1 _12783_ (.Y(_03725_),
    .A(_03724_),
    .B(net48));
 sg13g2_o21ai_1 _12784_ (.B1(_03725_),
    .Y(_03726_),
    .A1(net46),
    .A2(_03719_));
 sg13g2_xnor2_1 _12785_ (.Y(_03727_),
    .A(_03499_),
    .B(_03726_));
 sg13g2_xnor2_1 _12786_ (.Y(_03728_),
    .A(_03702_),
    .B(_03727_));
 sg13g2_buf_2 _12787_ (.A(_03728_),
    .X(_03729_));
 sg13g2_inv_1 _12788_ (.Y(_03730_),
    .A(_03729_));
 sg13g2_nand2_1 _12789_ (.Y(_03731_),
    .A(_03698_),
    .B(_03730_));
 sg13g2_nand3_1 _12790_ (.B(_03697_),
    .C(_03729_),
    .A(_03692_),
    .Y(_03732_));
 sg13g2_nand2_1 _12791_ (.Y(_03733_),
    .A(_03731_),
    .B(_03732_));
 sg13g2_nand2_1 _12792_ (.Y(_03734_),
    .A(_03669_),
    .B(_03733_));
 sg13g2_xnor2_1 _12793_ (.Y(_03735_),
    .A(_03729_),
    .B(_03698_));
 sg13g2_nand2_1 _12794_ (.Y(_03736_),
    .A(_03668_),
    .B(_03689_));
 sg13g2_nand3_1 _12795_ (.B(_03527_),
    .C(_03667_),
    .A(_03663_),
    .Y(_03737_));
 sg13g2_nand2_2 _12796_ (.Y(_03738_),
    .A(_03736_),
    .B(_03737_));
 sg13g2_nand2_1 _12797_ (.Y(_03739_),
    .A(_03735_),
    .B(_03738_));
 sg13g2_nand2_1 _12798_ (.Y(_03740_),
    .A(_03734_),
    .B(_03739_));
 sg13g2_nand3_1 _12799_ (.B(_03548_),
    .C(_03550_),
    .A(_03552_),
    .Y(_03741_));
 sg13g2_nor2b_1 _12800_ (.A(_03542_),
    .B_N(_03532_),
    .Y(_03742_));
 sg13g2_o21ai_1 _12801_ (.B1(_03544_),
    .Y(_03743_),
    .A1(_03741_),
    .A2(_03742_));
 sg13g2_nand2_1 _12802_ (.Y(_03744_),
    .A(_03568_),
    .B(_03572_));
 sg13g2_nor2_1 _12803_ (.A(_03588_),
    .B(_03744_),
    .Y(_03745_));
 sg13g2_nand2_1 _12804_ (.Y(_03746_),
    .A(_03743_),
    .B(_03745_));
 sg13g2_nand2_1 _12805_ (.Y(_03747_),
    .A(_03568_),
    .B(_03586_));
 sg13g2_nand2_1 _12806_ (.Y(_03748_),
    .A(_03747_),
    .B(_03587_));
 sg13g2_nand2_1 _12807_ (.Y(_03749_),
    .A(_03746_),
    .B(_03748_));
 sg13g2_inv_1 _12808_ (.Y(_03750_),
    .A(_03600_));
 sg13g2_nand2_1 _12809_ (.Y(_03751_),
    .A(_03621_),
    .B(_03750_));
 sg13g2_inv_1 _12810_ (.Y(_03752_),
    .A(_03751_));
 sg13g2_nand2_1 _12811_ (.Y(_03753_),
    .A(_03749_),
    .B(_03752_));
 sg13g2_nand2_1 _12812_ (.Y(_03754_),
    .A(_03605_),
    .B(_03620_));
 sg13g2_nand2b_1 _12813_ (.Y(_03755_),
    .B(_03754_),
    .A_N(_03619_));
 sg13g2_inv_1 _12814_ (.Y(_03756_),
    .A(_03755_));
 sg13g2_nand2_1 _12815_ (.Y(_03757_),
    .A(_03753_),
    .B(_03756_));
 sg13g2_nand2_1 _12816_ (.Y(_03758_),
    .A(_03635_),
    .B(_03665_));
 sg13g2_nand2_1 _12817_ (.Y(_03759_),
    .A(_03664_),
    .B(_03689_));
 sg13g2_nor2_1 _12818_ (.A(_03758_),
    .B(_03759_),
    .Y(_03760_));
 sg13g2_nand2_1 _12819_ (.Y(_03761_),
    .A(_03757_),
    .B(_03760_));
 sg13g2_a21o_1 _12820_ (.A2(_03659_),
    .A1(_03525_),
    .B1(_03694_),
    .X(_03762_));
 sg13g2_inv_1 _12821_ (.Y(_03763_),
    .A(_03633_));
 sg13g2_nor2b_1 _12822_ (.A(_03655_),
    .B_N(_03653_),
    .Y(_03764_));
 sg13g2_o21ai_1 _12823_ (.B1(_03656_),
    .Y(_03765_),
    .A1(_03763_),
    .A2(_03764_));
 sg13g2_nor2b_1 _12824_ (.A(_03759_),
    .B_N(_03765_),
    .Y(_03766_));
 sg13g2_nor2_1 _12825_ (.A(_03762_),
    .B(_03766_),
    .Y(_03767_));
 sg13g2_nand2_1 _12826_ (.Y(_03768_),
    .A(_03761_),
    .B(_03767_));
 sg13g2_inv_2 _12827_ (.Y(_03769_),
    .A(_03688_));
 sg13g2_nand2_1 _12828_ (.Y(_03770_),
    .A(_03768_),
    .B(_03769_));
 sg13g2_nand3_1 _12829_ (.B(_03688_),
    .C(_03767_),
    .A(_03761_),
    .Y(_03771_));
 sg13g2_nand2_2 _12830_ (.Y(_03772_),
    .A(_03770_),
    .B(_03771_));
 sg13g2_nor2_1 _12831_ (.A(_03751_),
    .B(_03758_),
    .Y(_03773_));
 sg13g2_nand2_1 _12832_ (.Y(_03774_),
    .A(_03749_),
    .B(_03773_));
 sg13g2_nor2_1 _12833_ (.A(_03756_),
    .B(_03758_),
    .Y(_03775_));
 sg13g2_nor2_1 _12834_ (.A(_03765_),
    .B(_03775_),
    .Y(_03776_));
 sg13g2_nand2_1 _12835_ (.Y(_03777_),
    .A(_03774_),
    .B(_03776_));
 sg13g2_xnor2_1 _12836_ (.Y(_03778_),
    .A(_03664_),
    .B(_03777_));
 sg13g2_inv_2 _12837_ (.Y(_03779_),
    .A(_03778_));
 sg13g2_nand2_1 _12838_ (.Y(_03780_),
    .A(_03772_),
    .B(_03779_));
 sg13g2_inv_1 _12839_ (.Y(_03781_),
    .A(_03780_));
 sg13g2_nand2_1 _12840_ (.Y(_03782_),
    .A(_03740_),
    .B(_03781_));
 sg13g2_inv_1 _12841_ (.Y(_03783_),
    .A(_03782_));
 sg13g2_nor2_1 _12842_ (.A(_03738_),
    .B(_03735_),
    .Y(_03784_));
 sg13g2_inv_1 _12843_ (.Y(_03785_),
    .A(_03772_));
 sg13g2_nand2_1 _12844_ (.Y(_03786_),
    .A(_03724_),
    .B(net47));
 sg13g2_o21ai_1 _12845_ (.B1(_03786_),
    .Y(_03787_),
    .A1(net47),
    .A2(_03719_));
 sg13g2_xnor2_1 _12846_ (.Y(_03788_),
    .A(_03573_),
    .B(_03787_));
 sg13g2_nand2_1 _12847_ (.Y(_03789_),
    .A(_03676_),
    .B(_03463_));
 sg13g2_nand2_1 _12848_ (.Y(_03790_),
    .A(_03789_),
    .B(_03472_));
 sg13g2_xnor2_1 _12849_ (.Y(_03791_),
    .A(_03476_),
    .B(_03790_));
 sg13g2_buf_1 _12850_ (.A(net47),
    .X(_03792_));
 sg13g2_nand2b_1 _12851_ (.Y(_03793_),
    .B(_03283_),
    .A_N(_03394_));
 sg13g2_nand2b_1 _12852_ (.Y(_03794_),
    .B(_03793_),
    .A_N(_03404_));
 sg13g2_xnor2_1 _12853_ (.Y(_03795_),
    .A(_03350_),
    .B(_03794_));
 sg13g2_nor2b_1 _12854_ (.A(net47),
    .B_N(_03795_),
    .Y(_03796_));
 sg13g2_a21oi_1 _12855_ (.A1(_03791_),
    .A2(_03792_),
    .Y(_03797_),
    .B1(_03796_));
 sg13g2_xnor2_1 _12856_ (.Y(_03798_),
    .A(net38),
    .B(_03797_));
 sg13g2_xnor2_1 _12857_ (.Y(_03799_),
    .A(_03788_),
    .B(_03798_));
 sg13g2_nor3_1 _12858_ (.A(_03769_),
    .B(_03729_),
    .C(_03759_),
    .Y(_03800_));
 sg13g2_nand2_1 _12859_ (.Y(_03801_),
    .A(_03777_),
    .B(_03800_));
 sg13g2_nor2_1 _12860_ (.A(_03769_),
    .B(_03729_),
    .Y(_03802_));
 sg13g2_o21ai_1 _12861_ (.B1(_03686_),
    .Y(_03803_),
    .A1(_03702_),
    .A2(_03727_));
 sg13g2_nand2_1 _12862_ (.Y(_03804_),
    .A(_03727_),
    .B(_03702_));
 sg13g2_nand2_1 _12863_ (.Y(_03805_),
    .A(_03803_),
    .B(_03804_));
 sg13g2_a21oi_1 _12864_ (.A1(_03802_),
    .A2(_03762_),
    .Y(_03806_),
    .B1(_03805_));
 sg13g2_nand2_1 _12865_ (.Y(_03807_),
    .A(_03801_),
    .B(_03806_));
 sg13g2_xnor2_1 _12866_ (.Y(_03808_),
    .A(_03799_),
    .B(_03807_));
 sg13g2_nand2_2 _12867_ (.Y(_03809_),
    .A(_03785_),
    .B(_03808_));
 sg13g2_inv_1 _12868_ (.Y(_03810_),
    .A(_03799_));
 sg13g2_nand2_1 _12869_ (.Y(_03811_),
    .A(_03807_),
    .B(_03810_));
 sg13g2_nand3_1 _12870_ (.B(_03806_),
    .C(_03799_),
    .A(_03801_),
    .Y(_03812_));
 sg13g2_nand2_1 _12871_ (.Y(_03813_),
    .A(_03811_),
    .B(_03812_));
 sg13g2_nand2_1 _12872_ (.Y(_03814_),
    .A(_03772_),
    .B(_03813_));
 sg13g2_nand3_1 _12873_ (.B(_03809_),
    .C(_03814_),
    .A(_03784_),
    .Y(_03815_));
 sg13g2_nand2_1 _12874_ (.Y(_03816_),
    .A(_03783_),
    .B(_03815_));
 sg13g2_nand2_1 _12875_ (.Y(_03817_),
    .A(_03809_),
    .B(_03814_));
 sg13g2_nand2_1 _12876_ (.Y(_03818_),
    .A(_03817_),
    .B(_03734_));
 sg13g2_nand2_1 _12877_ (.Y(_03819_),
    .A(_03816_),
    .B(_03818_));
 sg13g2_nand2_1 _12878_ (.Y(_03820_),
    .A(_03815_),
    .B(_03818_));
 sg13g2_nand3_1 _12879_ (.B(_03739_),
    .C(_03780_),
    .A(_03734_),
    .Y(_03821_));
 sg13g2_nand2_1 _12880_ (.Y(_03822_),
    .A(_03782_),
    .B(_03821_));
 sg13g2_nor2_1 _12881_ (.A(_03820_),
    .B(_03822_),
    .Y(_03823_));
 sg13g2_nand2_1 _12882_ (.Y(_03824_),
    .A(_03671_),
    .B(_03673_));
 sg13g2_inv_1 _12883_ (.Y(_03825_),
    .A(_03665_));
 sg13g2_nand2_1 _12884_ (.Y(_03826_),
    .A(_03824_),
    .B(_03825_));
 sg13g2_nand3_1 _12885_ (.B(_03665_),
    .C(_03673_),
    .A(_03671_),
    .Y(_03827_));
 sg13g2_nand2_1 _12886_ (.Y(_03828_),
    .A(_03826_),
    .B(_03827_));
 sg13g2_inv_1 _12887_ (.Y(_03829_),
    .A(_03828_));
 sg13g2_nand2_2 _12888_ (.Y(_03830_),
    .A(_03738_),
    .B(_03829_));
 sg13g2_nand3_1 _12889_ (.B(_03737_),
    .C(_03828_),
    .A(_03736_),
    .Y(_03831_));
 sg13g2_nand2_1 _12890_ (.Y(_03832_),
    .A(_03757_),
    .B(_03635_));
 sg13g2_nand3_1 _12891_ (.B(_03636_),
    .C(_03756_),
    .A(_03753_),
    .Y(_03833_));
 sg13g2_nand2_1 _12892_ (.Y(_03834_),
    .A(_03832_),
    .B(_03833_));
 sg13g2_nor2_1 _12893_ (.A(_03834_),
    .B(_03778_),
    .Y(_03835_));
 sg13g2_nand3_1 _12894_ (.B(_03831_),
    .C(_03835_),
    .A(_03830_),
    .Y(_03836_));
 sg13g2_buf_1 _12895_ (.A(_03836_),
    .X(_03837_));
 sg13g2_xnor2_1 _12896_ (.Y(_03838_),
    .A(_03778_),
    .B(_03772_));
 sg13g2_inv_2 _12897_ (.Y(_03839_),
    .A(_03830_));
 sg13g2_nand2_1 _12898_ (.Y(_03840_),
    .A(_03838_),
    .B(_03839_));
 sg13g2_xnor2_1 _12899_ (.Y(_03841_),
    .A(_03779_),
    .B(_03772_));
 sg13g2_nand2_1 _12900_ (.Y(_03842_),
    .A(_03841_),
    .B(_03830_));
 sg13g2_inv_1 _12901_ (.Y(_03843_),
    .A(_03842_));
 sg13g2_a21oi_1 _12902_ (.A1(_03837_),
    .A2(_03840_),
    .Y(_03844_),
    .B1(_03843_));
 sg13g2_nand2_1 _12903_ (.Y(_03845_),
    .A(_03823_),
    .B(_03844_));
 sg13g2_nand2b_1 _12904_ (.Y(_03846_),
    .B(_03845_),
    .A_N(_03819_));
 sg13g2_xnor2_1 _12905_ (.Y(_03847_),
    .A(_03600_),
    .B(_03749_));
 sg13g2_inv_1 _12906_ (.Y(_03848_),
    .A(_03847_));
 sg13g2_xnor2_1 _12907_ (.Y(_03849_),
    .A(_03744_),
    .B(_03743_));
 sg13g2_nor2b_1 _12908_ (.A(_03848_),
    .B_N(_03849_),
    .Y(_03850_));
 sg13g2_nand2_1 _12909_ (.Y(_03851_),
    .A(_03570_),
    .B(_03572_));
 sg13g2_xnor2_1 _12910_ (.Y(_03852_),
    .A(_03588_),
    .B(_03851_));
 sg13g2_nand2_1 _12911_ (.Y(_03853_),
    .A(_03607_),
    .B(_03621_));
 sg13g2_nand3_1 _12912_ (.B(_03606_),
    .C(_03622_),
    .A(_03603_),
    .Y(_03854_));
 sg13g2_nand3b_1 _12913_ (.B(_03853_),
    .C(_03854_),
    .Y(_03855_),
    .A_N(_03852_));
 sg13g2_buf_1 _12914_ (.A(_03855_),
    .X(_03856_));
 sg13g2_nand2_1 _12915_ (.Y(_03857_),
    .A(_03853_),
    .B(_03854_));
 sg13g2_nand2_1 _12916_ (.Y(_03858_),
    .A(_03857_),
    .B(_03852_));
 sg13g2_nand2_1 _12917_ (.Y(_03859_),
    .A(_03856_),
    .B(_03858_));
 sg13g2_nand2b_1 _12918_ (.Y(_03860_),
    .B(_03859_),
    .A_N(_03850_));
 sg13g2_nand3_1 _12919_ (.B(_03858_),
    .C(_03850_),
    .A(_03856_),
    .Y(_03861_));
 sg13g2_buf_1 _12920_ (.A(_03861_),
    .X(_03862_));
 sg13g2_a21oi_1 _12921_ (.A1(_03544_),
    .A2(_03554_),
    .Y(_03863_),
    .B1(_03553_));
 sg13g2_nor2b_1 _12922_ (.A(_03863_),
    .B_N(_03555_),
    .Y(_03864_));
 sg13g2_nand2b_1 _12923_ (.Y(_03865_),
    .B(_03864_),
    .A_N(_03852_));
 sg13g2_xnor2_1 _12924_ (.Y(_03866_),
    .A(_03849_),
    .B(_03847_));
 sg13g2_nor2_1 _12925_ (.A(_03865_),
    .B(_03866_),
    .Y(_03867_));
 sg13g2_nand3_1 _12926_ (.B(_03862_),
    .C(_03867_),
    .A(_03860_),
    .Y(_03868_));
 sg13g2_inv_1 _12927_ (.Y(_03869_),
    .A(_03862_));
 sg13g2_nand2_1 _12928_ (.Y(_03870_),
    .A(_03834_),
    .B(_03848_));
 sg13g2_nand3_1 _12929_ (.B(_03833_),
    .C(_03847_),
    .A(_03832_),
    .Y(_03871_));
 sg13g2_buf_1 _12930_ (.A(_03871_),
    .X(_03872_));
 sg13g2_nand2_1 _12931_ (.Y(_03873_),
    .A(_03870_),
    .B(_03872_));
 sg13g2_nor2_1 _12932_ (.A(_03856_),
    .B(_03873_),
    .Y(_03874_));
 sg13g2_nor2_1 _12933_ (.A(_03869_),
    .B(_03874_),
    .Y(_03875_));
 sg13g2_nand2_1 _12934_ (.Y(_03876_),
    .A(_03873_),
    .B(_03856_));
 sg13g2_inv_1 _12935_ (.Y(_03877_),
    .A(_03876_));
 sg13g2_a21oi_1 _12936_ (.A1(_03868_),
    .A2(_03875_),
    .Y(_03878_),
    .B1(_03877_));
 sg13g2_xnor2_1 _12937_ (.Y(_03879_),
    .A(_03622_),
    .B(_03607_));
 sg13g2_nand3_1 _12938_ (.B(_03826_),
    .C(_03827_),
    .A(_03879_),
    .Y(_03880_));
 sg13g2_buf_1 _12939_ (.A(_03880_),
    .X(_03881_));
 sg13g2_nand2_1 _12940_ (.Y(_03882_),
    .A(_03828_),
    .B(_03857_));
 sg13g2_nand2_1 _12941_ (.Y(_03883_),
    .A(_03881_),
    .B(_03882_));
 sg13g2_nand2_1 _12942_ (.Y(_03884_),
    .A(_03883_),
    .B(_03872_));
 sg13g2_inv_1 _12943_ (.Y(_03885_),
    .A(_03872_));
 sg13g2_nand3_1 _12944_ (.B(_03882_),
    .C(_03885_),
    .A(_03881_),
    .Y(_03886_));
 sg13g2_nand2_1 _12945_ (.Y(_03887_),
    .A(_03884_),
    .B(_03886_));
 sg13g2_xnor2_1 _12946_ (.Y(_03888_),
    .A(_03834_),
    .B(_03778_));
 sg13g2_nor2_1 _12947_ (.A(_03881_),
    .B(_03888_),
    .Y(_03889_));
 sg13g2_nand2_1 _12948_ (.Y(_03890_),
    .A(_03888_),
    .B(_03881_));
 sg13g2_nand2b_1 _12949_ (.Y(_03891_),
    .B(_03890_),
    .A_N(_03889_));
 sg13g2_nor2_1 _12950_ (.A(_03887_),
    .B(_03891_),
    .Y(_03892_));
 sg13g2_inv_1 _12951_ (.Y(_03893_),
    .A(_03886_));
 sg13g2_a21oi_1 _12952_ (.A1(_03893_),
    .A2(_03890_),
    .Y(_03894_),
    .B1(_03889_));
 sg13g2_inv_1 _12953_ (.Y(_03895_),
    .A(_03894_));
 sg13g2_a21oi_1 _12954_ (.A1(_03878_),
    .A2(_03892_),
    .Y(_03896_),
    .B1(_03895_));
 sg13g2_nand2_1 _12955_ (.Y(_03897_),
    .A(_03842_),
    .B(_03840_));
 sg13g2_nand2_1 _12956_ (.Y(_03898_),
    .A(_03830_),
    .B(_03831_));
 sg13g2_inv_1 _12957_ (.Y(_03899_),
    .A(_03835_));
 sg13g2_nand2_1 _12958_ (.Y(_03900_),
    .A(_03898_),
    .B(_03899_));
 sg13g2_nand2_1 _12959_ (.Y(_03901_),
    .A(_03900_),
    .B(_03837_));
 sg13g2_nor2_1 _12960_ (.A(_03897_),
    .B(_03901_),
    .Y(_03902_));
 sg13g2_nand2_1 _12961_ (.Y(_03903_),
    .A(_03823_),
    .B(_03902_));
 sg13g2_nor2_1 _12962_ (.A(_03896_),
    .B(_03903_),
    .Y(_03904_));
 sg13g2_nor2_1 _12963_ (.A(_03846_),
    .B(_03904_),
    .Y(_03905_));
 sg13g2_mux2_1 _12964_ (.A0(_03795_),
    .A1(_03791_),
    .S(net46),
    .X(_03906_));
 sg13g2_xnor2_1 _12965_ (.Y(_03907_),
    .A(_03518_),
    .B(_03906_));
 sg13g2_nand2b_1 _12966_ (.Y(_03908_),
    .B(_03384_),
    .A_N(_03723_));
 sg13g2_a21oi_1 _12967_ (.A1(_03908_),
    .A2(_03403_),
    .Y(_03909_),
    .B1(_03350_));
 sg13g2_nor2b_1 _12968_ (.A(_03909_),
    .B_N(_03406_),
    .Y(_03910_));
 sg13g2_xnor2_1 _12969_ (.Y(_03911_),
    .A(_03370_),
    .B(_03910_));
 sg13g2_nand2_1 _12970_ (.Y(_03912_),
    .A(_03717_),
    .B(_03462_));
 sg13g2_nand3_1 _12971_ (.B(_03382_),
    .C(_03474_),
    .A(_03912_),
    .Y(_03913_));
 sg13g2_nand2_1 _12972_ (.Y(_03914_),
    .A(_03913_),
    .B(_03475_));
 sg13g2_xnor2_1 _12973_ (.Y(_03915_),
    .A(_03478_),
    .B(_03914_));
 sg13g2_nor2b_1 _12974_ (.A(_03703_),
    .B_N(_03915_),
    .Y(_03916_));
 sg13g2_a21oi_1 _12975_ (.A1(_03911_),
    .A2(_03703_),
    .Y(_03917_),
    .B1(_03916_));
 sg13g2_xnor2_1 _12976_ (.Y(_03918_),
    .A(_03675_),
    .B(_03917_));
 sg13g2_or2_1 _12977_ (.X(_03919_),
    .B(_03918_),
    .A(_03907_));
 sg13g2_buf_1 _12978_ (.A(_03919_),
    .X(_03920_));
 sg13g2_nand2_1 _12979_ (.Y(_03921_),
    .A(_03918_),
    .B(_03907_));
 sg13g2_nand2_1 _12980_ (.Y(_03922_),
    .A(_03920_),
    .B(_03921_));
 sg13g2_nand3_1 _12981_ (.B(_03667_),
    .C(_03693_),
    .A(_03663_),
    .Y(_03923_));
 sg13g2_nand2_1 _12982_ (.Y(_03924_),
    .A(_03923_),
    .B(_03695_));
 sg13g2_nor2_1 _12983_ (.A(_03729_),
    .B(_03810_),
    .Y(_03925_));
 sg13g2_nand2_1 _12984_ (.Y(_03926_),
    .A(_03924_),
    .B(_03925_));
 sg13g2_inv_1 _12985_ (.Y(_03927_),
    .A(_03804_));
 sg13g2_nor2b_1 _12986_ (.A(_03798_),
    .B_N(_03788_),
    .Y(_03928_));
 sg13g2_a21oi_1 _12987_ (.A1(_03799_),
    .A2(_03927_),
    .Y(_03929_),
    .B1(_03928_));
 sg13g2_nand3b_1 _12988_ (.B(_03926_),
    .C(_03929_),
    .Y(_03930_),
    .A_N(_03922_));
 sg13g2_nand2_1 _12989_ (.Y(_03931_),
    .A(_03926_),
    .B(_03929_));
 sg13g2_nand2_1 _12990_ (.Y(_03932_),
    .A(_03931_),
    .B(_03922_));
 sg13g2_nand2_2 _12991_ (.Y(_03933_),
    .A(_03930_),
    .B(_03932_));
 sg13g2_nand2_1 _12992_ (.Y(_03934_),
    .A(_03933_),
    .B(_03735_));
 sg13g2_nand3_1 _12993_ (.B(_03932_),
    .C(_03733_),
    .A(_03930_),
    .Y(_03935_));
 sg13g2_buf_1 _12994_ (.A(_03935_),
    .X(_03936_));
 sg13g2_nand2_2 _12995_ (.Y(_03937_),
    .A(_03934_),
    .B(_03936_));
 sg13g2_xnor2_1 _12996_ (.Y(_03938_),
    .A(_03809_),
    .B(_03937_));
 sg13g2_nand2_1 _12997_ (.Y(_03939_),
    .A(_03905_),
    .B(_03938_));
 sg13g2_buf_8 _12998_ (.A(_03939_),
    .X(_03940_));
 sg13g2_xnor2_1 _12999_ (.Y(_03941_),
    .A(_03835_),
    .B(_03898_));
 sg13g2_xnor2_1 _13000_ (.Y(_03942_),
    .A(_03839_),
    .B(_03841_));
 sg13g2_nand2_1 _13001_ (.Y(_03943_),
    .A(_03941_),
    .B(_03942_));
 sg13g2_xnor2_1 _13002_ (.Y(_03944_),
    .A(_03733_),
    .B(_03738_));
 sg13g2_xnor2_1 _13003_ (.Y(_03945_),
    .A(_03781_),
    .B(_03944_));
 sg13g2_xnor2_1 _13004_ (.Y(_03946_),
    .A(_03784_),
    .B(_03817_));
 sg13g2_nand2_1 _13005_ (.Y(_03947_),
    .A(_03945_),
    .B(_03946_));
 sg13g2_nor2_1 _13006_ (.A(_03943_),
    .B(_03947_),
    .Y(_03948_));
 sg13g2_nand2_1 _13007_ (.Y(_03949_),
    .A(_03878_),
    .B(_03892_));
 sg13g2_nand2_1 _13008_ (.Y(_03950_),
    .A(_03949_),
    .B(_03894_));
 sg13g2_nand2_1 _13009_ (.Y(_03951_),
    .A(_03948_),
    .B(_03950_));
 sg13g2_a21oi_1 _13010_ (.A1(_03823_),
    .A2(_03844_),
    .Y(_03952_),
    .B1(_03819_));
 sg13g2_nand2_1 _13011_ (.Y(_03953_),
    .A(_03951_),
    .B(_03952_));
 sg13g2_inv_1 _13012_ (.Y(_03954_),
    .A(_03809_));
 sg13g2_xnor2_1 _13013_ (.Y(_03955_),
    .A(_03954_),
    .B(_03937_));
 sg13g2_nand2_1 _13014_ (.Y(_03956_),
    .A(_03953_),
    .B(_03955_));
 sg13g2_buf_8 _13015_ (.A(_03956_),
    .X(_03957_));
 sg13g2_nand2_1 _13016_ (.Y(_03958_),
    .A(_03940_),
    .B(_03957_));
 sg13g2_buf_8 _13017_ (.A(_03958_),
    .X(_03959_));
 sg13g2_buf_8 _13018_ (.A(_03959_),
    .X(_03960_));
 sg13g2_buf_8 _13019_ (.A(_03960_),
    .X(_03961_));
 sg13g2_buf_8 _13020_ (.A(_03961_),
    .X(_03962_));
 sg13g2_xnor2_1 _13021_ (.Y(_03963_),
    .A(\vgadonut.donut.donuthit.rx[13] ),
    .B(net35));
 sg13g2_buf_2 _13022_ (.A(_03963_),
    .X(_03964_));
 sg13g2_inv_1 _13023_ (.Y(_03965_),
    .A(_03964_));
 sg13g2_xnor2_1 _13024_ (.Y(_03966_),
    .A(_03856_),
    .B(_03873_));
 sg13g2_nor2_1 _13025_ (.A(_03966_),
    .B(_03887_),
    .Y(_03967_));
 sg13g2_a21oi_1 _13026_ (.A1(_03860_),
    .A2(_03867_),
    .Y(_03968_),
    .B1(_03869_));
 sg13g2_inv_1 _13027_ (.Y(_03969_),
    .A(_03968_));
 sg13g2_nand2_1 _13028_ (.Y(_03970_),
    .A(_03967_),
    .B(_03969_));
 sg13g2_a21oi_1 _13029_ (.A1(_03884_),
    .A2(_03874_),
    .Y(_03971_),
    .B1(_03893_));
 sg13g2_nand2_1 _13030_ (.Y(_03972_),
    .A(_03970_),
    .B(_03971_));
 sg13g2_xnor2_1 _13031_ (.Y(_03973_),
    .A(_03891_),
    .B(_03972_));
 sg13g2_buf_1 _13032_ (.A(_03973_),
    .X(_03974_));
 sg13g2_nand2b_1 _13033_ (.Y(_03975_),
    .B(net37),
    .A_N(_03974_));
 sg13g2_nand3_1 _13034_ (.B(_03957_),
    .C(_03974_),
    .A(_03940_),
    .Y(_03976_));
 sg13g2_nand2_1 _13035_ (.Y(_03977_),
    .A(_03975_),
    .B(_03976_));
 sg13g2_xnor2_1 _13036_ (.Y(_03978_),
    .A(_03887_),
    .B(_03878_));
 sg13g2_buf_1 _13037_ (.A(_03978_),
    .X(_03979_));
 sg13g2_inv_1 _13038_ (.Y(_03980_),
    .A(_03979_));
 sg13g2_nand2_1 _13039_ (.Y(_03981_),
    .A(net37),
    .B(_03980_));
 sg13g2_nand3_1 _13040_ (.B(_03957_),
    .C(_03979_),
    .A(_03940_),
    .Y(_03982_));
 sg13g2_nand2_1 _13041_ (.Y(_03983_),
    .A(_03981_),
    .B(_03982_));
 sg13g2_nand2_1 _13042_ (.Y(_03984_),
    .A(_03977_),
    .B(_03983_));
 sg13g2_xnor2_1 _13043_ (.Y(_03985_),
    .A(_03941_),
    .B(_03950_));
 sg13g2_xnor2_1 _13044_ (.Y(_03986_),
    .A(_03985_),
    .B(net37));
 sg13g2_nor2_1 _13045_ (.A(_03891_),
    .B(_03901_),
    .Y(_03987_));
 sg13g2_nand2_1 _13046_ (.Y(_03988_),
    .A(_03972_),
    .B(_03987_));
 sg13g2_inv_1 _13047_ (.Y(_03989_),
    .A(_03837_));
 sg13g2_a21oi_1 _13048_ (.A1(_03900_),
    .A2(_03889_),
    .Y(_03990_),
    .B1(_03989_));
 sg13g2_nand2_1 _13049_ (.Y(_03991_),
    .A(_03988_),
    .B(_03990_));
 sg13g2_xnor2_1 _13050_ (.Y(_03992_),
    .A(_03897_),
    .B(_03991_));
 sg13g2_inv_1 _13051_ (.Y(_03993_),
    .A(_03992_));
 sg13g2_nand2_1 _13052_ (.Y(_03994_),
    .A(net37),
    .B(_03993_));
 sg13g2_nand3_1 _13053_ (.B(_03957_),
    .C(_03992_),
    .A(_03940_),
    .Y(_03995_));
 sg13g2_nand2_1 _13054_ (.Y(_03996_),
    .A(_03994_),
    .B(_03995_));
 sg13g2_nand2_1 _13055_ (.Y(_03997_),
    .A(_03986_),
    .B(_03996_));
 sg13g2_nor2_1 _13056_ (.A(_03984_),
    .B(_03997_),
    .Y(_03998_));
 sg13g2_a21oi_1 _13057_ (.A1(_03950_),
    .A2(_03902_),
    .Y(_03999_),
    .B1(_03844_));
 sg13g2_xnor2_1 _13058_ (.Y(_04000_),
    .A(_03945_),
    .B(_03999_));
 sg13g2_xnor2_1 _13059_ (.Y(_04001_),
    .A(_04000_),
    .B(net37));
 sg13g2_nor2_1 _13060_ (.A(_03897_),
    .B(_03822_),
    .Y(_04002_));
 sg13g2_nand2_1 _13061_ (.Y(_04003_),
    .A(_03991_),
    .B(_04002_));
 sg13g2_inv_1 _13062_ (.Y(_04004_),
    .A(_03840_));
 sg13g2_a21oi_1 _13063_ (.A1(_04004_),
    .A2(_03821_),
    .Y(_04005_),
    .B1(_03783_));
 sg13g2_nand2_1 _13064_ (.Y(_04006_),
    .A(_04003_),
    .B(_04005_));
 sg13g2_xnor2_1 _13065_ (.Y(_04007_),
    .A(_03820_),
    .B(_04006_));
 sg13g2_nand2_1 _13066_ (.Y(_04008_),
    .A(_04007_),
    .B(_03959_));
 sg13g2_nand2_1 _13067_ (.Y(_04009_),
    .A(_04006_),
    .B(_03946_));
 sg13g2_nand3_1 _13068_ (.B(_03820_),
    .C(_04005_),
    .A(_04003_),
    .Y(_04010_));
 sg13g2_nand2_1 _13069_ (.Y(_04011_),
    .A(_04009_),
    .B(_04010_));
 sg13g2_xnor2_1 _13070_ (.Y(_04012_),
    .A(_03938_),
    .B(_03953_));
 sg13g2_nand2_1 _13071_ (.Y(_04013_),
    .A(_04011_),
    .B(_04012_));
 sg13g2_nand2_1 _13072_ (.Y(_04014_),
    .A(_04008_),
    .B(_04013_));
 sg13g2_buf_1 _13073_ (.A(_04014_),
    .X(_04015_));
 sg13g2_nor2_1 _13074_ (.A(_04001_),
    .B(net34),
    .Y(_04016_));
 sg13g2_buf_1 _13075_ (.A(_04016_),
    .X(_04017_));
 sg13g2_xor2_1 _13076_ (.B(_03968_),
    .A(_03966_),
    .X(_04018_));
 sg13g2_nand2_1 _13077_ (.Y(_04019_),
    .A(_03959_),
    .B(_04018_));
 sg13g2_inv_1 _13078_ (.Y(_04020_),
    .A(_04018_));
 sg13g2_nand3_1 _13079_ (.B(_03957_),
    .C(_04020_),
    .A(_03940_),
    .Y(_04021_));
 sg13g2_nand2_1 _13080_ (.Y(_04022_),
    .A(_04019_),
    .B(_04021_));
 sg13g2_nand3_1 _13081_ (.B(net30),
    .C(_04022_),
    .A(_03998_),
    .Y(_04023_));
 sg13g2_buf_1 _13082_ (.A(_04023_),
    .X(_04024_));
 sg13g2_nor2_1 _13083_ (.A(_03965_),
    .B(_04024_),
    .Y(_04025_));
 sg13g2_xnor2_1 _13084_ (.Y(_04026_),
    .A(_03959_),
    .B(_04011_));
 sg13g2_xor2_1 _13085_ (.B(_03959_),
    .A(_04000_),
    .X(_04027_));
 sg13g2_nand2_1 _13086_ (.Y(_04028_),
    .A(_04026_),
    .B(_04027_));
 sg13g2_buf_1 _13087_ (.A(_04028_),
    .X(_04029_));
 sg13g2_nor2_1 _13088_ (.A(_03997_),
    .B(_04029_),
    .Y(_04030_));
 sg13g2_buf_8 _13089_ (.A(_04030_),
    .X(_04031_));
 sg13g2_xnor2_1 _13090_ (.Y(_04032_),
    .A(_03974_),
    .B(_03959_));
 sg13g2_buf_2 _13091_ (.A(_04032_),
    .X(_04033_));
 sg13g2_xnor2_1 _13092_ (.Y(_04034_),
    .A(\vgadonut.donut.donuthit.rx[11] ),
    .B(net35));
 sg13g2_buf_1 _13093_ (.A(_04034_),
    .X(_04035_));
 sg13g2_nand3_1 _13094_ (.B(_04033_),
    .C(_04035_),
    .A(net26),
    .Y(_04036_));
 sg13g2_nor2b_1 _13095_ (.A(_04025_),
    .B_N(_04036_),
    .Y(_04037_));
 sg13g2_xnor2_1 _13096_ (.Y(_04038_),
    .A(\vgadonut.donut.donuthit.rx[12] ),
    .B(net35));
 sg13g2_buf_2 _13097_ (.A(_04038_),
    .X(_04039_));
 sg13g2_inv_1 _13098_ (.Y(_04040_),
    .A(_04039_));
 sg13g2_nor2_1 _13099_ (.A(_03983_),
    .B(_04033_),
    .Y(_04041_));
 sg13g2_buf_1 _13100_ (.A(_04041_),
    .X(_04042_));
 sg13g2_nand2_1 _13101_ (.Y(_04043_),
    .A(net26),
    .B(_04042_));
 sg13g2_buf_2 _13102_ (.A(_04043_),
    .X(_04044_));
 sg13g2_nor2_1 _13103_ (.A(_04040_),
    .B(_04044_),
    .Y(_04045_));
 sg13g2_xnor2_1 _13104_ (.Y(_04046_),
    .A(\vgadonut.donut.donuthit.rx[14] ),
    .B(_03962_));
 sg13g2_buf_2 _13105_ (.A(_04046_),
    .X(_04047_));
 sg13g2_inv_1 _13106_ (.Y(_04048_),
    .A(_04047_));
 sg13g2_inv_1 _13107_ (.Y(_04049_),
    .A(_04022_));
 sg13g2_a21oi_1 _13108_ (.A1(_03860_),
    .A2(_03862_),
    .Y(_04050_),
    .B1(_03867_));
 sg13g2_nand2b_1 _13109_ (.Y(_04051_),
    .B(_03868_),
    .A_N(_04050_));
 sg13g2_buf_1 _13110_ (.A(_04051_),
    .X(_04052_));
 sg13g2_nand2b_1 _13111_ (.Y(_04053_),
    .B(_03960_),
    .A_N(_04052_));
 sg13g2_nand3_1 _13112_ (.B(_03957_),
    .C(_04052_),
    .A(_03940_),
    .Y(_04054_));
 sg13g2_nand2_1 _13113_ (.Y(_04055_),
    .A(_04053_),
    .B(_04054_));
 sg13g2_nand2_1 _13114_ (.Y(_04056_),
    .A(_04049_),
    .B(_04055_));
 sg13g2_nor2_1 _13115_ (.A(_03984_),
    .B(_04056_),
    .Y(_04057_));
 sg13g2_nand2_1 _13116_ (.Y(_04058_),
    .A(_04030_),
    .B(_04057_));
 sg13g2_buf_2 _13117_ (.A(_04058_),
    .X(_04059_));
 sg13g2_nor2_1 _13118_ (.A(_04048_),
    .B(_04059_),
    .Y(_04060_));
 sg13g2_nor2_1 _13119_ (.A(_04045_),
    .B(_04060_),
    .Y(_04061_));
 sg13g2_nand2_1 _13120_ (.Y(_04062_),
    .A(_04037_),
    .B(_04061_));
 sg13g2_xnor2_1 _13121_ (.Y(_04063_),
    .A(_03979_),
    .B(net37));
 sg13g2_nor2_1 _13122_ (.A(_04033_),
    .B(_04063_),
    .Y(_04064_));
 sg13g2_buf_1 _13123_ (.A(_04064_),
    .X(_04065_));
 sg13g2_nor2_1 _13124_ (.A(_04022_),
    .B(_04055_),
    .Y(_04066_));
 sg13g2_nand2_1 _13125_ (.Y(_04067_),
    .A(_04065_),
    .B(_04066_));
 sg13g2_inv_1 _13126_ (.Y(_04068_),
    .A(_03985_));
 sg13g2_nand2_1 _13127_ (.Y(_04069_),
    .A(net37),
    .B(_04068_));
 sg13g2_nand3_1 _13128_ (.B(_03957_),
    .C(_03985_),
    .A(_03940_),
    .Y(_04070_));
 sg13g2_nand2_1 _13129_ (.Y(_04071_),
    .A(_04069_),
    .B(_04070_));
 sg13g2_xnor2_1 _13130_ (.Y(_04072_),
    .A(_03865_),
    .B(_03866_));
 sg13g2_buf_2 _13131_ (.A(_04072_),
    .X(_04073_));
 sg13g2_xnor2_1 _13132_ (.Y(_04074_),
    .A(_04073_),
    .B(net36));
 sg13g2_nor2_1 _13133_ (.A(_04071_),
    .B(_04074_),
    .Y(_04075_));
 sg13g2_nor2b_1 _13134_ (.A(_04067_),
    .B_N(_04075_),
    .Y(_04076_));
 sg13g2_xnor2_1 _13135_ (.Y(_04077_),
    .A(_03992_),
    .B(net37));
 sg13g2_nor2_1 _13136_ (.A(_04077_),
    .B(_04029_),
    .Y(_04078_));
 sg13g2_nand2_1 _13137_ (.Y(_04079_),
    .A(_04076_),
    .B(_04078_));
 sg13g2_xnor2_1 _13138_ (.Y(_04080_),
    .A(_03864_),
    .B(_03852_));
 sg13g2_nor3_1 _13139_ (.A(_04073_),
    .B(_04080_),
    .C(net36),
    .Y(_04081_));
 sg13g2_inv_1 _13140_ (.Y(_04082_),
    .A(_04080_));
 sg13g2_nand2_1 _13141_ (.Y(_04083_),
    .A(net36),
    .B(_04073_));
 sg13g2_nor2_1 _13142_ (.A(_04082_),
    .B(_04083_),
    .Y(_04084_));
 sg13g2_nor2_1 _13143_ (.A(_04081_),
    .B(_04084_),
    .Y(_04085_));
 sg13g2_xnor2_1 _13144_ (.Y(_04086_),
    .A(_04052_),
    .B(net36));
 sg13g2_nand2_1 _13145_ (.Y(_04087_),
    .A(_04049_),
    .B(_04086_));
 sg13g2_nor3_1 _13146_ (.A(_03984_),
    .B(_04085_),
    .C(_04087_),
    .Y(_04088_));
 sg13g2_nand2_1 _13147_ (.Y(_04089_),
    .A(_04088_),
    .B(_04031_));
 sg13g2_nand2_1 _13148_ (.Y(_04090_),
    .A(_04079_),
    .B(_04089_));
 sg13g2_buf_2 _13149_ (.A(_04090_),
    .X(_04091_));
 sg13g2_xor2_1 _13150_ (.B(net35),
    .A(\vgadonut.donut.donuthit.rx[15] ),
    .X(_04092_));
 sg13g2_inv_1 _13151_ (.Y(_04093_),
    .A(_04092_));
 sg13g2_buf_1 _13152_ (.A(_04093_),
    .X(_04094_));
 sg13g2_nand2_1 _13153_ (.Y(_04095_),
    .A(_04091_),
    .B(net25));
 sg13g2_nor2_1 _13154_ (.A(_04027_),
    .B(_04015_),
    .Y(_04096_));
 sg13g2_buf_1 _13155_ (.A(_04096_),
    .X(_04097_));
 sg13g2_buf_8 _13156_ (.A(_03961_),
    .X(_04098_));
 sg13g2_xnor2_1 _13157_ (.Y(_04099_),
    .A(\vgadonut.donut.donuthit.rx[8] ),
    .B(net33));
 sg13g2_nand2_1 _13158_ (.Y(_04100_),
    .A(net29),
    .B(_04099_));
 sg13g2_xnor2_1 _13159_ (.Y(_04101_),
    .A(\vgadonut.donut.donuthit.rx[7] ),
    .B(_04098_));
 sg13g2_nand2_1 _13160_ (.Y(_04102_),
    .A(net34),
    .B(_04101_));
 sg13g2_nand2_1 _13161_ (.Y(_04103_),
    .A(_04100_),
    .B(_04102_));
 sg13g2_xnor2_1 _13162_ (.Y(_04104_),
    .A(\vgadonut.donut.donuthit.rx[9] ),
    .B(_04098_));
 sg13g2_inv_1 _13163_ (.Y(_04105_),
    .A(_04104_));
 sg13g2_nand2_1 _13164_ (.Y(_04106_),
    .A(net30),
    .B(_04077_));
 sg13g2_buf_2 _13165_ (.A(_04106_),
    .X(_04107_));
 sg13g2_nor2_1 _13166_ (.A(_04105_),
    .B(_04107_),
    .Y(_04108_));
 sg13g2_nor2_1 _13167_ (.A(_04103_),
    .B(_04108_),
    .Y(_04109_));
 sg13g2_nand2_1 _13168_ (.Y(_04110_),
    .A(net30),
    .B(_03996_));
 sg13g2_buf_8 _13169_ (.A(_04110_),
    .X(_04111_));
 sg13g2_nor2_1 _13170_ (.A(_03986_),
    .B(_04111_),
    .Y(_04112_));
 sg13g2_buf_2 _13171_ (.A(_04112_),
    .X(_04113_));
 sg13g2_xnor2_1 _13172_ (.Y(_04114_),
    .A(\vgadonut.donut.donuthit.rx[10] ),
    .B(_03962_));
 sg13g2_buf_1 _13173_ (.A(_04114_),
    .X(_04115_));
 sg13g2_nand2_1 _13174_ (.Y(_04116_),
    .A(_04113_),
    .B(_04115_));
 sg13g2_nand2_1 _13175_ (.Y(_04117_),
    .A(_04109_),
    .B(_04116_));
 sg13g2_inv_1 _13176_ (.Y(_04118_),
    .A(_04117_));
 sg13g2_nand2_1 _13177_ (.Y(_04119_),
    .A(_04095_),
    .B(_04118_));
 sg13g2_nor2_1 _13178_ (.A(_04062_),
    .B(_04119_),
    .Y(_04120_));
 sg13g2_inv_1 _13179_ (.Y(_04121_),
    .A(_04115_));
 sg13g2_nor2_1 _13180_ (.A(_04121_),
    .B(_04044_),
    .Y(_04122_));
 sg13g2_nor2_1 _13181_ (.A(_04071_),
    .B(_04077_),
    .Y(_04123_));
 sg13g2_buf_8 _13182_ (.A(_04123_),
    .X(_04124_));
 sg13g2_nand2_1 _13183_ (.Y(_04125_),
    .A(net30),
    .B(_04124_));
 sg13g2_buf_8 _13184_ (.A(_04125_),
    .X(_04126_));
 sg13g2_nand3b_1 _13185_ (.B(_04012_),
    .C(_04082_),
    .Y(_04127_),
    .A_N(_04073_));
 sg13g2_nand3_1 _13186_ (.B(_04073_),
    .C(_04080_),
    .A(net36),
    .Y(_04128_));
 sg13g2_nand2_1 _13187_ (.Y(_04129_),
    .A(_04127_),
    .B(_04128_));
 sg13g2_nand3_1 _13188_ (.B(_04066_),
    .C(_04129_),
    .A(_04065_),
    .Y(_04130_));
 sg13g2_buf_2 _13189_ (.A(_04130_),
    .X(_04131_));
 sg13g2_nor3_1 _13190_ (.A(_04126_),
    .B(_04048_),
    .C(_04131_),
    .Y(_04132_));
 sg13g2_nor2_1 _13191_ (.A(_04122_),
    .B(_04132_),
    .Y(_04133_));
 sg13g2_inv_1 _13192_ (.Y(_04134_),
    .A(_04099_));
 sg13g2_nand2_1 _13193_ (.Y(_04135_),
    .A(_04078_),
    .B(_04071_));
 sg13g2_buf_1 _13194_ (.A(_04135_),
    .X(_04136_));
 sg13g2_nor2_1 _13195_ (.A(_04134_),
    .B(net24),
    .Y(_04137_));
 sg13g2_buf_1 _13196_ (.A(net29),
    .X(_04138_));
 sg13g2_buf_1 _13197_ (.A(net36),
    .X(_04139_));
 sg13g2_xnor2_1 _13198_ (.Y(_04140_),
    .A(\vgadonut.donut.donuthit.rx[6] ),
    .B(net32));
 sg13g2_nand2_1 _13199_ (.Y(_04141_),
    .A(_04008_),
    .B(\vgadonut.donut.donuthit.rx[5] ));
 sg13g2_nand2b_1 _13200_ (.Y(_04142_),
    .B(_04013_),
    .A_N(\vgadonut.donut.donuthit.rx[5] ));
 sg13g2_and2_1 _13201_ (.A(_04141_),
    .B(_04142_),
    .X(_04143_));
 sg13g2_a21oi_1 _13202_ (.A1(net23),
    .A2(_04140_),
    .Y(_04144_),
    .B1(_04143_));
 sg13g2_nor2_1 _13203_ (.A(_03996_),
    .B(_04029_),
    .Y(_04145_));
 sg13g2_buf_1 _13204_ (.A(_04145_),
    .X(_04146_));
 sg13g2_buf_1 _13205_ (.A(net28),
    .X(_04147_));
 sg13g2_nand2_1 _13206_ (.Y(_04148_),
    .A(_04147_),
    .B(_04101_));
 sg13g2_nand2_1 _13207_ (.Y(_04149_),
    .A(_04144_),
    .B(_04148_));
 sg13g2_nor2_1 _13208_ (.A(_04137_),
    .B(_04149_),
    .Y(_04150_));
 sg13g2_nand2_1 _13209_ (.Y(_04151_),
    .A(_04133_),
    .B(_04150_));
 sg13g2_nand2_1 _13210_ (.Y(_04152_),
    .A(net26),
    .B(_04033_));
 sg13g2_buf_2 _13211_ (.A(_04152_),
    .X(_04153_));
 sg13g2_nor2_1 _13212_ (.A(_04105_),
    .B(_04153_),
    .Y(_04154_));
 sg13g2_nand3_1 _13213_ (.B(_04075_),
    .C(_04066_),
    .A(_04065_),
    .Y(_04155_));
 sg13g2_buf_1 _13214_ (.A(_04155_),
    .X(_04156_));
 sg13g2_nor3_1 _13215_ (.A(_03965_),
    .B(_04111_),
    .C(_04156_),
    .Y(_04157_));
 sg13g2_nor2_1 _13216_ (.A(_04154_),
    .B(_04157_),
    .Y(_04158_));
 sg13g2_nor2_1 _13217_ (.A(_04040_),
    .B(_04059_),
    .Y(_04159_));
 sg13g2_inv_1 _13218_ (.Y(_04160_),
    .A(_04035_));
 sg13g2_nor2_1 _13219_ (.A(_04160_),
    .B(net18),
    .Y(_04161_));
 sg13g2_nor2_1 _13220_ (.A(_04159_),
    .B(_04161_),
    .Y(_04162_));
 sg13g2_nand2_1 _13221_ (.Y(_04163_),
    .A(_04158_),
    .B(_04162_));
 sg13g2_nor2_1 _13222_ (.A(_04151_),
    .B(_04163_),
    .Y(_04164_));
 sg13g2_nand2_1 _13223_ (.Y(_04165_),
    .A(_04120_),
    .B(_04164_));
 sg13g2_nor2_2 _13224_ (.A(_04126_),
    .B(_04131_),
    .Y(_04166_));
 sg13g2_nor2_1 _13225_ (.A(_04111_),
    .B(_04156_),
    .Y(_04167_));
 sg13g2_nor2_1 _13226_ (.A(_04166_),
    .B(_04167_),
    .Y(_04168_));
 sg13g2_inv_4 _13227_ (.A(_04059_),
    .Y(_04169_));
 sg13g2_nand2_1 _13228_ (.Y(_04170_),
    .A(_04065_),
    .B(_04124_));
 sg13g2_nor3_2 _13229_ (.A(_04029_),
    .B(_04049_),
    .C(_04170_),
    .Y(_04171_));
 sg13g2_nor2_1 _13230_ (.A(_04169_),
    .B(_04171_),
    .Y(_04172_));
 sg13g2_nor2_1 _13231_ (.A(_04029_),
    .B(_04170_),
    .Y(_04173_));
 sg13g2_nand3_1 _13232_ (.B(_04172_),
    .C(_04173_),
    .A(_04168_),
    .Y(_04174_));
 sg13g2_buf_2 _13233_ (.A(_04174_),
    .X(_04175_));
 sg13g2_buf_8 _13234_ (.A(_04175_),
    .X(_04176_));
 sg13g2_buf_8 _13235_ (.A(_04176_),
    .X(_04177_));
 sg13g2_buf_8 _13236_ (.A(_04177_),
    .X(_04178_));
 sg13g2_nand2_1 _13237_ (.Y(_04179_),
    .A(_04165_),
    .B(net10));
 sg13g2_a21oi_1 _13238_ (.A1(_04091_),
    .A2(net25),
    .Y(_04180_),
    .B1(_04117_));
 sg13g2_inv_1 _13239_ (.Y(_04181_),
    .A(_04060_));
 sg13g2_inv_1 _13240_ (.Y(_04182_),
    .A(_04045_));
 sg13g2_nand2_1 _13241_ (.Y(_04183_),
    .A(_04181_),
    .B(_04182_));
 sg13g2_o21ai_1 _13242_ (.B1(_04036_),
    .Y(_04184_),
    .A1(_03965_),
    .A2(net18));
 sg13g2_nor2_1 _13243_ (.A(_04183_),
    .B(_04184_),
    .Y(_04185_));
 sg13g2_nand2_1 _13244_ (.Y(_04186_),
    .A(_04180_),
    .B(_04185_));
 sg13g2_nand3b_1 _13245_ (.B(_04186_),
    .C(net10),
    .Y(_04187_),
    .A_N(_04164_));
 sg13g2_nand2b_1 _13246_ (.Y(_04188_),
    .B(_04187_),
    .A_N(_04179_));
 sg13g2_nand2b_1 _13247_ (.Y(_04189_),
    .B(_01959_),
    .A_N(_04188_));
 sg13g2_buf_1 _13248_ (.A(_09979_),
    .X(_04190_));
 sg13g2_buf_1 _13249_ (.A(net138),
    .X(_04191_));
 sg13g2_inv_1 _13250_ (.Y(_04192_),
    .A(_01959_));
 sg13g2_nand2_1 _13251_ (.Y(_04193_),
    .A(_04188_),
    .B(_04192_));
 sg13g2_nand3_1 _13252_ (.B(_04191_),
    .C(_04193_),
    .A(_04189_),
    .Y(_04194_));
 sg13g2_buf_1 _13253_ (.A(_09996_),
    .X(_04195_));
 sg13g2_inv_1 _13254_ (.Y(_04196_),
    .A(\vgadonut.donut.donuthit.rxin[5] ));
 sg13g2_buf_1 _13255_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[2] ),
    .X(_04197_));
 sg13g2_buf_1 _13256_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[4] ),
    .X(_04198_));
 sg13g2_nor2_1 _13257_ (.A(net252),
    .B(net251),
    .Y(_04199_));
 sg13g2_nand2_1 _13258_ (.Y(_04200_),
    .A(_04197_),
    .B(net251));
 sg13g2_nor2b_1 _13259_ (.A(_04199_),
    .B_N(_04200_),
    .Y(_04201_));
 sg13g2_buf_1 _13260_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[1] ),
    .X(_04202_));
 sg13g2_buf_1 _13261_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[3] ),
    .X(_04203_));
 sg13g2_nor2_1 _13262_ (.A(net250),
    .B(net249),
    .Y(_04204_));
 sg13g2_buf_2 _13263_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[0] ),
    .X(_04205_));
 sg13g2_buf_1 _13264_ (.A(\vgadonut.donut.sB[1] ),
    .X(_04206_));
 sg13g2_nand2_1 _13265_ (.Y(_04207_),
    .A(_04206_),
    .B(net250));
 sg13g2_buf_1 _13266_ (.A(\vgadonut.donut.sB[0] ),
    .X(_04208_));
 sg13g2_nand2_1 _13267_ (.Y(_04209_),
    .A(_04208_),
    .B(_04205_));
 sg13g2_nand2_1 _13268_ (.Y(_04210_),
    .A(_04207_),
    .B(_04209_));
 sg13g2_nor2_1 _13269_ (.A(_04205_),
    .B(net252),
    .Y(_04211_));
 sg13g2_nor2_1 _13270_ (.A(_04206_),
    .B(net250),
    .Y(_04212_));
 sg13g2_nor2_1 _13271_ (.A(_04211_),
    .B(_04212_),
    .Y(_04213_));
 sg13g2_a22oi_1 _13272_ (.Y(_04214_),
    .B1(_04210_),
    .B2(_04213_),
    .A2(net252),
    .A1(_04205_));
 sg13g2_nand2_1 _13273_ (.Y(_04215_),
    .A(net250),
    .B(net249));
 sg13g2_o21ai_1 _13274_ (.B1(_04215_),
    .Y(_04216_),
    .A1(_04204_),
    .A2(_04214_));
 sg13g2_xnor2_1 _13275_ (.Y(_04217_),
    .A(_04201_),
    .B(_04216_));
 sg13g2_nor2_1 _13276_ (.A(_04196_),
    .B(_04217_),
    .Y(_04218_));
 sg13g2_inv_1 _13277_ (.Y(_04219_),
    .A(_04218_));
 sg13g2_nand2_1 _13278_ (.Y(_04220_),
    .A(_04217_),
    .B(_04196_));
 sg13g2_nand3_1 _13279_ (.B(_04219_),
    .C(_04220_),
    .A(net112),
    .Y(_04221_));
 sg13g2_nand2_1 _13280_ (.Y(_00047_),
    .A(_04194_),
    .B(_04221_));
 sg13g2_buf_1 _13281_ (.A(\vgadonut.donut.donuthit.rxin[6] ),
    .X(_04222_));
 sg13g2_buf_1 _13282_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[5] ),
    .X(_04223_));
 sg13g2_nor2_1 _13283_ (.A(net249),
    .B(net248),
    .Y(_04224_));
 sg13g2_nand2_1 _13284_ (.Y(_04225_),
    .A(net249),
    .B(net248));
 sg13g2_nor2b_1 _13285_ (.A(_04224_),
    .B_N(_04225_),
    .Y(_04226_));
 sg13g2_inv_1 _13286_ (.Y(_04227_),
    .A(_04216_));
 sg13g2_a21oi_1 _13287_ (.A1(_04227_),
    .A2(_04200_),
    .Y(_04228_),
    .B1(_04199_));
 sg13g2_xnor2_1 _13288_ (.Y(_04229_),
    .A(_04226_),
    .B(_04228_));
 sg13g2_xnor2_1 _13289_ (.Y(_04230_),
    .A(_04222_),
    .B(_04229_));
 sg13g2_nor2b_1 _13290_ (.A(_04219_),
    .B_N(_04230_),
    .Y(_04231_));
 sg13g2_o21ai_1 _13291_ (.B1(net112),
    .Y(_04232_),
    .A1(_04218_),
    .A2(_04230_));
 sg13g2_a22oi_1 _13292_ (.Y(_04233_),
    .B1(_04104_),
    .B2(net29),
    .A2(_04099_),
    .A1(net34));
 sg13g2_nand2_1 _13293_ (.Y(_04234_),
    .A(net28),
    .B(_04115_));
 sg13g2_nand2_1 _13294_ (.Y(_04235_),
    .A(_04233_),
    .B(_04234_));
 sg13g2_nor2_1 _13295_ (.A(_04048_),
    .B(_04024_),
    .Y(_04236_));
 sg13g2_nor2_1 _13296_ (.A(_04235_),
    .B(_04236_),
    .Y(_04237_));
 sg13g2_nand2_1 _13297_ (.Y(_04238_),
    .A(_04095_),
    .B(_04237_));
 sg13g2_nand3_1 _13298_ (.B(_04057_),
    .C(_04093_),
    .A(_04031_),
    .Y(_04239_));
 sg13g2_nand4_1 _13299_ (.B(_04124_),
    .C(_04042_),
    .A(_04017_),
    .Y(_04240_),
    .D(_03964_));
 sg13g2_nand2_1 _13300_ (.Y(_04241_),
    .A(_04239_),
    .B(_04240_));
 sg13g2_nand2_1 _13301_ (.Y(_04242_),
    .A(_04113_),
    .B(_04035_));
 sg13g2_nand3_1 _13302_ (.B(_04033_),
    .C(_04039_),
    .A(net26),
    .Y(_04243_));
 sg13g2_nand2_1 _13303_ (.Y(_04244_),
    .A(_04242_),
    .B(_04243_));
 sg13g2_nor2_1 _13304_ (.A(_04241_),
    .B(_04244_),
    .Y(_04245_));
 sg13g2_nor2b_1 _13305_ (.A(_04238_),
    .B_N(_04245_),
    .Y(_04246_));
 sg13g2_nand2_1 _13306_ (.Y(_04247_),
    .A(net34),
    .B(_04140_));
 sg13g2_inv_1 _13307_ (.Y(_04248_),
    .A(_04247_));
 sg13g2_a21oi_1 _13308_ (.A1(net23),
    .A2(_04101_),
    .Y(_04249_),
    .B1(_04248_));
 sg13g2_nand2_1 _13309_ (.Y(_04250_),
    .A(net28),
    .B(_04099_));
 sg13g2_nand2_1 _13310_ (.Y(_04251_),
    .A(_04249_),
    .B(_04250_));
 sg13g2_nor2b_1 _13311_ (.A(net18),
    .B_N(_04039_),
    .Y(_04252_));
 sg13g2_nor2_1 _13312_ (.A(_04251_),
    .B(_04252_),
    .Y(_04253_));
 sg13g2_nor2_1 _13313_ (.A(_03965_),
    .B(_04059_),
    .Y(_04254_));
 sg13g2_nor2_1 _13314_ (.A(_04121_),
    .B(_04153_),
    .Y(_04255_));
 sg13g2_nor2_1 _13315_ (.A(_04254_),
    .B(_04255_),
    .Y(_04256_));
 sg13g2_nand2_1 _13316_ (.Y(_04257_),
    .A(_04253_),
    .B(_04256_));
 sg13g2_nor2_1 _13317_ (.A(_04160_),
    .B(_04044_),
    .Y(_04258_));
 sg13g2_nor3_1 _13318_ (.A(_04111_),
    .B(_04048_),
    .C(_04156_),
    .Y(_04259_));
 sg13g2_nor2_1 _13319_ (.A(_04258_),
    .B(_04259_),
    .Y(_04260_));
 sg13g2_nor2_1 _13320_ (.A(_04105_),
    .B(net24),
    .Y(_04261_));
 sg13g2_nor3_1 _13321_ (.A(_04126_),
    .B(_04092_),
    .C(_04131_),
    .Y(_04262_));
 sg13g2_nor2_1 _13322_ (.A(_04261_),
    .B(_04262_),
    .Y(_04263_));
 sg13g2_nand2_1 _13323_ (.Y(_04264_),
    .A(_04260_),
    .B(_04263_));
 sg13g2_nor2_1 _13324_ (.A(_04257_),
    .B(_04264_),
    .Y(_04265_));
 sg13g2_inv_2 _13325_ (.Y(_04266_),
    .A(net15));
 sg13g2_a21oi_1 _13326_ (.A1(_04246_),
    .A2(_04265_),
    .Y(_04267_),
    .B1(_04266_));
 sg13g2_nand3_1 _13327_ (.B(_04095_),
    .C(_04237_),
    .A(_04245_),
    .Y(_04268_));
 sg13g2_buf_1 _13328_ (.A(_04268_),
    .X(_04269_));
 sg13g2_nand2_1 _13329_ (.Y(_04270_),
    .A(_04166_),
    .B(_04094_));
 sg13g2_buf_8 _13330_ (.A(_04113_),
    .X(_04271_));
 sg13g2_nand2_1 _13331_ (.Y(_04272_),
    .A(net16),
    .B(_04104_));
 sg13g2_nand2_1 _13332_ (.Y(_04273_),
    .A(_04270_),
    .B(_04272_));
 sg13g2_nand2_1 _13333_ (.Y(_04274_),
    .A(_04167_),
    .B(_04047_));
 sg13g2_inv_1 _13334_ (.Y(_04275_),
    .A(_04258_));
 sg13g2_nand2_1 _13335_ (.Y(_04276_),
    .A(_04274_),
    .B(_04275_));
 sg13g2_nor2_1 _13336_ (.A(_04273_),
    .B(_04276_),
    .Y(_04277_));
 sg13g2_nand2_1 _13337_ (.Y(_04278_),
    .A(_04169_),
    .B(_03964_));
 sg13g2_nor2_1 _13338_ (.A(_03977_),
    .B(_04126_),
    .Y(_04279_));
 sg13g2_buf_2 _13339_ (.A(_04279_),
    .X(_04280_));
 sg13g2_nand2_1 _13340_ (.Y(_04281_),
    .A(_04280_),
    .B(_04115_));
 sg13g2_nand2_1 _13341_ (.Y(_04282_),
    .A(_04278_),
    .B(_04281_));
 sg13g2_nand2_1 _13342_ (.Y(_04283_),
    .A(_04171_),
    .B(_04039_));
 sg13g2_nand2_1 _13343_ (.Y(_04284_),
    .A(_04097_),
    .B(_04101_));
 sg13g2_nand2_1 _13344_ (.Y(_04285_),
    .A(_04284_),
    .B(_04247_));
 sg13g2_nor2_1 _13345_ (.A(_04134_),
    .B(_04107_),
    .Y(_04286_));
 sg13g2_nor2_1 _13346_ (.A(_04285_),
    .B(_04286_),
    .Y(_04287_));
 sg13g2_nand2_1 _13347_ (.Y(_04288_),
    .A(_04283_),
    .B(_04287_));
 sg13g2_nor2_1 _13348_ (.A(_04282_),
    .B(_04288_),
    .Y(_04289_));
 sg13g2_nand2_1 _13349_ (.Y(_04290_),
    .A(_04277_),
    .B(_04289_));
 sg13g2_buf_8 _13350_ (.A(_04175_),
    .X(_04291_));
 sg13g2_nand3_1 _13351_ (.B(_04290_),
    .C(net14),
    .A(_04269_),
    .Y(_04292_));
 sg13g2_buf_1 _13352_ (.A(_04292_),
    .X(_04293_));
 sg13g2_nand2_1 _13353_ (.Y(_04294_),
    .A(_04267_),
    .B(_04293_));
 sg13g2_inv_1 _13354_ (.Y(_04295_),
    .A(_01950_));
 sg13g2_nand2_1 _13355_ (.Y(_04296_),
    .A(_04294_),
    .B(_04295_));
 sg13g2_nand3_1 _13356_ (.B(_04293_),
    .C(_01950_),
    .A(_04267_),
    .Y(_04297_));
 sg13g2_nand2_1 _13357_ (.Y(_04298_),
    .A(_04296_),
    .B(_04297_));
 sg13g2_o21ai_1 _13358_ (.B1(_04187_),
    .Y(_04299_),
    .A1(_04192_),
    .A2(_04179_));
 sg13g2_nor2b_1 _13359_ (.A(_04298_),
    .B_N(_04299_),
    .Y(_04300_));
 sg13g2_inv_2 _13360_ (.Y(_04301_),
    .A(_04300_));
 sg13g2_nand2b_1 _13361_ (.Y(_04302_),
    .B(_04298_),
    .A_N(_04299_));
 sg13g2_buf_1 _13362_ (.A(net138),
    .X(_04303_));
 sg13g2_nand3_1 _13363_ (.B(_04302_),
    .C(_04303_),
    .A(_04301_),
    .Y(_04304_));
 sg13g2_o21ai_1 _13364_ (.B1(_04304_),
    .Y(_00054_),
    .A1(_04231_),
    .A2(_04232_));
 sg13g2_buf_8 _13365_ (.A(_09979_),
    .X(_04305_));
 sg13g2_buf_1 _13366_ (.A(net137),
    .X(_04306_));
 sg13g2_inv_1 _13367_ (.Y(_04307_),
    .A(_04222_));
 sg13g2_nor2_1 _13368_ (.A(_04307_),
    .B(_04229_),
    .Y(_04308_));
 sg13g2_nor2_1 _13369_ (.A(_04308_),
    .B(_04231_),
    .Y(_04309_));
 sg13g2_buf_1 _13370_ (.A(\vgadonut.donut.donuthit.rxin[7] ),
    .X(_04310_));
 sg13g2_buf_1 _13371_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[6] ),
    .X(_04311_));
 sg13g2_buf_1 _13372_ (.A(_04311_),
    .X(_04312_));
 sg13g2_nor2_1 _13373_ (.A(net251),
    .B(net213),
    .Y(_04313_));
 sg13g2_nand2_1 _13374_ (.Y(_04314_),
    .A(net251),
    .B(net213));
 sg13g2_inv_1 _13375_ (.Y(_04315_),
    .A(_04314_));
 sg13g2_nor2_1 _13376_ (.A(_04313_),
    .B(_04315_),
    .Y(_04316_));
 sg13g2_inv_1 _13377_ (.Y(_04317_),
    .A(_04228_));
 sg13g2_a21oi_1 _13378_ (.A1(_04317_),
    .A2(_04225_),
    .Y(_04318_),
    .B1(_04224_));
 sg13g2_xor2_1 _13379_ (.B(_04318_),
    .A(_04316_),
    .X(_04319_));
 sg13g2_nor2_1 _13380_ (.A(_04310_),
    .B(_04319_),
    .Y(_04320_));
 sg13g2_inv_1 _13381_ (.Y(_04321_),
    .A(_04310_));
 sg13g2_nor2b_1 _13382_ (.A(_04321_),
    .B_N(_04319_),
    .Y(_04322_));
 sg13g2_nor2_1 _13383_ (.A(_04320_),
    .B(_04322_),
    .Y(_04323_));
 sg13g2_xor2_1 _13384_ (.B(_04323_),
    .A(_04309_),
    .X(_04324_));
 sg13g2_buf_8 _13385_ (.A(net15),
    .X(_04325_));
 sg13g2_nand2_1 _13386_ (.Y(_04326_),
    .A(_04186_),
    .B(net12));
 sg13g2_nand2_1 _13387_ (.Y(_04327_),
    .A(_04168_),
    .B(_04172_));
 sg13g2_nand2_1 _13388_ (.Y(_04328_),
    .A(_04327_),
    .B(net25));
 sg13g2_buf_2 _13389_ (.A(_04328_),
    .X(_04329_));
 sg13g2_nand2_1 _13390_ (.Y(_04330_),
    .A(_04280_),
    .B(_03964_));
 sg13g2_nor2b_1 _13391_ (.A(_04126_),
    .B_N(_04042_),
    .Y(_04331_));
 sg13g2_buf_1 _13392_ (.A(_04331_),
    .X(_04332_));
 sg13g2_nand2_1 _13393_ (.Y(_04333_),
    .A(net17),
    .B(_04047_));
 sg13g2_nand2_1 _13394_ (.Y(_04334_),
    .A(_04330_),
    .B(_04333_));
 sg13g2_nor2_1 _13395_ (.A(_04160_),
    .B(_04107_),
    .Y(_04335_));
 sg13g2_nand2_2 _13396_ (.Y(_04336_),
    .A(_04026_),
    .B(_04001_));
 sg13g2_nand2_1 _13397_ (.Y(_04337_),
    .A(net34),
    .B(_04104_));
 sg13g2_o21ai_1 _13398_ (.B1(_04337_),
    .Y(_04338_),
    .A1(_04121_),
    .A2(_04336_));
 sg13g2_nor2_1 _13399_ (.A(_04335_),
    .B(_04338_),
    .Y(_04339_));
 sg13g2_nand2_1 _13400_ (.Y(_04340_),
    .A(_04113_),
    .B(_04039_));
 sg13g2_nand2_1 _13401_ (.Y(_04341_),
    .A(_04339_),
    .B(_04340_));
 sg13g2_nor2_1 _13402_ (.A(_04334_),
    .B(_04341_),
    .Y(_04342_));
 sg13g2_nand2_1 _13403_ (.Y(_04343_),
    .A(_04329_),
    .B(_04342_));
 sg13g2_nand2_1 _13404_ (.Y(_04344_),
    .A(_04343_),
    .B(net14));
 sg13g2_nand2_1 _13405_ (.Y(_04345_),
    .A(_04326_),
    .B(_04344_));
 sg13g2_nand3_1 _13406_ (.B(_04343_),
    .C(_04291_),
    .A(_04186_),
    .Y(_04346_));
 sg13g2_buf_1 _13407_ (.A(_04346_),
    .X(_04347_));
 sg13g2_nand2_1 _13408_ (.Y(_04348_),
    .A(_04345_),
    .B(_04347_));
 sg13g2_inv_1 _13409_ (.Y(_04349_),
    .A(net253));
 sg13g2_nand2_1 _13410_ (.Y(_04350_),
    .A(_04348_),
    .B(_04349_));
 sg13g2_nand3_1 _13411_ (.B(_04347_),
    .C(net253),
    .A(_04345_),
    .Y(_04351_));
 sg13g2_buf_1 _13412_ (.A(_04351_),
    .X(_04352_));
 sg13g2_nand2_1 _13413_ (.Y(_04353_),
    .A(_04246_),
    .B(_04265_));
 sg13g2_buf_8 _13414_ (.A(net14),
    .X(_04354_));
 sg13g2_nand2_1 _13415_ (.Y(_04355_),
    .A(_04353_),
    .B(_04354_));
 sg13g2_o21ai_1 _13416_ (.B1(_04293_),
    .Y(_04356_),
    .A1(_04295_),
    .A2(_04355_));
 sg13g2_a21oi_1 _13417_ (.A1(_04350_),
    .A2(_04352_),
    .Y(_04357_),
    .B1(_04356_));
 sg13g2_nand3_1 _13418_ (.B(_04350_),
    .C(_04352_),
    .A(_04356_),
    .Y(_04358_));
 sg13g2_buf_1 _13419_ (.A(_04358_),
    .X(_04359_));
 sg13g2_inv_1 _13420_ (.Y(_04360_),
    .A(_04359_));
 sg13g2_o21ai_1 _13421_ (.B1(_04301_),
    .Y(_04361_),
    .A1(_04357_),
    .A2(_04360_));
 sg13g2_buf_1 _13422_ (.A(net138),
    .X(_04362_));
 sg13g2_nand2_1 _13423_ (.Y(_04363_),
    .A(_04350_),
    .B(_04352_));
 sg13g2_inv_1 _13424_ (.Y(_04364_),
    .A(_04356_));
 sg13g2_nand2_1 _13425_ (.Y(_04365_),
    .A(_04363_),
    .B(_04364_));
 sg13g2_nand3_1 _13426_ (.B(_04300_),
    .C(_04365_),
    .A(_04359_),
    .Y(_04366_));
 sg13g2_nand3_1 _13427_ (.B(net123),
    .C(_04366_),
    .A(_04361_),
    .Y(_04367_));
 sg13g2_o21ai_1 _13428_ (.B1(_04367_),
    .Y(_00055_),
    .A1(net124),
    .A2(_04324_));
 sg13g2_nor2_1 _13429_ (.A(_04320_),
    .B(_04309_),
    .Y(_04368_));
 sg13g2_nor2_1 _13430_ (.A(_04322_),
    .B(_04368_),
    .Y(_04369_));
 sg13g2_buf_1 _13431_ (.A(\vgadonut.donut.donuthit.rxin[8] ),
    .X(_04370_));
 sg13g2_inv_1 _13432_ (.Y(_04371_),
    .A(_04370_));
 sg13g2_buf_1 _13433_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[7] ),
    .X(_04372_));
 sg13g2_buf_1 _13434_ (.A(_04372_),
    .X(_04373_));
 sg13g2_nor2_1 _13435_ (.A(net248),
    .B(net212),
    .Y(_04374_));
 sg13g2_nand2_1 _13436_ (.Y(_04375_),
    .A(net248),
    .B(net212));
 sg13g2_nor2b_1 _13437_ (.A(_04374_),
    .B_N(_04375_),
    .Y(_04376_));
 sg13g2_inv_1 _13438_ (.Y(_04377_),
    .A(_04313_));
 sg13g2_a21oi_1 _13439_ (.A1(_04318_),
    .A2(_04377_),
    .Y(_04378_),
    .B1(_04315_));
 sg13g2_xnor2_1 _13440_ (.Y(_04379_),
    .A(_04376_),
    .B(_04378_));
 sg13g2_inv_1 _13441_ (.Y(_04380_),
    .A(_04379_));
 sg13g2_nor2_1 _13442_ (.A(_04371_),
    .B(_04380_),
    .Y(_04381_));
 sg13g2_nand2_1 _13443_ (.Y(_04382_),
    .A(_04380_),
    .B(_04371_));
 sg13g2_nand2b_1 _13444_ (.Y(_04383_),
    .B(_04382_),
    .A_N(_04381_));
 sg13g2_xnor2_1 _13445_ (.Y(_04384_),
    .A(_04369_),
    .B(_04383_));
 sg13g2_o21ai_1 _13446_ (.B1(_04359_),
    .Y(_04385_),
    .A1(_04357_),
    .A2(_04301_));
 sg13g2_inv_1 _13447_ (.Y(_04386_),
    .A(_04385_));
 sg13g2_inv_1 _13448_ (.Y(_04387_),
    .A(_04347_));
 sg13g2_a21oi_2 _13449_ (.B1(_04387_),
    .Y(_04388_),
    .A2(_01956_),
    .A1(_04345_));
 sg13g2_a22oi_1 _13450_ (.Y(_04389_),
    .B1(_04280_),
    .B2(_04047_),
    .A2(_04094_),
    .A1(net17));
 sg13g2_nor2_1 _13451_ (.A(_03965_),
    .B(_04136_),
    .Y(_04390_));
 sg13g2_buf_8 _13452_ (.A(net34),
    .X(_04391_));
 sg13g2_a22oi_1 _13453_ (.Y(_04392_),
    .B1(_04035_),
    .B2(_04138_),
    .A2(_04115_),
    .A1(net31));
 sg13g2_nand2_1 _13454_ (.Y(_04393_),
    .A(_04146_),
    .B(_04039_));
 sg13g2_nand2_1 _13455_ (.Y(_04394_),
    .A(_04392_),
    .B(_04393_));
 sg13g2_nor2_1 _13456_ (.A(_04390_),
    .B(_04394_),
    .Y(_04395_));
 sg13g2_nand2_1 _13457_ (.Y(_04396_),
    .A(_04389_),
    .B(_04395_));
 sg13g2_inv_4 _13458_ (.A(_04329_),
    .Y(_04397_));
 sg13g2_a21oi_1 _13459_ (.A1(_04396_),
    .A2(_04291_),
    .Y(_04398_),
    .B1(_04397_));
 sg13g2_nand2_1 _13460_ (.Y(_04399_),
    .A(_04269_),
    .B(_04177_));
 sg13g2_nand2_1 _13461_ (.Y(_04400_),
    .A(_04398_),
    .B(_04399_));
 sg13g2_nand2_1 _13462_ (.Y(_04401_),
    .A(_04396_),
    .B(net15));
 sg13g2_nand2_1 _13463_ (.Y(_04402_),
    .A(_04401_),
    .B(_04329_));
 sg13g2_nand2_1 _13464_ (.Y(_04403_),
    .A(_04402_),
    .B(_04269_));
 sg13g2_nand2_1 _13465_ (.Y(_04404_),
    .A(_04400_),
    .B(_04403_));
 sg13g2_xnor2_1 _13466_ (.Y(_04405_),
    .A(_01974_),
    .B(_04404_));
 sg13g2_xnor2_1 _13467_ (.Y(_04406_),
    .A(_04388_),
    .B(_04405_));
 sg13g2_buf_1 _13468_ (.A(_09996_),
    .X(_04407_));
 sg13g2_a21oi_1 _13469_ (.A1(_04386_),
    .A2(_04406_),
    .Y(_04408_),
    .B1(net111));
 sg13g2_o21ai_1 _13470_ (.B1(_04408_),
    .Y(_04409_),
    .A1(_04386_),
    .A2(_04406_));
 sg13g2_o21ai_1 _13471_ (.B1(_04409_),
    .Y(_00056_),
    .A1(net124),
    .A2(_04384_));
 sg13g2_inv_1 _13472_ (.Y(_04410_),
    .A(_04369_));
 sg13g2_a21oi_1 _13473_ (.A1(_04410_),
    .A2(_04382_),
    .Y(_04411_),
    .B1(_04381_));
 sg13g2_buf_1 _13474_ (.A(\vgadonut.donut.donuthit.rxin[9] ),
    .X(_04412_));
 sg13g2_buf_1 _13475_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[8] ),
    .X(_04413_));
 sg13g2_buf_1 _13476_ (.A(_04413_),
    .X(_04414_));
 sg13g2_nor2_1 _13477_ (.A(net213),
    .B(net211),
    .Y(_04415_));
 sg13g2_nand2_1 _13478_ (.Y(_04416_),
    .A(net213),
    .B(net211));
 sg13g2_inv_1 _13479_ (.Y(_04417_),
    .A(_04416_));
 sg13g2_nor2_1 _13480_ (.A(_04415_),
    .B(_04417_),
    .Y(_04418_));
 sg13g2_o21ai_1 _13481_ (.B1(_04375_),
    .Y(_04419_),
    .A1(_04374_),
    .A2(_04378_));
 sg13g2_xor2_1 _13482_ (.B(_04419_),
    .A(_04418_),
    .X(_04420_));
 sg13g2_nor2_1 _13483_ (.A(_04412_),
    .B(_04420_),
    .Y(_04421_));
 sg13g2_inv_1 _13484_ (.Y(_04422_),
    .A(_04412_));
 sg13g2_nor2b_1 _13485_ (.A(_04422_),
    .B_N(_04420_),
    .Y(_04423_));
 sg13g2_nor2_1 _13486_ (.A(_04421_),
    .B(_04423_),
    .Y(_04424_));
 sg13g2_xor2_1 _13487_ (.B(_04424_),
    .A(_04411_),
    .X(_04425_));
 sg13g2_a22oi_1 _13488_ (.Y(_04426_),
    .B1(_01973_),
    .B2(_04400_),
    .A2(_04402_),
    .A1(_04269_));
 sg13g2_buf_1 _13489_ (.A(_04426_),
    .X(_04427_));
 sg13g2_nand2_1 _13490_ (.Y(_04428_),
    .A(_04391_),
    .B(_04035_));
 sg13g2_o21ai_1 _13491_ (.B1(_04428_),
    .Y(_04429_),
    .A1(_04040_),
    .A2(_04336_));
 sg13g2_a21oi_1 _13492_ (.A1(_03964_),
    .A2(_04147_),
    .Y(_04430_),
    .B1(_04429_));
 sg13g2_nor2_1 _13493_ (.A(_04065_),
    .B(_04126_),
    .Y(_04431_));
 sg13g2_nand2_1 _13494_ (.Y(_04432_),
    .A(_04431_),
    .B(_04093_));
 sg13g2_nand2_1 _13495_ (.Y(_04433_),
    .A(net16),
    .B(_04047_));
 sg13g2_nand3_1 _13496_ (.B(_04432_),
    .C(_04433_),
    .A(_04430_),
    .Y(_04434_));
 sg13g2_a21oi_1 _13497_ (.A1(_04434_),
    .A2(net15),
    .Y(_04435_),
    .B1(_04397_));
 sg13g2_nand2_1 _13498_ (.Y(_04436_),
    .A(_04435_),
    .B(_04344_));
 sg13g2_nand2_1 _13499_ (.Y(_04437_),
    .A(_04434_),
    .B(net15));
 sg13g2_nand2_1 _13500_ (.Y(_04438_),
    .A(_04437_),
    .B(_04329_));
 sg13g2_nand2_1 _13501_ (.Y(_04439_),
    .A(_04438_),
    .B(_04343_));
 sg13g2_nand2_1 _13502_ (.Y(_04440_),
    .A(_04436_),
    .B(_04439_));
 sg13g2_xnor2_1 _13503_ (.Y(_04441_),
    .A(_02046_),
    .B(_04440_));
 sg13g2_xnor2_1 _13504_ (.Y(_04442_),
    .A(_04427_),
    .B(_04441_));
 sg13g2_nor2_1 _13505_ (.A(_04388_),
    .B(_04405_),
    .Y(_04443_));
 sg13g2_nor2_1 _13506_ (.A(_04443_),
    .B(_04360_),
    .Y(_04444_));
 sg13g2_nand2_1 _13507_ (.Y(_04445_),
    .A(_04366_),
    .B(_04444_));
 sg13g2_nand2_1 _13508_ (.Y(_04446_),
    .A(_04405_),
    .B(_04388_));
 sg13g2_nand2_1 _13509_ (.Y(_04447_),
    .A(_04445_),
    .B(_04446_));
 sg13g2_a21oi_1 _13510_ (.A1(_04447_),
    .A2(_04442_),
    .Y(_04448_),
    .B1(net111));
 sg13g2_o21ai_1 _13511_ (.B1(_04448_),
    .Y(_04449_),
    .A1(_04442_),
    .A2(_04447_));
 sg13g2_o21ai_1 _13512_ (.B1(_04449_),
    .Y(_00057_),
    .A1(net124),
    .A2(_04425_));
 sg13g2_buf_1 _13513_ (.A(\vgadonut.donut.donuthit.rxin[10] ),
    .X(_04450_));
 sg13g2_inv_1 _13514_ (.Y(_04451_),
    .A(_04450_));
 sg13g2_buf_1 _13515_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[9] ),
    .X(_04452_));
 sg13g2_nor2_1 _13516_ (.A(_04373_),
    .B(net247),
    .Y(_04453_));
 sg13g2_nand2_1 _13517_ (.Y(_04454_),
    .A(_04373_),
    .B(net247));
 sg13g2_nand2b_1 _13518_ (.Y(_04455_),
    .B(_04454_),
    .A_N(_04453_));
 sg13g2_inv_1 _13519_ (.Y(_04456_),
    .A(_04415_));
 sg13g2_a21oi_1 _13520_ (.A1(_04419_),
    .A2(_04456_),
    .Y(_04457_),
    .B1(_04417_));
 sg13g2_xnor2_1 _13521_ (.Y(_04458_),
    .A(_04455_),
    .B(_04457_));
 sg13g2_nor2_1 _13522_ (.A(_04451_),
    .B(_04458_),
    .Y(_04459_));
 sg13g2_nand2_1 _13523_ (.Y(_04460_),
    .A(_04458_),
    .B(_04451_));
 sg13g2_inv_1 _13524_ (.Y(_04461_),
    .A(_04460_));
 sg13g2_nor2_1 _13525_ (.A(_04459_),
    .B(_04461_),
    .Y(_04462_));
 sg13g2_inv_1 _13526_ (.Y(_04463_),
    .A(_04462_));
 sg13g2_nor2_1 _13527_ (.A(_04421_),
    .B(_04411_),
    .Y(_04464_));
 sg13g2_nor2_1 _13528_ (.A(_04423_),
    .B(_04464_),
    .Y(_04465_));
 sg13g2_xnor2_1 _13529_ (.Y(_04466_),
    .A(_04463_),
    .B(_04465_));
 sg13g2_nor2_1 _13530_ (.A(_04442_),
    .B(_04406_),
    .Y(_04467_));
 sg13g2_nand2_1 _13531_ (.Y(_04468_),
    .A(_04385_),
    .B(_04467_));
 sg13g2_nand2_1 _13532_ (.Y(_04469_),
    .A(_04441_),
    .B(_04427_));
 sg13g2_nor2_1 _13533_ (.A(_04427_),
    .B(_04441_),
    .Y(_04470_));
 sg13g2_a21oi_1 _13534_ (.A1(_04443_),
    .A2(_04469_),
    .Y(_04471_),
    .B1(_04470_));
 sg13g2_nand2_1 _13535_ (.Y(_04472_),
    .A(_04468_),
    .B(_04471_));
 sg13g2_a22oi_1 _13536_ (.Y(_04473_),
    .B1(_01969_),
    .B2(_04436_),
    .A2(_04438_),
    .A1(_04343_));
 sg13g2_nor2_1 _13537_ (.A(_04092_),
    .B(_04136_),
    .Y(_04474_));
 sg13g2_nand2_1 _13538_ (.Y(_04475_),
    .A(net22),
    .B(_04047_));
 sg13g2_a22oi_1 _13539_ (.Y(_04476_),
    .B1(_03964_),
    .B2(net23),
    .A2(_04039_),
    .A1(net31));
 sg13g2_nand3_1 _13540_ (.B(_04475_),
    .C(_04476_),
    .A(_04432_),
    .Y(_04477_));
 sg13g2_nor2_1 _13541_ (.A(_04474_),
    .B(_04477_),
    .Y(_04478_));
 sg13g2_nand2_1 _13542_ (.Y(_04479_),
    .A(_04478_),
    .B(_04329_));
 sg13g2_nand2_1 _13543_ (.Y(_04480_),
    .A(_04479_),
    .B(net12));
 sg13g2_nand2_1 _13544_ (.Y(_04481_),
    .A(_04398_),
    .B(_04480_));
 sg13g2_nand2_1 _13545_ (.Y(_04482_),
    .A(_04402_),
    .B(_04479_));
 sg13g2_nand2_1 _13546_ (.Y(_04483_),
    .A(_04481_),
    .B(_04482_));
 sg13g2_xnor2_1 _13547_ (.Y(_04484_),
    .A(_01982_),
    .B(_04483_));
 sg13g2_nand2b_1 _13548_ (.Y(_04485_),
    .B(_04484_),
    .A_N(_04473_));
 sg13g2_xnor2_1 _13549_ (.Y(_04486_),
    .A(_02052_),
    .B(_04483_));
 sg13g2_nand2_1 _13550_ (.Y(_04487_),
    .A(_04486_),
    .B(_04473_));
 sg13g2_nand2_1 _13551_ (.Y(_04488_),
    .A(_04485_),
    .B(_04487_));
 sg13g2_inv_1 _13552_ (.Y(_04489_),
    .A(_04488_));
 sg13g2_nand2_1 _13553_ (.Y(_04490_),
    .A(_04472_),
    .B(_04489_));
 sg13g2_nand3_1 _13554_ (.B(_04471_),
    .C(_04488_),
    .A(_04468_),
    .Y(_04491_));
 sg13g2_nand3_1 _13555_ (.B(_04491_),
    .C(net125),
    .A(_04490_),
    .Y(_04492_));
 sg13g2_o21ai_1 _13556_ (.B1(_04492_),
    .Y(_00058_),
    .A1(_04306_),
    .A2(_04466_));
 sg13g2_buf_1 _13557_ (.A(\vgadonut.donut.donuthit.rxin[11] ),
    .X(_04493_));
 sg13g2_inv_1 _13558_ (.Y(_04494_),
    .A(_04493_));
 sg13g2_buf_1 _13559_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[10] ),
    .X(_04495_));
 sg13g2_buf_1 _13560_ (.A(_04495_),
    .X(_04496_));
 sg13g2_nor2_1 _13561_ (.A(_04414_),
    .B(net210),
    .Y(_04497_));
 sg13g2_nand2_1 _13562_ (.Y(_04498_),
    .A(_04414_),
    .B(net210));
 sg13g2_inv_1 _13563_ (.Y(_04499_),
    .A(_04498_));
 sg13g2_nor2_1 _13564_ (.A(_04497_),
    .B(_04499_),
    .Y(_04500_));
 sg13g2_o21ai_1 _13565_ (.B1(_04454_),
    .Y(_04501_),
    .A1(_04453_),
    .A2(_04457_));
 sg13g2_xnor2_1 _13566_ (.Y(_04502_),
    .A(_04500_),
    .B(_04501_));
 sg13g2_nor2_1 _13567_ (.A(_04494_),
    .B(_04502_),
    .Y(_04503_));
 sg13g2_nand2_1 _13568_ (.Y(_04504_),
    .A(_04502_),
    .B(_04494_));
 sg13g2_nand2b_1 _13569_ (.Y(_04505_),
    .B(_04504_),
    .A_N(_04503_));
 sg13g2_inv_1 _13570_ (.Y(_04506_),
    .A(_04459_));
 sg13g2_o21ai_1 _13571_ (.B1(_04506_),
    .Y(_04507_),
    .A1(_04461_),
    .A2(_04465_));
 sg13g2_xor2_1 _13572_ (.B(_04507_),
    .A(_04505_),
    .X(_04508_));
 sg13g2_nor2_1 _13573_ (.A(_04442_),
    .B(_04488_),
    .Y(_04509_));
 sg13g2_nand3_1 _13574_ (.B(_04446_),
    .C(_04509_),
    .A(_04445_),
    .Y(_04510_));
 sg13g2_nor2_1 _13575_ (.A(_04473_),
    .B(_04486_),
    .Y(_04511_));
 sg13g2_o21ai_1 _13576_ (.B1(_04487_),
    .Y(_04512_),
    .A1(_04470_),
    .A2(_04511_));
 sg13g2_nand2_1 _13577_ (.Y(_04513_),
    .A(_04510_),
    .B(_04512_));
 sg13g2_a22oi_1 _13578_ (.Y(_04514_),
    .B1(_01982_),
    .B2(_04481_),
    .A2(_04479_),
    .A1(_04402_));
 sg13g2_nand2_1 _13579_ (.Y(_04515_),
    .A(_04170_),
    .B(net30));
 sg13g2_nand3_1 _13580_ (.B(_04172_),
    .C(_04515_),
    .A(_04168_),
    .Y(_04516_));
 sg13g2_buf_1 _13581_ (.A(_04516_),
    .X(_04517_));
 sg13g2_nand2_1 _13582_ (.Y(_04518_),
    .A(_04517_),
    .B(net25));
 sg13g2_buf_1 _13583_ (.A(net31),
    .X(_04519_));
 sg13g2_buf_1 _13584_ (.A(net29),
    .X(_04520_));
 sg13g2_a22oi_1 _13585_ (.Y(_04521_),
    .B1(_04047_),
    .B2(net21),
    .A2(_03964_),
    .A1(net27));
 sg13g2_nand2_1 _13586_ (.Y(_04522_),
    .A(_04518_),
    .B(_04521_));
 sg13g2_nand2_1 _13587_ (.Y(_04523_),
    .A(_04522_),
    .B(net13));
 sg13g2_nand2_1 _13588_ (.Y(_04524_),
    .A(_04523_),
    .B(_04435_));
 sg13g2_nand2_1 _13589_ (.Y(_04525_),
    .A(_04438_),
    .B(_04522_));
 sg13g2_nand2_1 _13590_ (.Y(_04526_),
    .A(_04524_),
    .B(_04525_));
 sg13g2_xnor2_1 _13591_ (.Y(_04527_),
    .A(_01987_),
    .B(_04526_));
 sg13g2_xnor2_1 _13592_ (.Y(_04528_),
    .A(_04514_),
    .B(_04527_));
 sg13g2_a21oi_1 _13593_ (.A1(_04513_),
    .A2(_04528_),
    .Y(_04529_),
    .B1(net111));
 sg13g2_o21ai_1 _13594_ (.B1(_04529_),
    .Y(_04530_),
    .A1(_04513_),
    .A2(_04528_));
 sg13g2_o21ai_1 _13595_ (.B1(_04530_),
    .Y(_00059_),
    .A1(_04306_),
    .A2(_04508_));
 sg13g2_buf_1 _13596_ (.A(net137),
    .X(_04531_));
 sg13g2_buf_2 _13597_ (.A(\vgadonut.donut.donuthit.rxin[12] ),
    .X(_04532_));
 sg13g2_buf_1 _13598_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[11] ),
    .X(_04533_));
 sg13g2_buf_1 _13599_ (.A(_04533_),
    .X(_04534_));
 sg13g2_nor2_1 _13600_ (.A(_04452_),
    .B(net209),
    .Y(_04535_));
 sg13g2_nand2_1 _13601_ (.Y(_04536_),
    .A(_04452_),
    .B(net209));
 sg13g2_nor2b_1 _13602_ (.A(_04535_),
    .B_N(_04536_),
    .Y(_04537_));
 sg13g2_inv_1 _13603_ (.Y(_04538_),
    .A(_04497_));
 sg13g2_a21oi_1 _13604_ (.A1(_04501_),
    .A2(_04538_),
    .Y(_04539_),
    .B1(_04499_));
 sg13g2_xnor2_1 _13605_ (.Y(_04540_),
    .A(_04537_),
    .B(_04539_));
 sg13g2_nor2_1 _13606_ (.A(_04532_),
    .B(_04540_),
    .Y(_04541_));
 sg13g2_nand2_1 _13607_ (.Y(_04542_),
    .A(_04540_),
    .B(_04532_));
 sg13g2_nand2b_1 _13608_ (.Y(_04543_),
    .B(_04542_),
    .A_N(_04541_));
 sg13g2_a21oi_1 _13609_ (.A1(_04507_),
    .A2(_04504_),
    .Y(_04544_),
    .B1(_04503_));
 sg13g2_xnor2_1 _13610_ (.Y(_04545_),
    .A(_04543_),
    .B(_04544_));
 sg13g2_inv_1 _13611_ (.Y(_04546_),
    .A(_04471_));
 sg13g2_nand2b_1 _13612_ (.Y(_04547_),
    .B(_04527_),
    .A_N(_04514_));
 sg13g2_nor2b_1 _13613_ (.A(_04527_),
    .B_N(_04514_),
    .Y(_04548_));
 sg13g2_a21oi_1 _13614_ (.A1(_04547_),
    .A2(_04485_),
    .Y(_04549_),
    .B1(_04548_));
 sg13g2_nor2_1 _13615_ (.A(_04546_),
    .B(_04549_),
    .Y(_04550_));
 sg13g2_nand2_1 _13616_ (.Y(_04551_),
    .A(_04550_),
    .B(_04468_));
 sg13g2_inv_1 _13617_ (.Y(_04552_),
    .A(_04549_));
 sg13g2_nand2_1 _13618_ (.Y(_04553_),
    .A(_04528_),
    .B(_04489_));
 sg13g2_nand2_1 _13619_ (.Y(_04554_),
    .A(_04552_),
    .B(_04553_));
 sg13g2_a22oi_1 _13620_ (.Y(_04555_),
    .B1(_01987_),
    .B2(_04524_),
    .A2(_04522_),
    .A1(_04438_));
 sg13g2_a22oi_1 _13621_ (.Y(_04556_),
    .B1(net25),
    .B2(net21),
    .A2(_04047_),
    .A1(net27));
 sg13g2_nand2_1 _13622_ (.Y(_04557_),
    .A(_04518_),
    .B(_04556_));
 sg13g2_nand2_1 _13623_ (.Y(_04558_),
    .A(_04557_),
    .B(net13));
 sg13g2_nand2_1 _13624_ (.Y(_04559_),
    .A(_04558_),
    .B(_04480_));
 sg13g2_nand3_1 _13625_ (.B(_04354_),
    .C(_04479_),
    .A(_04557_),
    .Y(_04560_));
 sg13g2_nand2_1 _13626_ (.Y(_04561_),
    .A(_04559_),
    .B(_04560_));
 sg13g2_xnor2_1 _13627_ (.Y(_04562_),
    .A(_02070_),
    .B(_04561_));
 sg13g2_nor2_1 _13628_ (.A(_04555_),
    .B(_04562_),
    .Y(_04563_));
 sg13g2_inv_1 _13629_ (.Y(_04564_),
    .A(_04555_));
 sg13g2_xnor2_1 _13630_ (.Y(_04565_),
    .A(_01895_),
    .B(_04561_));
 sg13g2_nor2_1 _13631_ (.A(_04564_),
    .B(_04565_),
    .Y(_04566_));
 sg13g2_nor2_1 _13632_ (.A(_04563_),
    .B(_04566_),
    .Y(_04567_));
 sg13g2_a21oi_1 _13633_ (.A1(_04551_),
    .A2(_04554_),
    .Y(_04568_),
    .B1(_04567_));
 sg13g2_nand3_1 _13634_ (.B(_04567_),
    .C(_04554_),
    .A(_04551_),
    .Y(_04569_));
 sg13g2_nand3b_1 _13635_ (.B(net123),
    .C(_04569_),
    .Y(_04570_),
    .A_N(_04568_));
 sg13g2_o21ai_1 _13636_ (.B1(_04570_),
    .Y(_00060_),
    .A1(_04531_),
    .A2(_04545_));
 sg13g2_buf_1 _13637_ (.A(\vgadonut.donut.donuthit.rxin[13] ),
    .X(_04571_));
 sg13g2_inv_1 _13638_ (.Y(_04572_),
    .A(_04571_));
 sg13g2_buf_1 _13639_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[12] ),
    .X(_04573_));
 sg13g2_nor2_1 _13640_ (.A(net210),
    .B(net246),
    .Y(_04574_));
 sg13g2_nand2_1 _13641_ (.Y(_04575_),
    .A(net210),
    .B(net246));
 sg13g2_inv_1 _13642_ (.Y(_04576_),
    .A(_04575_));
 sg13g2_nor2_1 _13643_ (.A(_04574_),
    .B(_04576_),
    .Y(_04577_));
 sg13g2_o21ai_1 _13644_ (.B1(_04536_),
    .Y(_04578_),
    .A1(_04535_),
    .A2(_04539_));
 sg13g2_xnor2_1 _13645_ (.Y(_04579_),
    .A(_04577_),
    .B(_04578_));
 sg13g2_xnor2_1 _13646_ (.Y(_04580_),
    .A(_04572_),
    .B(_04579_));
 sg13g2_o21ai_1 _13647_ (.B1(_04542_),
    .Y(_04581_),
    .A1(_04541_),
    .A2(_04544_));
 sg13g2_xor2_1 _13648_ (.B(_04581_),
    .A(_04580_),
    .X(_04582_));
 sg13g2_nand2_1 _13649_ (.Y(_04583_),
    .A(_04565_),
    .B(_04564_));
 sg13g2_a21oi_1 _13650_ (.A1(_04547_),
    .A2(_04583_),
    .Y(_04584_),
    .B1(_04566_));
 sg13g2_nor2b_1 _13651_ (.A(_04584_),
    .B_N(_04512_),
    .Y(_04585_));
 sg13g2_nand2_1 _13652_ (.Y(_04586_),
    .A(_04510_),
    .B(_04585_));
 sg13g2_nand2_1 _13653_ (.Y(_04587_),
    .A(_04567_),
    .B(_04528_));
 sg13g2_nand2b_1 _13654_ (.Y(_04588_),
    .B(_04587_),
    .A_N(_04584_));
 sg13g2_inv_1 _13655_ (.Y(_04589_),
    .A(_04560_));
 sg13g2_a21oi_2 _13656_ (.B1(_04589_),
    .Y(_04590_),
    .A2(_01895_),
    .A1(_04559_));
 sg13g2_nand2_1 _13657_ (.Y(_04591_),
    .A(net12),
    .B(net25));
 sg13g2_buf_2 _13658_ (.A(_04591_),
    .X(_04592_));
 sg13g2_nand2_1 _13659_ (.Y(_04593_),
    .A(_04523_),
    .B(_04592_));
 sg13g2_nand3_1 _13660_ (.B(net25),
    .C(_04178_),
    .A(_04522_),
    .Y(_04594_));
 sg13g2_nand2_1 _13661_ (.Y(_04595_),
    .A(_04593_),
    .B(_04594_));
 sg13g2_xnor2_1 _13662_ (.Y(_04596_),
    .A(_02011_),
    .B(_04595_));
 sg13g2_xor2_1 _13663_ (.B(_04596_),
    .A(_04590_),
    .X(_04597_));
 sg13g2_a21oi_1 _13664_ (.A1(_04586_),
    .A2(_04588_),
    .Y(_04598_),
    .B1(_04597_));
 sg13g2_nand3_1 _13665_ (.B(_04597_),
    .C(_04588_),
    .A(_04586_),
    .Y(_04599_));
 sg13g2_nand3b_1 _13666_ (.B(_04362_),
    .C(_04599_),
    .Y(_04600_),
    .A_N(_04598_));
 sg13g2_o21ai_1 _13667_ (.B1(_04600_),
    .Y(_00061_),
    .A1(net122),
    .A2(_04582_));
 sg13g2_inv_1 _13668_ (.Y(_04601_),
    .A(\vgadonut.donut.donuthit.rxin[14] ));
 sg13g2_buf_1 _13669_ (.A(\vgadonut.donut.donuthit.cordicxy.x2in[13] ),
    .X(_04602_));
 sg13g2_buf_1 _13670_ (.A(_04602_),
    .X(_04603_));
 sg13g2_nor2_1 _13671_ (.A(net209),
    .B(net208),
    .Y(_04604_));
 sg13g2_nand2_1 _13672_ (.Y(_04605_),
    .A(_04534_),
    .B(net208));
 sg13g2_nor2b_1 _13673_ (.A(_04604_),
    .B_N(_04605_),
    .Y(_04606_));
 sg13g2_inv_1 _13674_ (.Y(_04607_),
    .A(_04574_));
 sg13g2_a21oi_1 _13675_ (.A1(_04578_),
    .A2(_04607_),
    .Y(_04608_),
    .B1(_04576_));
 sg13g2_xor2_1 _13676_ (.B(_04608_),
    .A(_04606_),
    .X(_04609_));
 sg13g2_xnor2_1 _13677_ (.Y(_04610_),
    .A(_04601_),
    .B(_04609_));
 sg13g2_inv_1 _13678_ (.Y(_04611_),
    .A(_04580_));
 sg13g2_nor2_1 _13679_ (.A(_04572_),
    .B(_04579_),
    .Y(_04612_));
 sg13g2_a21oi_1 _13680_ (.A1(_04611_),
    .A2(_04581_),
    .Y(_04613_),
    .B1(_04612_));
 sg13g2_nor2_1 _13681_ (.A(_04610_),
    .B(_04613_),
    .Y(_04614_));
 sg13g2_a21o_1 _13682_ (.A2(_04610_),
    .A1(_04613_),
    .B1(net137),
    .X(_04615_));
 sg13g2_nand2_1 _13683_ (.Y(_04616_),
    .A(_04597_),
    .B(_04567_));
 sg13g2_nor2_1 _13684_ (.A(_04553_),
    .B(_04616_),
    .Y(_04617_));
 sg13g2_nand2_1 _13685_ (.Y(_04618_),
    .A(_04472_),
    .B(_04617_));
 sg13g2_nor2_1 _13686_ (.A(_04590_),
    .B(_04596_),
    .Y(_04619_));
 sg13g2_nor2_1 _13687_ (.A(_04563_),
    .B(_04619_),
    .Y(_04620_));
 sg13g2_nand2_1 _13688_ (.Y(_04621_),
    .A(_04596_),
    .B(_04590_));
 sg13g2_nor2b_1 _13689_ (.A(_04620_),
    .B_N(_04621_),
    .Y(_04622_));
 sg13g2_nor2_1 _13690_ (.A(_04616_),
    .B(_04552_),
    .Y(_04623_));
 sg13g2_nor2_1 _13691_ (.A(_04622_),
    .B(_04623_),
    .Y(_04624_));
 sg13g2_nand2_1 _13692_ (.Y(_04625_),
    .A(_04618_),
    .B(_04624_));
 sg13g2_inv_1 _13693_ (.Y(_04626_),
    .A(_04594_));
 sg13g2_a21oi_2 _13694_ (.B1(_04626_),
    .Y(_04627_),
    .A2(_01891_),
    .A1(_04593_));
 sg13g2_nand2_1 _13695_ (.Y(_04628_),
    .A(_04558_),
    .B(_04592_));
 sg13g2_nand3_1 _13696_ (.B(net25),
    .C(_04178_),
    .A(_04557_),
    .Y(_04629_));
 sg13g2_nand2_1 _13697_ (.Y(_04630_),
    .A(_04628_),
    .B(_04629_));
 sg13g2_xor2_1 _13698_ (.B(_04630_),
    .A(_01902_),
    .X(_04631_));
 sg13g2_xor2_1 _13699_ (.B(_04631_),
    .A(_04627_),
    .X(_04632_));
 sg13g2_nand2_1 _13700_ (.Y(_04633_),
    .A(_04625_),
    .B(_04632_));
 sg13g2_xnor2_1 _13701_ (.Y(_04634_),
    .A(_04627_),
    .B(_04631_));
 sg13g2_nand3_1 _13702_ (.B(_04624_),
    .C(_04634_),
    .A(_04618_),
    .Y(_04635_));
 sg13g2_nand3_1 _13703_ (.B(_04635_),
    .C(net125),
    .A(_04633_),
    .Y(_04636_));
 sg13g2_o21ai_1 _13704_ (.B1(_04636_),
    .Y(_00062_),
    .A1(_04614_),
    .A2(_04615_));
 sg13g2_xnor2_1 _13705_ (.Y(_04637_),
    .A(_04590_),
    .B(_04596_));
 sg13g2_nor2_1 _13706_ (.A(_04637_),
    .B(_04634_),
    .Y(_04638_));
 sg13g2_nand2_1 _13707_ (.Y(_04639_),
    .A(_04638_),
    .B(_04584_));
 sg13g2_nor2_1 _13708_ (.A(_04627_),
    .B(_04631_),
    .Y(_04640_));
 sg13g2_nand2_1 _13709_ (.Y(_04641_),
    .A(_04631_),
    .B(_04627_));
 sg13g2_o21ai_1 _13710_ (.B1(_04641_),
    .Y(_04642_),
    .A1(_04619_),
    .A2(_04640_));
 sg13g2_nand2_1 _13711_ (.Y(_04643_),
    .A(_04639_),
    .B(_04642_));
 sg13g2_inv_1 _13712_ (.Y(_04644_),
    .A(_04638_));
 sg13g2_nor2_1 _13713_ (.A(_04587_),
    .B(_04644_),
    .Y(_04645_));
 sg13g2_nand2_1 _13714_ (.Y(_04646_),
    .A(_04513_),
    .B(_04645_));
 sg13g2_nand2b_1 _13715_ (.Y(_04647_),
    .B(_04646_),
    .A_N(_04643_));
 sg13g2_inv_1 _13716_ (.Y(_04648_),
    .A(_04629_));
 sg13g2_a21oi_1 _13717_ (.A1(_04628_),
    .A2(_01902_),
    .Y(_04649_),
    .B1(_04648_));
 sg13g2_nor2_1 _13718_ (.A(_01905_),
    .B(_04649_),
    .Y(_04650_));
 sg13g2_inv_2 _13719_ (.Y(_04651_),
    .A(_04650_));
 sg13g2_nand2_1 _13720_ (.Y(_04652_),
    .A(_04649_),
    .B(_01905_));
 sg13g2_nand2_1 _13721_ (.Y(_04653_),
    .A(_04651_),
    .B(_04652_));
 sg13g2_nand2b_1 _13722_ (.Y(_04654_),
    .B(_04653_),
    .A_N(_04647_));
 sg13g2_inv_1 _13723_ (.Y(_04655_),
    .A(_04653_));
 sg13g2_nand2_1 _13724_ (.Y(_04656_),
    .A(_04647_),
    .B(_04655_));
 sg13g2_nand3_1 _13725_ (.B(net126),
    .C(_04656_),
    .A(_04654_),
    .Y(_04657_));
 sg13g2_inv_1 _13726_ (.Y(_04658_),
    .A(_04614_));
 sg13g2_o21ai_1 _13727_ (.B1(_04658_),
    .Y(_04659_),
    .A1(_04601_),
    .A2(_04609_));
 sg13g2_buf_1 _13728_ (.A(\vgadonut.donut.donuthit.rxin[15] ),
    .X(_04660_));
 sg13g2_xor2_1 _13729_ (.B(net208),
    .A(_04573_),
    .X(_04661_));
 sg13g2_o21ai_1 _13730_ (.B1(_04605_),
    .Y(_04662_),
    .A1(_04604_),
    .A2(_04608_));
 sg13g2_xnor2_1 _13731_ (.Y(_04663_),
    .A(_04661_),
    .B(_04662_));
 sg13g2_xnor2_1 _13732_ (.Y(_04664_),
    .A(_04660_),
    .B(_04663_));
 sg13g2_a21oi_1 _13733_ (.A1(_04659_),
    .A2(_04664_),
    .Y(_04665_),
    .B1(net137));
 sg13g2_o21ai_1 _13734_ (.B1(_04665_),
    .Y(_04666_),
    .A1(_04659_),
    .A2(_04664_));
 sg13g2_nand2_1 _13735_ (.Y(_00048_),
    .A(_04657_),
    .B(_04666_));
 sg13g2_buf_1 _13736_ (.A(_09996_),
    .X(_04667_));
 sg13g2_xnor2_1 _13737_ (.Y(_04668_),
    .A(_02083_),
    .B(_04592_));
 sg13g2_inv_1 _13738_ (.Y(_04669_),
    .A(_04668_));
 sg13g2_nor2_1 _13739_ (.A(_04653_),
    .B(_04634_),
    .Y(_04670_));
 sg13g2_nand2_1 _13740_ (.Y(_04671_),
    .A(_04670_),
    .B(_04622_));
 sg13g2_o21ai_1 _13741_ (.B1(_04652_),
    .Y(_04672_),
    .A1(_04650_),
    .A2(_04640_));
 sg13g2_nand2_1 _13742_ (.Y(_04673_),
    .A(_04671_),
    .B(_04672_));
 sg13g2_nand2_1 _13743_ (.Y(_04674_),
    .A(_04632_),
    .B(_04655_));
 sg13g2_nor2_1 _13744_ (.A(_04616_),
    .B(_04674_),
    .Y(_04675_));
 sg13g2_nand3_1 _13745_ (.B(_04554_),
    .C(_04675_),
    .A(_04551_),
    .Y(_04676_));
 sg13g2_nand2b_1 _13746_ (.Y(_04677_),
    .B(_04676_),
    .A_N(_04673_));
 sg13g2_xnor2_1 _13747_ (.Y(_04678_),
    .A(_04669_),
    .B(_04677_));
 sg13g2_nand3b_1 _13748_ (.B(_04606_),
    .C(_04661_),
    .Y(_04679_),
    .A_N(_04608_));
 sg13g2_o21ai_1 _13749_ (.B1(net208),
    .Y(_04680_),
    .A1(_04534_),
    .A2(net246));
 sg13g2_nand2_1 _13750_ (.Y(_04681_),
    .A(_04679_),
    .B(_04680_));
 sg13g2_xnor2_1 _13751_ (.Y(_04682_),
    .A(_04660_),
    .B(_04681_));
 sg13g2_nand2_1 _13752_ (.Y(_04683_),
    .A(_04659_),
    .B(_04664_));
 sg13g2_o21ai_1 _13753_ (.B1(_04683_),
    .Y(_04684_),
    .A1(_00174_),
    .A2(_04663_));
 sg13g2_nor2_1 _13754_ (.A(_04682_),
    .B(_04684_),
    .Y(_04685_));
 sg13g2_and2_1 _13755_ (.A(_04684_),
    .B(_04682_),
    .X(_04686_));
 sg13g2_o21ai_1 _13756_ (.B1(net112),
    .Y(_04687_),
    .A1(_04685_),
    .A2(_04686_));
 sg13g2_o21ai_1 _13757_ (.B1(_04687_),
    .Y(_00049_),
    .A1(_04667_),
    .A2(_04678_));
 sg13g2_nor2_1 _13758_ (.A(_04668_),
    .B(_04653_),
    .Y(_04688_));
 sg13g2_inv_1 _13759_ (.Y(_04689_),
    .A(_04688_));
 sg13g2_nor2_1 _13760_ (.A(_04689_),
    .B(_04644_),
    .Y(_04690_));
 sg13g2_nand3_1 _13761_ (.B(_04588_),
    .C(_04690_),
    .A(_04586_),
    .Y(_04691_));
 sg13g2_inv_1 _13762_ (.Y(_04692_),
    .A(_04642_));
 sg13g2_nor2_1 _13763_ (.A(_04668_),
    .B(_04651_),
    .Y(_04693_));
 sg13g2_a21oi_1 _13764_ (.A1(_04692_),
    .A2(_04688_),
    .Y(_04694_),
    .B1(_04693_));
 sg13g2_nand2_1 _13765_ (.Y(_04695_),
    .A(_04691_),
    .B(_04694_));
 sg13g2_inv_1 _13766_ (.Y(_04696_),
    .A(_04592_));
 sg13g2_nand2_1 _13767_ (.Y(_04697_),
    .A(_04696_),
    .B(_02083_));
 sg13g2_xnor2_1 _13768_ (.Y(_04698_),
    .A(_02081_),
    .B(_04697_));
 sg13g2_inv_1 _13769_ (.Y(_04699_),
    .A(_04698_));
 sg13g2_nand2_1 _13770_ (.Y(_04700_),
    .A(_04695_),
    .B(_04699_));
 sg13g2_nand3_1 _13771_ (.B(_04694_),
    .C(_04698_),
    .A(_04691_),
    .Y(_04701_));
 sg13g2_nand3_1 _13772_ (.B(_04701_),
    .C(net126),
    .A(_04700_),
    .Y(_04702_));
 sg13g2_a21oi_1 _13773_ (.A1(_04679_),
    .A2(_04680_),
    .Y(_04703_),
    .B1(_00174_));
 sg13g2_inv_1 _13774_ (.Y(_04704_),
    .A(_04660_));
 sg13g2_a21oi_1 _13775_ (.A1(_04703_),
    .A2(_04704_),
    .Y(_04705_),
    .B1(_09979_));
 sg13g2_o21ai_1 _13776_ (.B1(_04705_),
    .Y(_04706_),
    .A1(_04703_),
    .A2(_04685_));
 sg13g2_buf_1 _13777_ (.A(_04706_),
    .X(_04707_));
 sg13g2_nand2_1 _13778_ (.Y(_00050_),
    .A(_04702_),
    .B(_04707_));
 sg13g2_nand2_1 _13779_ (.Y(_04708_),
    .A(_04699_),
    .B(_04669_));
 sg13g2_nor2_1 _13780_ (.A(_04708_),
    .B(_04674_),
    .Y(_04709_));
 sg13g2_nand2_1 _13781_ (.Y(_04710_),
    .A(_04625_),
    .B(_04709_));
 sg13g2_nand2_1 _13782_ (.Y(_04711_),
    .A(_04696_),
    .B(_02081_));
 sg13g2_nor2_1 _13783_ (.A(_02083_),
    .B(_04711_),
    .Y(_04712_));
 sg13g2_nor2_1 _13784_ (.A(_04708_),
    .B(_04672_),
    .Y(_04713_));
 sg13g2_nor2_1 _13785_ (.A(_04712_),
    .B(_04713_),
    .Y(_04714_));
 sg13g2_nand2_1 _13786_ (.Y(_04715_),
    .A(_04710_),
    .B(_04714_));
 sg13g2_inv_1 _13787_ (.Y(_04716_),
    .A(_00175_));
 sg13g2_nor2_1 _13788_ (.A(_01918_),
    .B(_04716_),
    .Y(_04717_));
 sg13g2_a22oi_1 _13789_ (.Y(_04718_),
    .B1(_04716_),
    .B2(_04711_),
    .A2(_04717_),
    .A1(_04696_));
 sg13g2_buf_1 _13790_ (.A(_04718_),
    .X(_04719_));
 sg13g2_inv_1 _13791_ (.Y(_04720_),
    .A(_04719_));
 sg13g2_nand2_1 _13792_ (.Y(_04721_),
    .A(_04715_),
    .B(_04720_));
 sg13g2_nand3_1 _13793_ (.B(_04714_),
    .C(_04719_),
    .A(_04710_),
    .Y(_04722_));
 sg13g2_nand3_1 _13794_ (.B(_04722_),
    .C(net126),
    .A(_04721_),
    .Y(_04723_));
 sg13g2_nand2_1 _13795_ (.Y(_00051_),
    .A(_04723_),
    .B(_04707_));
 sg13g2_nand2_1 _13796_ (.Y(_04724_),
    .A(_04720_),
    .B(_04699_));
 sg13g2_nor2_1 _13797_ (.A(_04724_),
    .B(_04689_),
    .Y(_04725_));
 sg13g2_nand3_1 _13798_ (.B(_04645_),
    .C(_04725_),
    .A(_04513_),
    .Y(_04726_));
 sg13g2_inv_1 _13799_ (.Y(_04727_),
    .A(_04693_));
 sg13g2_nor2_1 _13800_ (.A(_04716_),
    .B(_04592_),
    .Y(_04728_));
 sg13g2_o21ai_1 _13801_ (.B1(_04728_),
    .Y(_04729_),
    .A1(_01918_),
    .A2(_01922_));
 sg13g2_o21ai_1 _13802_ (.B1(_04729_),
    .Y(_04730_),
    .A1(_04724_),
    .A2(_04727_));
 sg13g2_a21oi_1 _13803_ (.A1(_04643_),
    .A2(_04725_),
    .Y(_04731_),
    .B1(_04730_));
 sg13g2_nand2_1 _13804_ (.Y(_04732_),
    .A(_04726_),
    .B(_04731_));
 sg13g2_inv_1 _13805_ (.Y(_04733_),
    .A(_00176_));
 sg13g2_nor2_1 _13806_ (.A(_04733_),
    .B(_04592_),
    .Y(_04734_));
 sg13g2_inv_1 _13807_ (.Y(_04735_),
    .A(_04728_));
 sg13g2_a22oi_1 _13808_ (.Y(_04736_),
    .B1(_04733_),
    .B2(_04735_),
    .A2(_00175_),
    .A1(_04734_));
 sg13g2_nand2_1 _13809_ (.Y(_04737_),
    .A(_04732_),
    .B(_04736_));
 sg13g2_inv_1 _13810_ (.Y(_04738_),
    .A(_04736_));
 sg13g2_nand3_1 _13811_ (.B(_04731_),
    .C(_04738_),
    .A(_04726_),
    .Y(_04739_));
 sg13g2_nand2_1 _13812_ (.Y(_04740_),
    .A(_04737_),
    .B(_04739_));
 sg13g2_buf_8 _13813_ (.A(net137),
    .X(_04741_));
 sg13g2_nand2_1 _13814_ (.Y(_04742_),
    .A(_04740_),
    .B(_04741_));
 sg13g2_nand2_1 _13815_ (.Y(_00052_),
    .A(_04742_),
    .B(_04707_));
 sg13g2_nor3_1 _13816_ (.A(_04719_),
    .B(_04736_),
    .C(_04708_),
    .Y(_04743_));
 sg13g2_nand4_1 _13817_ (.B(_04554_),
    .C(_04675_),
    .A(_04551_),
    .Y(_04744_),
    .D(_04743_));
 sg13g2_inv_1 _13818_ (.Y(_04745_),
    .A(_04734_));
 sg13g2_nand3_1 _13819_ (.B(_04720_),
    .C(_04712_),
    .A(_04738_),
    .Y(_04746_));
 sg13g2_o21ai_1 _13820_ (.B1(_04746_),
    .Y(_04747_),
    .A1(_04717_),
    .A2(_04745_));
 sg13g2_a21oi_1 _13821_ (.A1(_04673_),
    .A2(_04743_),
    .Y(_04748_),
    .B1(_04747_));
 sg13g2_nand2_1 _13822_ (.Y(_04749_),
    .A(_04744_),
    .B(_04748_));
 sg13g2_xor2_1 _13823_ (.B(_04734_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[15] ),
    .X(_04750_));
 sg13g2_nand2_1 _13824_ (.Y(_04751_),
    .A(_04749_),
    .B(_04750_));
 sg13g2_inv_1 _13825_ (.Y(_04752_),
    .A(_04750_));
 sg13g2_nand3_1 _13826_ (.B(_04748_),
    .C(_04752_),
    .A(_04744_),
    .Y(_04753_));
 sg13g2_nand3_1 _13827_ (.B(_04753_),
    .C(net126),
    .A(_04751_),
    .Y(_04754_));
 sg13g2_nand2_1 _13828_ (.Y(_00053_),
    .A(_04754_),
    .B(_04707_));
 sg13g2_xor2_1 _13829_ (.B(net33),
    .A(\vgadonut.donut.donuthit.ry[15] ),
    .X(_04755_));
 sg13g2_inv_1 _13830_ (.Y(_04756_),
    .A(_04755_));
 sg13g2_buf_1 _13831_ (.A(_04756_),
    .X(_04757_));
 sg13g2_xnor2_1 _13832_ (.Y(_04758_),
    .A(\vgadonut.donut.donuthit.ry[8] ),
    .B(net33));
 sg13g2_nand2_1 _13833_ (.Y(_04759_),
    .A(net29),
    .B(_04758_));
 sg13g2_xnor2_1 _13834_ (.Y(_04760_),
    .A(\vgadonut.donut.donuthit.ry[7] ),
    .B(net32));
 sg13g2_nand2_1 _13835_ (.Y(_04761_),
    .A(net34),
    .B(_04760_));
 sg13g2_nand2_1 _13836_ (.Y(_04762_),
    .A(_04759_),
    .B(_04761_));
 sg13g2_xor2_1 _13837_ (.B(net33),
    .A(\vgadonut.donut.donuthit.ry[9] ),
    .X(_04763_));
 sg13g2_nor2_1 _13838_ (.A(_04763_),
    .B(_04107_),
    .Y(_04764_));
 sg13g2_nor2_1 _13839_ (.A(_04762_),
    .B(_04764_),
    .Y(_04765_));
 sg13g2_xnor2_1 _13840_ (.Y(_04766_),
    .A(\vgadonut.donut.donuthit.ry[10] ),
    .B(net32));
 sg13g2_buf_1 _13841_ (.A(_04766_),
    .X(_04767_));
 sg13g2_nand2_1 _13842_ (.Y(_04768_),
    .A(net16),
    .B(_04767_));
 sg13g2_nand2_1 _13843_ (.Y(_04769_),
    .A(_04765_),
    .B(_04768_));
 sg13g2_a21oi_1 _13844_ (.A1(_04091_),
    .A2(net20),
    .Y(_04770_),
    .B1(_04769_));
 sg13g2_xor2_1 _13845_ (.B(net32),
    .A(\vgadonut.donut.donuthit.ry[14] ),
    .X(_04771_));
 sg13g2_buf_2 _13846_ (.A(_04771_),
    .X(_04772_));
 sg13g2_inv_1 _13847_ (.Y(_04773_),
    .A(_04772_));
 sg13g2_nand2_1 _13848_ (.Y(_04774_),
    .A(_04169_),
    .B(_04773_));
 sg13g2_xnor2_1 _13849_ (.Y(_04775_),
    .A(\vgadonut.donut.donuthit.ry[12] ),
    .B(net32));
 sg13g2_buf_2 _13850_ (.A(_04775_),
    .X(_04776_));
 sg13g2_nand2_1 _13851_ (.Y(_04777_),
    .A(net17),
    .B(_04776_));
 sg13g2_nand2_1 _13852_ (.Y(_04778_),
    .A(_04774_),
    .B(_04777_));
 sg13g2_xor2_1 _13853_ (.B(net35),
    .A(\vgadonut.donut.donuthit.ry[13] ),
    .X(_04779_));
 sg13g2_inv_2 _13854_ (.Y(_04780_),
    .A(_04779_));
 sg13g2_nand2_1 _13855_ (.Y(_04781_),
    .A(_04171_),
    .B(_04780_));
 sg13g2_xor2_1 _13856_ (.B(net33),
    .A(\vgadonut.donut.donuthit.ry[11] ),
    .X(_04782_));
 sg13g2_inv_2 _13857_ (.Y(_04783_),
    .A(_04782_));
 sg13g2_nand2_1 _13858_ (.Y(_04784_),
    .A(_04280_),
    .B(_04783_));
 sg13g2_nand2_1 _13859_ (.Y(_04785_),
    .A(_04781_),
    .B(_04784_));
 sg13g2_nor2_1 _13860_ (.A(_04778_),
    .B(_04785_),
    .Y(_04786_));
 sg13g2_nand2_1 _13861_ (.Y(_04787_),
    .A(_04770_),
    .B(_04786_));
 sg13g2_nand2_1 _13862_ (.Y(_04788_),
    .A(_04787_),
    .B(net14));
 sg13g2_inv_1 _13863_ (.Y(_04789_),
    .A(_04763_));
 sg13g2_nand2_1 _13864_ (.Y(_04790_),
    .A(_04280_),
    .B(_04789_));
 sg13g2_o21ai_1 _13865_ (.B1(_04790_),
    .Y(_04791_),
    .A1(_04779_),
    .A2(_04079_));
 sg13g2_xnor2_1 _13866_ (.Y(_04792_),
    .A(\vgadonut.donut.donuthit.ry[6] ),
    .B(net32));
 sg13g2_inv_1 _13867_ (.Y(_04793_),
    .A(_04792_));
 sg13g2_inv_1 _13868_ (.Y(_04794_),
    .A(_04013_));
 sg13g2_nand2_1 _13869_ (.Y(_04795_),
    .A(_04008_),
    .B(\vgadonut.donut.donuthit.ry[5] ));
 sg13g2_o21ai_1 _13870_ (.B1(_04795_),
    .Y(_04796_),
    .A1(\vgadonut.donut.donuthit.ry[5] ),
    .A2(_04794_));
 sg13g2_o21ai_1 _13871_ (.B1(_04796_),
    .Y(_04797_),
    .A1(_04793_),
    .A2(_04336_));
 sg13g2_a21oi_1 _13872_ (.A1(net22),
    .A2(_04760_),
    .Y(_04798_),
    .B1(_04797_));
 sg13g2_nand2_1 _13873_ (.Y(_04799_),
    .A(net17),
    .B(_04767_));
 sg13g2_nand2_1 _13874_ (.Y(_04800_),
    .A(_04798_),
    .B(_04799_));
 sg13g2_nor2_1 _13875_ (.A(_04791_),
    .B(_04800_),
    .Y(_04801_));
 sg13g2_nand2_1 _13876_ (.Y(_04802_),
    .A(net16),
    .B(_04758_));
 sg13g2_o21ai_1 _13877_ (.B1(_04802_),
    .Y(_04803_),
    .A1(_04782_),
    .A2(net18));
 sg13g2_nand2_1 _13878_ (.Y(_04804_),
    .A(_04169_),
    .B(_04776_));
 sg13g2_o21ai_1 _13879_ (.B1(_04804_),
    .Y(_04805_),
    .A1(_04772_),
    .A2(_04089_));
 sg13g2_nor2_1 _13880_ (.A(_04803_),
    .B(_04805_),
    .Y(_04806_));
 sg13g2_nand2_1 _13881_ (.Y(_04807_),
    .A(_04801_),
    .B(_04806_));
 sg13g2_nor2b_1 _13882_ (.A(_04788_),
    .B_N(_04807_),
    .Y(_04808_));
 sg13g2_nor2_1 _13883_ (.A(_04787_),
    .B(_04807_),
    .Y(_04809_));
 sg13g2_nor2_1 _13884_ (.A(_04266_),
    .B(_04809_),
    .Y(_04810_));
 sg13g2_nand2b_1 _13885_ (.Y(_04811_),
    .B(_04810_),
    .A_N(_04808_));
 sg13g2_nand2b_1 _13886_ (.Y(_04812_),
    .B(_01958_),
    .A_N(_04811_));
 sg13g2_nand2_1 _13887_ (.Y(_04813_),
    .A(_04811_),
    .B(_02029_));
 sg13g2_nand3_1 _13888_ (.B(net126),
    .C(_04813_),
    .A(_04812_),
    .Y(_04814_));
 sg13g2_buf_2 _13889_ (.A(\vgadonut.donut.sAcB[4] ),
    .X(_04815_));
 sg13g2_buf_1 _13890_ (.A(\vgadonut.donut.sAcB[6] ),
    .X(_04816_));
 sg13g2_nor2_1 _13891_ (.A(_04815_),
    .B(net244),
    .Y(_04817_));
 sg13g2_nand2_1 _13892_ (.Y(_04818_),
    .A(_04815_),
    .B(net244));
 sg13g2_nor2b_1 _13893_ (.A(_04817_),
    .B_N(_04818_),
    .Y(_04819_));
 sg13g2_buf_2 _13894_ (.A(\vgadonut.donut.sAcB[3] ),
    .X(_04820_));
 sg13g2_buf_1 _13895_ (.A(\vgadonut.donut.sAcB[5] ),
    .X(_04821_));
 sg13g2_nor2_1 _13896_ (.A(_04820_),
    .B(_04821_),
    .Y(_04822_));
 sg13g2_buf_2 _13897_ (.A(\vgadonut.donut.sAcB[2] ),
    .X(_04823_));
 sg13g2_buf_2 _13898_ (.A(\vgadonut.donut.sAcB[1] ),
    .X(_04824_));
 sg13g2_nand2_1 _13899_ (.Y(_04825_),
    .A(_04824_),
    .B(_04820_));
 sg13g2_buf_2 _13900_ (.A(\vgadonut.donut.sAcB[0] ),
    .X(_04826_));
 sg13g2_nand2_1 _13901_ (.Y(_04827_),
    .A(_04826_),
    .B(_04823_));
 sg13g2_nand2_1 _13902_ (.Y(_04828_),
    .A(_04825_),
    .B(_04827_));
 sg13g2_nor2_1 _13903_ (.A(_04823_),
    .B(_04815_),
    .Y(_04829_));
 sg13g2_nor2_1 _13904_ (.A(_04824_),
    .B(_04820_),
    .Y(_04830_));
 sg13g2_nor2_1 _13905_ (.A(_04829_),
    .B(_04830_),
    .Y(_04831_));
 sg13g2_a22oi_1 _13906_ (.Y(_04832_),
    .B1(_04828_),
    .B2(_04831_),
    .A2(_04815_),
    .A1(_04823_));
 sg13g2_nand2_1 _13907_ (.Y(_04833_),
    .A(_04820_),
    .B(_04821_));
 sg13g2_o21ai_1 _13908_ (.B1(_04833_),
    .Y(_04834_),
    .A1(_04822_),
    .A2(_04832_));
 sg13g2_xnor2_1 _13909_ (.Y(_04835_),
    .A(_04819_),
    .B(_04834_));
 sg13g2_nor2b_1 _13910_ (.A(_04835_),
    .B_N(_00123_),
    .Y(_04836_));
 sg13g2_nor2b_1 _13911_ (.A(_00123_),
    .B_N(_04835_),
    .Y(_04837_));
 sg13g2_o21ai_1 _13912_ (.B1(_04195_),
    .Y(_04838_),
    .A1(_04836_),
    .A2(_04837_));
 sg13g2_nand2_1 _13913_ (.Y(_00063_),
    .A(_04814_),
    .B(_04838_));
 sg13g2_inv_1 _13914_ (.Y(_04839_),
    .A(\vgadonut.donut.donuthit.ryin[5] ));
 sg13g2_nor2_1 _13915_ (.A(_04839_),
    .B(_04835_),
    .Y(_04840_));
 sg13g2_inv_1 _13916_ (.Y(_04841_),
    .A(_04840_));
 sg13g2_buf_1 _13917_ (.A(\vgadonut.donut.sAcB[7] ),
    .X(_04842_));
 sg13g2_nor2_1 _13918_ (.A(net243),
    .B(net242),
    .Y(_04843_));
 sg13g2_nand2_1 _13919_ (.Y(_04844_),
    .A(net243),
    .B(net242));
 sg13g2_nor2b_1 _13920_ (.A(_04843_),
    .B_N(_04844_),
    .Y(_04845_));
 sg13g2_inv_1 _13921_ (.Y(_04846_),
    .A(_04834_));
 sg13g2_a21oi_1 _13922_ (.A1(_04846_),
    .A2(_04818_),
    .Y(_04847_),
    .B1(_04817_));
 sg13g2_xnor2_1 _13923_ (.Y(_04848_),
    .A(_04845_),
    .B(_04847_));
 sg13g2_xnor2_1 _13924_ (.Y(_04849_),
    .A(\vgadonut.donut.donuthit.ryin[6] ),
    .B(_04848_));
 sg13g2_inv_1 _13925_ (.Y(_04850_),
    .A(_04849_));
 sg13g2_nor2_1 _13926_ (.A(_04841_),
    .B(_04850_),
    .Y(_04851_));
 sg13g2_o21ai_1 _13927_ (.B1(_04195_),
    .Y(_04852_),
    .A1(_04840_),
    .A2(_04849_));
 sg13g2_nand2_1 _13928_ (.Y(_04853_),
    .A(_04091_),
    .B(net20));
 sg13g2_a22oi_1 _13929_ (.Y(_04854_),
    .B1(_04789_),
    .B2(net23),
    .A2(_04758_),
    .A1(net31));
 sg13g2_nand2_1 _13930_ (.Y(_04855_),
    .A(net28),
    .B(_04767_));
 sg13g2_nand2_1 _13931_ (.Y(_04856_),
    .A(_04854_),
    .B(_04855_));
 sg13g2_nor2_1 _13932_ (.A(_04772_),
    .B(net18),
    .Y(_04857_));
 sg13g2_nor2_1 _13933_ (.A(_04856_),
    .B(_04857_),
    .Y(_04858_));
 sg13g2_nand2_1 _13934_ (.Y(_04859_),
    .A(_04853_),
    .B(_04858_));
 sg13g2_nand3_1 _13935_ (.B(_04057_),
    .C(_04756_),
    .A(net26),
    .Y(_04860_));
 sg13g2_nand4_1 _13936_ (.B(_04124_),
    .C(_04042_),
    .A(net30),
    .Y(_04861_),
    .D(_04780_));
 sg13g2_nand2_1 _13937_ (.Y(_04862_),
    .A(_04860_),
    .B(_04861_));
 sg13g2_nand3_1 _13938_ (.B(_04071_),
    .C(_04783_),
    .A(_04078_),
    .Y(_04863_));
 sg13g2_nand3_1 _13939_ (.B(_04033_),
    .C(_04776_),
    .A(net26),
    .Y(_04864_));
 sg13g2_nand2_1 _13940_ (.Y(_04865_),
    .A(_04863_),
    .B(_04864_));
 sg13g2_nor2_1 _13941_ (.A(_04862_),
    .B(_04865_),
    .Y(_04866_));
 sg13g2_nor2b_1 _13942_ (.A(_04859_),
    .B_N(_04866_),
    .Y(_04867_));
 sg13g2_nor2b_1 _13943_ (.A(net18),
    .B_N(_04776_),
    .Y(_04868_));
 sg13g2_nand4_1 _13944_ (.B(_04124_),
    .C(_04042_),
    .A(net30),
    .Y(_04869_),
    .D(_04783_));
 sg13g2_nor2b_1 _13945_ (.A(_04868_),
    .B_N(_04869_),
    .Y(_04870_));
 sg13g2_nor2_1 _13946_ (.A(_04763_),
    .B(net24),
    .Y(_04871_));
 sg13g2_nor2_1 _13947_ (.A(_04793_),
    .B(_04026_),
    .Y(_04872_));
 sg13g2_a21oi_1 _13948_ (.A1(net23),
    .A2(_04760_),
    .Y(_04873_),
    .B1(_04872_));
 sg13g2_nand2_1 _13949_ (.Y(_04874_),
    .A(net28),
    .B(_04758_));
 sg13g2_nand2_1 _13950_ (.Y(_04875_),
    .A(_04873_),
    .B(_04874_));
 sg13g2_nor2_1 _13951_ (.A(_04871_),
    .B(_04875_),
    .Y(_04876_));
 sg13g2_nand2_1 _13952_ (.Y(_04877_),
    .A(_04870_),
    .B(_04876_));
 sg13g2_nor2b_1 _13953_ (.A(_04153_),
    .B_N(_04767_),
    .Y(_04878_));
 sg13g2_nor3_1 _13954_ (.A(_04111_),
    .B(_04772_),
    .C(_04156_),
    .Y(_04879_));
 sg13g2_nor2_1 _13955_ (.A(_04878_),
    .B(_04879_),
    .Y(_04880_));
 sg13g2_nor2_1 _13956_ (.A(_04779_),
    .B(_04059_),
    .Y(_04881_));
 sg13g2_nor3_1 _13957_ (.A(_04126_),
    .B(_04755_),
    .C(_04131_),
    .Y(_04882_));
 sg13g2_nor2_1 _13958_ (.A(_04881_),
    .B(_04882_),
    .Y(_04883_));
 sg13g2_nand2_1 _13959_ (.Y(_04884_),
    .A(_04880_),
    .B(_04883_));
 sg13g2_nor2_1 _13960_ (.A(_04877_),
    .B(_04884_),
    .Y(_04885_));
 sg13g2_a21oi_1 _13961_ (.A1(_04867_),
    .A2(_04885_),
    .Y(_04886_),
    .B1(_04266_));
 sg13g2_inv_1 _13962_ (.Y(_04887_),
    .A(_04877_));
 sg13g2_nand2_1 _13963_ (.Y(_04888_),
    .A(_04166_),
    .B(net20));
 sg13g2_inv_1 _13964_ (.Y(_04889_),
    .A(_04881_));
 sg13g2_nand2_1 _13965_ (.Y(_04890_),
    .A(_04888_),
    .B(_04889_));
 sg13g2_nand2_1 _13966_ (.Y(_04891_),
    .A(_04167_),
    .B(_04773_));
 sg13g2_nand2b_1 _13967_ (.Y(_04892_),
    .B(_04891_),
    .A_N(_04878_));
 sg13g2_nor2_1 _13968_ (.A(_04890_),
    .B(_04892_),
    .Y(_04893_));
 sg13g2_nand2_1 _13969_ (.Y(_04894_),
    .A(_04887_),
    .B(_04893_));
 sg13g2_nand3_1 _13970_ (.B(_04853_),
    .C(_04858_),
    .A(_04866_),
    .Y(_04895_));
 sg13g2_buf_1 _13971_ (.A(_04895_),
    .X(_04896_));
 sg13g2_nand3_1 _13972_ (.B(_04896_),
    .C(net12),
    .A(_04894_),
    .Y(_04897_));
 sg13g2_buf_1 _13973_ (.A(_04897_),
    .X(_04898_));
 sg13g2_nand2_1 _13974_ (.Y(_04899_),
    .A(_04886_),
    .B(_04898_));
 sg13g2_nand2_1 _13975_ (.Y(_04900_),
    .A(_04899_),
    .B(_02032_));
 sg13g2_nand3_1 _13976_ (.B(_04898_),
    .C(_01949_),
    .A(_04886_),
    .Y(_04901_));
 sg13g2_nand2_1 _13977_ (.Y(_04902_),
    .A(_04900_),
    .B(_04901_));
 sg13g2_a21oi_1 _13978_ (.A1(_04810_),
    .A2(_01958_),
    .Y(_04903_),
    .B1(_04808_));
 sg13g2_a21oi_1 _13979_ (.A1(_04902_),
    .A2(_04903_),
    .Y(_04904_),
    .B1(_04407_));
 sg13g2_xnor2_1 _13980_ (.Y(_04905_),
    .A(_01949_),
    .B(_04899_));
 sg13g2_nand2b_1 _13981_ (.Y(_04906_),
    .B(_04905_),
    .A_N(_04903_));
 sg13g2_nand2_1 _13982_ (.Y(_04907_),
    .A(_04904_),
    .B(_04906_));
 sg13g2_o21ai_1 _13983_ (.B1(_04907_),
    .Y(_00070_),
    .A1(_04851_),
    .A2(_04852_));
 sg13g2_nor2b_1 _13984_ (.A(net24),
    .B_N(_04776_),
    .Y(_04908_));
 sg13g2_a22oi_1 _13985_ (.Y(_04909_),
    .B1(_04767_),
    .B2(net29),
    .A2(_04789_),
    .A1(net31));
 sg13g2_nand2_1 _13986_ (.Y(_04910_),
    .A(net28),
    .B(_04783_));
 sg13g2_nand2_1 _13987_ (.Y(_04911_),
    .A(_04909_),
    .B(_04910_));
 sg13g2_nor2_1 _13988_ (.A(_04908_),
    .B(_04911_),
    .Y(_04912_));
 sg13g2_nor2_1 _13989_ (.A(_04779_),
    .B(_04153_),
    .Y(_04913_));
 sg13g2_nor2_1 _13990_ (.A(_04772_),
    .B(_04044_),
    .Y(_04914_));
 sg13g2_nor2_1 _13991_ (.A(_04913_),
    .B(_04914_),
    .Y(_04915_));
 sg13g2_nand2_1 _13992_ (.Y(_04916_),
    .A(_04912_),
    .B(_04915_));
 sg13g2_nand2_1 _13993_ (.Y(_04917_),
    .A(_04327_),
    .B(net20));
 sg13g2_buf_1 _13994_ (.A(_04917_),
    .X(_04918_));
 sg13g2_inv_1 _13995_ (.Y(_04919_),
    .A(_04918_));
 sg13g2_a21oi_1 _13996_ (.A1(net15),
    .A2(_04916_),
    .Y(_04920_),
    .B1(_04919_));
 sg13g2_nand2_1 _13997_ (.Y(_04921_),
    .A(_04788_),
    .B(_04920_));
 sg13g2_nand2_1 _13998_ (.Y(_04922_),
    .A(net15),
    .B(_04916_));
 sg13g2_nand2_1 _13999_ (.Y(_04923_),
    .A(_04922_),
    .B(_04918_));
 sg13g2_nand2_1 _14000_ (.Y(_04924_),
    .A(_04923_),
    .B(_04787_));
 sg13g2_nand2_1 _14001_ (.Y(_04925_),
    .A(_04921_),
    .B(_04924_));
 sg13g2_nand2_1 _14002_ (.Y(_04926_),
    .A(_04925_),
    .B(_02034_));
 sg13g2_nand3_1 _14003_ (.B(_04924_),
    .C(_01955_),
    .A(_04921_),
    .Y(_04927_));
 sg13g2_buf_1 _14004_ (.A(_04927_),
    .X(_04928_));
 sg13g2_nand2_1 _14005_ (.Y(_04929_),
    .A(_04867_),
    .B(_04885_));
 sg13g2_nand2_1 _14006_ (.Y(_04930_),
    .A(_04929_),
    .B(net11));
 sg13g2_o21ai_1 _14007_ (.B1(_04898_),
    .Y(_04931_),
    .A1(_02032_),
    .A2(_04930_));
 sg13g2_a21oi_1 _14008_ (.A1(_04926_),
    .A2(_04928_),
    .Y(_04932_),
    .B1(_04931_));
 sg13g2_nand3_1 _14009_ (.B(_04926_),
    .C(_04928_),
    .A(_04931_),
    .Y(_04933_));
 sg13g2_buf_1 _14010_ (.A(_04933_),
    .X(_04934_));
 sg13g2_inv_1 _14011_ (.Y(_04935_),
    .A(_04934_));
 sg13g2_o21ai_1 _14012_ (.B1(_04906_),
    .Y(_04936_),
    .A1(_04932_),
    .A2(_04935_));
 sg13g2_nor2_1 _14013_ (.A(_04903_),
    .B(_04902_),
    .Y(_04937_));
 sg13g2_nand2_1 _14014_ (.Y(_04938_),
    .A(_04926_),
    .B(_04928_));
 sg13g2_inv_1 _14015_ (.Y(_04939_),
    .A(_04931_));
 sg13g2_nand2_1 _14016_ (.Y(_04940_),
    .A(_04938_),
    .B(_04939_));
 sg13g2_nand3_1 _14017_ (.B(_04934_),
    .C(_04940_),
    .A(_04937_),
    .Y(_04941_));
 sg13g2_nand3_1 _14018_ (.B(net126),
    .C(_04941_),
    .A(_04936_),
    .Y(_04942_));
 sg13g2_nor2_1 _14019_ (.A(_00124_),
    .B(_04848_),
    .Y(_04943_));
 sg13g2_buf_1 _14020_ (.A(\vgadonut.donut.sAcB[8] ),
    .X(_04944_));
 sg13g2_nor2_1 _14021_ (.A(net244),
    .B(net241),
    .Y(_04945_));
 sg13g2_nand2_1 _14022_ (.Y(_04946_),
    .A(_04816_),
    .B(net241));
 sg13g2_inv_1 _14023_ (.Y(_04947_),
    .A(_04946_));
 sg13g2_nor2_1 _14024_ (.A(_04945_),
    .B(_04947_),
    .Y(_04948_));
 sg13g2_inv_1 _14025_ (.Y(_04949_),
    .A(_04847_));
 sg13g2_a21oi_1 _14026_ (.A1(_04949_),
    .A2(_04844_),
    .Y(_04950_),
    .B1(_04843_));
 sg13g2_xnor2_1 _14027_ (.Y(_04951_),
    .A(_04948_),
    .B(_04950_));
 sg13g2_xnor2_1 _14028_ (.Y(_04952_),
    .A(\vgadonut.donut.donuthit.ryin[7] ),
    .B(_04951_));
 sg13g2_o21ai_1 _14029_ (.B1(_04952_),
    .Y(_04953_),
    .A1(_04851_),
    .A2(_04943_));
 sg13g2_nor2_1 _14030_ (.A(_04943_),
    .B(_04851_),
    .Y(_04954_));
 sg13g2_nand2b_1 _14031_ (.Y(_04955_),
    .B(_04954_),
    .A_N(_04952_));
 sg13g2_nand3_1 _14032_ (.B(_04955_),
    .C(net112),
    .A(_04953_),
    .Y(_04956_));
 sg13g2_nand2_1 _14033_ (.Y(_00071_),
    .A(_04942_),
    .B(_04956_));
 sg13g2_inv_1 _14034_ (.Y(_04957_),
    .A(\vgadonut.donut.donuthit.ryin[8] ));
 sg13g2_buf_1 _14035_ (.A(\vgadonut.donut.sAcB[9] ),
    .X(_04958_));
 sg13g2_buf_1 _14036_ (.A(_04958_),
    .X(_04959_));
 sg13g2_nor2_1 _14037_ (.A(net242),
    .B(net207),
    .Y(_04960_));
 sg13g2_nand2_1 _14038_ (.Y(_04961_),
    .A(net242),
    .B(net207));
 sg13g2_nor2b_1 _14039_ (.A(_04960_),
    .B_N(_04961_),
    .Y(_04962_));
 sg13g2_inv_1 _14040_ (.Y(_04963_),
    .A(_04950_));
 sg13g2_a21oi_1 _14041_ (.A1(_04963_),
    .A2(_04946_),
    .Y(_04964_),
    .B1(_04945_));
 sg13g2_xor2_1 _14042_ (.B(_04964_),
    .A(_04962_),
    .X(_04965_));
 sg13g2_xnor2_1 _14043_ (.Y(_04966_),
    .A(_04957_),
    .B(_04965_));
 sg13g2_o21ai_1 _14044_ (.B1(_04953_),
    .Y(_04967_),
    .A1(_00125_),
    .A2(_04951_));
 sg13g2_xor2_1 _14045_ (.B(_04967_),
    .A(_04966_),
    .X(_04968_));
 sg13g2_o21ai_1 _14046_ (.B1(_04934_),
    .Y(_04969_),
    .A1(_04932_),
    .A2(_04906_));
 sg13g2_inv_1 _14047_ (.Y(_04970_),
    .A(_04969_));
 sg13g2_a22oi_1 _14048_ (.Y(_04971_),
    .B1(_01955_),
    .B2(_04921_),
    .A2(_04923_),
    .A1(_04787_));
 sg13g2_buf_1 _14049_ (.A(_04971_),
    .X(_04972_));
 sg13g2_nand2_1 _14050_ (.Y(_04973_),
    .A(net17),
    .B(_04757_));
 sg13g2_o21ai_1 _14051_ (.B1(_04973_),
    .Y(_04974_),
    .A1(_04153_),
    .A2(_04772_));
 sg13g2_nand2_1 _14052_ (.Y(_04975_),
    .A(net16),
    .B(_04780_));
 sg13g2_nand2_1 _14053_ (.Y(_04976_),
    .A(net22),
    .B(_04776_));
 sg13g2_a22oi_1 _14054_ (.Y(_04977_),
    .B1(_04783_),
    .B2(net21),
    .A2(_04767_),
    .A1(net27));
 sg13g2_nand3_1 _14055_ (.B(_04976_),
    .C(_04977_),
    .A(_04975_),
    .Y(_04978_));
 sg13g2_nor2_1 _14056_ (.A(_04974_),
    .B(_04978_),
    .Y(_04979_));
 sg13g2_nand2_1 _14057_ (.Y(_04980_),
    .A(_04979_),
    .B(_04918_));
 sg13g2_nand2_1 _14058_ (.Y(_04981_),
    .A(_04980_),
    .B(net13));
 sg13g2_nand2_1 _14059_ (.Y(_04982_),
    .A(_04896_),
    .B(net11));
 sg13g2_nand2_1 _14060_ (.Y(_04983_),
    .A(_04981_),
    .B(_04982_));
 sg13g2_nand3_1 _14061_ (.B(_04896_),
    .C(net10),
    .A(_04980_),
    .Y(_04984_));
 sg13g2_nand2_1 _14062_ (.Y(_04985_),
    .A(_04983_),
    .B(_04984_));
 sg13g2_xnor2_1 _14063_ (.Y(_04986_),
    .A(_01977_),
    .B(_04985_));
 sg13g2_xnor2_1 _14064_ (.Y(_04987_),
    .A(_04972_),
    .B(_04986_));
 sg13g2_o21ai_1 _14065_ (.B1(net138),
    .Y(_04988_),
    .A1(_04987_),
    .A2(_04970_));
 sg13g2_a21oi_1 _14066_ (.A1(_04970_),
    .A2(_04987_),
    .Y(_04989_),
    .B1(_04988_));
 sg13g2_a21o_1 _14067_ (.A2(_04968_),
    .A1(net110),
    .B1(_04989_),
    .X(_00072_));
 sg13g2_buf_1 _14068_ (.A(\vgadonut.donut.sAcB[10] ),
    .X(_04990_));
 sg13g2_nor2_1 _14069_ (.A(net241),
    .B(net240),
    .Y(_04991_));
 sg13g2_nand2_1 _14070_ (.Y(_04992_),
    .A(net241),
    .B(net240));
 sg13g2_nor2b_1 _14071_ (.A(_04991_),
    .B_N(_04992_),
    .Y(_04993_));
 sg13g2_inv_1 _14072_ (.Y(_04994_),
    .A(_04964_));
 sg13g2_a21oi_1 _14073_ (.A1(_04994_),
    .A2(_04961_),
    .Y(_04995_),
    .B1(_04960_));
 sg13g2_xor2_1 _14074_ (.B(_04995_),
    .A(_04993_),
    .X(_04996_));
 sg13g2_xnor2_1 _14075_ (.Y(_04997_),
    .A(\vgadonut.donut.donuthit.ryin[9] ),
    .B(_04996_));
 sg13g2_inv_1 _14076_ (.Y(_04998_),
    .A(_00126_));
 sg13g2_a22oi_1 _14077_ (.Y(_04999_),
    .B1(_04966_),
    .B2(_04967_),
    .A2(_04965_),
    .A1(_04998_));
 sg13g2_nor2_1 _14078_ (.A(_04997_),
    .B(_04999_),
    .Y(_05000_));
 sg13g2_inv_1 _14079_ (.Y(_05001_),
    .A(_05000_));
 sg13g2_a21oi_1 _14080_ (.A1(_04999_),
    .A2(_04997_),
    .Y(_05002_),
    .B1(net125));
 sg13g2_inv_1 _14081_ (.Y(_05003_),
    .A(_04984_));
 sg13g2_a21oi_2 _14082_ (.B1(_05003_),
    .Y(_05004_),
    .A2(_01975_),
    .A1(_04983_));
 sg13g2_nand2_1 _14083_ (.Y(_05005_),
    .A(net16),
    .B(_04773_));
 sg13g2_nand2_1 _14084_ (.Y(_05006_),
    .A(net22),
    .B(_04780_));
 sg13g2_a22oi_1 _14085_ (.Y(_05007_),
    .B1(_04776_),
    .B2(net21),
    .A2(_04783_),
    .A1(net27));
 sg13g2_nand3_1 _14086_ (.B(_05006_),
    .C(_05007_),
    .A(_05005_),
    .Y(_05008_));
 sg13g2_nand2_1 _14087_ (.Y(_05009_),
    .A(_04431_),
    .B(_04756_));
 sg13g2_nor2b_1 _14088_ (.A(_05008_),
    .B_N(_05009_),
    .Y(_05010_));
 sg13g2_nand2_1 _14089_ (.Y(_05011_),
    .A(_05010_),
    .B(_04918_));
 sg13g2_nand2_1 _14090_ (.Y(_05012_),
    .A(_05011_),
    .B(net12));
 sg13g2_nand2_1 _14091_ (.Y(_05013_),
    .A(_05012_),
    .B(_04920_));
 sg13g2_nand2_1 _14092_ (.Y(_05014_),
    .A(_04923_),
    .B(_05011_));
 sg13g2_nand2_1 _14093_ (.Y(_05015_),
    .A(_05013_),
    .B(_05014_));
 sg13g2_xnor2_1 _14094_ (.Y(_05016_),
    .A(_02048_),
    .B(_05015_));
 sg13g2_xnor2_1 _14095_ (.Y(_05017_),
    .A(_05004_),
    .B(_05016_));
 sg13g2_nor2_1 _14096_ (.A(_04972_),
    .B(_04986_),
    .Y(_05018_));
 sg13g2_nor2_1 _14097_ (.A(_05018_),
    .B(_04935_),
    .Y(_05019_));
 sg13g2_nand2_1 _14098_ (.Y(_05020_),
    .A(_04941_),
    .B(_05019_));
 sg13g2_nand2_1 _14099_ (.Y(_05021_),
    .A(_04986_),
    .B(_04972_));
 sg13g2_nand2_1 _14100_ (.Y(_05022_),
    .A(_05020_),
    .B(_05021_));
 sg13g2_o21ai_1 _14101_ (.B1(net138),
    .Y(_05023_),
    .A1(_05017_),
    .A2(_05022_));
 sg13g2_a21oi_1 _14102_ (.A1(_05017_),
    .A2(_05022_),
    .Y(_05024_),
    .B1(_05023_));
 sg13g2_a21o_1 _14103_ (.A2(_05002_),
    .A1(_05001_),
    .B1(_05024_),
    .X(_00073_));
 sg13g2_buf_1 _14104_ (.A(\vgadonut.donut.sAcB[11] ),
    .X(_05025_));
 sg13g2_nor2_1 _14105_ (.A(net207),
    .B(net239),
    .Y(_05026_));
 sg13g2_nand2_1 _14106_ (.Y(_05027_),
    .A(net207),
    .B(net239));
 sg13g2_nor2b_1 _14107_ (.A(_05026_),
    .B_N(_05027_),
    .Y(_05028_));
 sg13g2_inv_1 _14108_ (.Y(_05029_),
    .A(_04995_));
 sg13g2_a21oi_1 _14109_ (.A1(_05029_),
    .A2(_04992_),
    .Y(_05030_),
    .B1(_04991_));
 sg13g2_xor2_1 _14110_ (.B(_05030_),
    .A(_05028_),
    .X(_05031_));
 sg13g2_xnor2_1 _14111_ (.Y(_05032_),
    .A(\vgadonut.donut.donuthit.ryin[10] ),
    .B(_05031_));
 sg13g2_inv_1 _14112_ (.Y(_05033_),
    .A(_00127_));
 sg13g2_a21oi_1 _14113_ (.A1(_05033_),
    .A2(_04996_),
    .Y(_05034_),
    .B1(_05000_));
 sg13g2_nor2_1 _14114_ (.A(_05032_),
    .B(_05034_),
    .Y(_05035_));
 sg13g2_a21o_1 _14115_ (.A2(_05032_),
    .A1(_05034_),
    .B1(net137),
    .X(_05036_));
 sg13g2_nor2_1 _14116_ (.A(_05017_),
    .B(_04987_),
    .Y(_05037_));
 sg13g2_nand2_1 _14117_ (.Y(_05038_),
    .A(_04969_),
    .B(_05037_));
 sg13g2_nand2_1 _14118_ (.Y(_05039_),
    .A(_05016_),
    .B(_05004_));
 sg13g2_nor2_1 _14119_ (.A(_05004_),
    .B(_05016_),
    .Y(_05040_));
 sg13g2_a21oi_1 _14120_ (.A1(_05018_),
    .A2(_05039_),
    .Y(_05041_),
    .B1(_05040_));
 sg13g2_nand2_1 _14121_ (.Y(_05042_),
    .A(_05038_),
    .B(_05041_));
 sg13g2_nor2_1 _14122_ (.A(_04755_),
    .B(net24),
    .Y(_05043_));
 sg13g2_nand2_1 _14123_ (.Y(_05044_),
    .A(net22),
    .B(_04773_));
 sg13g2_a22oi_1 _14124_ (.Y(_05045_),
    .B1(_04780_),
    .B2(net21),
    .A2(_04776_),
    .A1(net27));
 sg13g2_nand3_1 _14125_ (.B(_05044_),
    .C(_05045_),
    .A(_05009_),
    .Y(_05046_));
 sg13g2_nor2_1 _14126_ (.A(_05043_),
    .B(_05046_),
    .Y(_05047_));
 sg13g2_nand2_1 _14127_ (.Y(_05048_),
    .A(_05047_),
    .B(_04918_));
 sg13g2_nand2_1 _14128_ (.Y(_05049_),
    .A(_05048_),
    .B(net13));
 sg13g2_nand2_1 _14129_ (.Y(_05050_),
    .A(_04981_),
    .B(_05049_));
 sg13g2_nand3_1 _14130_ (.B(_05048_),
    .C(net10),
    .A(_04980_),
    .Y(_05051_));
 sg13g2_nand2_1 _14131_ (.Y(_05052_),
    .A(_05050_),
    .B(_05051_));
 sg13g2_xor2_1 _14132_ (.B(_05052_),
    .A(_01981_),
    .X(_05053_));
 sg13g2_a22oi_1 _14133_ (.Y(_05054_),
    .B1(_01968_),
    .B2(_05013_),
    .A2(_05011_),
    .A1(_04923_));
 sg13g2_nand2_1 _14134_ (.Y(_05055_),
    .A(_05053_),
    .B(_05054_));
 sg13g2_xnor2_1 _14135_ (.Y(_05056_),
    .A(_01981_),
    .B(_05052_));
 sg13g2_nand2b_1 _14136_ (.Y(_05057_),
    .B(_05056_),
    .A_N(_05054_));
 sg13g2_nand2_1 _14137_ (.Y(_05058_),
    .A(_05055_),
    .B(_05057_));
 sg13g2_inv_1 _14138_ (.Y(_05059_),
    .A(_05058_));
 sg13g2_a21oi_1 _14139_ (.A1(_05042_),
    .A2(_05059_),
    .Y(_05060_),
    .B1(net111));
 sg13g2_o21ai_1 _14140_ (.B1(_05060_),
    .Y(_05061_),
    .A1(_05042_),
    .A2(_05059_));
 sg13g2_o21ai_1 _14141_ (.B1(_05061_),
    .Y(_00074_),
    .A1(_05035_),
    .A2(_05036_));
 sg13g2_buf_1 _14142_ (.A(\vgadonut.donut.sAcB[12] ),
    .X(_05062_));
 sg13g2_nor2_1 _14143_ (.A(net240),
    .B(net238),
    .Y(_05063_));
 sg13g2_nand2_1 _14144_ (.Y(_05064_),
    .A(net240),
    .B(net238));
 sg13g2_inv_1 _14145_ (.Y(_05065_),
    .A(_05064_));
 sg13g2_nor2_1 _14146_ (.A(_05063_),
    .B(_05065_),
    .Y(_05066_));
 sg13g2_inv_1 _14147_ (.Y(_05067_),
    .A(_05030_));
 sg13g2_a21oi_1 _14148_ (.A1(_05067_),
    .A2(_05027_),
    .Y(_05068_),
    .B1(_05026_));
 sg13g2_xor2_1 _14149_ (.B(_05068_),
    .A(_05066_),
    .X(_05069_));
 sg13g2_xnor2_1 _14150_ (.Y(_05070_),
    .A(\vgadonut.donut.donuthit.ryin[11] ),
    .B(_05069_));
 sg13g2_inv_1 _14151_ (.Y(_05071_),
    .A(_00128_));
 sg13g2_a21oi_1 _14152_ (.A1(_05071_),
    .A2(_05031_),
    .Y(_05072_),
    .B1(_05035_));
 sg13g2_or2_1 _14153_ (.X(_05073_),
    .B(_05072_),
    .A(_05070_));
 sg13g2_a21oi_1 _14154_ (.A1(_05072_),
    .A2(_05070_),
    .Y(_05074_),
    .B1(net125));
 sg13g2_nor2_1 _14155_ (.A(_05017_),
    .B(_05058_),
    .Y(_05075_));
 sg13g2_nand3_1 _14156_ (.B(_05021_),
    .C(_05075_),
    .A(_05020_),
    .Y(_05076_));
 sg13g2_inv_1 _14157_ (.Y(_05077_),
    .A(_05057_));
 sg13g2_a21oi_1 _14158_ (.A1(_05055_),
    .A2(_05040_),
    .Y(_05078_),
    .B1(_05077_));
 sg13g2_nand2_1 _14159_ (.Y(_05079_),
    .A(_05076_),
    .B(_05078_));
 sg13g2_inv_1 _14160_ (.Y(_05080_),
    .A(_05051_));
 sg13g2_a21oi_1 _14161_ (.A1(_05050_),
    .A2(_01981_),
    .Y(_05081_),
    .B1(_05080_));
 sg13g2_nand2_1 _14162_ (.Y(_05082_),
    .A(_04517_),
    .B(net20));
 sg13g2_a22oi_1 _14163_ (.Y(_05083_),
    .B1(_04773_),
    .B2(net21),
    .A2(_04780_),
    .A1(net27));
 sg13g2_nand2_1 _14164_ (.Y(_05084_),
    .A(_05082_),
    .B(_05083_));
 sg13g2_nand2_1 _14165_ (.Y(_05085_),
    .A(_05084_),
    .B(net11));
 sg13g2_nand2_1 _14166_ (.Y(_05086_),
    .A(_05085_),
    .B(_05012_));
 sg13g2_nand3_1 _14167_ (.B(net11),
    .C(_05011_),
    .A(_05084_),
    .Y(_05087_));
 sg13g2_nand2_1 _14168_ (.Y(_05088_),
    .A(_05086_),
    .B(_05087_));
 sg13g2_xnor2_1 _14169_ (.Y(_05089_),
    .A(_01986_),
    .B(_05088_));
 sg13g2_xnor2_1 _14170_ (.Y(_05090_),
    .A(_05081_),
    .B(_05089_));
 sg13g2_o21ai_1 _14171_ (.B1(net138),
    .Y(_05091_),
    .A1(_05090_),
    .A2(_05079_));
 sg13g2_a21oi_1 _14172_ (.A1(_05079_),
    .A2(_05090_),
    .Y(_05092_),
    .B1(_05091_));
 sg13g2_a21o_1 _14173_ (.A2(_05074_),
    .A1(_05073_),
    .B1(_05092_),
    .X(_00075_));
 sg13g2_inv_1 _14174_ (.Y(_05093_),
    .A(\vgadonut.donut.donuthit.ryin[12] ));
 sg13g2_buf_1 _14175_ (.A(\vgadonut.donut.sAcB[13] ),
    .X(_05094_));
 sg13g2_buf_1 _14176_ (.A(_05094_),
    .X(_05095_));
 sg13g2_nor2_1 _14177_ (.A(net239),
    .B(net206),
    .Y(_05096_));
 sg13g2_nand2_1 _14178_ (.Y(_05097_),
    .A(net239),
    .B(net206));
 sg13g2_nor2b_1 _14179_ (.A(_05096_),
    .B_N(_05097_),
    .Y(_05098_));
 sg13g2_inv_1 _14180_ (.Y(_05099_),
    .A(_05063_));
 sg13g2_a21oi_1 _14181_ (.A1(_05068_),
    .A2(_05099_),
    .Y(_05100_),
    .B1(_05065_));
 sg13g2_xnor2_1 _14182_ (.Y(_05101_),
    .A(_05098_),
    .B(_05100_));
 sg13g2_xnor2_1 _14183_ (.Y(_05102_),
    .A(_05093_),
    .B(_05101_));
 sg13g2_inv_1 _14184_ (.Y(_05103_),
    .A(_05069_));
 sg13g2_o21ai_1 _14185_ (.B1(_05073_),
    .Y(_05104_),
    .A1(_00129_),
    .A2(_05103_));
 sg13g2_xnor2_1 _14186_ (.Y(_05105_),
    .A(_05102_),
    .B(_05104_));
 sg13g2_inv_1 _14187_ (.Y(_05106_),
    .A(_05041_));
 sg13g2_inv_1 _14188_ (.Y(_05107_),
    .A(_05081_));
 sg13g2_nand2_1 _14189_ (.Y(_05108_),
    .A(_05089_),
    .B(_05107_));
 sg13g2_nor2_1 _14190_ (.A(_05107_),
    .B(_05089_),
    .Y(_05109_));
 sg13g2_a21oi_1 _14191_ (.A1(_05108_),
    .A2(_05057_),
    .Y(_05110_),
    .B1(_05109_));
 sg13g2_nor2_1 _14192_ (.A(_05106_),
    .B(_05110_),
    .Y(_05111_));
 sg13g2_nand2_1 _14193_ (.Y(_05112_),
    .A(_05111_),
    .B(_05038_));
 sg13g2_inv_1 _14194_ (.Y(_05113_),
    .A(_05110_));
 sg13g2_nand2_1 _14195_ (.Y(_05114_),
    .A(_05090_),
    .B(_05059_));
 sg13g2_nand2_1 _14196_ (.Y(_05115_),
    .A(_05113_),
    .B(_05114_));
 sg13g2_inv_1 _14197_ (.Y(_05116_),
    .A(_05087_));
 sg13g2_a21oi_1 _14198_ (.A1(_05086_),
    .A2(_01986_),
    .Y(_05117_),
    .B1(_05116_));
 sg13g2_inv_1 _14199_ (.Y(_05118_),
    .A(_05117_));
 sg13g2_a22oi_1 _14200_ (.Y(_05119_),
    .B1(_04757_),
    .B2(net21),
    .A2(_04773_),
    .A1(net27));
 sg13g2_nand2_1 _14201_ (.Y(_05120_),
    .A(_05082_),
    .B(_05119_));
 sg13g2_nand2_1 _14202_ (.Y(_05121_),
    .A(_05120_),
    .B(net13));
 sg13g2_nand2_1 _14203_ (.Y(_05122_),
    .A(_05121_),
    .B(_05049_));
 sg13g2_nand3_1 _14204_ (.B(net11),
    .C(_05048_),
    .A(_05120_),
    .Y(_05123_));
 sg13g2_nand2_1 _14205_ (.Y(_05124_),
    .A(_05122_),
    .B(_05123_));
 sg13g2_xnor2_1 _14206_ (.Y(_05125_),
    .A(_01894_),
    .B(_05124_));
 sg13g2_nor2_1 _14207_ (.A(_05118_),
    .B(_05125_),
    .Y(_05126_));
 sg13g2_nand2_1 _14208_ (.Y(_05127_),
    .A(_05125_),
    .B(_05118_));
 sg13g2_inv_1 _14209_ (.Y(_05128_),
    .A(_05127_));
 sg13g2_nor2_1 _14210_ (.A(_05126_),
    .B(_05128_),
    .Y(_05129_));
 sg13g2_a21oi_1 _14211_ (.A1(_05112_),
    .A2(_05115_),
    .Y(_05130_),
    .B1(_05129_));
 sg13g2_nand3_1 _14212_ (.B(_05129_),
    .C(_05115_),
    .A(_05112_),
    .Y(_05131_));
 sg13g2_nand3b_1 _14213_ (.B(net123),
    .C(_05131_),
    .Y(_05132_),
    .A_N(_05130_));
 sg13g2_o21ai_1 _14214_ (.B1(_05132_),
    .Y(_00076_),
    .A1(net122),
    .A2(_05105_));
 sg13g2_inv_1 _14215_ (.Y(_05133_),
    .A(\vgadonut.donut.donuthit.ryin[13] ));
 sg13g2_buf_1 _14216_ (.A(\vgadonut.donut.sAcB[14] ),
    .X(_05134_));
 sg13g2_buf_1 _14217_ (.A(_05134_),
    .X(_05135_));
 sg13g2_nor2_1 _14218_ (.A(net238),
    .B(net205),
    .Y(_05136_));
 sg13g2_nand2_1 _14219_ (.Y(_05137_),
    .A(net238),
    .B(net205));
 sg13g2_inv_1 _14220_ (.Y(_05138_),
    .A(_05137_));
 sg13g2_nor2_1 _14221_ (.A(_05136_),
    .B(_05138_),
    .Y(_05139_));
 sg13g2_o21ai_1 _14222_ (.B1(_05097_),
    .Y(_05140_),
    .A1(_05096_),
    .A2(_05100_));
 sg13g2_xor2_1 _14223_ (.B(_05140_),
    .A(_05139_),
    .X(_05141_));
 sg13g2_xnor2_1 _14224_ (.Y(_05142_),
    .A(_05133_),
    .B(_05141_));
 sg13g2_inv_1 _14225_ (.Y(_05143_),
    .A(_05101_));
 sg13g2_nand2_1 _14226_ (.Y(_05144_),
    .A(_05104_),
    .B(_05102_));
 sg13g2_o21ai_1 _14227_ (.B1(_05144_),
    .Y(_05145_),
    .A1(_00130_),
    .A2(_05143_));
 sg13g2_xnor2_1 _14228_ (.Y(_05146_),
    .A(_05142_),
    .B(_05145_));
 sg13g2_a21oi_1 _14229_ (.A1(_05108_),
    .A2(_05127_),
    .Y(_05147_),
    .B1(_05126_));
 sg13g2_nor2b_1 _14230_ (.A(_05147_),
    .B_N(_05078_),
    .Y(_05148_));
 sg13g2_nand2_1 _14231_ (.Y(_05149_),
    .A(_05076_),
    .B(_05148_));
 sg13g2_nand2_1 _14232_ (.Y(_05150_),
    .A(_05129_),
    .B(_05090_));
 sg13g2_nand2b_1 _14233_ (.Y(_05151_),
    .B(_05150_),
    .A_N(_05147_));
 sg13g2_inv_1 _14234_ (.Y(_05152_),
    .A(_05123_));
 sg13g2_a21oi_2 _14235_ (.B1(_05152_),
    .Y(_05153_),
    .A2(_01894_),
    .A1(_05122_));
 sg13g2_nand2_1 _14236_ (.Y(_05154_),
    .A(net12),
    .B(net20));
 sg13g2_buf_2 _14237_ (.A(_05154_),
    .X(_05155_));
 sg13g2_nand2_1 _14238_ (.Y(_05156_),
    .A(_05085_),
    .B(_05155_));
 sg13g2_nand3_1 _14239_ (.B(net10),
    .C(net20),
    .A(_05084_),
    .Y(_05157_));
 sg13g2_nand2_1 _14240_ (.Y(_05158_),
    .A(_05156_),
    .B(_05157_));
 sg13g2_xnor2_1 _14241_ (.Y(_05159_),
    .A(_02013_),
    .B(_05158_));
 sg13g2_xnor2_1 _14242_ (.Y(_05160_),
    .A(_05153_),
    .B(_05159_));
 sg13g2_inv_2 _14243_ (.Y(_05161_),
    .A(_05160_));
 sg13g2_a21oi_1 _14244_ (.A1(_05149_),
    .A2(_05151_),
    .Y(_05162_),
    .B1(_05161_));
 sg13g2_nand3_1 _14245_ (.B(_05161_),
    .C(_05151_),
    .A(_05149_),
    .Y(_05163_));
 sg13g2_nand3b_1 _14246_ (.B(net123),
    .C(_05163_),
    .Y(_05164_),
    .A_N(_05162_));
 sg13g2_o21ai_1 _14247_ (.B1(_05164_),
    .Y(_00077_),
    .A1(net122),
    .A2(_05146_));
 sg13g2_nor2b_1 _14248_ (.A(_00131_),
    .B_N(_05141_),
    .Y(_05165_));
 sg13g2_a21oi_1 _14249_ (.A1(_05145_),
    .A2(_05142_),
    .Y(_05166_),
    .B1(_05165_));
 sg13g2_inv_2 _14250_ (.Y(_05167_),
    .A(\vgadonut.donut.donuthit.ryin[14] ));
 sg13g2_buf_2 _14251_ (.A(\vgadonut.donut.sAcB[15] ),
    .X(_05168_));
 sg13g2_buf_1 _14252_ (.A(_05168_),
    .X(_05169_));
 sg13g2_nor2_1 _14253_ (.A(net206),
    .B(net204),
    .Y(_05170_));
 sg13g2_nand2_1 _14254_ (.Y(_05171_),
    .A(net206),
    .B(net204));
 sg13g2_nor2b_1 _14255_ (.A(_05170_),
    .B_N(_05171_),
    .Y(_05172_));
 sg13g2_inv_1 _14256_ (.Y(_05173_),
    .A(_05136_));
 sg13g2_a21oi_1 _14257_ (.A1(_05140_),
    .A2(_05173_),
    .Y(_05174_),
    .B1(_05138_));
 sg13g2_xnor2_1 _14258_ (.Y(_05175_),
    .A(_05172_),
    .B(_05174_));
 sg13g2_xnor2_1 _14259_ (.Y(_05176_),
    .A(_05167_),
    .B(_05175_));
 sg13g2_nor2b_1 _14260_ (.A(_05166_),
    .B_N(_05176_),
    .Y(_05177_));
 sg13g2_inv_1 _14261_ (.Y(_05178_),
    .A(_05166_));
 sg13g2_o21ai_1 _14262_ (.B1(net112),
    .Y(_05179_),
    .A1(_05176_),
    .A2(_05178_));
 sg13g2_nand2_1 _14263_ (.Y(_05180_),
    .A(_05161_),
    .B(_05129_));
 sg13g2_nor2_1 _14264_ (.A(_05114_),
    .B(_05180_),
    .Y(_05181_));
 sg13g2_nand2_1 _14265_ (.Y(_05182_),
    .A(_05042_),
    .B(_05181_));
 sg13g2_nor2_1 _14266_ (.A(_05153_),
    .B(_05159_),
    .Y(_05183_));
 sg13g2_nor2_1 _14267_ (.A(_05183_),
    .B(_05128_),
    .Y(_05184_));
 sg13g2_nand2_1 _14268_ (.Y(_05185_),
    .A(_05159_),
    .B(_05153_));
 sg13g2_nor2b_1 _14269_ (.A(_05184_),
    .B_N(_05185_),
    .Y(_05186_));
 sg13g2_nor2_1 _14270_ (.A(_05113_),
    .B(_05180_),
    .Y(_05187_));
 sg13g2_nor2_1 _14271_ (.A(_05186_),
    .B(_05187_),
    .Y(_05188_));
 sg13g2_nand2_1 _14272_ (.Y(_05189_),
    .A(_05182_),
    .B(_05188_));
 sg13g2_inv_1 _14273_ (.Y(_05190_),
    .A(_05157_));
 sg13g2_a21oi_2 _14274_ (.B1(_05190_),
    .Y(_05191_),
    .A2(_01890_),
    .A1(_05156_));
 sg13g2_nand2_1 _14275_ (.Y(_05192_),
    .A(_05121_),
    .B(_05155_));
 sg13g2_nand3_1 _14276_ (.B(net10),
    .C(net20),
    .A(_05120_),
    .Y(_05193_));
 sg13g2_nand2_1 _14277_ (.Y(_05194_),
    .A(_05192_),
    .B(_05193_));
 sg13g2_xnor2_1 _14278_ (.Y(_05195_),
    .A(_02074_),
    .B(_05194_));
 sg13g2_xor2_1 _14279_ (.B(_05195_),
    .A(_05191_),
    .X(_05196_));
 sg13g2_a21oi_1 _14280_ (.A1(_05189_),
    .A2(_05196_),
    .Y(_05197_),
    .B1(net111));
 sg13g2_o21ai_1 _14281_ (.B1(_05197_),
    .Y(_05198_),
    .A1(_05189_),
    .A2(_05196_));
 sg13g2_o21ai_1 _14282_ (.B1(_05198_),
    .Y(_00078_),
    .A1(_05177_),
    .A2(_05179_));
 sg13g2_inv_1 _14283_ (.Y(_05199_),
    .A(_05193_));
 sg13g2_a21oi_1 _14284_ (.A1(_05192_),
    .A2(_01901_),
    .Y(_05200_),
    .B1(_05199_));
 sg13g2_nor2_1 _14285_ (.A(_01904_),
    .B(_05200_),
    .Y(_05201_));
 sg13g2_inv_1 _14286_ (.Y(_05202_),
    .A(_05201_));
 sg13g2_nand2_1 _14287_ (.Y(_05203_),
    .A(_05200_),
    .B(_01904_));
 sg13g2_nand2_1 _14288_ (.Y(_05204_),
    .A(_05202_),
    .B(_05203_));
 sg13g2_inv_1 _14289_ (.Y(_05205_),
    .A(_05204_));
 sg13g2_xnor2_1 _14290_ (.Y(_05206_),
    .A(_05191_),
    .B(_05195_));
 sg13g2_nor2_1 _14291_ (.A(_05160_),
    .B(_05206_),
    .Y(_05207_));
 sg13g2_nand2_1 _14292_ (.Y(_05208_),
    .A(_05207_),
    .B(_05147_));
 sg13g2_nor2_1 _14293_ (.A(_05191_),
    .B(_05195_),
    .Y(_05209_));
 sg13g2_nand2_1 _14294_ (.Y(_05210_),
    .A(_05195_),
    .B(_05191_));
 sg13g2_o21ai_1 _14295_ (.B1(_05210_),
    .Y(_05211_),
    .A1(_05183_),
    .A2(_05209_));
 sg13g2_nand2_1 _14296_ (.Y(_05212_),
    .A(_05208_),
    .B(_05211_));
 sg13g2_inv_1 _14297_ (.Y(_05213_),
    .A(_05207_));
 sg13g2_nor2_1 _14298_ (.A(_05150_),
    .B(_05213_),
    .Y(_05214_));
 sg13g2_nand2_1 _14299_ (.Y(_05215_),
    .A(_05079_),
    .B(_05214_));
 sg13g2_nand2b_1 _14300_ (.Y(_05216_),
    .B(_05215_),
    .A_N(_05212_));
 sg13g2_nor2_1 _14301_ (.A(_05205_),
    .B(_05216_),
    .Y(_05217_));
 sg13g2_nand2_1 _14302_ (.Y(_05218_),
    .A(_05216_),
    .B(_05205_));
 sg13g2_nand2_1 _14303_ (.Y(_05219_),
    .A(_05218_),
    .B(net125));
 sg13g2_inv_1 _14304_ (.Y(_05220_),
    .A(_00132_));
 sg13g2_a21oi_1 _14305_ (.A1(_05220_),
    .A2(_05175_),
    .Y(_05221_),
    .B1(_05177_));
 sg13g2_inv_2 _14306_ (.Y(_05222_),
    .A(\vgadonut.donut.donuthit.ryin[15] ));
 sg13g2_xor2_1 _14307_ (.B(net204),
    .A(net205),
    .X(_05223_));
 sg13g2_o21ai_1 _14308_ (.B1(_05171_),
    .Y(_05224_),
    .A1(_05170_),
    .A2(_05174_));
 sg13g2_xnor2_1 _14309_ (.Y(_05225_),
    .A(_05223_),
    .B(_05224_));
 sg13g2_xnor2_1 _14310_ (.Y(_05226_),
    .A(_05222_),
    .B(_05225_));
 sg13g2_a21oi_1 _14311_ (.A1(_05221_),
    .A2(_05226_),
    .Y(_05227_),
    .B1(net137));
 sg13g2_or2_1 _14312_ (.X(_05228_),
    .B(_05221_),
    .A(_05226_));
 sg13g2_nand2_1 _14313_ (.Y(_05229_),
    .A(_05227_),
    .B(_05228_));
 sg13g2_o21ai_1 _14314_ (.B1(_05229_),
    .Y(_00064_),
    .A1(_05217_),
    .A2(_05219_));
 sg13g2_inv_1 _14315_ (.Y(_05230_),
    .A(_01921_));
 sg13g2_xnor2_1 _14316_ (.Y(_05231_),
    .A(_05230_),
    .B(_05155_));
 sg13g2_inv_1 _14317_ (.Y(_05232_),
    .A(_05231_));
 sg13g2_nor2_1 _14318_ (.A(_05204_),
    .B(_05206_),
    .Y(_05233_));
 sg13g2_nand2_1 _14319_ (.Y(_05234_),
    .A(_05186_),
    .B(_05233_));
 sg13g2_o21ai_1 _14320_ (.B1(_05203_),
    .Y(_05235_),
    .A1(_05201_),
    .A2(_05209_));
 sg13g2_nand2_1 _14321_ (.Y(_05236_),
    .A(_05234_),
    .B(_05235_));
 sg13g2_nand2_1 _14322_ (.Y(_05237_),
    .A(_05196_),
    .B(_05205_));
 sg13g2_nor2_1 _14323_ (.A(_05237_),
    .B(_05180_),
    .Y(_05238_));
 sg13g2_nand3_1 _14324_ (.B(_05115_),
    .C(_05238_),
    .A(_05112_),
    .Y(_05239_));
 sg13g2_nand2b_1 _14325_ (.Y(_05240_),
    .B(_05239_),
    .A_N(_05236_));
 sg13g2_xnor2_1 _14326_ (.Y(_05241_),
    .A(_05232_),
    .B(_05240_));
 sg13g2_o21ai_1 _14327_ (.B1(_05228_),
    .Y(_05242_),
    .A1(_00181_),
    .A2(_05225_));
 sg13g2_nand3b_1 _14328_ (.B(_05172_),
    .C(_05223_),
    .Y(_05243_),
    .A_N(_05174_));
 sg13g2_o21ai_1 _14329_ (.B1(_05169_),
    .Y(_05244_),
    .A1(net206),
    .A2(net205));
 sg13g2_nand2_1 _14330_ (.Y(_05245_),
    .A(_05243_),
    .B(_05244_));
 sg13g2_xnor2_1 _14331_ (.Y(_05246_),
    .A(_05222_),
    .B(_05245_));
 sg13g2_nor2b_1 _14332_ (.A(_05242_),
    .B_N(_05246_),
    .Y(_05247_));
 sg13g2_nor2b_1 _14333_ (.A(_05246_),
    .B_N(_05242_),
    .Y(_05248_));
 sg13g2_o21ai_1 _14334_ (.B1(net112),
    .Y(_05249_),
    .A1(_05247_),
    .A2(_05248_));
 sg13g2_o21ai_1 _14335_ (.B1(_05249_),
    .Y(_00065_),
    .A1(net110),
    .A2(_05241_));
 sg13g2_nor2_1 _14336_ (.A(_05231_),
    .B(_05204_),
    .Y(_05250_));
 sg13g2_inv_1 _14337_ (.Y(_05251_),
    .A(_05250_));
 sg13g2_nor2_1 _14338_ (.A(_05251_),
    .B(_05213_),
    .Y(_05252_));
 sg13g2_nand3_1 _14339_ (.B(_05151_),
    .C(_05252_),
    .A(_05149_),
    .Y(_05253_));
 sg13g2_inv_1 _14340_ (.Y(_05254_),
    .A(_05211_));
 sg13g2_nor2_1 _14341_ (.A(_05231_),
    .B(_05202_),
    .Y(_05255_));
 sg13g2_a21oi_1 _14342_ (.A1(_05254_),
    .A2(_05250_),
    .Y(_05256_),
    .B1(_05255_));
 sg13g2_nand2_1 _14343_ (.Y(_05257_),
    .A(_05253_),
    .B(_05256_));
 sg13g2_inv_1 _14344_ (.Y(_05258_),
    .A(_01917_));
 sg13g2_inv_1 _14345_ (.Y(_05259_),
    .A(_05155_));
 sg13g2_nand2_1 _14346_ (.Y(_05260_),
    .A(_05259_),
    .B(_05230_));
 sg13g2_xnor2_1 _14347_ (.Y(_05261_),
    .A(_05258_),
    .B(_05260_));
 sg13g2_nand2_1 _14348_ (.Y(_05262_),
    .A(_05257_),
    .B(_05261_));
 sg13g2_inv_1 _14349_ (.Y(_05263_),
    .A(_05261_));
 sg13g2_nand3_1 _14350_ (.B(_05256_),
    .C(_05263_),
    .A(_05253_),
    .Y(_05264_));
 sg13g2_nand2_1 _14351_ (.Y(_05265_),
    .A(_05262_),
    .B(_05264_));
 sg13g2_nand2_1 _14352_ (.Y(_05266_),
    .A(_05265_),
    .B(net121));
 sg13g2_nand2b_1 _14353_ (.Y(_05267_),
    .B(_05245_),
    .A_N(_00181_));
 sg13g2_nand2_1 _14354_ (.Y(_05268_),
    .A(_05247_),
    .B(_05267_));
 sg13g2_o21ai_1 _14355_ (.B1(_05268_),
    .Y(_05269_),
    .A1(_05222_),
    .A2(_05267_));
 sg13g2_nand2_1 _14356_ (.Y(_05270_),
    .A(_05269_),
    .B(net111));
 sg13g2_nand2_1 _14357_ (.Y(_00066_),
    .A(_05266_),
    .B(_05270_));
 sg13g2_nand2_1 _14358_ (.Y(_05271_),
    .A(_05263_),
    .B(_05232_));
 sg13g2_nor2_1 _14359_ (.A(_05271_),
    .B(_05237_),
    .Y(_05272_));
 sg13g2_nand2_1 _14360_ (.Y(_05273_),
    .A(_05189_),
    .B(_05272_));
 sg13g2_nand2_1 _14361_ (.Y(_05274_),
    .A(_05259_),
    .B(_05258_));
 sg13g2_nor2_1 _14362_ (.A(_05230_),
    .B(_05274_),
    .Y(_05275_));
 sg13g2_nor2_1 _14363_ (.A(_05271_),
    .B(_05235_),
    .Y(_05276_));
 sg13g2_nor2_1 _14364_ (.A(_05275_),
    .B(_05276_),
    .Y(_05277_));
 sg13g2_nand2_1 _14365_ (.Y(_05278_),
    .A(_05273_),
    .B(_05277_));
 sg13g2_inv_1 _14366_ (.Y(_05279_),
    .A(_00182_));
 sg13g2_nor2_1 _14367_ (.A(_01917_),
    .B(_05279_),
    .Y(_05280_));
 sg13g2_a22oi_1 _14368_ (.Y(_05281_),
    .B1(_05279_),
    .B2(_05274_),
    .A2(_05280_),
    .A1(_05259_));
 sg13g2_buf_1 _14369_ (.A(_05281_),
    .X(_05282_));
 sg13g2_inv_1 _14370_ (.Y(_05283_),
    .A(_05282_));
 sg13g2_nand2_1 _14371_ (.Y(_05284_),
    .A(_05278_),
    .B(_05283_));
 sg13g2_nand3_1 _14372_ (.B(_05277_),
    .C(_05282_),
    .A(_05273_),
    .Y(_05285_));
 sg13g2_nand3_1 _14373_ (.B(_05285_),
    .C(net123),
    .A(_05284_),
    .Y(_05286_));
 sg13g2_nand2_1 _14374_ (.Y(_00067_),
    .A(_05286_),
    .B(_05270_));
 sg13g2_nand2_1 _14375_ (.Y(_05287_),
    .A(_05283_),
    .B(_05263_));
 sg13g2_nor2_1 _14376_ (.A(_05287_),
    .B(_05251_),
    .Y(_05288_));
 sg13g2_nand3_1 _14377_ (.B(_05214_),
    .C(_05288_),
    .A(_05079_),
    .Y(_05289_));
 sg13g2_inv_1 _14378_ (.Y(_05290_),
    .A(_05255_));
 sg13g2_nor2_1 _14379_ (.A(_05279_),
    .B(_05155_),
    .Y(_05291_));
 sg13g2_o21ai_1 _14380_ (.B1(_05291_),
    .Y(_05292_),
    .A1(_01917_),
    .A2(_01921_));
 sg13g2_o21ai_1 _14381_ (.B1(_05292_),
    .Y(_05293_),
    .A1(_05287_),
    .A2(_05290_));
 sg13g2_a21oi_1 _14382_ (.A1(_05212_),
    .A2(_05288_),
    .Y(_05294_),
    .B1(_05293_));
 sg13g2_nand2_1 _14383_ (.Y(_05295_),
    .A(_05289_),
    .B(_05294_));
 sg13g2_inv_1 _14384_ (.Y(_05296_),
    .A(_00183_));
 sg13g2_nor2_1 _14385_ (.A(_05296_),
    .B(_05155_),
    .Y(_05297_));
 sg13g2_inv_1 _14386_ (.Y(_05298_),
    .A(_05291_));
 sg13g2_a22oi_1 _14387_ (.Y(_05299_),
    .B1(_05296_),
    .B2(_05298_),
    .A2(_00182_),
    .A1(_05297_));
 sg13g2_nand2_1 _14388_ (.Y(_05300_),
    .A(_05295_),
    .B(_05299_));
 sg13g2_inv_1 _14389_ (.Y(_05301_),
    .A(_05299_));
 sg13g2_nand3_1 _14390_ (.B(_05294_),
    .C(_05301_),
    .A(_05289_),
    .Y(_05302_));
 sg13g2_nand2_1 _14391_ (.Y(_05303_),
    .A(_05300_),
    .B(_05302_));
 sg13g2_nand2_1 _14392_ (.Y(_05304_),
    .A(_05303_),
    .B(net121));
 sg13g2_nand2_1 _14393_ (.Y(_00068_),
    .A(_05304_),
    .B(_05270_));
 sg13g2_nor3_1 _14394_ (.A(_05282_),
    .B(_05299_),
    .C(_05271_),
    .Y(_05305_));
 sg13g2_nand4_1 _14395_ (.B(_05115_),
    .C(_05238_),
    .A(_05112_),
    .Y(_05306_),
    .D(_05305_));
 sg13g2_inv_1 _14396_ (.Y(_05307_),
    .A(_05297_));
 sg13g2_nand3_1 _14397_ (.B(_05283_),
    .C(_05275_),
    .A(_05301_),
    .Y(_05308_));
 sg13g2_o21ai_1 _14398_ (.B1(_05308_),
    .Y(_05309_),
    .A1(_05280_),
    .A2(_05307_));
 sg13g2_a21oi_1 _14399_ (.A1(_05236_),
    .A2(_05305_),
    .Y(_05310_),
    .B1(_05309_));
 sg13g2_nand2_1 _14400_ (.Y(_05311_),
    .A(_05306_),
    .B(_05310_));
 sg13g2_xnor2_1 _14401_ (.Y(_05312_),
    .A(_03228_),
    .B(_05297_));
 sg13g2_nand2_1 _14402_ (.Y(_05313_),
    .A(_05311_),
    .B(_05312_));
 sg13g2_inv_1 _14403_ (.Y(_05314_),
    .A(_05312_));
 sg13g2_nand3_1 _14404_ (.B(_05310_),
    .C(_05314_),
    .A(_05306_),
    .Y(_05315_));
 sg13g2_nand3_1 _14405_ (.B(_05315_),
    .C(net123),
    .A(_05313_),
    .Y(_05316_));
 sg13g2_nand2_1 _14406_ (.Y(_00069_),
    .A(_05316_),
    .B(_05270_));
 sg13g2_xor2_1 _14407_ (.B(net32),
    .A(\vgadonut.donut.donuthit.rz[14] ),
    .X(_05317_));
 sg13g2_buf_2 _14408_ (.A(_05317_),
    .X(_05318_));
 sg13g2_inv_2 _14409_ (.Y(_05319_),
    .A(_05318_));
 sg13g2_nand2_1 _14410_ (.Y(_05320_),
    .A(_04166_),
    .B(_05319_));
 sg13g2_xor2_1 _14411_ (.B(net35),
    .A(\vgadonut.donut.donuthit.rz[9] ),
    .X(_05321_));
 sg13g2_inv_1 _14412_ (.Y(_05322_),
    .A(_05321_));
 sg13g2_nand2_1 _14413_ (.Y(_05323_),
    .A(_04280_),
    .B(_05322_));
 sg13g2_nand2_1 _14414_ (.Y(_05324_),
    .A(_05320_),
    .B(_05323_));
 sg13g2_xor2_1 _14415_ (.B(net36),
    .A(\vgadonut.donut.donuthit.rz[13] ),
    .X(_05325_));
 sg13g2_buf_1 _14416_ (.A(_05325_),
    .X(_05326_));
 sg13g2_xnor2_1 _14417_ (.Y(_05327_),
    .A(\vgadonut.donut.donuthit.rz[8] ),
    .B(net33));
 sg13g2_nand2_1 _14418_ (.Y(_05328_),
    .A(net16),
    .B(_05327_));
 sg13g2_o21ai_1 _14419_ (.B1(_05328_),
    .Y(_05329_),
    .A1(_05326_),
    .A2(_04079_));
 sg13g2_nor2_1 _14420_ (.A(_05324_),
    .B(_05329_),
    .Y(_05330_));
 sg13g2_xor2_1 _14421_ (.B(net35),
    .A(\vgadonut.donut.donuthit.rz[11] ),
    .X(_05331_));
 sg13g2_inv_2 _14422_ (.Y(_05332_),
    .A(_05331_));
 sg13g2_nand2_1 _14423_ (.Y(_05333_),
    .A(_04171_),
    .B(_05332_));
 sg13g2_xnor2_1 _14424_ (.Y(_05334_),
    .A(\vgadonut.donut.donuthit.rz[7] ),
    .B(net33));
 sg13g2_nor2b_1 _14425_ (.A(_04107_),
    .B_N(_05334_),
    .Y(_05335_));
 sg13g2_xnor2_1 _14426_ (.Y(_05336_),
    .A(\vgadonut.donut.donuthit.rz[6] ),
    .B(net32));
 sg13g2_inv_1 _14427_ (.Y(_05337_),
    .A(_05336_));
 sg13g2_nand2_1 _14428_ (.Y(_05338_),
    .A(_04008_),
    .B(\vgadonut.donut.donuthit.rz[5] ));
 sg13g2_o21ai_1 _14429_ (.B1(_05338_),
    .Y(_05339_),
    .A1(\vgadonut.donut.donuthit.rz[5] ),
    .A2(_04794_));
 sg13g2_o21ai_1 _14430_ (.B1(_05339_),
    .Y(_05340_),
    .A1(_05337_),
    .A2(_04336_));
 sg13g2_nor2_1 _14431_ (.A(_05335_),
    .B(_05340_),
    .Y(_05341_));
 sg13g2_nand2_1 _14432_ (.Y(_05342_),
    .A(_05333_),
    .B(_05341_));
 sg13g2_xnor2_1 _14433_ (.Y(_05343_),
    .A(\vgadonut.donut.donuthit.rz[12] ),
    .B(net36));
 sg13g2_buf_1 _14434_ (.A(_05343_),
    .X(_05344_));
 sg13g2_inv_1 _14435_ (.Y(_05345_),
    .A(_05344_));
 sg13g2_xnor2_1 _14436_ (.Y(_05346_),
    .A(\vgadonut.donut.donuthit.rz[10] ),
    .B(net33));
 sg13g2_buf_2 _14437_ (.A(_05346_),
    .X(_05347_));
 sg13g2_nand2_1 _14438_ (.Y(_05348_),
    .A(_04332_),
    .B(_05347_));
 sg13g2_o21ai_1 _14439_ (.B1(_05348_),
    .Y(_05349_),
    .A1(_04059_),
    .A2(_05345_));
 sg13g2_nor2_1 _14440_ (.A(_05342_),
    .B(_05349_),
    .Y(_05350_));
 sg13g2_nand2_1 _14441_ (.Y(_05351_),
    .A(_05330_),
    .B(_05350_));
 sg13g2_nand2_1 _14442_ (.Y(_05352_),
    .A(_05351_),
    .B(_04325_));
 sg13g2_xor2_1 _14443_ (.B(net35),
    .A(\vgadonut.donut.donuthit.rz[15] ),
    .X(_05353_));
 sg13g2_inv_2 _14444_ (.Y(_05354_),
    .A(_05353_));
 sg13g2_buf_8 _14445_ (.A(_05354_),
    .X(_05355_));
 sg13g2_nand2_1 _14446_ (.Y(_05356_),
    .A(net29),
    .B(_05327_));
 sg13g2_nand2_1 _14447_ (.Y(_05357_),
    .A(_04391_),
    .B(_05334_));
 sg13g2_nand2_1 _14448_ (.Y(_05358_),
    .A(_05356_),
    .B(_05357_));
 sg13g2_nor2_1 _14449_ (.A(_05321_),
    .B(_04107_),
    .Y(_05359_));
 sg13g2_nor2_1 _14450_ (.A(_05358_),
    .B(_05359_),
    .Y(_05360_));
 sg13g2_nand2_1 _14451_ (.Y(_05361_),
    .A(_04271_),
    .B(_05347_));
 sg13g2_nand2_1 _14452_ (.Y(_05362_),
    .A(_05360_),
    .B(_05361_));
 sg13g2_a21oi_1 _14453_ (.A1(_04091_),
    .A2(net19),
    .Y(_05363_),
    .B1(_05362_));
 sg13g2_nand2_1 _14454_ (.Y(_05364_),
    .A(_04169_),
    .B(_05319_));
 sg13g2_nand2_1 _14455_ (.Y(_05365_),
    .A(net17),
    .B(_05344_));
 sg13g2_nand2_1 _14456_ (.Y(_05366_),
    .A(_05364_),
    .B(_05365_));
 sg13g2_inv_1 _14457_ (.Y(_05367_),
    .A(_05326_));
 sg13g2_nand2_1 _14458_ (.Y(_05368_),
    .A(_04171_),
    .B(_05367_));
 sg13g2_nand2_1 _14459_ (.Y(_05369_),
    .A(_04280_),
    .B(_05332_));
 sg13g2_nand2_1 _14460_ (.Y(_05370_),
    .A(_05368_),
    .B(_05369_));
 sg13g2_nor2_1 _14461_ (.A(_05366_),
    .B(_05370_),
    .Y(_05371_));
 sg13g2_nand2_1 _14462_ (.Y(_05372_),
    .A(_05363_),
    .B(_05371_));
 sg13g2_nand2_1 _14463_ (.Y(_05373_),
    .A(_05372_),
    .B(net14));
 sg13g2_nand2_1 _14464_ (.Y(_05374_),
    .A(_05352_),
    .B(_05373_));
 sg13g2_nand3_1 _14465_ (.B(_05372_),
    .C(net11),
    .A(_05351_),
    .Y(_05375_));
 sg13g2_buf_1 _14466_ (.A(_05375_),
    .X(_05376_));
 sg13g2_a21oi_1 _14467_ (.A1(_05374_),
    .A2(_05376_),
    .Y(_05377_),
    .B1(_03008_));
 sg13g2_nand3_1 _14468_ (.B(_05376_),
    .C(_03008_),
    .A(_05374_),
    .Y(_05378_));
 sg13g2_nand3b_1 _14469_ (.B(net126),
    .C(_05378_),
    .Y(_05379_),
    .A_N(_05377_));
 sg13g2_buf_2 _14470_ (.A(\vgadonut.donut.cAcB[3] ),
    .X(_05380_));
 sg13g2_buf_1 _14471_ (.A(\vgadonut.donut.cAcB[5] ),
    .X(_05381_));
 sg13g2_nor2_1 _14472_ (.A(_05380_),
    .B(net237),
    .Y(_05382_));
 sg13g2_inv_1 _14473_ (.Y(_05383_),
    .A(_05382_));
 sg13g2_buf_1 _14474_ (.A(\vgadonut.donut.cAcB[4] ),
    .X(_05384_));
 sg13g2_buf_1 _14475_ (.A(\vgadonut.donut.cAcB[6] ),
    .X(_05385_));
 sg13g2_nor2_1 _14476_ (.A(net236),
    .B(net235),
    .Y(_05386_));
 sg13g2_nand2_1 _14477_ (.Y(_05387_),
    .A(net236),
    .B(net235));
 sg13g2_nor2b_1 _14478_ (.A(_05386_),
    .B_N(_05387_),
    .Y(_05388_));
 sg13g2_xnor2_1 _14479_ (.Y(_05389_),
    .A(_05383_),
    .B(_05388_));
 sg13g2_buf_2 _14480_ (.A(\vgadonut.donut.cAcB[2] ),
    .X(_05390_));
 sg13g2_nor2_1 _14481_ (.A(_05390_),
    .B(net236),
    .Y(_05391_));
 sg13g2_inv_1 _14482_ (.Y(_05392_),
    .A(_05391_));
 sg13g2_xor2_1 _14483_ (.B(net237),
    .A(_05380_),
    .X(_05393_));
 sg13g2_inv_1 _14484_ (.Y(_05394_),
    .A(_05393_));
 sg13g2_nor2_1 _14485_ (.A(_05392_),
    .B(_05394_),
    .Y(_05395_));
 sg13g2_buf_2 _14486_ (.A(\vgadonut.donut.cAcB[1] ),
    .X(_05396_));
 sg13g2_nand2_1 _14487_ (.Y(_05397_),
    .A(_05396_),
    .B(_05380_));
 sg13g2_xnor2_1 _14488_ (.Y(_05398_),
    .A(_05390_),
    .B(net236));
 sg13g2_xnor2_1 _14489_ (.Y(_05399_),
    .A(_05397_),
    .B(_05398_));
 sg13g2_inv_1 _14490_ (.Y(_05400_),
    .A(_05396_));
 sg13g2_inv_1 _14491_ (.Y(_05401_),
    .A(_05380_));
 sg13g2_nand2_1 _14492_ (.Y(_05402_),
    .A(_05400_),
    .B(_05401_));
 sg13g2_buf_2 _14493_ (.A(\vgadonut.donut.cAcB[0] ),
    .X(_05403_));
 sg13g2_inv_1 _14494_ (.Y(_05404_),
    .A(_05403_));
 sg13g2_inv_1 _14495_ (.Y(_05405_),
    .A(_05390_));
 sg13g2_nand2_1 _14496_ (.Y(_05406_),
    .A(_05404_),
    .B(_05405_));
 sg13g2_a21oi_1 _14497_ (.A1(_05402_),
    .A2(_05397_),
    .Y(_05407_),
    .B1(_05406_));
 sg13g2_nor2b_1 _14498_ (.A(_05398_),
    .B_N(_05397_),
    .Y(_05408_));
 sg13g2_a21oi_1 _14499_ (.A1(_05399_),
    .A2(_05407_),
    .Y(_05409_),
    .B1(_05408_));
 sg13g2_inv_1 _14500_ (.Y(_05410_),
    .A(_05409_));
 sg13g2_nand2_1 _14501_ (.Y(_05411_),
    .A(_05394_),
    .B(_05392_));
 sg13g2_o21ai_1 _14502_ (.B1(_05411_),
    .Y(_05412_),
    .A1(_05395_),
    .A2(_05410_));
 sg13g2_xnor2_1 _14503_ (.Y(_05413_),
    .A(_05389_),
    .B(_05412_));
 sg13g2_inv_1 _14504_ (.Y(_05414_),
    .A(_05413_));
 sg13g2_inv_1 _14505_ (.Y(_05415_),
    .A(\vgadonut.donut.donuthit.rzin[5] ));
 sg13g2_a21oi_1 _14506_ (.A1(_05414_),
    .A2(_05415_),
    .Y(_05416_),
    .B1(_04305_));
 sg13g2_nor2_1 _14507_ (.A(_05415_),
    .B(_05414_),
    .Y(_05417_));
 sg13g2_inv_1 _14508_ (.Y(_05418_),
    .A(_05417_));
 sg13g2_nand2_1 _14509_ (.Y(_05419_),
    .A(_05416_),
    .B(_05418_));
 sg13g2_nand2_1 _14510_ (.Y(_00079_),
    .A(_05379_),
    .B(_05419_));
 sg13g2_inv_1 _14511_ (.Y(_05420_),
    .A(\vgadonut.donut.donuthit.rzin[6] ));
 sg13g2_buf_1 _14512_ (.A(\vgadonut.donut.cAcB[7] ),
    .X(_05421_));
 sg13g2_xor2_1 _14513_ (.B(net234),
    .A(net237),
    .X(_05422_));
 sg13g2_xor2_1 _14514_ (.B(_05422_),
    .A(_05386_),
    .X(_05423_));
 sg13g2_inv_1 _14515_ (.Y(_05424_),
    .A(_05423_));
 sg13g2_inv_1 _14516_ (.Y(_05425_),
    .A(_05395_));
 sg13g2_and3_1 _14517_ (.X(_05426_),
    .A(_05389_),
    .B(_05411_),
    .C(_05425_));
 sg13g2_o21ai_1 _14518_ (.B1(_05388_),
    .Y(_05427_),
    .A1(_05382_),
    .A2(_05395_));
 sg13g2_inv_1 _14519_ (.Y(_05428_),
    .A(_05427_));
 sg13g2_a21oi_1 _14520_ (.A1(_05426_),
    .A2(_05410_),
    .Y(_05429_),
    .B1(_05428_));
 sg13g2_xnor2_1 _14521_ (.Y(_05430_),
    .A(_05424_),
    .B(_05429_));
 sg13g2_nor2_1 _14522_ (.A(_05420_),
    .B(_05430_),
    .Y(_05431_));
 sg13g2_nand2_1 _14523_ (.Y(_05432_),
    .A(_05430_),
    .B(_05420_));
 sg13g2_nor2b_1 _14524_ (.A(_05431_),
    .B_N(_05432_),
    .Y(_05433_));
 sg13g2_nor2b_1 _14525_ (.A(_05418_),
    .B_N(_05433_),
    .Y(_05434_));
 sg13g2_o21ai_1 _14526_ (.B1(net112),
    .Y(_05435_),
    .A1(_05417_),
    .A2(_05433_));
 sg13g2_nand2_1 _14527_ (.Y(_05436_),
    .A(_05374_),
    .B(\vgadonut.donut.donuthit.cordicxz.xin[0] ));
 sg13g2_nand2_1 _14528_ (.Y(_05437_),
    .A(_05436_),
    .B(_05376_));
 sg13g2_nand2_1 _14529_ (.Y(_05438_),
    .A(_04091_),
    .B(net19));
 sg13g2_a22oi_1 _14530_ (.Y(_05439_),
    .B1(_05322_),
    .B2(net23),
    .A2(_05327_),
    .A1(net31));
 sg13g2_nand2_1 _14531_ (.Y(_05440_),
    .A(net28),
    .B(_05347_));
 sg13g2_nand2_1 _14532_ (.Y(_05441_),
    .A(_05439_),
    .B(_05440_));
 sg13g2_nor2_1 _14533_ (.A(_05318_),
    .B(net18),
    .Y(_05442_));
 sg13g2_nor2_1 _14534_ (.A(_05441_),
    .B(_05442_),
    .Y(_05443_));
 sg13g2_nand2_1 _14535_ (.Y(_05444_),
    .A(_05438_),
    .B(_05443_));
 sg13g2_nand3_1 _14536_ (.B(_04057_),
    .C(_05354_),
    .A(net26),
    .Y(_05445_));
 sg13g2_nand4_1 _14537_ (.B(_04124_),
    .C(_04042_),
    .A(net30),
    .Y(_05446_),
    .D(_05367_));
 sg13g2_nand2_1 _14538_ (.Y(_05447_),
    .A(_05445_),
    .B(_05446_));
 sg13g2_nand2_1 _14539_ (.Y(_05448_),
    .A(_04113_),
    .B(_05332_));
 sg13g2_nand3_1 _14540_ (.B(_04033_),
    .C(_05344_),
    .A(net26),
    .Y(_05449_));
 sg13g2_nand2_1 _14541_ (.Y(_05450_),
    .A(_05448_),
    .B(_05449_));
 sg13g2_nor2_1 _14542_ (.A(_05447_),
    .B(_05450_),
    .Y(_05451_));
 sg13g2_nor2b_1 _14543_ (.A(_05444_),
    .B_N(_05451_),
    .Y(_05452_));
 sg13g2_nor2_1 _14544_ (.A(_05321_),
    .B(net24),
    .Y(_05453_));
 sg13g2_nor3_1 _14545_ (.A(_04126_),
    .B(_05353_),
    .C(_04131_),
    .Y(_05454_));
 sg13g2_nor2_1 _14546_ (.A(_05453_),
    .B(_05454_),
    .Y(_05455_));
 sg13g2_nor2_1 _14547_ (.A(_05331_),
    .B(_04044_),
    .Y(_05456_));
 sg13g2_nor2_1 _14548_ (.A(_05337_),
    .B(_04026_),
    .Y(_05457_));
 sg13g2_a21oi_1 _14549_ (.A1(_04520_),
    .A2(_05334_),
    .Y(_05458_),
    .B1(_05457_));
 sg13g2_nand2_1 _14550_ (.Y(_05459_),
    .A(net22),
    .B(_05327_));
 sg13g2_nand2_1 _14551_ (.Y(_05460_),
    .A(_05458_),
    .B(_05459_));
 sg13g2_nor2_1 _14552_ (.A(_05456_),
    .B(_05460_),
    .Y(_05461_));
 sg13g2_nand2_1 _14553_ (.Y(_05462_),
    .A(_05455_),
    .B(_05461_));
 sg13g2_nor2_1 _14554_ (.A(_05326_),
    .B(_04059_),
    .Y(_05463_));
 sg13g2_nor3_1 _14555_ (.A(_04111_),
    .B(_05318_),
    .C(_04156_),
    .Y(_05464_));
 sg13g2_nor2_1 _14556_ (.A(_05463_),
    .B(_05464_),
    .Y(_05465_));
 sg13g2_nor2b_1 _14557_ (.A(_04153_),
    .B_N(_05347_),
    .Y(_05466_));
 sg13g2_nor2_1 _14558_ (.A(_05345_),
    .B(net18),
    .Y(_05467_));
 sg13g2_nor2_1 _14559_ (.A(_05466_),
    .B(_05467_),
    .Y(_05468_));
 sg13g2_nand2_1 _14560_ (.Y(_05469_),
    .A(_05465_),
    .B(_05468_));
 sg13g2_nor2_1 _14561_ (.A(_05462_),
    .B(_05469_),
    .Y(_05470_));
 sg13g2_a21oi_1 _14562_ (.A1(_05452_),
    .A2(_05470_),
    .Y(_05471_),
    .B1(_04266_));
 sg13g2_nand3_1 _14563_ (.B(_05438_),
    .C(_05443_),
    .A(_05451_),
    .Y(_05472_));
 sg13g2_buf_1 _14564_ (.A(_05472_),
    .X(_05473_));
 sg13g2_nand3_1 _14565_ (.B(_04022_),
    .C(_05344_),
    .A(_04173_),
    .Y(_05474_));
 sg13g2_nand2_1 _14566_ (.Y(_05475_),
    .A(_04280_),
    .B(_05347_));
 sg13g2_nand2_1 _14567_ (.Y(_05476_),
    .A(_05474_),
    .B(_05475_));
 sg13g2_nand2_1 _14568_ (.Y(_05477_),
    .A(_04167_),
    .B(_05319_));
 sg13g2_inv_1 _14569_ (.Y(_05478_),
    .A(_05463_));
 sg13g2_nand2_1 _14570_ (.Y(_05479_),
    .A(_05477_),
    .B(_05478_));
 sg13g2_nor2_1 _14571_ (.A(_05476_),
    .B(_05479_),
    .Y(_05480_));
 sg13g2_nand2_1 _14572_ (.Y(_05481_),
    .A(_04138_),
    .B(_05334_));
 sg13g2_nand2b_1 _14573_ (.Y(_05482_),
    .B(_05481_),
    .A_N(_05457_));
 sg13g2_nor2b_1 _14574_ (.A(_04107_),
    .B_N(_05327_),
    .Y(_05483_));
 sg13g2_nor2_1 _14575_ (.A(_05482_),
    .B(_05483_),
    .Y(_05484_));
 sg13g2_nand2_1 _14576_ (.Y(_05485_),
    .A(net17),
    .B(_05332_));
 sg13g2_nand2_1 _14577_ (.Y(_05486_),
    .A(_05484_),
    .B(_05485_));
 sg13g2_nand2_1 _14578_ (.Y(_05487_),
    .A(_04166_),
    .B(net19));
 sg13g2_nand2_1 _14579_ (.Y(_05488_),
    .A(_04271_),
    .B(_05322_));
 sg13g2_nand2_1 _14580_ (.Y(_05489_),
    .A(_05487_),
    .B(_05488_));
 sg13g2_nor2_1 _14581_ (.A(_05486_),
    .B(_05489_),
    .Y(_05490_));
 sg13g2_nand2_1 _14582_ (.Y(_05491_),
    .A(_05480_),
    .B(_05490_));
 sg13g2_nand3_1 _14583_ (.B(_05491_),
    .C(_04325_),
    .A(_05473_),
    .Y(_05492_));
 sg13g2_buf_1 _14584_ (.A(_05492_),
    .X(_05493_));
 sg13g2_nand2_1 _14585_ (.Y(_05494_),
    .A(_05471_),
    .B(_05493_));
 sg13g2_nand2_1 _14586_ (.Y(_05495_),
    .A(_05494_),
    .B(_03001_));
 sg13g2_nand3_1 _14587_ (.B(_05493_),
    .C(_03000_),
    .A(_05471_),
    .Y(_05496_));
 sg13g2_nand2_1 _14588_ (.Y(_05497_),
    .A(_05495_),
    .B(_05496_));
 sg13g2_nand2b_1 _14589_ (.Y(_05498_),
    .B(_05497_),
    .A_N(_05437_));
 sg13g2_nand3_1 _14590_ (.B(_05495_),
    .C(_05496_),
    .A(_05437_),
    .Y(_05499_));
 sg13g2_buf_1 _14591_ (.A(_05499_),
    .X(_05500_));
 sg13g2_nand3_1 _14592_ (.B(_05500_),
    .C(net125),
    .A(_05498_),
    .Y(_05501_));
 sg13g2_o21ai_1 _14593_ (.B1(_05501_),
    .Y(_00086_),
    .A1(_05434_),
    .A2(_05435_));
 sg13g2_buf_1 _14594_ (.A(\vgadonut.donut.donuthit.rzin[7] ),
    .X(_05502_));
 sg13g2_inv_1 _14595_ (.Y(_05503_),
    .A(_05502_));
 sg13g2_nor2_1 _14596_ (.A(net237),
    .B(net234),
    .Y(_05504_));
 sg13g2_buf_1 _14597_ (.A(\vgadonut.donut.cAcB[8] ),
    .X(_05505_));
 sg13g2_xor2_1 _14598_ (.B(net233),
    .A(net235),
    .X(_05506_));
 sg13g2_xor2_1 _14599_ (.B(_05506_),
    .A(_05504_),
    .X(_05507_));
 sg13g2_nand2_1 _14600_ (.Y(_05508_),
    .A(_05389_),
    .B(_05423_));
 sg13g2_nor2b_1 _14601_ (.A(_05383_),
    .B_N(_05388_),
    .Y(_05509_));
 sg13g2_nand2_1 _14602_ (.Y(_05510_),
    .A(_05422_),
    .B(_05386_));
 sg13g2_inv_1 _14603_ (.Y(_05511_),
    .A(_05510_));
 sg13g2_a21oi_1 _14604_ (.A1(_05509_),
    .A2(net234),
    .Y(_05512_),
    .B1(_05511_));
 sg13g2_o21ai_1 _14605_ (.B1(_05512_),
    .Y(_05513_),
    .A1(_05508_),
    .A2(_05412_));
 sg13g2_xnor2_1 _14606_ (.Y(_05514_),
    .A(_05507_),
    .B(_05513_));
 sg13g2_nor2_1 _14607_ (.A(_05503_),
    .B(_05514_),
    .Y(_05515_));
 sg13g2_nand2_1 _14608_ (.Y(_05516_),
    .A(_05514_),
    .B(_05503_));
 sg13g2_nor2b_1 _14609_ (.A(_05515_),
    .B_N(_05516_),
    .Y(_05517_));
 sg13g2_nor2_1 _14610_ (.A(_05431_),
    .B(_05434_),
    .Y(_05518_));
 sg13g2_xor2_1 _14611_ (.B(_05518_),
    .A(_05517_),
    .X(_05519_));
 sg13g2_nor2_1 _14612_ (.A(_05345_),
    .B(net24),
    .Y(_05520_));
 sg13g2_a22oi_1 _14613_ (.Y(_05521_),
    .B1(_05347_),
    .B2(net29),
    .A2(_05322_),
    .A1(net31));
 sg13g2_nand2_1 _14614_ (.Y(_05522_),
    .A(net28),
    .B(_05332_));
 sg13g2_nand2_1 _14615_ (.Y(_05523_),
    .A(_05521_),
    .B(_05522_));
 sg13g2_nor2_1 _14616_ (.A(_05520_),
    .B(_05523_),
    .Y(_05524_));
 sg13g2_nor2_1 _14617_ (.A(_05326_),
    .B(_04153_),
    .Y(_05525_));
 sg13g2_nor2_1 _14618_ (.A(_05318_),
    .B(_04044_),
    .Y(_05526_));
 sg13g2_nor2_1 _14619_ (.A(_05525_),
    .B(_05526_),
    .Y(_05527_));
 sg13g2_nand2_1 _14620_ (.Y(_05528_),
    .A(_05524_),
    .B(_05527_));
 sg13g2_a21oi_1 _14621_ (.A1(_04168_),
    .A2(_04172_),
    .Y(_05529_),
    .B1(_05353_));
 sg13g2_a21oi_1 _14622_ (.A1(_04176_),
    .A2(_05528_),
    .Y(_05530_),
    .B1(_05529_));
 sg13g2_nand2_1 _14623_ (.Y(_05531_),
    .A(_05373_),
    .B(_05530_));
 sg13g2_nand2_1 _14624_ (.Y(_05532_),
    .A(_04175_),
    .B(_05528_));
 sg13g2_nand2_1 _14625_ (.Y(_05533_),
    .A(_04327_),
    .B(net19));
 sg13g2_nand2_1 _14626_ (.Y(_05534_),
    .A(_05532_),
    .B(_05533_));
 sg13g2_nand2_1 _14627_ (.Y(_05535_),
    .A(_05534_),
    .B(_05372_));
 sg13g2_nand2_1 _14628_ (.Y(_05536_),
    .A(_05531_),
    .B(_05535_));
 sg13g2_xnor2_1 _14629_ (.Y(_05537_),
    .A(_02994_),
    .B(_05536_));
 sg13g2_inv_1 _14630_ (.Y(_05538_),
    .A(_05493_));
 sg13g2_a21oi_1 _14631_ (.A1(_05471_),
    .A2(_03000_),
    .Y(_05539_),
    .B1(_05538_));
 sg13g2_nor2b_1 _14632_ (.A(_05537_),
    .B_N(_05539_),
    .Y(_05540_));
 sg13g2_nand2b_1 _14633_ (.Y(_05541_),
    .B(_05537_),
    .A_N(_05539_));
 sg13g2_inv_2 _14634_ (.Y(_05542_),
    .A(_05541_));
 sg13g2_o21ai_1 _14635_ (.B1(_05500_),
    .Y(_05543_),
    .A1(_05540_),
    .A2(_05542_));
 sg13g2_nor2b_1 _14636_ (.A(_05497_),
    .B_N(_05437_),
    .Y(_05544_));
 sg13g2_nand2b_1 _14637_ (.Y(_05545_),
    .B(_05536_),
    .A_N(_02994_));
 sg13g2_nand3_1 _14638_ (.B(_05535_),
    .C(_02994_),
    .A(_05531_),
    .Y(_05546_));
 sg13g2_nand2_1 _14639_ (.Y(_05547_),
    .A(_05545_),
    .B(_05546_));
 sg13g2_nand2_1 _14640_ (.Y(_05548_),
    .A(_05547_),
    .B(_05539_));
 sg13g2_nand3_1 _14641_ (.B(_05544_),
    .C(_05548_),
    .A(_05541_),
    .Y(_05549_));
 sg13g2_nand3_1 _14642_ (.B(_04362_),
    .C(_05549_),
    .A(_05543_),
    .Y(_05550_));
 sg13g2_o21ai_1 _14643_ (.B1(_05550_),
    .Y(_00087_),
    .A1(net122),
    .A2(_05519_));
 sg13g2_buf_1 _14644_ (.A(\vgadonut.donut.donuthit.rzin[8] ),
    .X(_05551_));
 sg13g2_nor2_1 _14645_ (.A(net235),
    .B(net233),
    .Y(_05552_));
 sg13g2_buf_1 _14646_ (.A(\vgadonut.donut.cAcB[9] ),
    .X(_05553_));
 sg13g2_xor2_1 _14647_ (.B(net232),
    .A(net234),
    .X(_05554_));
 sg13g2_xor2_1 _14648_ (.B(_05554_),
    .A(_05552_),
    .X(_05555_));
 sg13g2_inv_1 _14649_ (.Y(_05556_),
    .A(_05429_));
 sg13g2_inv_1 _14650_ (.Y(_05557_),
    .A(_05507_));
 sg13g2_nor2_1 _14651_ (.A(_05424_),
    .B(_05557_),
    .Y(_05558_));
 sg13g2_nand2_1 _14652_ (.Y(_05559_),
    .A(_05506_),
    .B(_05504_));
 sg13g2_inv_1 _14653_ (.Y(_05560_),
    .A(_05559_));
 sg13g2_a21oi_1 _14654_ (.A1(_05511_),
    .A2(net233),
    .Y(_05561_),
    .B1(_05560_));
 sg13g2_inv_1 _14655_ (.Y(_05562_),
    .A(_05561_));
 sg13g2_a21oi_1 _14656_ (.A1(_05556_),
    .A2(_05558_),
    .Y(_05563_),
    .B1(_05562_));
 sg13g2_xnor2_1 _14657_ (.Y(_05564_),
    .A(_05555_),
    .B(_05563_));
 sg13g2_nor2_1 _14658_ (.A(_05551_),
    .B(_05564_),
    .Y(_05565_));
 sg13g2_nand2_1 _14659_ (.Y(_05566_),
    .A(_05564_),
    .B(_05551_));
 sg13g2_nand2b_1 _14660_ (.Y(_05567_),
    .B(_05566_),
    .A_N(_05565_));
 sg13g2_inv_1 _14661_ (.Y(_05568_),
    .A(_05518_));
 sg13g2_a21oi_1 _14662_ (.A1(_05568_),
    .A2(_05516_),
    .Y(_05569_),
    .B1(_05515_));
 sg13g2_xnor2_1 _14663_ (.Y(_05570_),
    .A(_05567_),
    .B(_05569_));
 sg13g2_o21ai_1 _14664_ (.B1(_05541_),
    .Y(_05571_),
    .A1(_05500_),
    .A2(_05540_));
 sg13g2_inv_1 _14665_ (.Y(_05572_),
    .A(_05571_));
 sg13g2_a22oi_1 _14666_ (.Y(_05573_),
    .B1(_02994_),
    .B2(_05531_),
    .A2(_05534_),
    .A1(_05372_));
 sg13g2_buf_1 _14667_ (.A(_05573_),
    .X(_05574_));
 sg13g2_nand2_1 _14668_ (.Y(_05575_),
    .A(net17),
    .B(_05355_));
 sg13g2_o21ai_1 _14669_ (.B1(_05575_),
    .Y(_05576_),
    .A1(_04153_),
    .A2(_05318_));
 sg13g2_nand2_1 _14670_ (.Y(_05577_),
    .A(net16),
    .B(_05367_));
 sg13g2_nand2_1 _14671_ (.Y(_05578_),
    .A(net22),
    .B(_05344_));
 sg13g2_a22oi_1 _14672_ (.Y(_05579_),
    .B1(_05332_),
    .B2(net23),
    .A2(_05347_),
    .A1(net31));
 sg13g2_nand3_1 _14673_ (.B(_05578_),
    .C(_05579_),
    .A(_05577_),
    .Y(_05580_));
 sg13g2_nor2_1 _14674_ (.A(_05576_),
    .B(_05580_),
    .Y(_05581_));
 sg13g2_nand2_1 _14675_ (.Y(_05582_),
    .A(_05581_),
    .B(_05533_));
 sg13g2_nand2_1 _14676_ (.Y(_05583_),
    .A(_05582_),
    .B(net14));
 sg13g2_nand2_1 _14677_ (.Y(_05584_),
    .A(_05473_),
    .B(net13));
 sg13g2_nand2_1 _14678_ (.Y(_05585_),
    .A(_05583_),
    .B(_05584_));
 sg13g2_nand3_1 _14679_ (.B(_05473_),
    .C(net13),
    .A(_05582_),
    .Y(_05586_));
 sg13g2_buf_1 _14680_ (.A(_05586_),
    .X(_05587_));
 sg13g2_nand2_1 _14681_ (.Y(_05588_),
    .A(_05585_),
    .B(_05587_));
 sg13g2_nand2_1 _14682_ (.Y(_05589_),
    .A(_05588_),
    .B(_02984_));
 sg13g2_nand3_1 _14683_ (.B(_05587_),
    .C(_02983_),
    .A(_05585_),
    .Y(_05590_));
 sg13g2_nand2_1 _14684_ (.Y(_05591_),
    .A(_05589_),
    .B(_05590_));
 sg13g2_xnor2_1 _14685_ (.Y(_05592_),
    .A(_05574_),
    .B(_05591_));
 sg13g2_a21oi_1 _14686_ (.A1(_05572_),
    .A2(_05592_),
    .Y(_05593_),
    .B1(_04407_));
 sg13g2_o21ai_1 _14687_ (.B1(_05593_),
    .Y(_05594_),
    .A1(_05572_),
    .A2(_05592_));
 sg13g2_o21ai_1 _14688_ (.B1(_05594_),
    .Y(_00088_),
    .A1(net122),
    .A2(_05570_));
 sg13g2_buf_1 _14689_ (.A(\vgadonut.donut.donuthit.rzin[9] ),
    .X(_05595_));
 sg13g2_nor2_1 _14690_ (.A(net234),
    .B(net232),
    .Y(_05596_));
 sg13g2_buf_1 _14691_ (.A(\vgadonut.donut.cAcB[10] ),
    .X(_05597_));
 sg13g2_buf_1 _14692_ (.A(_05597_),
    .X(_05598_));
 sg13g2_xor2_1 _14693_ (.B(net203),
    .A(net233),
    .X(_05599_));
 sg13g2_xor2_1 _14694_ (.B(_05599_),
    .A(_05596_),
    .X(_05600_));
 sg13g2_inv_1 _14695_ (.Y(_05601_),
    .A(_05555_));
 sg13g2_nor2_1 _14696_ (.A(_05557_),
    .B(_05601_),
    .Y(_05602_));
 sg13g2_nand2_1 _14697_ (.Y(_05603_),
    .A(_05554_),
    .B(_05552_));
 sg13g2_inv_1 _14698_ (.Y(_05604_),
    .A(_05603_));
 sg13g2_a21oi_1 _14699_ (.A1(_05560_),
    .A2(net232),
    .Y(_05605_),
    .B1(_05604_));
 sg13g2_inv_1 _14700_ (.Y(_05606_),
    .A(_05605_));
 sg13g2_a21oi_1 _14701_ (.A1(_05513_),
    .A2(_05602_),
    .Y(_05607_),
    .B1(_05606_));
 sg13g2_xnor2_1 _14702_ (.Y(_05608_),
    .A(_05600_),
    .B(_05607_));
 sg13g2_nor2_1 _14703_ (.A(_05595_),
    .B(_05608_),
    .Y(_05609_));
 sg13g2_nand2_1 _14704_ (.Y(_05610_),
    .A(_05608_),
    .B(_05595_));
 sg13g2_nor2b_1 _14705_ (.A(_05609_),
    .B_N(_05610_),
    .Y(_05611_));
 sg13g2_a21oi_1 _14706_ (.A1(_05569_),
    .A2(_05566_),
    .Y(_05612_),
    .B1(_05565_));
 sg13g2_xnor2_1 _14707_ (.Y(_05613_),
    .A(_05611_),
    .B(_05612_));
 sg13g2_inv_1 _14708_ (.Y(_05614_),
    .A(_05587_));
 sg13g2_a21oi_2 _14709_ (.B1(_05614_),
    .Y(_05615_),
    .A2(_02983_),
    .A1(_05585_));
 sg13g2_nor2_1 _14710_ (.A(_05326_),
    .B(_04107_),
    .Y(_05616_));
 sg13g2_nand2_1 _14711_ (.Y(_05617_),
    .A(net34),
    .B(_05332_));
 sg13g2_o21ai_1 _14712_ (.B1(_05617_),
    .Y(_05618_),
    .A1(_05345_),
    .A2(_04336_));
 sg13g2_nor2_1 _14713_ (.A(_05616_),
    .B(_05618_),
    .Y(_05619_));
 sg13g2_nand2_1 _14714_ (.Y(_05620_),
    .A(_04113_),
    .B(_05319_));
 sg13g2_nand2_1 _14715_ (.Y(_05621_),
    .A(_04431_),
    .B(_05354_));
 sg13g2_nand3_1 _14716_ (.B(_05620_),
    .C(_05621_),
    .A(_05619_),
    .Y(_05622_));
 sg13g2_nand2b_1 _14717_ (.Y(_05623_),
    .B(_05533_),
    .A_N(_05622_));
 sg13g2_nand2_1 _14718_ (.Y(_05624_),
    .A(_05623_),
    .B(net15));
 sg13g2_nand2_1 _14719_ (.Y(_05625_),
    .A(_05624_),
    .B(_05530_));
 sg13g2_nand2_1 _14720_ (.Y(_05626_),
    .A(_05534_),
    .B(_05623_));
 sg13g2_nand2_1 _14721_ (.Y(_05627_),
    .A(_05625_),
    .B(_05626_));
 sg13g2_nand2_1 _14722_ (.Y(_05628_),
    .A(_05627_),
    .B(_02977_));
 sg13g2_nand3_1 _14723_ (.B(_05626_),
    .C(\vgadonut.donut.donuthit.cordicxz.xin[4] ),
    .A(_05625_),
    .Y(_05629_));
 sg13g2_nand2_1 _14724_ (.Y(_05630_),
    .A(_05628_),
    .B(_05629_));
 sg13g2_xnor2_1 _14725_ (.Y(_05631_),
    .A(_05615_),
    .B(_05630_));
 sg13g2_nor2_1 _14726_ (.A(_05574_),
    .B(_05591_),
    .Y(_05632_));
 sg13g2_nor2_1 _14727_ (.A(_05632_),
    .B(_05542_),
    .Y(_05633_));
 sg13g2_nand2_1 _14728_ (.Y(_05634_),
    .A(_05549_),
    .B(_05633_));
 sg13g2_nand2_1 _14729_ (.Y(_05635_),
    .A(_05591_),
    .B(_05574_));
 sg13g2_nand2_1 _14730_ (.Y(_05636_),
    .A(_05634_),
    .B(_05635_));
 sg13g2_xor2_1 _14731_ (.B(_05636_),
    .A(_05631_),
    .X(_05637_));
 sg13g2_nand2_1 _14732_ (.Y(_05638_),
    .A(_05637_),
    .B(net126));
 sg13g2_o21ai_1 _14733_ (.B1(_05638_),
    .Y(_00089_),
    .A1(net122),
    .A2(_05613_));
 sg13g2_buf_1 _14734_ (.A(\vgadonut.donut.donuthit.rzin[10] ),
    .X(_05639_));
 sg13g2_inv_1 _14735_ (.Y(_05640_),
    .A(_05639_));
 sg13g2_nor2_1 _14736_ (.A(_05505_),
    .B(net203),
    .Y(_05641_));
 sg13g2_buf_1 _14737_ (.A(\vgadonut.donut.cAcB[11] ),
    .X(_05642_));
 sg13g2_buf_1 _14738_ (.A(_05642_),
    .X(_05643_));
 sg13g2_xor2_1 _14739_ (.B(net202),
    .A(net232),
    .X(_05644_));
 sg13g2_xor2_1 _14740_ (.B(_05644_),
    .A(_05641_),
    .X(_05645_));
 sg13g2_inv_1 _14741_ (.Y(_05646_),
    .A(_05645_));
 sg13g2_inv_1 _14742_ (.Y(_05647_),
    .A(_05563_));
 sg13g2_inv_1 _14743_ (.Y(_05648_),
    .A(_05600_));
 sg13g2_nor2_1 _14744_ (.A(_05601_),
    .B(_05648_),
    .Y(_05649_));
 sg13g2_nand2_1 _14745_ (.Y(_05650_),
    .A(_05599_),
    .B(_05596_));
 sg13g2_inv_1 _14746_ (.Y(_05651_),
    .A(_05650_));
 sg13g2_a221oi_1 _14747_ (.B2(_05649_),
    .C1(_05651_),
    .B1(_05647_),
    .A1(net203),
    .Y(_05652_),
    .A2(_05604_));
 sg13g2_xnor2_1 _14748_ (.Y(_05653_),
    .A(_05646_),
    .B(_05652_));
 sg13g2_nor2_1 _14749_ (.A(_05640_),
    .B(_05653_),
    .Y(_05654_));
 sg13g2_inv_1 _14750_ (.Y(_05655_),
    .A(_05654_));
 sg13g2_nand2_1 _14751_ (.Y(_05656_),
    .A(_05653_),
    .B(_05640_));
 sg13g2_nand2_1 _14752_ (.Y(_05657_),
    .A(_05655_),
    .B(_05656_));
 sg13g2_inv_1 _14753_ (.Y(_05658_),
    .A(_05612_));
 sg13g2_a21oi_1 _14754_ (.A1(_05658_),
    .A2(_05610_),
    .Y(_05659_),
    .B1(_05609_));
 sg13g2_xor2_1 _14755_ (.B(_05659_),
    .A(_05657_),
    .X(_05660_));
 sg13g2_nor2_1 _14756_ (.A(_05615_),
    .B(_05630_),
    .Y(_05661_));
 sg13g2_nor2_1 _14757_ (.A(_05661_),
    .B(_05632_),
    .Y(_05662_));
 sg13g2_nand2_1 _14758_ (.Y(_05663_),
    .A(_05630_),
    .B(_05615_));
 sg13g2_nor2b_1 _14759_ (.A(_05662_),
    .B_N(_05663_),
    .Y(_05664_));
 sg13g2_nor2_1 _14760_ (.A(_05631_),
    .B(_05592_),
    .Y(_05665_));
 sg13g2_nand2_1 _14761_ (.Y(_05666_),
    .A(_05571_),
    .B(_05665_));
 sg13g2_nand2b_1 _14762_ (.Y(_05667_),
    .B(_05666_),
    .A_N(_05664_));
 sg13g2_nand2_1 _14763_ (.Y(_05668_),
    .A(_05629_),
    .B(_05626_));
 sg13g2_nor2_1 _14764_ (.A(_05353_),
    .B(net24),
    .Y(_05669_));
 sg13g2_nand2_1 _14765_ (.Y(_05670_),
    .A(net22),
    .B(_05319_));
 sg13g2_a22oi_1 _14766_ (.Y(_05671_),
    .B1(_05367_),
    .B2(net23),
    .A2(_05344_),
    .A1(net27));
 sg13g2_nand3_1 _14767_ (.B(_05670_),
    .C(_05671_),
    .A(_05621_),
    .Y(_05672_));
 sg13g2_nor2_1 _14768_ (.A(_05669_),
    .B(_05672_),
    .Y(_05673_));
 sg13g2_nand2_1 _14769_ (.Y(_05674_),
    .A(_05673_),
    .B(_05533_));
 sg13g2_nand2_1 _14770_ (.Y(_05675_),
    .A(_05674_),
    .B(net14));
 sg13g2_nand2_1 _14771_ (.Y(_05676_),
    .A(_05583_),
    .B(_05675_));
 sg13g2_nand3_1 _14772_ (.B(_05674_),
    .C(net12),
    .A(_05582_),
    .Y(_05677_));
 sg13g2_buf_1 _14773_ (.A(_05677_),
    .X(_05678_));
 sg13g2_nand2_1 _14774_ (.Y(_05679_),
    .A(_05676_),
    .B(_05678_));
 sg13g2_nand2_1 _14775_ (.Y(_05680_),
    .A(_05679_),
    .B(_03441_));
 sg13g2_nand3_1 _14776_ (.B(_05678_),
    .C(_02964_),
    .A(_05676_),
    .Y(_05681_));
 sg13g2_nand3_1 _14777_ (.B(_05680_),
    .C(_05681_),
    .A(_05668_),
    .Y(_05682_));
 sg13g2_buf_1 _14778_ (.A(_05682_),
    .X(_05683_));
 sg13g2_nand2_1 _14779_ (.Y(_05684_),
    .A(_05680_),
    .B(_05681_));
 sg13g2_inv_1 _14780_ (.Y(_05685_),
    .A(_05668_));
 sg13g2_nand2_1 _14781_ (.Y(_05686_),
    .A(_05684_),
    .B(_05685_));
 sg13g2_nand2_1 _14782_ (.Y(_05687_),
    .A(_05683_),
    .B(_05686_));
 sg13g2_inv_1 _14783_ (.Y(_05688_),
    .A(_05687_));
 sg13g2_a21oi_1 _14784_ (.A1(_05667_),
    .A2(_05688_),
    .Y(_05689_),
    .B1(net111));
 sg13g2_o21ai_1 _14785_ (.B1(_05689_),
    .Y(_05690_),
    .A1(_05667_),
    .A2(_05688_));
 sg13g2_o21ai_1 _14786_ (.B1(_05690_),
    .Y(_00090_),
    .A1(net122),
    .A2(_05660_));
 sg13g2_buf_2 _14787_ (.A(\vgadonut.donut.donuthit.rzin[11] ),
    .X(_05691_));
 sg13g2_nor2_1 _14788_ (.A(net232),
    .B(net202),
    .Y(_05692_));
 sg13g2_buf_1 _14789_ (.A(\vgadonut.donut.cAcB[12] ),
    .X(_05693_));
 sg13g2_buf_1 _14790_ (.A(_05693_),
    .X(_05694_));
 sg13g2_xor2_1 _14791_ (.B(net201),
    .A(_05598_),
    .X(_05695_));
 sg13g2_xor2_1 _14792_ (.B(_05695_),
    .A(_05692_),
    .X(_05696_));
 sg13g2_inv_1 _14793_ (.Y(_05697_),
    .A(_05607_));
 sg13g2_nor2_1 _14794_ (.A(_05648_),
    .B(_05646_),
    .Y(_05698_));
 sg13g2_nand2_1 _14795_ (.Y(_05699_),
    .A(_05644_),
    .B(_05641_));
 sg13g2_inv_1 _14796_ (.Y(_05700_),
    .A(_05699_));
 sg13g2_a221oi_1 _14797_ (.B2(_05698_),
    .C1(_05700_),
    .B1(_05697_),
    .A1(net202),
    .Y(_05701_),
    .A2(_05651_));
 sg13g2_xnor2_1 _14798_ (.Y(_05702_),
    .A(_05696_),
    .B(_05701_));
 sg13g2_nor2_1 _14799_ (.A(_05691_),
    .B(_05702_),
    .Y(_05703_));
 sg13g2_nand2_1 _14800_ (.Y(_05704_),
    .A(_05702_),
    .B(_05691_));
 sg13g2_inv_1 _14801_ (.Y(_05705_),
    .A(_05704_));
 sg13g2_nor2_1 _14802_ (.A(_05703_),
    .B(_05705_),
    .Y(_05706_));
 sg13g2_a21o_1 _14803_ (.A2(_05656_),
    .A1(_05659_),
    .B1(_05654_),
    .X(_05707_));
 sg13g2_xnor2_1 _14804_ (.Y(_05708_),
    .A(_05706_),
    .B(_05707_));
 sg13g2_nor2_1 _14805_ (.A(_05631_),
    .B(_05687_),
    .Y(_05709_));
 sg13g2_nand3_1 _14806_ (.B(_05635_),
    .C(_05709_),
    .A(_05634_),
    .Y(_05710_));
 sg13g2_inv_1 _14807_ (.Y(_05711_),
    .A(_05683_));
 sg13g2_a21oi_1 _14808_ (.A1(_05686_),
    .A2(_05661_),
    .Y(_05712_),
    .B1(_05711_));
 sg13g2_nand2_1 _14809_ (.Y(_05713_),
    .A(_05710_),
    .B(_05712_));
 sg13g2_inv_1 _14810_ (.Y(_05714_),
    .A(_05678_));
 sg13g2_a21oi_1 _14811_ (.A1(_05676_),
    .A2(_02964_),
    .Y(_05715_),
    .B1(_05714_));
 sg13g2_nand2_1 _14812_ (.Y(_05716_),
    .A(_04517_),
    .B(net19));
 sg13g2_a22oi_1 _14813_ (.Y(_05717_),
    .B1(_05319_),
    .B2(net21),
    .A2(_05367_),
    .A1(_04519_));
 sg13g2_nand2_1 _14814_ (.Y(_05718_),
    .A(_05716_),
    .B(_05717_));
 sg13g2_nand2_1 _14815_ (.Y(_05719_),
    .A(_05718_),
    .B(net13));
 sg13g2_nand2_1 _14816_ (.Y(_05720_),
    .A(_05719_),
    .B(_05624_));
 sg13g2_nand3_1 _14817_ (.B(net11),
    .C(_05623_),
    .A(_05718_),
    .Y(_05721_));
 sg13g2_nand2_1 _14818_ (.Y(_05722_),
    .A(_05720_),
    .B(_05721_));
 sg13g2_xnor2_1 _14819_ (.Y(_05723_),
    .A(_02957_),
    .B(_05722_));
 sg13g2_xnor2_1 _14820_ (.Y(_05724_),
    .A(_05715_),
    .B(_05723_));
 sg13g2_a21oi_1 _14821_ (.A1(_05713_),
    .A2(_05724_),
    .Y(_05725_),
    .B1(net111));
 sg13g2_o21ai_1 _14822_ (.B1(_05725_),
    .Y(_05726_),
    .A1(_05713_),
    .A2(_05724_));
 sg13g2_o21ai_1 _14823_ (.B1(_05726_),
    .Y(_00091_),
    .A1(net122),
    .A2(_05708_));
 sg13g2_buf_1 _14824_ (.A(\vgadonut.donut.donuthit.rzin[12] ),
    .X(_05727_));
 sg13g2_nor2_1 _14825_ (.A(net203),
    .B(net201),
    .Y(_05728_));
 sg13g2_buf_1 _14826_ (.A(\vgadonut.donut.cAcB[13] ),
    .X(_05729_));
 sg13g2_buf_1 _14827_ (.A(_05729_),
    .X(_05730_));
 sg13g2_xnor2_1 _14828_ (.Y(_05731_),
    .A(net202),
    .B(net200));
 sg13g2_xnor2_1 _14829_ (.Y(_05732_),
    .A(_05728_),
    .B(_05731_));
 sg13g2_nand2_1 _14830_ (.Y(_05733_),
    .A(_05645_),
    .B(_05696_));
 sg13g2_and2_1 _14831_ (.A(_05695_),
    .B(_05692_),
    .X(_05734_));
 sg13g2_a21oi_1 _14832_ (.A1(_05700_),
    .A2(net201),
    .Y(_05735_),
    .B1(_05734_));
 sg13g2_o21ai_1 _14833_ (.B1(_05735_),
    .Y(_05736_),
    .A1(_05733_),
    .A2(_05652_));
 sg13g2_xor2_1 _14834_ (.B(_05736_),
    .A(_05732_),
    .X(_05737_));
 sg13g2_nor2_1 _14835_ (.A(_05727_),
    .B(_05737_),
    .Y(_05738_));
 sg13g2_nand2_1 _14836_ (.Y(_05739_),
    .A(_05737_),
    .B(_05727_));
 sg13g2_inv_1 _14837_ (.Y(_05740_),
    .A(_05739_));
 sg13g2_nor2_1 _14838_ (.A(_05738_),
    .B(_05740_),
    .Y(_05741_));
 sg13g2_inv_1 _14839_ (.Y(_05742_),
    .A(_05703_));
 sg13g2_a21oi_1 _14840_ (.A1(_05707_),
    .A2(_05742_),
    .Y(_05743_),
    .B1(_05705_));
 sg13g2_xor2_1 _14841_ (.B(_05743_),
    .A(_05741_),
    .X(_05744_));
 sg13g2_inv_1 _14842_ (.Y(_05745_),
    .A(_05721_));
 sg13g2_a21oi_1 _14843_ (.A1(_05720_),
    .A2(_02957_),
    .Y(_05746_),
    .B1(_05745_));
 sg13g2_a22oi_1 _14844_ (.Y(_05747_),
    .B1(_05355_),
    .B2(_04520_),
    .A2(_05319_),
    .A1(_04519_));
 sg13g2_nand2_1 _14845_ (.Y(_05748_),
    .A(_05716_),
    .B(_05747_));
 sg13g2_nand2_1 _14846_ (.Y(_05749_),
    .A(_05748_),
    .B(net12));
 sg13g2_nand2_1 _14847_ (.Y(_05750_),
    .A(_05749_),
    .B(_05675_));
 sg13g2_nand3_1 _14848_ (.B(net11),
    .C(_05674_),
    .A(_05748_),
    .Y(_05751_));
 sg13g2_nand2_1 _14849_ (.Y(_05752_),
    .A(_05750_),
    .B(_05751_));
 sg13g2_xnor2_1 _14850_ (.Y(_05753_),
    .A(_03449_),
    .B(_05752_));
 sg13g2_nor2_1 _14851_ (.A(_05746_),
    .B(_05753_),
    .Y(_05754_));
 sg13g2_inv_1 _14852_ (.Y(_05755_),
    .A(_05746_));
 sg13g2_xnor2_1 _14853_ (.Y(_05756_),
    .A(_03275_),
    .B(_05752_));
 sg13g2_nor2_1 _14854_ (.A(_05755_),
    .B(_05756_),
    .Y(_05757_));
 sg13g2_nor2_1 _14855_ (.A(_05754_),
    .B(_05757_),
    .Y(_05758_));
 sg13g2_nand2_1 _14856_ (.Y(_05759_),
    .A(_05724_),
    .B(_05688_));
 sg13g2_inv_1 _14857_ (.Y(_05760_),
    .A(_05715_));
 sg13g2_nor2_1 _14858_ (.A(_05760_),
    .B(_05723_),
    .Y(_05761_));
 sg13g2_nand2_1 _14859_ (.Y(_05762_),
    .A(_05723_),
    .B(_05760_));
 sg13g2_nand2_1 _14860_ (.Y(_05763_),
    .A(_05762_),
    .B(_05683_));
 sg13g2_nand2b_1 _14861_ (.Y(_05764_),
    .B(_05763_),
    .A_N(_05761_));
 sg13g2_a21oi_1 _14862_ (.A1(_05762_),
    .A2(_05683_),
    .Y(_05765_),
    .B1(_05761_));
 sg13g2_nor2_1 _14863_ (.A(_05664_),
    .B(_05765_),
    .Y(_05766_));
 sg13g2_a22oi_1 _14864_ (.Y(_05767_),
    .B1(_05666_),
    .B2(_05766_),
    .A2(_05764_),
    .A1(_05759_));
 sg13g2_a21oi_1 _14865_ (.A1(_05767_),
    .A2(_05758_),
    .Y(_05768_),
    .B1(_09996_));
 sg13g2_o21ai_1 _14866_ (.B1(_05768_),
    .Y(_05769_),
    .A1(_05758_),
    .A2(_05767_));
 sg13g2_o21ai_1 _14867_ (.B1(_05769_),
    .Y(_00092_),
    .A1(_04531_),
    .A2(_05744_));
 sg13g2_buf_1 _14868_ (.A(\vgadonut.donut.donuthit.rzin[13] ),
    .X(_05770_));
 sg13g2_nor2_1 _14869_ (.A(net202),
    .B(net200),
    .Y(_05771_));
 sg13g2_buf_1 _14870_ (.A(\vgadonut.donut.cAcB[14] ),
    .X(_05772_));
 sg13g2_buf_1 _14871_ (.A(_05772_),
    .X(_05773_));
 sg13g2_xnor2_1 _14872_ (.Y(_05774_),
    .A(net201),
    .B(_05773_));
 sg13g2_xnor2_1 _14873_ (.Y(_05775_),
    .A(_05771_),
    .B(_05774_));
 sg13g2_nand2_1 _14874_ (.Y(_05776_),
    .A(_05696_),
    .B(_05732_));
 sg13g2_nor2b_1 _14875_ (.A(_05731_),
    .B_N(_05728_),
    .Y(_05777_));
 sg13g2_a21oi_1 _14876_ (.A1(_05734_),
    .A2(net200),
    .Y(_05778_),
    .B1(_05777_));
 sg13g2_o21ai_1 _14877_ (.B1(_05778_),
    .Y(_05779_),
    .A1(_05776_),
    .A2(_05701_));
 sg13g2_xor2_1 _14878_ (.B(_05779_),
    .A(_05775_),
    .X(_05780_));
 sg13g2_nor2_1 _14879_ (.A(_05770_),
    .B(_05780_),
    .Y(_05781_));
 sg13g2_nand2_1 _14880_ (.Y(_05782_),
    .A(_05780_),
    .B(_05770_));
 sg13g2_inv_1 _14881_ (.Y(_05783_),
    .A(_05782_));
 sg13g2_nor2_1 _14882_ (.A(_05781_),
    .B(_05783_),
    .Y(_05784_));
 sg13g2_a21oi_1 _14883_ (.A1(_05743_),
    .A2(_05739_),
    .Y(_05785_),
    .B1(_05738_));
 sg13g2_xnor2_1 _14884_ (.Y(_05786_),
    .A(_05784_),
    .B(_05785_));
 sg13g2_nand2_1 _14885_ (.Y(_05787_),
    .A(_05756_),
    .B(_05755_));
 sg13g2_a21oi_1 _14886_ (.A1(_05762_),
    .A2(_05787_),
    .Y(_05788_),
    .B1(_05757_));
 sg13g2_nor2b_1 _14887_ (.A(_05788_),
    .B_N(_05712_),
    .Y(_05789_));
 sg13g2_nand2_1 _14888_ (.Y(_05790_),
    .A(_05710_),
    .B(_05789_));
 sg13g2_nand2_1 _14889_ (.Y(_05791_),
    .A(_05758_),
    .B(_05724_));
 sg13g2_nand2b_1 _14890_ (.Y(_05792_),
    .B(_05791_),
    .A_N(_05788_));
 sg13g2_inv_1 _14891_ (.Y(_05793_),
    .A(_05751_));
 sg13g2_a21oi_2 _14892_ (.B1(_05793_),
    .Y(_05794_),
    .A2(_03275_),
    .A1(_05750_));
 sg13g2_nand2_1 _14893_ (.Y(_05795_),
    .A(net14),
    .B(net19));
 sg13g2_buf_2 _14894_ (.A(_05795_),
    .X(_05796_));
 sg13g2_nand2_1 _14895_ (.Y(_05797_),
    .A(_05719_),
    .B(_05796_));
 sg13g2_nand3_1 _14896_ (.B(net10),
    .C(net19),
    .A(_05718_),
    .Y(_05798_));
 sg13g2_nand2_1 _14897_ (.Y(_05799_),
    .A(_05797_),
    .B(_05798_));
 sg13g2_xnor2_1 _14898_ (.Y(_05800_),
    .A(_03146_),
    .B(_05799_));
 sg13g2_xor2_1 _14899_ (.B(_05800_),
    .A(_05794_),
    .X(_05801_));
 sg13g2_a21oi_1 _14900_ (.A1(_05790_),
    .A2(_05792_),
    .Y(_05802_),
    .B1(_05801_));
 sg13g2_nand3_1 _14901_ (.B(_05801_),
    .C(_05792_),
    .A(_05790_),
    .Y(_05803_));
 sg13g2_nand3b_1 _14902_ (.B(net123),
    .C(_05803_),
    .Y(_05804_),
    .A_N(_05802_));
 sg13g2_o21ai_1 _14903_ (.B1(_05804_),
    .Y(_00093_),
    .A1(net121),
    .A2(_05786_));
 sg13g2_inv_1 _14904_ (.Y(_05805_),
    .A(\vgadonut.donut.donuthit.rzin[14] ));
 sg13g2_nor2_1 _14905_ (.A(_05694_),
    .B(net199),
    .Y(_05806_));
 sg13g2_buf_4 _14906_ (.X(_05807_),
    .A(\vgadonut.donut.cAcB[15] ));
 sg13g2_xnor2_1 _14907_ (.Y(_05808_),
    .A(net200),
    .B(_05807_));
 sg13g2_xnor2_1 _14908_ (.Y(_05809_),
    .A(_05806_),
    .B(_05808_));
 sg13g2_nand3_1 _14909_ (.B(_05732_),
    .C(_05775_),
    .A(_05736_),
    .Y(_05810_));
 sg13g2_nor2b_1 _14910_ (.A(_05774_),
    .B_N(_05771_),
    .Y(_05811_));
 sg13g2_a21oi_1 _14911_ (.A1(_05777_),
    .A2(_05773_),
    .Y(_05812_),
    .B1(_05811_));
 sg13g2_nand2_1 _14912_ (.Y(_05813_),
    .A(_05810_),
    .B(_05812_));
 sg13g2_xor2_1 _14913_ (.B(_05813_),
    .A(_05809_),
    .X(_05814_));
 sg13g2_inv_1 _14914_ (.Y(_05815_),
    .A(_05814_));
 sg13g2_nor2_1 _14915_ (.A(_05805_),
    .B(_05815_),
    .Y(_05816_));
 sg13g2_nand2_1 _14916_ (.Y(_05817_),
    .A(_05815_),
    .B(_05805_));
 sg13g2_nand2b_1 _14917_ (.Y(_05818_),
    .B(_05817_),
    .A_N(_05816_));
 sg13g2_nand2b_1 _14918_ (.Y(_05819_),
    .B(_05741_),
    .A_N(_05743_));
 sg13g2_nor2_1 _14919_ (.A(_05740_),
    .B(_05783_),
    .Y(_05820_));
 sg13g2_a21oi_1 _14920_ (.A1(_05819_),
    .A2(_05820_),
    .Y(_05821_),
    .B1(_05781_));
 sg13g2_xor2_1 _14921_ (.B(_05821_),
    .A(_05818_),
    .X(_05822_));
 sg13g2_nand2_1 _14922_ (.Y(_05823_),
    .A(_05801_),
    .B(_05758_));
 sg13g2_nor2_1 _14923_ (.A(_05759_),
    .B(_05823_),
    .Y(_05824_));
 sg13g2_nand2_1 _14924_ (.Y(_05825_),
    .A(_05667_),
    .B(_05824_));
 sg13g2_nor2_1 _14925_ (.A(_05794_),
    .B(_05800_),
    .Y(_05826_));
 sg13g2_nor2_1 _14926_ (.A(_05754_),
    .B(_05826_),
    .Y(_05827_));
 sg13g2_nand2_1 _14927_ (.Y(_05828_),
    .A(_05800_),
    .B(_05794_));
 sg13g2_nor2b_1 _14928_ (.A(_05827_),
    .B_N(_05828_),
    .Y(_05829_));
 sg13g2_nor2_1 _14929_ (.A(_05764_),
    .B(_05823_),
    .Y(_05830_));
 sg13g2_nor2_1 _14930_ (.A(_05829_),
    .B(_05830_),
    .Y(_05831_));
 sg13g2_nand2_1 _14931_ (.Y(_05832_),
    .A(_05825_),
    .B(_05831_));
 sg13g2_inv_1 _14932_ (.Y(_05833_),
    .A(_05798_));
 sg13g2_a21oi_2 _14933_ (.B1(_05833_),
    .Y(_05834_),
    .A2(\vgadonut.donut.donuthit.cordicxz.xin[8] ),
    .A1(_05797_));
 sg13g2_nand2_1 _14934_ (.Y(_05835_),
    .A(_05749_),
    .B(_05796_));
 sg13g2_nand3_1 _14935_ (.B(net10),
    .C(net19),
    .A(_05748_),
    .Y(_05836_));
 sg13g2_nand2_1 _14936_ (.Y(_05837_),
    .A(_05835_),
    .B(_05836_));
 sg13g2_xnor2_1 _14937_ (.Y(_05838_),
    .A(_03270_),
    .B(_05837_));
 sg13g2_xor2_1 _14938_ (.B(_05838_),
    .A(_05834_),
    .X(_05839_));
 sg13g2_a21oi_1 _14939_ (.A1(_05832_),
    .A2(_05839_),
    .Y(_05840_),
    .B1(_09996_));
 sg13g2_o21ai_1 _14940_ (.B1(_05840_),
    .Y(_05841_),
    .A1(_05832_),
    .A2(_05839_));
 sg13g2_o21ai_1 _14941_ (.B1(_05841_),
    .Y(_00094_),
    .A1(net121),
    .A2(_05822_));
 sg13g2_inv_1 _14942_ (.Y(_05842_),
    .A(_05836_));
 sg13g2_a21oi_1 _14943_ (.A1(_05835_),
    .A2(\vgadonut.donut.donuthit.cordicxz.xin[9] ),
    .Y(_05843_),
    .B1(_05842_));
 sg13g2_xnor2_1 _14944_ (.Y(_05844_),
    .A(_03258_),
    .B(_05843_));
 sg13g2_inv_2 _14945_ (.Y(_05845_),
    .A(_05844_));
 sg13g2_xnor2_1 _14946_ (.Y(_05846_),
    .A(_05794_),
    .B(_05800_));
 sg13g2_xnor2_1 _14947_ (.Y(_05847_),
    .A(_05834_),
    .B(_05838_));
 sg13g2_nor2_1 _14948_ (.A(_05846_),
    .B(_05847_),
    .Y(_05848_));
 sg13g2_nand2_1 _14949_ (.Y(_05849_),
    .A(_05848_),
    .B(_05788_));
 sg13g2_nor2_1 _14950_ (.A(_05834_),
    .B(_05838_),
    .Y(_05850_));
 sg13g2_nand2_1 _14951_ (.Y(_05851_),
    .A(_05838_),
    .B(_05834_));
 sg13g2_o21ai_1 _14952_ (.B1(_05851_),
    .Y(_05852_),
    .A1(_05850_),
    .A2(_05826_));
 sg13g2_nand2_1 _14953_ (.Y(_05853_),
    .A(_05849_),
    .B(_05852_));
 sg13g2_inv_1 _14954_ (.Y(_05854_),
    .A(_05848_));
 sg13g2_nor2_1 _14955_ (.A(_05791_),
    .B(_05854_),
    .Y(_05855_));
 sg13g2_nand2_1 _14956_ (.Y(_05856_),
    .A(_05713_),
    .B(_05855_));
 sg13g2_nand2b_1 _14957_ (.Y(_05857_),
    .B(_05856_),
    .A_N(_05853_));
 sg13g2_nor2_1 _14958_ (.A(_05845_),
    .B(_05857_),
    .Y(_05858_));
 sg13g2_nand2_1 _14959_ (.Y(_05859_),
    .A(_05857_),
    .B(_05845_));
 sg13g2_nand2_1 _14960_ (.Y(_05860_),
    .A(_05859_),
    .B(net125));
 sg13g2_buf_1 _14961_ (.A(\vgadonut.donut.donuthit.rzin[15] ),
    .X(_05861_));
 sg13g2_nor2_1 _14962_ (.A(net200),
    .B(_05807_),
    .Y(_05862_));
 sg13g2_xor2_1 _14963_ (.B(_05807_),
    .A(net199),
    .X(_05863_));
 sg13g2_nor2_1 _14964_ (.A(_05862_),
    .B(_05863_),
    .Y(_05864_));
 sg13g2_a21o_1 _14965_ (.A2(_05862_),
    .A1(net199),
    .B1(_05864_),
    .X(_05865_));
 sg13g2_nor2_1 _14966_ (.A(_05806_),
    .B(_05811_),
    .Y(_05866_));
 sg13g2_nand3_1 _14967_ (.B(_05775_),
    .C(_05809_),
    .A(_05779_),
    .Y(_05867_));
 sg13g2_o21ai_1 _14968_ (.B1(_05867_),
    .Y(_05868_),
    .A1(_05808_),
    .A2(_05866_));
 sg13g2_xnor2_1 _14969_ (.Y(_05869_),
    .A(_05865_),
    .B(_05868_));
 sg13g2_xnor2_1 _14970_ (.Y(_05870_),
    .A(_05861_),
    .B(_05869_));
 sg13g2_a21oi_1 _14971_ (.A1(_05821_),
    .A2(_05817_),
    .Y(_05871_),
    .B1(_05816_));
 sg13g2_or2_1 _14972_ (.X(_05872_),
    .B(_05871_),
    .A(_05870_));
 sg13g2_nand2_1 _14973_ (.Y(_05873_),
    .A(_05871_),
    .B(_05870_));
 sg13g2_nand3_1 _14974_ (.B(net112),
    .C(_05873_),
    .A(_05872_),
    .Y(_05874_));
 sg13g2_o21ai_1 _14975_ (.B1(_05874_),
    .Y(_00080_),
    .A1(_05858_),
    .A2(_05860_));
 sg13g2_xor2_1 _14976_ (.B(_05796_),
    .A(_00158_),
    .X(_05875_));
 sg13g2_inv_1 _14977_ (.Y(_05876_),
    .A(_05875_));
 sg13g2_nand2_1 _14978_ (.Y(_05877_),
    .A(_05839_),
    .B(_05845_));
 sg13g2_nor2_1 _14979_ (.A(_05877_),
    .B(_05823_),
    .Y(_05878_));
 sg13g2_nand2_1 _14980_ (.Y(_05879_),
    .A(_05767_),
    .B(_05878_));
 sg13g2_nor2_1 _14981_ (.A(_05844_),
    .B(_05847_),
    .Y(_05880_));
 sg13g2_nand2_1 _14982_ (.Y(_05881_),
    .A(_05829_),
    .B(_05880_));
 sg13g2_nor2_1 _14983_ (.A(_00164_),
    .B(_05843_),
    .Y(_05882_));
 sg13g2_a21oi_1 _14984_ (.A1(_05845_),
    .A2(_05850_),
    .Y(_05883_),
    .B1(_05882_));
 sg13g2_nand2_1 _14985_ (.Y(_05884_),
    .A(_05881_),
    .B(_05883_));
 sg13g2_inv_1 _14986_ (.Y(_05885_),
    .A(_05884_));
 sg13g2_nand2_1 _14987_ (.Y(_05886_),
    .A(_05879_),
    .B(_05885_));
 sg13g2_xnor2_1 _14988_ (.Y(_05887_),
    .A(_05876_),
    .B(_05886_));
 sg13g2_nand2_1 _14989_ (.Y(_05888_),
    .A(_05887_),
    .B(net121));
 sg13g2_inv_1 _14990_ (.Y(_05889_),
    .A(_05861_));
 sg13g2_nor2_1 _14991_ (.A(net199),
    .B(_05807_),
    .Y(_05890_));
 sg13g2_nand2_1 _14992_ (.Y(_05891_),
    .A(_05813_),
    .B(_05809_));
 sg13g2_nor4_1 _14993_ (.A(net201),
    .B(net199),
    .C(_05808_),
    .D(_05865_),
    .Y(_05892_));
 sg13g2_a21oi_1 _14994_ (.A1(net199),
    .A2(_05862_),
    .Y(_05893_),
    .B1(_05892_));
 sg13g2_o21ai_1 _14995_ (.B1(_05893_),
    .Y(_05894_),
    .A1(_05864_),
    .A2(_05891_));
 sg13g2_xnor2_1 _14996_ (.Y(_05895_),
    .A(_05890_),
    .B(_05894_));
 sg13g2_xnor2_1 _14997_ (.Y(_05896_),
    .A(_05889_),
    .B(_05895_));
 sg13g2_inv_1 _14998_ (.Y(_05897_),
    .A(_05869_));
 sg13g2_o21ai_1 _14999_ (.B1(_05872_),
    .Y(_05898_),
    .A1(_00095_),
    .A2(_05897_));
 sg13g2_xnor2_1 _15000_ (.Y(_05899_),
    .A(_05896_),
    .B(_05898_));
 sg13g2_nand2_1 _15001_ (.Y(_05900_),
    .A(_05899_),
    .B(net110));
 sg13g2_nand2_1 _15002_ (.Y(_00081_),
    .A(_05888_),
    .B(_05900_));
 sg13g2_nor2_1 _15003_ (.A(_05876_),
    .B(_05844_),
    .Y(_05901_));
 sg13g2_nor2b_1 _15004_ (.A(_05854_),
    .B_N(_05901_),
    .Y(_05902_));
 sg13g2_nand3_1 _15005_ (.B(_05792_),
    .C(_05902_),
    .A(_05790_),
    .Y(_05903_));
 sg13g2_inv_1 _15006_ (.Y(_05904_),
    .A(_05852_));
 sg13g2_nor3_1 _15007_ (.A(_00164_),
    .B(_05876_),
    .C(_05843_),
    .Y(_05905_));
 sg13g2_a21oi_1 _15008_ (.A1(_05904_),
    .A2(_05901_),
    .Y(_05906_),
    .B1(_05905_));
 sg13g2_nand2_1 _15009_ (.Y(_05907_),
    .A(_05903_),
    .B(_05906_));
 sg13g2_inv_1 _15010_ (.Y(_05908_),
    .A(_05796_));
 sg13g2_nand2_1 _15011_ (.Y(_05909_),
    .A(_05908_),
    .B(_03456_));
 sg13g2_xnor2_1 _15012_ (.Y(_05910_),
    .A(_03381_),
    .B(_05909_));
 sg13g2_inv_2 _15013_ (.Y(_05911_),
    .A(_05910_));
 sg13g2_nand2_1 _15014_ (.Y(_05912_),
    .A(_05907_),
    .B(_05911_));
 sg13g2_nand3_1 _15015_ (.B(_05906_),
    .C(_05910_),
    .A(_05903_),
    .Y(_05913_));
 sg13g2_nand2_1 _15016_ (.Y(_05914_),
    .A(_05912_),
    .B(_05913_));
 sg13g2_nand2_1 _15017_ (.Y(_05915_),
    .A(_05914_),
    .B(net121));
 sg13g2_nor3_1 _15018_ (.A(_05889_),
    .B(_00095_),
    .C(_05895_),
    .Y(_05916_));
 sg13g2_nor2_1 _15019_ (.A(_00095_),
    .B(_05895_),
    .Y(_05917_));
 sg13g2_nor3_1 _15020_ (.A(_05896_),
    .B(_05917_),
    .C(_05898_),
    .Y(_05918_));
 sg13g2_o21ai_1 _15021_ (.B1(_09996_),
    .Y(_05919_),
    .A1(_05916_),
    .A2(_05918_));
 sg13g2_buf_1 _15022_ (.A(_05919_),
    .X(_05920_));
 sg13g2_nand2_1 _15023_ (.Y(_00082_),
    .A(_05915_),
    .B(_05920_));
 sg13g2_nor2_1 _15024_ (.A(_03398_),
    .B(_05796_),
    .Y(_05921_));
 sg13g2_xnor2_1 _15025_ (.Y(_05922_),
    .A(_03346_),
    .B(_05921_));
 sg13g2_nor2_1 _15026_ (.A(_05876_),
    .B(_05911_),
    .Y(_05923_));
 sg13g2_nor2b_1 _15027_ (.A(_05877_),
    .B_N(_05923_),
    .Y(_05924_));
 sg13g2_nand2_1 _15028_ (.Y(_05925_),
    .A(_05832_),
    .B(_05924_));
 sg13g2_inv_1 _15029_ (.Y(_05926_),
    .A(_05883_));
 sg13g2_nor3_1 _15030_ (.A(_03456_),
    .B(_03381_),
    .C(_05796_),
    .Y(_05927_));
 sg13g2_a21oi_1 _15031_ (.A1(_05926_),
    .A2(_05923_),
    .Y(_05928_),
    .B1(_05927_));
 sg13g2_nand2_1 _15032_ (.Y(_05929_),
    .A(_05925_),
    .B(_05928_));
 sg13g2_nand2b_1 _15033_ (.Y(_05930_),
    .B(_05929_),
    .A_N(_05922_));
 sg13g2_nand3_1 _15034_ (.B(_05928_),
    .C(_05922_),
    .A(_05925_),
    .Y(_05931_));
 sg13g2_nand2_1 _15035_ (.Y(_05932_),
    .A(_05930_),
    .B(_05931_));
 sg13g2_nand2_1 _15036_ (.Y(_05933_),
    .A(_05932_),
    .B(net121));
 sg13g2_nand2_1 _15037_ (.Y(_00083_),
    .A(_05933_),
    .B(_05920_));
 sg13g2_nand2_1 _15038_ (.Y(_05934_),
    .A(_05923_),
    .B(_05922_));
 sg13g2_nor2_1 _15039_ (.A(_05934_),
    .B(_05844_),
    .Y(_05935_));
 sg13g2_nand3_1 _15040_ (.B(_05855_),
    .C(_05935_),
    .A(_05713_),
    .Y(_05936_));
 sg13g2_nand3_1 _15041_ (.B(_05910_),
    .C(_05922_),
    .A(_05905_),
    .Y(_05937_));
 sg13g2_nand2_1 _15042_ (.Y(_05938_),
    .A(_05922_),
    .B(_05927_));
 sg13g2_nand3_1 _15043_ (.B(_03398_),
    .C(_03346_),
    .A(_05908_),
    .Y(_05939_));
 sg13g2_nand3_1 _15044_ (.B(_05938_),
    .C(_05939_),
    .A(_05937_),
    .Y(_05940_));
 sg13g2_a21oi_1 _15045_ (.A1(_05853_),
    .A2(_05935_),
    .Y(_05941_),
    .B1(_05940_));
 sg13g2_nand2_1 _15046_ (.Y(_05942_),
    .A(_05936_),
    .B(_05941_));
 sg13g2_nor2_1 _15047_ (.A(_03477_),
    .B(_05796_),
    .Y(_05943_));
 sg13g2_nand2_1 _15048_ (.Y(_05944_),
    .A(_05908_),
    .B(_03346_));
 sg13g2_a22oi_1 _15049_ (.Y(_05945_),
    .B1(_03477_),
    .B2(_05944_),
    .A2(_03346_),
    .A1(_05943_));
 sg13g2_buf_1 _15050_ (.A(_05945_),
    .X(_05946_));
 sg13g2_nand2_1 _15051_ (.Y(_05947_),
    .A(_05942_),
    .B(_05946_));
 sg13g2_inv_1 _15052_ (.Y(_05948_),
    .A(_05946_));
 sg13g2_nand3_1 _15053_ (.B(_05941_),
    .C(_05948_),
    .A(_05936_),
    .Y(_05949_));
 sg13g2_nand2_1 _15054_ (.Y(_05950_),
    .A(_05947_),
    .B(_05949_));
 sg13g2_nand2_1 _15055_ (.Y(_05951_),
    .A(_05950_),
    .B(net121));
 sg13g2_nand2_1 _15056_ (.Y(_00084_),
    .A(_05951_),
    .B(_05920_));
 sg13g2_nand2_1 _15057_ (.Y(_05952_),
    .A(_05766_),
    .B(_05666_));
 sg13g2_nand2_1 _15058_ (.Y(_05953_),
    .A(_05759_),
    .B(_05764_));
 sg13g2_nor2_1 _15059_ (.A(_05946_),
    .B(_05934_),
    .Y(_05954_));
 sg13g2_nand4_1 _15060_ (.B(_05953_),
    .C(_05878_),
    .A(_05952_),
    .Y(_05955_),
    .D(_05954_));
 sg13g2_o21ai_1 _15061_ (.B1(_05943_),
    .Y(_05956_),
    .A1(_03398_),
    .A2(_03348_));
 sg13g2_o21ai_1 _15062_ (.B1(_05956_),
    .Y(_05957_),
    .A1(_05946_),
    .A2(_05938_));
 sg13g2_a21oi_1 _15063_ (.A1(_05884_),
    .A2(_05954_),
    .Y(_05958_),
    .B1(_05957_));
 sg13g2_nand2_1 _15064_ (.Y(_05959_),
    .A(_05955_),
    .B(_05958_));
 sg13g2_xnor2_1 _15065_ (.Y(_05960_),
    .A(_00165_),
    .B(_05943_));
 sg13g2_nand2_1 _15066_ (.Y(_05961_),
    .A(_05959_),
    .B(_05960_));
 sg13g2_inv_1 _15067_ (.Y(_05962_),
    .A(_05960_));
 sg13g2_nand3_1 _15068_ (.B(_05958_),
    .C(_05962_),
    .A(_05955_),
    .Y(_05963_));
 sg13g2_nand3_1 _15069_ (.B(_05963_),
    .C(net123),
    .A(_05961_),
    .Y(_05964_));
 sg13g2_nand2_1 _15070_ (.Y(_00085_),
    .A(_05964_),
    .B(_05920_));
 sg13g2_nand2_1 _15071_ (.Y(_05965_),
    .A(\vgadonut.donut.h_count[7] ),
    .B(net255));
 sg13g2_nor2_1 _15072_ (.A(_09905_),
    .B(_09884_),
    .Y(_05966_));
 sg13g2_inv_1 _15073_ (.Y(_05967_),
    .A(_05966_));
 sg13g2_nand3_1 _15074_ (.B(_09726_),
    .C(_09694_),
    .A(net254),
    .Y(_05968_));
 sg13g2_nor3_1 _15075_ (.A(_05965_),
    .B(_05967_),
    .C(_05968_),
    .Y(_05969_));
 sg13g2_nand2_2 _15076_ (.Y(_05970_),
    .A(_10040_),
    .B(_05969_));
 sg13g2_inv_2 _15077_ (.Y(_05971_),
    .A(_05970_));
 sg13g2_nor2_1 _15078_ (.A(_09884_),
    .B(_05971_),
    .Y(_00015_));
 sg13g2_nand2_2 _15079_ (.Y(_05972_),
    .A(_09905_),
    .B(_09884_));
 sg13g2_nor2b_1 _15080_ (.A(_05966_),
    .B_N(_05972_),
    .Y(_00017_));
 sg13g2_nor2_1 _15081_ (.A(_00171_),
    .B(_05972_),
    .Y(_05973_));
 sg13g2_inv_1 _15082_ (.Y(_05974_),
    .A(_09726_));
 sg13g2_nor3_1 _15083_ (.A(_05974_),
    .B(_09705_),
    .C(_05965_),
    .Y(_05975_));
 sg13g2_nand4_1 _15084_ (.B(net254),
    .C(_05966_),
    .A(_10040_),
    .Y(_05976_),
    .D(_05975_));
 sg13g2_inv_1 _15085_ (.Y(_05977_),
    .A(_05976_));
 sg13g2_a21oi_1 _15086_ (.A1(_00171_),
    .A2(_05972_),
    .Y(_05978_),
    .B1(_05977_));
 sg13g2_nor2b_1 _15087_ (.A(_05973_),
    .B_N(_05978_),
    .Y(_00018_));
 sg13g2_nor2_1 _15088_ (.A(_09853_),
    .B(_05972_),
    .Y(_05979_));
 sg13g2_xor2_1 _15089_ (.B(_05979_),
    .A(_00170_),
    .X(_05980_));
 sg13g2_nor2_1 _15090_ (.A(_05980_),
    .B(_05971_),
    .Y(_00019_));
 sg13g2_nand2_1 _15091_ (.Y(_05981_),
    .A(_05979_),
    .B(_09716_));
 sg13g2_nor2_1 _15092_ (.A(_05974_),
    .B(_05981_),
    .Y(_05982_));
 sg13g2_inv_1 _15093_ (.Y(_05983_),
    .A(_05982_));
 sg13g2_nand2_1 _15094_ (.Y(_05984_),
    .A(_05970_),
    .B(_05983_));
 sg13g2_a21oi_1 _15095_ (.A1(_05974_),
    .A2(_05981_),
    .Y(_00020_),
    .B1(_05984_));
 sg13g2_nor2_1 _15096_ (.A(_09694_),
    .B(_05982_),
    .Y(_05985_));
 sg13g2_nor2_1 _15097_ (.A(_09705_),
    .B(_05983_),
    .Y(_05986_));
 sg13g2_nor3_1 _15098_ (.A(_05985_),
    .B(_05971_),
    .C(_05986_),
    .Y(_00021_));
 sg13g2_nor2_1 _15099_ (.A(net255),
    .B(_05986_),
    .Y(_05987_));
 sg13g2_nand2_1 _15100_ (.Y(_05988_),
    .A(_05986_),
    .B(net255));
 sg13g2_inv_1 _15101_ (.Y(_05989_),
    .A(_05988_));
 sg13g2_nor3_1 _15102_ (.A(_05971_),
    .B(_05987_),
    .C(_05989_),
    .Y(_00022_));
 sg13g2_nor2_2 _15103_ (.A(_09663_),
    .B(_05988_),
    .Y(_05990_));
 sg13g2_nor2_1 _15104_ (.A(\vgadonut.donut.h_count[7] ),
    .B(_05989_),
    .Y(_05991_));
 sg13g2_nor3_1 _15105_ (.A(_05977_),
    .B(_05990_),
    .C(_05991_),
    .Y(_00023_));
 sg13g2_nand2b_1 _15106_ (.Y(_05992_),
    .B(net254),
    .A_N(_09716_));
 sg13g2_nor2_1 _15107_ (.A(_05967_),
    .B(_05992_),
    .Y(_05993_));
 sg13g2_and3_1 _15108_ (.X(_05994_),
    .A(_05975_),
    .B(_10029_),
    .C(_05993_));
 sg13g2_xor2_1 _15109_ (.B(_05990_),
    .A(_00172_),
    .X(_05995_));
 sg13g2_nor2_1 _15110_ (.A(_05994_),
    .B(_05995_),
    .Y(_00024_));
 sg13g2_a21oi_1 _15111_ (.A1(_05990_),
    .A2(_09654_),
    .Y(_05996_),
    .B1(_09645_));
 sg13g2_nand3_1 _15112_ (.B(_09645_),
    .C(_09654_),
    .A(_05990_),
    .Y(_05997_));
 sg13g2_buf_1 _15113_ (.A(_05997_),
    .X(_05998_));
 sg13g2_nor2b_1 _15114_ (.A(_05996_),
    .B_N(_05998_),
    .Y(_00025_));
 sg13g2_o21ai_1 _15115_ (.B1(_05970_),
    .Y(_05999_),
    .A1(_10011_),
    .A2(_05998_));
 sg13g2_a21oi_1 _15116_ (.A1(_10011_),
    .A2(_05998_),
    .Y(_00016_),
    .B1(_05999_));
 sg13g2_buf_1 _15117_ (.A(\vgadonut.donut.v_count[2] ),
    .X(_06000_));
 sg13g2_inv_1 _15118_ (.Y(_06001_),
    .A(_09894_));
 sg13g2_buf_1 _15119_ (.A(\vgadonut.donut.v_count[3] ),
    .X(_06002_));
 sg13g2_inv_1 _15120_ (.Y(_06003_),
    .A(_06002_));
 sg13g2_buf_2 _15121_ (.A(\vgadonut.donut.v_count[5] ),
    .X(_06004_));
 sg13g2_inv_1 _15122_ (.Y(_06005_),
    .A(_06004_));
 sg13g2_nor4_1 _15123_ (.A(_06000_),
    .B(_06001_),
    .C(_06003_),
    .D(_06005_),
    .Y(_06006_));
 sg13g2_buf_1 _15124_ (.A(\vgadonut.donut.v_count[7] ),
    .X(_06007_));
 sg13g2_buf_1 _15125_ (.A(\vgadonut.donut.v_count[6] ),
    .X(_06008_));
 sg13g2_buf_1 _15126_ (.A(\vgadonut.donut.v_count[4] ),
    .X(_06009_));
 sg13g2_inv_1 _15127_ (.Y(_06010_),
    .A(\vgadonut.donut.v_count[8] ));
 sg13g2_nor3_1 _15128_ (.A(_06009_),
    .B(\vgadonut.donut.v_count[9] ),
    .C(_06010_),
    .Y(_06011_));
 sg13g2_nand4_1 _15129_ (.B(_06007_),
    .C(_06008_),
    .A(_06006_),
    .Y(_00027_),
    .D(_06011_));
 sg13g2_nor2_1 _15130_ (.A(_09769_),
    .B(_05972_),
    .Y(_06012_));
 sg13g2_nor2_1 _15131_ (.A(_09716_),
    .B(_09726_),
    .Y(_06013_));
 sg13g2_nand2_1 _15132_ (.Y(_06014_),
    .A(_06013_),
    .B(_00171_));
 sg13g2_nor2_1 _15133_ (.A(_06012_),
    .B(_06014_),
    .Y(_06015_));
 sg13g2_nor3_1 _15134_ (.A(_10051_),
    .B(_06015_),
    .C(_09748_),
    .Y(_06016_));
 sg13g2_nor3_1 _15135_ (.A(_09716_),
    .B(_09645_),
    .C(_09654_),
    .Y(_06017_));
 sg13g2_nand3_1 _15136_ (.B(_06012_),
    .C(_06017_),
    .A(_10062_),
    .Y(_06018_));
 sg13g2_inv_1 _15137_ (.Y(_06019_),
    .A(_09790_));
 sg13g2_o21ai_1 _15138_ (.B1(_06019_),
    .Y(_06020_),
    .A1(_10011_),
    .A2(_06018_));
 sg13g2_nor2_1 _15139_ (.A(_09905_),
    .B(_09769_),
    .Y(_06021_));
 sg13g2_nor2_1 _15140_ (.A(_09694_),
    .B(net255),
    .Y(_06022_));
 sg13g2_o21ai_1 _15141_ (.B1(_06022_),
    .Y(_06023_),
    .A1(_09737_),
    .A2(_06021_));
 sg13g2_nor4_1 _15142_ (.A(_09645_),
    .B(_09663_),
    .C(_10020_),
    .D(_09672_),
    .Y(_06024_));
 sg13g2_a22oi_1 _15143_ (.Y(_06025_),
    .B1(_06023_),
    .B2(_06024_),
    .A2(\vgadonut.donut.h_count[10] ),
    .A1(_09645_));
 sg13g2_o21ai_1 _15144_ (.B1(_06025_),
    .Y(_00026_),
    .A1(_06016_),
    .A2(_06020_));
 sg13g2_buf_1 _15145_ (.A(\vgadonut.donut.sA[5] ),
    .X(_06026_));
 sg13g2_buf_1 _15146_ (.A(_06026_),
    .X(_06027_));
 sg13g2_xor2_1 _15147_ (.B(\vgadonut.donut.cA[0] ),
    .A(net198),
    .X(_06028_));
 sg13g2_buf_1 _15148_ (.A(\vgadonut.donut.cB[15] ),
    .X(_06029_));
 sg13g2_buf_1 _15149_ (.A(_06029_),
    .X(_06030_));
 sg13g2_buf_2 _15150_ (.A(\vgadonut.donut.cB[12] ),
    .X(_06031_));
 sg13g2_inv_1 _15151_ (.Y(_06032_),
    .A(_06031_));
 sg13g2_buf_2 _15152_ (.A(\vgadonut.donut.cB[11] ),
    .X(_06033_));
 sg13g2_inv_1 _15153_ (.Y(_06034_),
    .A(_06033_));
 sg13g2_buf_2 _15154_ (.A(\vgadonut.donut.cB[10] ),
    .X(_06035_));
 sg13g2_inv_1 _15155_ (.Y(_06036_),
    .A(net245));
 sg13g2_nor2_1 _15156_ (.A(_06035_),
    .B(_06036_),
    .Y(_06037_));
 sg13g2_buf_1 _15157_ (.A(\vgadonut.donut.cB[1] ),
    .X(_06038_));
 sg13g2_inv_1 _15158_ (.Y(_06039_),
    .A(net248));
 sg13g2_buf_1 _15159_ (.A(\vgadonut.donut.cB[0] ),
    .X(_06040_));
 sg13g2_inv_1 _15160_ (.Y(_06041_),
    .A(net251));
 sg13g2_nor2_1 _15161_ (.A(net230),
    .B(_06041_),
    .Y(_06042_));
 sg13g2_xnor2_1 _15162_ (.Y(_06043_),
    .A(net231),
    .B(net248));
 sg13g2_nor2b_1 _15163_ (.A(_06042_),
    .B_N(_06043_),
    .Y(_06044_));
 sg13g2_a21oi_1 _15164_ (.A1(net231),
    .A2(_06039_),
    .Y(_06045_),
    .B1(_06044_));
 sg13g2_inv_1 _15165_ (.Y(_06046_),
    .A(_06045_));
 sg13g2_buf_1 _15166_ (.A(\vgadonut.donut.cB[2] ),
    .X(_06047_));
 sg13g2_inv_1 _15167_ (.Y(_06048_),
    .A(net213));
 sg13g2_nor2_1 _15168_ (.A(_06047_),
    .B(_06048_),
    .Y(_06049_));
 sg13g2_inv_1 _15169_ (.Y(_06050_),
    .A(_06049_));
 sg13g2_nor2b_1 _15170_ (.A(net213),
    .B_N(_06047_),
    .Y(_06051_));
 sg13g2_a21oi_2 _15171_ (.B1(_06051_),
    .Y(_06052_),
    .A2(_06050_),
    .A1(_06046_));
 sg13g2_inv_1 _15172_ (.Y(_06053_),
    .A(_06052_));
 sg13g2_buf_1 _15173_ (.A(\vgadonut.donut.cB[3] ),
    .X(_06054_));
 sg13g2_inv_1 _15174_ (.Y(_06055_),
    .A(net229));
 sg13g2_nor2_1 _15175_ (.A(net212),
    .B(_06055_),
    .Y(_06056_));
 sg13g2_nor2b_1 _15176_ (.A(net229),
    .B_N(net212),
    .Y(_06057_));
 sg13g2_nor2_1 _15177_ (.A(_06056_),
    .B(_06057_),
    .Y(_06058_));
 sg13g2_nand2_1 _15178_ (.Y(_06059_),
    .A(_06053_),
    .B(_06058_));
 sg13g2_buf_2 _15179_ (.A(\vgadonut.donut.cB[4] ),
    .X(_06060_));
 sg13g2_inv_1 _15180_ (.Y(_06061_),
    .A(_06060_));
 sg13g2_nor2_1 _15181_ (.A(net211),
    .B(_06061_),
    .Y(_06062_));
 sg13g2_nor2_1 _15182_ (.A(_06062_),
    .B(_06056_),
    .Y(_06063_));
 sg13g2_nor2b_1 _15183_ (.A(_06060_),
    .B_N(net211),
    .Y(_06064_));
 sg13g2_a21oi_1 _15184_ (.A1(_06059_),
    .A2(_06063_),
    .Y(_06065_),
    .B1(_06064_));
 sg13g2_buf_2 _15185_ (.A(\vgadonut.donut.cB[5] ),
    .X(_06066_));
 sg13g2_inv_1 _15186_ (.Y(_06067_),
    .A(net247));
 sg13g2_nor2_1 _15187_ (.A(_06066_),
    .B(_06067_),
    .Y(_06068_));
 sg13g2_nor2b_1 _15188_ (.A(net247),
    .B_N(_06066_),
    .Y(_06069_));
 sg13g2_nor2_1 _15189_ (.A(_06068_),
    .B(_06069_),
    .Y(_06070_));
 sg13g2_nand2_1 _15190_ (.Y(_06071_),
    .A(_06065_),
    .B(_06070_));
 sg13g2_buf_2 _15191_ (.A(\vgadonut.donut.cB[6] ),
    .X(_06072_));
 sg13g2_nor2b_1 _15192_ (.A(_04496_),
    .B_N(_06072_),
    .Y(_06073_));
 sg13g2_nor2_1 _15193_ (.A(_06073_),
    .B(_06069_),
    .Y(_06074_));
 sg13g2_inv_1 _15194_ (.Y(_06075_),
    .A(_04495_));
 sg13g2_nor2_1 _15195_ (.A(_06072_),
    .B(_06075_),
    .Y(_06076_));
 sg13g2_a21oi_1 _15196_ (.A1(_06071_),
    .A2(_06074_),
    .Y(_06077_),
    .B1(_06076_));
 sg13g2_buf_2 _15197_ (.A(\vgadonut.donut.cB[7] ),
    .X(_06078_));
 sg13g2_inv_1 _15198_ (.Y(_06079_),
    .A(_06078_));
 sg13g2_nor2_1 _15199_ (.A(_04533_),
    .B(_06079_),
    .Y(_06080_));
 sg13g2_inv_1 _15200_ (.Y(_06081_),
    .A(_04533_));
 sg13g2_nor2_1 _15201_ (.A(_06078_),
    .B(_06081_),
    .Y(_06082_));
 sg13g2_nor2_1 _15202_ (.A(_06080_),
    .B(_06082_),
    .Y(_06083_));
 sg13g2_nand2_1 _15203_ (.Y(_06084_),
    .A(_06077_),
    .B(_06083_));
 sg13g2_buf_2 _15204_ (.A(\vgadonut.donut.cB[8] ),
    .X(_06085_));
 sg13g2_inv_1 _15205_ (.Y(_06086_),
    .A(_06085_));
 sg13g2_nor2_1 _15206_ (.A(net246),
    .B(_06086_),
    .Y(_06087_));
 sg13g2_nor2_1 _15207_ (.A(_06080_),
    .B(_06087_),
    .Y(_06088_));
 sg13g2_nor2b_1 _15208_ (.A(_06085_),
    .B_N(net246),
    .Y(_06089_));
 sg13g2_a21oi_1 _15209_ (.A1(_06084_),
    .A2(_06088_),
    .Y(_06090_),
    .B1(_06089_));
 sg13g2_buf_2 _15210_ (.A(\vgadonut.donut.cB[9] ),
    .X(_06091_));
 sg13g2_xnor2_1 _15211_ (.Y(_06092_),
    .A(_06091_),
    .B(net245));
 sg13g2_nand2_1 _15212_ (.Y(_06093_),
    .A(_06090_),
    .B(_06092_));
 sg13g2_o21ai_1 _15213_ (.B1(_06036_),
    .Y(_06094_),
    .A1(_06091_),
    .A2(_06035_));
 sg13g2_o21ai_1 _15214_ (.B1(_06094_),
    .Y(_06095_),
    .A1(_06037_),
    .A2(_06093_));
 sg13g2_xnor2_1 _15215_ (.Y(_06096_),
    .A(_06033_),
    .B(net245));
 sg13g2_nand2_1 _15216_ (.Y(_06097_),
    .A(_06095_),
    .B(_06096_));
 sg13g2_o21ai_1 _15217_ (.B1(_06097_),
    .Y(_06098_),
    .A1(_06034_),
    .A2(net245));
 sg13g2_xnor2_1 _15218_ (.Y(_06099_),
    .A(_06031_),
    .B(net245));
 sg13g2_nand2_1 _15219_ (.Y(_06100_),
    .A(_06098_),
    .B(_06099_));
 sg13g2_o21ai_1 _15220_ (.B1(_06100_),
    .Y(_06101_),
    .A1(_06032_),
    .A2(net208));
 sg13g2_buf_2 _15221_ (.A(\vgadonut.donut.cB[13] ),
    .X(_06102_));
 sg13g2_xnor2_1 _15222_ (.Y(_06103_),
    .A(_06102_),
    .B(net245));
 sg13g2_inv_1 _15223_ (.Y(_06104_),
    .A(_06102_));
 sg13g2_nor2_1 _15224_ (.A(net208),
    .B(_06104_),
    .Y(_06105_));
 sg13g2_a21oi_1 _15225_ (.A1(_06101_),
    .A2(_06103_),
    .Y(_06106_),
    .B1(_06105_));
 sg13g2_inv_1 _15226_ (.Y(_06107_),
    .A(_06106_));
 sg13g2_buf_1 _15227_ (.A(\vgadonut.donut.cB[14] ),
    .X(_06108_));
 sg13g2_nor2_1 _15228_ (.A(net228),
    .B(_06036_),
    .Y(_06109_));
 sg13g2_inv_1 _15229_ (.Y(_06110_),
    .A(_06109_));
 sg13g2_inv_1 _15230_ (.Y(_06111_),
    .A(net228));
 sg13g2_nor2_1 _15231_ (.A(net208),
    .B(_06111_),
    .Y(_06112_));
 sg13g2_a21oi_1 _15232_ (.A1(_06107_),
    .A2(_06110_),
    .Y(_06113_),
    .B1(_06112_));
 sg13g2_xnor2_1 _15233_ (.Y(_06114_),
    .A(net197),
    .B(_06113_));
 sg13g2_buf_1 _15234_ (.A(_00146_),
    .X(_06115_));
 sg13g2_xnor2_1 _15235_ (.Y(_06116_),
    .A(_06029_),
    .B(_04603_));
 sg13g2_inv_1 _15236_ (.Y(_06117_),
    .A(_06116_));
 sg13g2_xnor2_1 _15237_ (.Y(_06118_),
    .A(_06117_),
    .B(_06113_));
 sg13g2_buf_1 _15238_ (.A(_06118_),
    .X(_06119_));
 sg13g2_buf_1 _15239_ (.A(_06119_),
    .X(_06120_));
 sg13g2_a21oi_1 _15240_ (.A1(_00145_),
    .A2(_06115_),
    .Y(_06121_),
    .B1(net76));
 sg13g2_xnor2_1 _15241_ (.Y(_06122_),
    .A(net210),
    .B(_06120_));
 sg13g2_inv_1 _15242_ (.Y(_06123_),
    .A(_06122_));
 sg13g2_nor2_1 _15243_ (.A(_06112_),
    .B(_06109_),
    .Y(_06124_));
 sg13g2_xor2_1 _15244_ (.B(_06106_),
    .A(_06124_),
    .X(_06125_));
 sg13g2_nor2_1 _15245_ (.A(_00151_),
    .B(_06125_),
    .Y(_06126_));
 sg13g2_xnor2_1 _15246_ (.Y(_06127_),
    .A(_04312_),
    .B(_06125_));
 sg13g2_inv_1 _15247_ (.Y(_06128_),
    .A(_06127_));
 sg13g2_inv_1 _15248_ (.Y(_06129_),
    .A(_00152_));
 sg13g2_xor2_1 _15249_ (.B(_06101_),
    .A(_06103_),
    .X(_06130_));
 sg13g2_xnor2_1 _15250_ (.Y(_06131_),
    .A(_06039_),
    .B(_06130_));
 sg13g2_buf_1 _15251_ (.A(_00156_),
    .X(_06132_));
 sg13g2_xor2_1 _15252_ (.B(_06090_),
    .A(_06092_),
    .X(_06133_));
 sg13g2_nor2b_1 _15253_ (.A(_06132_),
    .B_N(_06133_),
    .Y(_06134_));
 sg13g2_xnor2_1 _15254_ (.Y(_06135_),
    .A(net250),
    .B(_06133_));
 sg13g2_inv_1 _15255_ (.Y(_06136_),
    .A(_00157_));
 sg13g2_nor2_1 _15256_ (.A(_06087_),
    .B(_06089_),
    .Y(_06137_));
 sg13g2_inv_1 _15257_ (.Y(_06138_),
    .A(_06056_));
 sg13g2_o21ai_1 _15258_ (.B1(_06138_),
    .Y(_06139_),
    .A1(_06057_),
    .A2(_06052_));
 sg13g2_nor2_1 _15259_ (.A(_06062_),
    .B(_06064_),
    .Y(_06140_));
 sg13g2_nand2_1 _15260_ (.Y(_06141_),
    .A(_06139_),
    .B(_06140_));
 sg13g2_nor2_1 _15261_ (.A(_06062_),
    .B(_06069_),
    .Y(_06142_));
 sg13g2_a21oi_1 _15262_ (.A1(_06141_),
    .A2(_06142_),
    .Y(_06143_),
    .B1(_06068_));
 sg13g2_nor2_1 _15263_ (.A(_06076_),
    .B(_06073_),
    .Y(_06144_));
 sg13g2_a221oi_1 _15264_ (.B2(_06144_),
    .C1(_06073_),
    .B1(_06143_),
    .A1(_06078_),
    .Y(_06145_),
    .A2(_06081_));
 sg13g2_nor2_1 _15265_ (.A(_06082_),
    .B(_06145_),
    .Y(_06146_));
 sg13g2_xor2_1 _15266_ (.B(_06146_),
    .A(_06137_),
    .X(_06147_));
 sg13g2_inv_1 _15267_ (.Y(_06148_),
    .A(_04206_));
 sg13g2_xor2_1 _15268_ (.B(_06077_),
    .A(_06083_),
    .X(_06149_));
 sg13g2_xnor2_1 _15269_ (.Y(_06150_),
    .A(_06148_),
    .B(_06149_));
 sg13g2_inv_1 _15270_ (.Y(_06151_),
    .A(_04208_));
 sg13g2_xnor2_1 _15271_ (.Y(_06152_),
    .A(_06144_),
    .B(_06143_));
 sg13g2_nor2_1 _15272_ (.A(_06151_),
    .B(_06152_),
    .Y(_06153_));
 sg13g2_nor2b_1 _15273_ (.A(_06148_),
    .B_N(_06149_),
    .Y(_06154_));
 sg13g2_a21oi_1 _15274_ (.A1(_06150_),
    .A2(_06153_),
    .Y(_06155_),
    .B1(_06154_));
 sg13g2_inv_1 _15275_ (.Y(_06156_),
    .A(_06155_));
 sg13g2_inv_1 _15276_ (.Y(_06157_),
    .A(_04205_));
 sg13g2_xnor2_1 _15277_ (.Y(_06158_),
    .A(_06157_),
    .B(_06147_));
 sg13g2_a22oi_1 _15278_ (.Y(_06159_),
    .B1(_06156_),
    .B2(_06158_),
    .A2(_06147_),
    .A1(_06136_));
 sg13g2_nor2_1 _15279_ (.A(_06135_),
    .B(_06159_),
    .Y(_06160_));
 sg13g2_nor2_1 _15280_ (.A(_06134_),
    .B(_06160_),
    .Y(_06161_));
 sg13g2_inv_1 _15281_ (.Y(_06162_),
    .A(_06161_));
 sg13g2_xor2_1 _15282_ (.B(net245),
    .A(_06035_),
    .X(_06163_));
 sg13g2_nand3_1 _15283_ (.B(_06092_),
    .C(_06137_),
    .A(_06146_),
    .Y(_06164_));
 sg13g2_inv_1 _15284_ (.Y(_06165_),
    .A(_06091_));
 sg13g2_nor2_1 _15285_ (.A(net245),
    .B(_06165_),
    .Y(_06166_));
 sg13g2_a21oi_1 _15286_ (.A1(_06092_),
    .A2(_06087_),
    .Y(_06167_),
    .B1(_06166_));
 sg13g2_nand2_1 _15287_ (.Y(_06168_),
    .A(_06164_),
    .B(_06167_));
 sg13g2_xnor2_1 _15288_ (.Y(_06169_),
    .A(_06163_),
    .B(_06168_));
 sg13g2_xnor2_1 _15289_ (.Y(_06170_),
    .A(net252),
    .B(_06169_));
 sg13g2_inv_1 _15290_ (.Y(_06171_),
    .A(_06170_));
 sg13g2_buf_1 _15291_ (.A(_00155_),
    .X(_06172_));
 sg13g2_nor2b_1 _15292_ (.A(_06172_),
    .B_N(_06169_),
    .Y(_06173_));
 sg13g2_a21oi_1 _15293_ (.A1(_06162_),
    .A2(_06171_),
    .Y(_06174_),
    .B1(_06173_));
 sg13g2_inv_1 _15294_ (.Y(_06175_),
    .A(_06174_));
 sg13g2_xor2_1 _15295_ (.B(_06095_),
    .A(_06096_),
    .X(_06176_));
 sg13g2_xor2_1 _15296_ (.B(_06176_),
    .A(net249),
    .X(_06177_));
 sg13g2_buf_1 _15297_ (.A(_00154_),
    .X(_06178_));
 sg13g2_nor2b_1 _15298_ (.A(_06178_),
    .B_N(_06176_),
    .Y(_06179_));
 sg13g2_a21oi_1 _15299_ (.A1(_06175_),
    .A2(_06177_),
    .Y(_06180_),
    .B1(_06179_));
 sg13g2_inv_1 _15300_ (.Y(_06181_),
    .A(_06180_));
 sg13g2_xor2_1 _15301_ (.B(_06098_),
    .A(_06099_),
    .X(_06182_));
 sg13g2_xnor2_1 _15302_ (.Y(_06183_),
    .A(_06041_),
    .B(_06182_));
 sg13g2_nor2b_1 _15303_ (.A(_00153_),
    .B_N(_06182_),
    .Y(_06184_));
 sg13g2_a21oi_1 _15304_ (.A1(_06181_),
    .A2(_06183_),
    .Y(_06185_),
    .B1(_06184_));
 sg13g2_inv_1 _15305_ (.Y(_06186_),
    .A(_06185_));
 sg13g2_a22oi_1 _15306_ (.Y(_06187_),
    .B1(_06131_),
    .B2(_06186_),
    .A2(_06130_),
    .A1(_06129_));
 sg13g2_nor2_1 _15307_ (.A(_06128_),
    .B(_06187_),
    .Y(_06188_));
 sg13g2_nor2_1 _15308_ (.A(_06126_),
    .B(_06188_),
    .Y(_06189_));
 sg13g2_inv_1 _15309_ (.Y(_06190_),
    .A(_06189_));
 sg13g2_xnor2_1 _15310_ (.Y(_06191_),
    .A(net212),
    .B(_06119_));
 sg13g2_buf_1 _15311_ (.A(_00150_),
    .X(_06192_));
 sg13g2_nor2_1 _15312_ (.A(_06192_),
    .B(_06119_),
    .Y(_06193_));
 sg13g2_a21oi_1 _15313_ (.A1(_06190_),
    .A2(_06191_),
    .Y(_06194_),
    .B1(_06193_));
 sg13g2_xnor2_1 _15314_ (.Y(_06195_),
    .A(net211),
    .B(_06119_));
 sg13g2_nand2b_1 _15315_ (.Y(_06196_),
    .B(_06195_),
    .A_N(_06194_));
 sg13g2_o21ai_1 _15316_ (.B1(_06196_),
    .Y(_06197_),
    .A1(_00149_),
    .A2(net76));
 sg13g2_xnor2_1 _15317_ (.Y(_06198_),
    .A(net247),
    .B(net76));
 sg13g2_nand2_1 _15318_ (.Y(_06199_),
    .A(_06197_),
    .B(_06198_));
 sg13g2_buf_1 _15319_ (.A(_00148_),
    .X(_06200_));
 sg13g2_nor2_1 _15320_ (.A(_06200_),
    .B(net76),
    .Y(_06201_));
 sg13g2_buf_1 _15321_ (.A(_00147_),
    .X(_06202_));
 sg13g2_nor2_1 _15322_ (.A(_06202_),
    .B(net76),
    .Y(_06203_));
 sg13g2_a21oi_1 _15323_ (.A1(_06201_),
    .A2(_06075_),
    .Y(_06204_),
    .B1(_06203_));
 sg13g2_o21ai_1 _15324_ (.B1(_06204_),
    .Y(_06205_),
    .A1(_06123_),
    .A2(_06199_));
 sg13g2_inv_1 _15325_ (.Y(_06206_),
    .A(_00145_));
 sg13g2_xnor2_1 _15326_ (.Y(_06207_),
    .A(_06206_),
    .B(_06120_));
 sg13g2_xnor2_1 _15327_ (.Y(_06208_),
    .A(net209),
    .B(net76));
 sg13g2_nand3_1 _15328_ (.B(_06207_),
    .C(_06208_),
    .A(_06205_),
    .Y(_06209_));
 sg13g2_nand2b_1 _15329_ (.Y(_06210_),
    .B(_06209_),
    .A_N(_06121_));
 sg13g2_xor2_1 _15330_ (.B(_06210_),
    .A(_06114_),
    .X(_06211_));
 sg13g2_nand2_1 _15331_ (.Y(_06212_),
    .A(_06010_),
    .B(\vgadonut.donut.v_count[9] ));
 sg13g2_nor3_1 _15332_ (.A(_06007_),
    .B(_06008_),
    .C(_06212_),
    .Y(_06213_));
 sg13g2_inv_1 _15333_ (.Y(_06214_),
    .A(_06009_));
 sg13g2_nand2_1 _15334_ (.Y(_06215_),
    .A(_06002_),
    .B(_06000_));
 sg13g2_inv_1 _15335_ (.Y(_06216_),
    .A(_06215_));
 sg13g2_nor2_1 _15336_ (.A(_09894_),
    .B(_09832_),
    .Y(_06217_));
 sg13g2_inv_1 _15337_ (.Y(_06218_),
    .A(_06217_));
 sg13g2_nor2_1 _15338_ (.A(_06004_),
    .B(_06218_),
    .Y(_06219_));
 sg13g2_nand4_1 _15339_ (.B(_06214_),
    .C(_06216_),
    .A(_06213_),
    .Y(_06220_),
    .D(_06219_));
 sg13g2_buf_2 _15340_ (.A(_06220_),
    .X(_06221_));
 sg13g2_nor2_2 _15341_ (.A(_10106_),
    .B(_06221_),
    .Y(_06222_));
 sg13g2_inv_1 _15342_ (.Y(_06223_),
    .A(_06222_));
 sg13g2_a21oi_1 _15343_ (.A1(_06211_),
    .A2(net208),
    .Y(_06224_),
    .B1(_06223_));
 sg13g2_buf_1 _15344_ (.A(_06224_),
    .X(_06225_));
 sg13g2_inv_1 _15345_ (.Y(_06226_),
    .A(_06225_));
 sg13g2_buf_1 _15346_ (.A(_06226_),
    .X(_06227_));
 sg13g2_buf_1 _15347_ (.A(net65),
    .X(_06228_));
 sg13g2_buf_2 _15348_ (.A(_06223_),
    .X(_06229_));
 sg13g2_buf_1 _15349_ (.A(_06229_),
    .X(_06230_));
 sg13g2_nand2_1 _15350_ (.Y(_06231_),
    .A(net136),
    .B(_00185_));
 sg13g2_o21ai_1 _15351_ (.B1(_06231_),
    .Y(_00232_),
    .A1(_06028_),
    .A2(net61));
 sg13g2_buf_2 _15352_ (.A(\vgadonut.donut.sA[15] ),
    .X(_06232_));
 sg13g2_buf_1 _15353_ (.A(\vgadonut.donut.cA[10] ),
    .X(_06233_));
 sg13g2_xor2_1 _15354_ (.B(net227),
    .A(_06232_),
    .X(_06234_));
 sg13g2_buf_2 _15355_ (.A(\vgadonut.donut.cA[9] ),
    .X(_06235_));
 sg13g2_buf_1 _15356_ (.A(\vgadonut.donut.sA[14] ),
    .X(_06236_));
 sg13g2_buf_1 _15357_ (.A(_06236_),
    .X(_06237_));
 sg13g2_inv_1 _15358_ (.Y(_06238_),
    .A(net196));
 sg13g2_nor2_1 _15359_ (.A(_06235_),
    .B(_06238_),
    .Y(_06239_));
 sg13g2_inv_1 _15360_ (.Y(_06240_),
    .A(_06235_));
 sg13g2_nor2_1 _15361_ (.A(net196),
    .B(_06240_),
    .Y(_06241_));
 sg13g2_nor2_1 _15362_ (.A(_06239_),
    .B(_06241_),
    .Y(_06242_));
 sg13g2_inv_1 _15363_ (.Y(_06243_),
    .A(_06242_));
 sg13g2_buf_1 _15364_ (.A(\vgadonut.donut.sA[13] ),
    .X(_06244_));
 sg13g2_buf_2 _15365_ (.A(\vgadonut.donut.cA[8] ),
    .X(_06245_));
 sg13g2_xor2_1 _15366_ (.B(_06245_),
    .A(net226),
    .X(_06246_));
 sg13g2_buf_1 _15367_ (.A(\vgadonut.donut.cA[7] ),
    .X(_06247_));
 sg13g2_buf_1 _15368_ (.A(\vgadonut.donut.sA[12] ),
    .X(_06248_));
 sg13g2_inv_2 _15369_ (.Y(_06249_),
    .A(net224));
 sg13g2_nor2_1 _15370_ (.A(net225),
    .B(_06249_),
    .Y(_06250_));
 sg13g2_buf_1 _15371_ (.A(\vgadonut.donut.sA[8] ),
    .X(_06251_));
 sg13g2_buf_2 _15372_ (.A(\vgadonut.donut.cA[3] ),
    .X(_06252_));
 sg13g2_inv_1 _15373_ (.Y(_06253_),
    .A(_06252_));
 sg13g2_nor2_1 _15374_ (.A(net223),
    .B(_06253_),
    .Y(_06254_));
 sg13g2_inv_1 _15375_ (.Y(_06255_),
    .A(net223));
 sg13g2_nor2_1 _15376_ (.A(_06252_),
    .B(_06255_),
    .Y(_06256_));
 sg13g2_buf_1 _15377_ (.A(\vgadonut.donut.sA[7] ),
    .X(_06257_));
 sg13g2_buf_1 _15378_ (.A(_06257_),
    .X(_06258_));
 sg13g2_inv_1 _15379_ (.Y(_06259_),
    .A(net195));
 sg13g2_buf_2 _15380_ (.A(\vgadonut.donut.cA[2] ),
    .X(_06260_));
 sg13g2_buf_1 _15381_ (.A(\vgadonut.donut.sA[6] ),
    .X(_06261_));
 sg13g2_buf_1 _15382_ (.A(_06261_),
    .X(_06262_));
 sg13g2_inv_2 _15383_ (.Y(_06263_),
    .A(net194));
 sg13g2_inv_1 _15384_ (.Y(_06264_),
    .A(net198));
 sg13g2_nor2_1 _15385_ (.A(\vgadonut.donut.cA[0] ),
    .B(_06264_),
    .Y(_06265_));
 sg13g2_xnor2_1 _15386_ (.Y(_06266_),
    .A(net194),
    .B(\vgadonut.donut.cA[1] ));
 sg13g2_nor2b_1 _15387_ (.A(_06265_),
    .B_N(_06266_),
    .Y(_06267_));
 sg13g2_a21oi_1 _15388_ (.A1(_06263_),
    .A2(\vgadonut.donut.cA[1] ),
    .Y(_06268_),
    .B1(_06267_));
 sg13g2_xnor2_1 _15389_ (.Y(_06269_),
    .A(net195),
    .B(_06260_));
 sg13g2_nor2b_1 _15390_ (.A(_06268_),
    .B_N(_06269_),
    .Y(_06270_));
 sg13g2_a21oi_1 _15391_ (.A1(_06259_),
    .A2(_06260_),
    .Y(_06271_),
    .B1(_06270_));
 sg13g2_nor2_1 _15392_ (.A(_06256_),
    .B(_06271_),
    .Y(_06272_));
 sg13g2_or2_1 _15393_ (.X(_06273_),
    .B(_06272_),
    .A(_06254_));
 sg13g2_buf_1 _15394_ (.A(\vgadonut.donut.sA[9] ),
    .X(_06274_));
 sg13g2_buf_1 _15395_ (.A(_06274_),
    .X(_06275_));
 sg13g2_buf_2 _15396_ (.A(\vgadonut.donut.cA[4] ),
    .X(_06276_));
 sg13g2_inv_1 _15397_ (.Y(_06277_),
    .A(_06276_));
 sg13g2_nor2_1 _15398_ (.A(net193),
    .B(_06277_),
    .Y(_06278_));
 sg13g2_inv_1 _15399_ (.Y(_06279_),
    .A(net193));
 sg13g2_nor2_1 _15400_ (.A(_06276_),
    .B(_06279_),
    .Y(_06280_));
 sg13g2_nor2_1 _15401_ (.A(_06278_),
    .B(_06280_),
    .Y(_06281_));
 sg13g2_nand2_1 _15402_ (.Y(_06282_),
    .A(_06273_),
    .B(_06281_));
 sg13g2_buf_1 _15403_ (.A(\vgadonut.donut.sA[10] ),
    .X(_06283_));
 sg13g2_buf_2 _15404_ (.A(\vgadonut.donut.cA[5] ),
    .X(_06284_));
 sg13g2_inv_1 _15405_ (.Y(_06285_),
    .A(_06284_));
 sg13g2_nor2_1 _15406_ (.A(net222),
    .B(_06285_),
    .Y(_06286_));
 sg13g2_nor2_1 _15407_ (.A(_06278_),
    .B(_06286_),
    .Y(_06287_));
 sg13g2_inv_1 _15408_ (.Y(_06288_),
    .A(net222));
 sg13g2_nor2_1 _15409_ (.A(_06284_),
    .B(_06288_),
    .Y(_06289_));
 sg13g2_a21oi_1 _15410_ (.A1(_06282_),
    .A2(_06287_),
    .Y(_06290_),
    .B1(_06289_));
 sg13g2_buf_1 _15411_ (.A(\vgadonut.donut.sA[11] ),
    .X(_06291_));
 sg13g2_buf_2 _15412_ (.A(\vgadonut.donut.cA[6] ),
    .X(_06292_));
 sg13g2_inv_1 _15413_ (.Y(_06293_),
    .A(_06292_));
 sg13g2_nor2_1 _15414_ (.A(net221),
    .B(_06293_),
    .Y(_06294_));
 sg13g2_inv_1 _15415_ (.Y(_06295_),
    .A(net221));
 sg13g2_nor2_1 _15416_ (.A(_06292_),
    .B(_06295_),
    .Y(_06296_));
 sg13g2_nor2_1 _15417_ (.A(_06294_),
    .B(_06296_),
    .Y(_06297_));
 sg13g2_a221oi_1 _15418_ (.B2(_06297_),
    .C1(_06294_),
    .B1(_06290_),
    .A1(_06249_),
    .Y(_06298_),
    .A2(net225));
 sg13g2_nor2_1 _15419_ (.A(_06250_),
    .B(_06298_),
    .Y(_06299_));
 sg13g2_nand2b_1 _15420_ (.Y(_06300_),
    .B(_06299_),
    .A_N(_06246_));
 sg13g2_inv_1 _15421_ (.Y(_06301_),
    .A(_06245_));
 sg13g2_nor2_1 _15422_ (.A(net226),
    .B(_06301_),
    .Y(_06302_));
 sg13g2_a21oi_1 _15423_ (.A1(_06242_),
    .A2(_06302_),
    .Y(_06303_),
    .B1(_06241_));
 sg13g2_o21ai_1 _15424_ (.B1(_06303_),
    .Y(_06304_),
    .A1(_06243_),
    .A2(_06300_));
 sg13g2_xnor2_1 _15425_ (.Y(_06305_),
    .A(_06234_),
    .B(_06304_));
 sg13g2_nand2_1 _15426_ (.Y(_06306_),
    .A(net136),
    .B(_00186_));
 sg13g2_o21ai_1 _15427_ (.B1(_06306_),
    .Y(_00233_),
    .A1(_06305_),
    .A2(_06228_));
 sg13g2_buf_1 _15428_ (.A(\vgadonut.donut.cA[11] ),
    .X(_06307_));
 sg13g2_xnor2_1 _15429_ (.Y(_06308_),
    .A(_06232_),
    .B(net220));
 sg13g2_inv_1 _15430_ (.Y(_06309_),
    .A(_06308_));
 sg13g2_buf_1 _15431_ (.A(_06232_),
    .X(_06310_));
 sg13g2_inv_1 _15432_ (.Y(_06311_),
    .A(net227));
 sg13g2_inv_2 _15433_ (.Y(_06312_),
    .A(_06232_));
 sg13g2_a21oi_1 _15434_ (.A1(_06312_),
    .A2(net227),
    .Y(_06313_),
    .B1(_06241_));
 sg13g2_inv_1 _15435_ (.Y(_06314_),
    .A(net225));
 sg13g2_nor2_1 _15436_ (.A(net224),
    .B(_06314_),
    .Y(_06315_));
 sg13g2_nor2_1 _15437_ (.A(_06302_),
    .B(_06315_),
    .Y(_06316_));
 sg13g2_nor3_1 _15438_ (.A(_06278_),
    .B(_06254_),
    .C(_06272_),
    .Y(_06317_));
 sg13g2_nor2_1 _15439_ (.A(_06280_),
    .B(_06317_),
    .Y(_06318_));
 sg13g2_nor2_1 _15440_ (.A(_06289_),
    .B(_06286_),
    .Y(_06319_));
 sg13g2_nand2_1 _15441_ (.Y(_06320_),
    .A(_06318_),
    .B(_06319_));
 sg13g2_nor2_1 _15442_ (.A(_06294_),
    .B(_06286_),
    .Y(_06321_));
 sg13g2_a21oi_1 _15443_ (.A1(_06320_),
    .A2(_06321_),
    .Y(_06322_),
    .B1(_06296_));
 sg13g2_nor2_1 _15444_ (.A(_06250_),
    .B(_06315_),
    .Y(_06323_));
 sg13g2_nand2_1 _15445_ (.Y(_06324_),
    .A(_06322_),
    .B(_06323_));
 sg13g2_a22oi_1 _15446_ (.Y(_06325_),
    .B1(_06316_),
    .B2(_06324_),
    .A2(_06301_),
    .A1(net226));
 sg13g2_nand2_1 _15447_ (.Y(_06326_),
    .A(_06325_),
    .B(_06242_));
 sg13g2_a22oi_1 _15448_ (.Y(_06327_),
    .B1(_06313_),
    .B2(_06326_),
    .A2(_06311_),
    .A1(net192));
 sg13g2_xnor2_1 _15449_ (.Y(_06328_),
    .A(_06309_),
    .B(_06327_));
 sg13g2_nand2_1 _15450_ (.Y(_06329_),
    .A(net136),
    .B(_00187_));
 sg13g2_o21ai_1 _15451_ (.B1(_06329_),
    .Y(_00234_),
    .A1(_06328_),
    .A2(_06228_));
 sg13g2_buf_2 _15452_ (.A(\vgadonut.donut.cA[12] ),
    .X(_06330_));
 sg13g2_inv_1 _15453_ (.Y(_06331_),
    .A(_06330_));
 sg13g2_nor3_1 _15454_ (.A(_10073_),
    .B(_09884_),
    .C(_05992_),
    .Y(_06332_));
 sg13g2_nand3_1 _15455_ (.B(_10062_),
    .C(_10029_),
    .A(_06332_),
    .Y(_06333_));
 sg13g2_buf_1 _15456_ (.A(_06333_),
    .X(_06334_));
 sg13g2_nor2_1 _15457_ (.A(_06004_),
    .B(_06009_),
    .Y(_06335_));
 sg13g2_inv_1 _15458_ (.Y(_06336_),
    .A(_06007_));
 sg13g2_inv_1 _15459_ (.Y(_06337_),
    .A(_06008_));
 sg13g2_nand3_1 _15460_ (.B(_06336_),
    .C(_06337_),
    .A(_06335_),
    .Y(_06338_));
 sg13g2_nor4_1 _15461_ (.A(_06212_),
    .B(_06218_),
    .C(_06215_),
    .D(_06338_),
    .Y(_06339_));
 sg13g2_inv_2 _15462_ (.Y(_06340_),
    .A(_06339_));
 sg13g2_nor2_1 _15463_ (.A(_06334_),
    .B(_06340_),
    .Y(_06341_));
 sg13g2_buf_1 _15464_ (.A(_06341_),
    .X(_06342_));
 sg13g2_buf_1 _15465_ (.A(_06342_),
    .X(_06343_));
 sg13g2_buf_1 _15466_ (.A(_06225_),
    .X(_06344_));
 sg13g2_buf_1 _15467_ (.A(net67),
    .X(_06345_));
 sg13g2_xnor2_1 _15468_ (.Y(_06346_),
    .A(net192),
    .B(_06330_));
 sg13g2_nand3b_1 _15469_ (.B(_06304_),
    .C(_06308_),
    .Y(_06347_),
    .A_N(_06234_));
 sg13g2_o21ai_1 _15470_ (.B1(_06312_),
    .Y(_06348_),
    .A1(net227),
    .A2(net220));
 sg13g2_nand2_1 _15471_ (.Y(_06349_),
    .A(_06347_),
    .B(_06348_));
 sg13g2_xor2_1 _15472_ (.B(_06349_),
    .A(_06346_),
    .X(_06350_));
 sg13g2_nand2_1 _15473_ (.Y(_06351_),
    .A(net64),
    .B(_06350_));
 sg13g2_o21ai_1 _15474_ (.B1(_06351_),
    .Y(_00235_),
    .A1(_06331_),
    .A2(net154));
 sg13g2_buf_1 _15475_ (.A(\vgadonut.donut.cA[13] ),
    .X(_06352_));
 sg13g2_xnor2_1 _15476_ (.Y(_06353_),
    .A(_06232_),
    .B(net219));
 sg13g2_nand3_1 _15477_ (.B(_06308_),
    .C(_06346_),
    .A(_06327_),
    .Y(_06354_));
 sg13g2_o21ai_1 _15478_ (.B1(_06312_),
    .Y(_06355_),
    .A1(net220),
    .A2(_06330_));
 sg13g2_nand2_1 _15479_ (.Y(_06356_),
    .A(_06354_),
    .B(_06355_));
 sg13g2_xnor2_1 _15480_ (.Y(_06357_),
    .A(_06353_),
    .B(_06356_));
 sg13g2_inv_1 _15481_ (.Y(_06358_),
    .A(_06357_));
 sg13g2_nand2_1 _15482_ (.Y(_06359_),
    .A(net136),
    .B(_00188_));
 sg13g2_o21ai_1 _15483_ (.B1(_06359_),
    .Y(_00236_),
    .A1(_06358_),
    .A2(net61));
 sg13g2_buf_1 _15484_ (.A(\vgadonut.donut.cA[14] ),
    .X(_06360_));
 sg13g2_inv_1 _15485_ (.Y(_06361_),
    .A(net218));
 sg13g2_xnor2_1 _15486_ (.Y(_06362_),
    .A(_06232_),
    .B(net218));
 sg13g2_nand2_1 _15487_ (.Y(_06363_),
    .A(_06346_),
    .B(_06353_));
 sg13g2_inv_1 _15488_ (.Y(_06364_),
    .A(net219));
 sg13g2_a21oi_1 _15489_ (.A1(_06331_),
    .A2(_06364_),
    .Y(_06365_),
    .B1(net192));
 sg13g2_nor2_1 _15490_ (.A(_06348_),
    .B(_06363_),
    .Y(_06366_));
 sg13g2_nor2_1 _15491_ (.A(_06365_),
    .B(_06366_),
    .Y(_06367_));
 sg13g2_o21ai_1 _15492_ (.B1(_06367_),
    .Y(_06368_),
    .A1(_06363_),
    .A2(_06347_));
 sg13g2_xor2_1 _15493_ (.B(_06368_),
    .A(_06362_),
    .X(_06369_));
 sg13g2_nand2_1 _15494_ (.Y(_06370_),
    .A(net64),
    .B(_06369_));
 sg13g2_o21ai_1 _15495_ (.B1(_06370_),
    .Y(_00237_),
    .A1(_06361_),
    .A2(net154));
 sg13g2_buf_2 _15496_ (.A(\vgadonut.donut.cA[15] ),
    .X(_06371_));
 sg13g2_inv_2 _15497_ (.Y(_06372_),
    .A(_06371_));
 sg13g2_xor2_1 _15498_ (.B(_06371_),
    .A(net192),
    .X(_06373_));
 sg13g2_nand2_1 _15499_ (.Y(_06374_),
    .A(_06353_),
    .B(_06362_));
 sg13g2_a21oi_1 _15500_ (.A1(_06364_),
    .A2(_06361_),
    .Y(_06375_),
    .B1(net192));
 sg13g2_nor2_1 _15501_ (.A(_06355_),
    .B(_06374_),
    .Y(_06376_));
 sg13g2_nor2_1 _15502_ (.A(_06375_),
    .B(_06376_),
    .Y(_06377_));
 sg13g2_o21ai_1 _15503_ (.B1(_06377_),
    .Y(_06378_),
    .A1(_06374_),
    .A2(_06354_));
 sg13g2_or2_1 _15504_ (.X(_06379_),
    .B(_06378_),
    .A(_06373_));
 sg13g2_nand2_1 _15505_ (.Y(_06380_),
    .A(_06378_),
    .B(_06373_));
 sg13g2_nand2_1 _15506_ (.Y(_06381_),
    .A(_06379_),
    .B(_06380_));
 sg13g2_buf_2 _15507_ (.A(_06381_),
    .X(_06382_));
 sg13g2_nand2_1 _15508_ (.Y(_06383_),
    .A(net64),
    .B(_06382_));
 sg13g2_o21ai_1 _15509_ (.B1(_06383_),
    .Y(_00238_),
    .A1(_06372_),
    .A2(net154));
 sg13g2_xnor2_1 _15510_ (.Y(_06384_),
    .A(_06265_),
    .B(_06266_));
 sg13g2_nand2_1 _15511_ (.Y(_06385_),
    .A(net136),
    .B(_00189_));
 sg13g2_o21ai_1 _15512_ (.B1(_06385_),
    .Y(_00239_),
    .A1(_06384_),
    .A2(net61));
 sg13g2_xnor2_1 _15513_ (.Y(_06386_),
    .A(_06269_),
    .B(_06268_));
 sg13g2_nand2_1 _15514_ (.Y(_06387_),
    .A(net136),
    .B(_00190_));
 sg13g2_o21ai_1 _15515_ (.B1(_06387_),
    .Y(_00240_),
    .A1(_06386_),
    .A2(net61));
 sg13g2_nor2_1 _15516_ (.A(_06254_),
    .B(_06256_),
    .Y(_06388_));
 sg13g2_xnor2_1 _15517_ (.Y(_06389_),
    .A(_06388_),
    .B(_06271_));
 sg13g2_nand2_1 _15518_ (.Y(_06390_),
    .A(_06230_),
    .B(_00191_));
 sg13g2_o21ai_1 _15519_ (.B1(_06390_),
    .Y(_00241_),
    .A1(_06389_),
    .A2(net61));
 sg13g2_xor2_1 _15520_ (.B(_06273_),
    .A(_06281_),
    .X(_06391_));
 sg13g2_nand2_1 _15521_ (.Y(_06392_),
    .A(_06230_),
    .B(_00192_));
 sg13g2_o21ai_1 _15522_ (.B1(_06392_),
    .Y(_00242_),
    .A1(_06391_),
    .A2(net61));
 sg13g2_xor2_1 _15523_ (.B(_06318_),
    .A(_06319_),
    .X(_06393_));
 sg13g2_buf_1 _15524_ (.A(_06229_),
    .X(_06394_));
 sg13g2_nand2_1 _15525_ (.Y(_06395_),
    .A(net135),
    .B(_00193_));
 sg13g2_o21ai_1 _15526_ (.B1(_06395_),
    .Y(_00243_),
    .A1(_06393_),
    .A2(net61));
 sg13g2_xor2_1 _15527_ (.B(_06290_),
    .A(_06297_),
    .X(_06396_));
 sg13g2_nand2_1 _15528_ (.Y(_06397_),
    .A(net64),
    .B(_06396_));
 sg13g2_o21ai_1 _15529_ (.B1(_06397_),
    .Y(_00244_),
    .A1(_06293_),
    .A2(net154));
 sg13g2_xor2_1 _15530_ (.B(_06322_),
    .A(_06323_),
    .X(_06398_));
 sg13g2_nand2_1 _15531_ (.Y(_06399_),
    .A(net64),
    .B(_06398_));
 sg13g2_o21ai_1 _15532_ (.B1(_06399_),
    .Y(_00245_),
    .A1(_06314_),
    .A2(net154));
 sg13g2_xnor2_1 _15533_ (.Y(_06400_),
    .A(_06246_),
    .B(_06299_));
 sg13g2_nand2_1 _15534_ (.Y(_06401_),
    .A(net135),
    .B(_00194_));
 sg13g2_o21ai_1 _15535_ (.B1(_06401_),
    .Y(_00246_),
    .A1(_06400_),
    .A2(net61));
 sg13g2_xnor2_1 _15536_ (.Y(_06402_),
    .A(_06243_),
    .B(_06325_));
 sg13g2_nand2_1 _15537_ (.Y(_06403_),
    .A(net64),
    .B(_06402_));
 sg13g2_o21ai_1 _15538_ (.B1(_06403_),
    .Y(_00247_),
    .A1(_06240_),
    .A2(net154));
 sg13g2_xnor2_1 _15539_ (.Y(_06404_),
    .A(_05403_),
    .B(net243));
 sg13g2_buf_1 _15540_ (.A(\vgadonut.donut.cAsB[6] ),
    .X(_06405_));
 sg13g2_buf_2 _15541_ (.A(\vgadonut.donut.sAsB[11] ),
    .X(_06406_));
 sg13g2_inv_1 _15542_ (.Y(_06407_),
    .A(_06406_));
 sg13g2_nor2_1 _15543_ (.A(_06405_),
    .B(_06407_),
    .Y(_06408_));
 sg13g2_nor2b_1 _15544_ (.A(_06406_),
    .B_N(_06405_),
    .Y(_06409_));
 sg13g2_inv_1 _15545_ (.Y(_06410_),
    .A(_06409_));
 sg13g2_nand2b_1 _15546_ (.Y(_06411_),
    .B(_06410_),
    .A_N(_06408_));
 sg13g2_buf_2 _15547_ (.A(\vgadonut.donut.cAsB[2] ),
    .X(_06412_));
 sg13g2_inv_1 _15548_ (.Y(_06413_),
    .A(_06412_));
 sg13g2_buf_2 _15549_ (.A(\vgadonut.donut.sAsB[7] ),
    .X(_06414_));
 sg13g2_buf_2 _15550_ (.A(\vgadonut.donut.cAsB[1] ),
    .X(_06415_));
 sg13g2_inv_1 _15551_ (.Y(_06416_),
    .A(_06415_));
 sg13g2_buf_2 _15552_ (.A(\vgadonut.donut.sAsB[6] ),
    .X(_06417_));
 sg13g2_xnor2_1 _15553_ (.Y(_06418_),
    .A(_06415_),
    .B(_06417_));
 sg13g2_buf_1 _15554_ (.A(\vgadonut.donut.cAsB[0] ),
    .X(_06419_));
 sg13g2_buf_2 _15555_ (.A(\vgadonut.donut.sAsB[5] ),
    .X(_06420_));
 sg13g2_nand2b_1 _15556_ (.Y(_06421_),
    .B(_06420_),
    .A_N(net217));
 sg13g2_nand2_1 _15557_ (.Y(_06422_),
    .A(_06418_),
    .B(_06421_));
 sg13g2_o21ai_1 _15558_ (.B1(_06422_),
    .Y(_06423_),
    .A1(_06416_),
    .A2(_06417_));
 sg13g2_xnor2_1 _15559_ (.Y(_06424_),
    .A(_06412_),
    .B(_06414_));
 sg13g2_nand2_1 _15560_ (.Y(_06425_),
    .A(_06423_),
    .B(_06424_));
 sg13g2_o21ai_1 _15561_ (.B1(_06425_),
    .Y(_06426_),
    .A1(_06413_),
    .A2(_06414_));
 sg13g2_buf_1 _15562_ (.A(\vgadonut.donut.cAsB[3] ),
    .X(_06427_));
 sg13g2_buf_2 _15563_ (.A(\vgadonut.donut.sAsB[8] ),
    .X(_06428_));
 sg13g2_xnor2_1 _15564_ (.Y(_06429_),
    .A(_06427_),
    .B(_06428_));
 sg13g2_nor2b_1 _15565_ (.A(_06428_),
    .B_N(_06427_),
    .Y(_06430_));
 sg13g2_a21oi_1 _15566_ (.A1(_06426_),
    .A2(_06429_),
    .Y(_06431_),
    .B1(_06430_));
 sg13g2_inv_1 _15567_ (.Y(_06432_),
    .A(_06431_));
 sg13g2_buf_1 _15568_ (.A(\vgadonut.donut.cAsB[4] ),
    .X(_06433_));
 sg13g2_buf_2 _15569_ (.A(\vgadonut.donut.sAsB[9] ),
    .X(_06434_));
 sg13g2_inv_1 _15570_ (.Y(_06435_),
    .A(_06434_));
 sg13g2_nor2_1 _15571_ (.A(_06433_),
    .B(_06435_),
    .Y(_06436_));
 sg13g2_inv_1 _15572_ (.Y(_06437_),
    .A(_06436_));
 sg13g2_nor2b_1 _15573_ (.A(_06434_),
    .B_N(_06433_),
    .Y(_06438_));
 sg13g2_a21oi_1 _15574_ (.A1(_06432_),
    .A2(_06437_),
    .Y(_06439_),
    .B1(_06438_));
 sg13g2_inv_1 _15575_ (.Y(_06440_),
    .A(_06439_));
 sg13g2_buf_1 _15576_ (.A(\vgadonut.donut.cAsB[5] ),
    .X(_06441_));
 sg13g2_buf_1 _15577_ (.A(\vgadonut.donut.sAsB[10] ),
    .X(_06442_));
 sg13g2_inv_1 _15578_ (.Y(_06443_),
    .A(_06442_));
 sg13g2_nor2_1 _15579_ (.A(_06441_),
    .B(_06443_),
    .Y(_06444_));
 sg13g2_inv_1 _15580_ (.Y(_06445_),
    .A(_06444_));
 sg13g2_inv_1 _15581_ (.Y(_06446_),
    .A(_06441_));
 sg13g2_nor2_1 _15582_ (.A(_06442_),
    .B(_06446_),
    .Y(_06447_));
 sg13g2_a21oi_1 _15583_ (.A1(_06440_),
    .A2(_06445_),
    .Y(_06448_),
    .B1(_06447_));
 sg13g2_xor2_1 _15584_ (.B(_06448_),
    .A(_06411_),
    .X(_06449_));
 sg13g2_buf_1 _15585_ (.A(_06449_),
    .X(_06450_));
 sg13g2_xnor2_1 _15586_ (.Y(_06451_),
    .A(_06404_),
    .B(_06450_));
 sg13g2_buf_1 _15587_ (.A(net65),
    .X(_06452_));
 sg13g2_nand2_1 _15588_ (.Y(_06453_),
    .A(net135),
    .B(_00195_));
 sg13g2_o21ai_1 _15589_ (.B1(_06453_),
    .Y(_00248_),
    .A1(_06451_),
    .A2(_06452_));
 sg13g2_inv_1 _15590_ (.Y(_06454_),
    .A(_05597_));
 sg13g2_nor2_1 _15591_ (.A(_05168_),
    .B(_06454_),
    .Y(_06455_));
 sg13g2_inv_1 _15592_ (.Y(_06456_),
    .A(_05168_));
 sg13g2_nor2_1 _15593_ (.A(_05597_),
    .B(_06456_),
    .Y(_06457_));
 sg13g2_nor2_1 _15594_ (.A(_06455_),
    .B(_06457_),
    .Y(_06458_));
 sg13g2_inv_1 _15595_ (.Y(_06459_),
    .A(_06458_));
 sg13g2_inv_1 _15596_ (.Y(_06460_),
    .A(net234));
 sg13g2_nor2_1 _15597_ (.A(net238),
    .B(_06460_),
    .Y(_06461_));
 sg13g2_inv_1 _15598_ (.Y(_06462_),
    .A(net237));
 sg13g2_nor2_1 _15599_ (.A(net240),
    .B(_06462_),
    .Y(_06463_));
 sg13g2_inv_1 _15600_ (.Y(_06464_),
    .A(net236));
 sg13g2_xnor2_1 _15601_ (.Y(_06465_),
    .A(_05396_),
    .B(net244));
 sg13g2_nand2_1 _15602_ (.Y(_06466_),
    .A(_05404_),
    .B(net243));
 sg13g2_nand2_1 _15603_ (.Y(_06467_),
    .A(_06465_),
    .B(_06466_));
 sg13g2_o21ai_1 _15604_ (.B1(_06467_),
    .Y(_06468_),
    .A1(_05400_),
    .A2(net244));
 sg13g2_xnor2_1 _15605_ (.Y(_06469_),
    .A(_05390_),
    .B(net242));
 sg13g2_nand2_1 _15606_ (.Y(_06470_),
    .A(_06468_),
    .B(_06469_));
 sg13g2_o21ai_1 _15607_ (.B1(_06470_),
    .Y(_06471_),
    .A1(_05405_),
    .A2(net242));
 sg13g2_xnor2_1 _15608_ (.Y(_06472_),
    .A(_05380_),
    .B(net241));
 sg13g2_nand2_1 _15609_ (.Y(_06473_),
    .A(_06471_),
    .B(_06472_));
 sg13g2_o21ai_1 _15610_ (.B1(_06473_),
    .Y(_06474_),
    .A1(_05401_),
    .A2(net241));
 sg13g2_xnor2_1 _15611_ (.Y(_06475_),
    .A(net236),
    .B(net207));
 sg13g2_nand2_1 _15612_ (.Y(_06476_),
    .A(_06474_),
    .B(_06475_));
 sg13g2_o21ai_1 _15613_ (.B1(_06476_),
    .Y(_06477_),
    .A1(_06464_),
    .A2(net207));
 sg13g2_inv_1 _15614_ (.Y(_06478_),
    .A(net240));
 sg13g2_nor2_1 _15615_ (.A(net237),
    .B(_06478_),
    .Y(_06479_));
 sg13g2_inv_1 _15616_ (.Y(_06480_),
    .A(_06479_));
 sg13g2_o21ai_1 _15617_ (.B1(_06480_),
    .Y(_06481_),
    .A1(_06463_),
    .A2(_06477_));
 sg13g2_inv_1 _15618_ (.Y(_06482_),
    .A(net235));
 sg13g2_nor2_1 _15619_ (.A(net239),
    .B(_06482_),
    .Y(_06483_));
 sg13g2_inv_1 _15620_ (.Y(_06484_),
    .A(_06483_));
 sg13g2_inv_1 _15621_ (.Y(_06485_),
    .A(net239));
 sg13g2_nor2_1 _15622_ (.A(net235),
    .B(_06485_),
    .Y(_06486_));
 sg13g2_a21oi_1 _15623_ (.A1(_06481_),
    .A2(_06484_),
    .Y(_06487_),
    .B1(_06486_));
 sg13g2_inv_1 _15624_ (.Y(_06488_),
    .A(net238));
 sg13g2_nor2_1 _15625_ (.A(net234),
    .B(_06488_),
    .Y(_06489_));
 sg13g2_inv_1 _15626_ (.Y(_06490_),
    .A(_06489_));
 sg13g2_o21ai_1 _15627_ (.B1(_06490_),
    .Y(_06491_),
    .A1(_06461_),
    .A2(_06487_));
 sg13g2_inv_1 _15628_ (.Y(_06492_),
    .A(_06491_));
 sg13g2_xnor2_1 _15629_ (.Y(_06493_),
    .A(_05553_),
    .B(_05134_));
 sg13g2_inv_1 _15630_ (.Y(_06494_),
    .A(\vgadonut.donut.cAcB[8] ));
 sg13g2_nor2_1 _15631_ (.A(net206),
    .B(_06494_),
    .Y(_06495_));
 sg13g2_inv_1 _15632_ (.Y(_06496_),
    .A(net206));
 sg13g2_nor2_1 _15633_ (.A(_05505_),
    .B(_06496_),
    .Y(_06497_));
 sg13g2_nor2_1 _15634_ (.A(_06495_),
    .B(_06497_),
    .Y(_06498_));
 sg13g2_nand3_1 _15635_ (.B(_06493_),
    .C(_06498_),
    .A(_06492_),
    .Y(_06499_));
 sg13g2_inv_1 _15636_ (.Y(_06500_),
    .A(_05553_));
 sg13g2_nor2_1 _15637_ (.A(net205),
    .B(_06500_),
    .Y(_06501_));
 sg13g2_a21oi_1 _15638_ (.A1(_06493_),
    .A2(_06495_),
    .Y(_06502_),
    .B1(_06501_));
 sg13g2_nand2_1 _15639_ (.Y(_06503_),
    .A(_06499_),
    .B(_06502_));
 sg13g2_xnor2_1 _15640_ (.Y(_06504_),
    .A(_06459_),
    .B(_06503_));
 sg13g2_buf_2 _15641_ (.A(\vgadonut.donut.cAsB[15] ),
    .X(_06505_));
 sg13g2_inv_1 _15642_ (.Y(_06506_),
    .A(_06505_));
 sg13g2_buf_1 _15643_ (.A(_06506_),
    .X(_06507_));
 sg13g2_buf_1 _15644_ (.A(\vgadonut.donut.cAsB[14] ),
    .X(_06508_));
 sg13g2_buf_1 _15645_ (.A(\vgadonut.donut.sAsB[15] ),
    .X(_06509_));
 sg13g2_buf_1 _15646_ (.A(_06509_),
    .X(_06510_));
 sg13g2_nand2_1 _15647_ (.Y(_06511_),
    .A(_06508_),
    .B(net191));
 sg13g2_inv_1 _15648_ (.Y(_06512_),
    .A(_06511_));
 sg13g2_buf_1 _15649_ (.A(\vgadonut.donut.cAsB[13] ),
    .X(_06513_));
 sg13g2_inv_1 _15650_ (.Y(_06514_),
    .A(_06513_));
 sg13g2_buf_1 _15651_ (.A(\vgadonut.donut.cAsB[10] ),
    .X(_06515_));
 sg13g2_inv_1 _15652_ (.Y(_06516_),
    .A(_06515_));
 sg13g2_inv_1 _15653_ (.Y(_06517_),
    .A(_06509_));
 sg13g2_buf_1 _15654_ (.A(\vgadonut.donut.sAsB[14] ),
    .X(_06518_));
 sg13g2_buf_1 _15655_ (.A(\vgadonut.donut.cAsB[9] ),
    .X(_06519_));
 sg13g2_inv_1 _15656_ (.Y(_06520_),
    .A(_06519_));
 sg13g2_nor2_1 _15657_ (.A(_06518_),
    .B(_06520_),
    .Y(_06521_));
 sg13g2_a21oi_1 _15658_ (.A1(_06515_),
    .A2(_06517_),
    .Y(_06522_),
    .B1(_06521_));
 sg13g2_o21ai_1 _15659_ (.B1(_06410_),
    .Y(_06523_),
    .A1(_06408_),
    .A2(_06448_));
 sg13g2_buf_1 _15660_ (.A(_06523_),
    .X(_06524_));
 sg13g2_buf_1 _15661_ (.A(\vgadonut.donut.sAsB[12] ),
    .X(_06525_));
 sg13g2_buf_1 _15662_ (.A(\vgadonut.donut.cAsB[7] ),
    .X(_06526_));
 sg13g2_inv_1 _15663_ (.Y(_06527_),
    .A(_06526_));
 sg13g2_nor2_1 _15664_ (.A(_06525_),
    .B(_06527_),
    .Y(_06528_));
 sg13g2_inv_1 _15665_ (.Y(_06529_),
    .A(_06525_));
 sg13g2_nor2_1 _15666_ (.A(_06526_),
    .B(_06529_),
    .Y(_06530_));
 sg13g2_nor2_1 _15667_ (.A(_06528_),
    .B(_06530_),
    .Y(_06531_));
 sg13g2_nand2_1 _15668_ (.Y(_06532_),
    .A(_06524_),
    .B(_06531_));
 sg13g2_buf_1 _15669_ (.A(\vgadonut.donut.sAsB[13] ),
    .X(_06533_));
 sg13g2_buf_1 _15670_ (.A(\vgadonut.donut.cAsB[8] ),
    .X(_06534_));
 sg13g2_inv_1 _15671_ (.Y(_06535_),
    .A(_06534_));
 sg13g2_nor2_1 _15672_ (.A(_06533_),
    .B(_06535_),
    .Y(_06536_));
 sg13g2_nor2_1 _15673_ (.A(_06528_),
    .B(_06536_),
    .Y(_06537_));
 sg13g2_inv_1 _15674_ (.Y(_06538_),
    .A(_06533_));
 sg13g2_nor2_1 _15675_ (.A(_06534_),
    .B(_06538_),
    .Y(_06539_));
 sg13g2_a21oi_1 _15676_ (.A1(_06532_),
    .A2(_06537_),
    .Y(_06540_),
    .B1(_06539_));
 sg13g2_inv_1 _15677_ (.Y(_06541_),
    .A(_06518_));
 sg13g2_nor2_1 _15678_ (.A(_06519_),
    .B(_06541_),
    .Y(_06542_));
 sg13g2_nor2_1 _15679_ (.A(_06521_),
    .B(_06542_),
    .Y(_06543_));
 sg13g2_nand2_1 _15680_ (.Y(_06544_),
    .A(_06540_),
    .B(_06543_));
 sg13g2_a22oi_1 _15681_ (.Y(_06545_),
    .B1(_06522_),
    .B2(_06544_),
    .A2(_06510_),
    .A1(_06516_));
 sg13g2_buf_1 _15682_ (.A(\vgadonut.donut.cAsB[11] ),
    .X(_06546_));
 sg13g2_xnor2_1 _15683_ (.Y(_06547_),
    .A(_06546_),
    .B(_06509_));
 sg13g2_inv_1 _15684_ (.Y(_06548_),
    .A(_06546_));
 sg13g2_nor2_1 _15685_ (.A(net191),
    .B(_06548_),
    .Y(_06549_));
 sg13g2_a21oi_1 _15686_ (.A1(_06545_),
    .A2(_06547_),
    .Y(_06550_),
    .B1(_06549_));
 sg13g2_inv_1 _15687_ (.Y(_06551_),
    .A(_06550_));
 sg13g2_buf_1 _15688_ (.A(\vgadonut.donut.cAsB[12] ),
    .X(_06552_));
 sg13g2_nor2_1 _15689_ (.A(_06552_),
    .B(_06517_),
    .Y(_06553_));
 sg13g2_inv_1 _15690_ (.Y(_06554_),
    .A(_06553_));
 sg13g2_inv_1 _15691_ (.Y(_06555_),
    .A(_06552_));
 sg13g2_nor2_1 _15692_ (.A(net191),
    .B(_06555_),
    .Y(_06556_));
 sg13g2_a21oi_1 _15693_ (.A1(_06551_),
    .A2(_06554_),
    .Y(_06557_),
    .B1(_06556_));
 sg13g2_xnor2_1 _15694_ (.Y(_06558_),
    .A(_06513_),
    .B(net191));
 sg13g2_nand2b_1 _15695_ (.Y(_06559_),
    .B(_06558_),
    .A_N(_06557_));
 sg13g2_o21ai_1 _15696_ (.B1(_06559_),
    .Y(_06560_),
    .A1(_06514_),
    .A2(net191));
 sg13g2_buf_1 _15697_ (.A(_06560_),
    .X(_06561_));
 sg13g2_nor2_1 _15698_ (.A(_06508_),
    .B(_06510_),
    .Y(_06562_));
 sg13g2_nor2b_1 _15699_ (.A(_06561_),
    .B_N(_06562_),
    .Y(_06563_));
 sg13g2_a21oi_1 _15700_ (.A1(_06512_),
    .A2(_06561_),
    .Y(_06564_),
    .B1(_06563_));
 sg13g2_xnor2_1 _15701_ (.Y(_06565_),
    .A(net184),
    .B(_06564_));
 sg13g2_buf_1 _15702_ (.A(_06565_),
    .X(_06566_));
 sg13g2_buf_1 _15703_ (.A(_06566_),
    .X(_06567_));
 sg13g2_nor2_1 _15704_ (.A(_06504_),
    .B(net75),
    .Y(_06568_));
 sg13g2_inv_1 _15705_ (.Y(_06569_),
    .A(_06504_));
 sg13g2_inv_1 _15706_ (.Y(_06570_),
    .A(_06566_));
 sg13g2_buf_1 _15707_ (.A(_06570_),
    .X(_06571_));
 sg13g2_nor2_1 _15708_ (.A(_06569_),
    .B(net74),
    .Y(_06572_));
 sg13g2_nor2_1 _15709_ (.A(_06568_),
    .B(_06572_),
    .Y(_06573_));
 sg13g2_xnor2_1 _15710_ (.Y(_06574_),
    .A(_06558_),
    .B(_06557_));
 sg13g2_buf_2 _15711_ (.A(_06574_),
    .X(_06575_));
 sg13g2_nand2b_1 _15712_ (.Y(_06576_),
    .B(_06490_),
    .A_N(_06461_));
 sg13g2_xor2_1 _15713_ (.B(_06487_),
    .A(_06576_),
    .X(_06577_));
 sg13g2_inv_1 _15714_ (.Y(_06578_),
    .A(_06575_));
 sg13g2_inv_1 _15715_ (.Y(_06579_),
    .A(_06577_));
 sg13g2_nor2_1 _15716_ (.A(_06479_),
    .B(_06463_),
    .Y(_06580_));
 sg13g2_xnor2_1 _15717_ (.Y(_06581_),
    .A(_06580_),
    .B(_06477_));
 sg13g2_inv_1 _15718_ (.Y(_06582_),
    .A(_06581_));
 sg13g2_xnor2_1 _15719_ (.Y(_06583_),
    .A(_06547_),
    .B(_06545_));
 sg13g2_buf_2 _15720_ (.A(_06583_),
    .X(_06584_));
 sg13g2_nor2_1 _15721_ (.A(_06582_),
    .B(_06584_),
    .Y(_06585_));
 sg13g2_xor2_1 _15722_ (.B(_06524_),
    .A(_06531_),
    .X(_06586_));
 sg13g2_buf_2 _15723_ (.A(_06586_),
    .X(_06587_));
 sg13g2_xnor2_1 _15724_ (.Y(_06588_),
    .A(_06466_),
    .B(_06465_));
 sg13g2_nand2_1 _15725_ (.Y(_06589_),
    .A(_06587_),
    .B(_06588_));
 sg13g2_nand2_1 _15726_ (.Y(_06590_),
    .A(_06450_),
    .B(_06404_));
 sg13g2_nor2_1 _15727_ (.A(_06588_),
    .B(_06587_),
    .Y(_06591_));
 sg13g2_a21oi_1 _15728_ (.A1(_06589_),
    .A2(_06590_),
    .Y(_06592_),
    .B1(_06591_));
 sg13g2_inv_1 _15729_ (.Y(_06593_),
    .A(_06592_));
 sg13g2_xnor2_1 _15730_ (.Y(_06594_),
    .A(_06469_),
    .B(_06468_));
 sg13g2_nor2_1 _15731_ (.A(_06539_),
    .B(_06536_),
    .Y(_06595_));
 sg13g2_inv_1 _15732_ (.Y(_06596_),
    .A(_06530_));
 sg13g2_a21oi_1 _15733_ (.A1(_06524_),
    .A2(_06596_),
    .Y(_06597_),
    .B1(_06528_));
 sg13g2_xnor2_1 _15734_ (.Y(_06598_),
    .A(_06595_),
    .B(_06597_));
 sg13g2_buf_2 _15735_ (.A(_06598_),
    .X(_06599_));
 sg13g2_xor2_1 _15736_ (.B(_06599_),
    .A(_06594_),
    .X(_06600_));
 sg13g2_nor2_1 _15737_ (.A(_06594_),
    .B(_06599_),
    .Y(_06601_));
 sg13g2_a21oi_1 _15738_ (.A1(_06593_),
    .A2(_06600_),
    .Y(_06602_),
    .B1(_06601_));
 sg13g2_xor2_1 _15739_ (.B(_06540_),
    .A(_06543_),
    .X(_06603_));
 sg13g2_xnor2_1 _15740_ (.Y(_06604_),
    .A(_06472_),
    .B(_06471_));
 sg13g2_nand2_1 _15741_ (.Y(_06605_),
    .A(_06603_),
    .B(_06604_));
 sg13g2_nand2b_1 _15742_ (.Y(_06606_),
    .B(_06605_),
    .A_N(_06602_));
 sg13g2_nor2_1 _15743_ (.A(_06604_),
    .B(_06603_),
    .Y(_06607_));
 sg13g2_inv_1 _15744_ (.Y(_06608_),
    .A(_06607_));
 sg13g2_nand2_1 _15745_ (.Y(_06609_),
    .A(_06606_),
    .B(_06608_));
 sg13g2_xor2_1 _15746_ (.B(net191),
    .A(_06515_),
    .X(_06610_));
 sg13g2_nand2b_1 _15747_ (.Y(_06611_),
    .B(_06595_),
    .A_N(_06597_));
 sg13g2_nor2_1 _15748_ (.A(_06521_),
    .B(_06536_),
    .Y(_06612_));
 sg13g2_a21oi_1 _15749_ (.A1(_06611_),
    .A2(_06612_),
    .Y(_06613_),
    .B1(_06542_));
 sg13g2_xor2_1 _15750_ (.B(_06613_),
    .A(_06610_),
    .X(_06614_));
 sg13g2_inv_1 _15751_ (.Y(_06615_),
    .A(_06614_));
 sg13g2_xor2_1 _15752_ (.B(_06474_),
    .A(_06475_),
    .X(_06616_));
 sg13g2_inv_1 _15753_ (.Y(_06617_),
    .A(_06616_));
 sg13g2_nand2_1 _15754_ (.Y(_06618_),
    .A(_06615_),
    .B(_06617_));
 sg13g2_nor2_1 _15755_ (.A(_06617_),
    .B(_06615_),
    .Y(_06619_));
 sg13g2_a221oi_1 _15756_ (.B2(_06618_),
    .C1(_06619_),
    .B1(_06609_),
    .A1(_06584_),
    .Y(_06620_),
    .A2(_06582_));
 sg13g2_nor2_1 _15757_ (.A(_06585_),
    .B(_06620_),
    .Y(_06621_));
 sg13g2_nand2b_1 _15758_ (.Y(_06622_),
    .B(_06484_),
    .A_N(_06486_));
 sg13g2_xnor2_1 _15759_ (.Y(_06623_),
    .A(_06622_),
    .B(_06481_));
 sg13g2_inv_1 _15760_ (.Y(_06624_),
    .A(_06623_));
 sg13g2_nand2b_1 _15761_ (.Y(_06625_),
    .B(_06554_),
    .A_N(_06556_));
 sg13g2_xnor2_1 _15762_ (.Y(_06626_),
    .A(_06625_),
    .B(_06550_));
 sg13g2_nor2_1 _15763_ (.A(_06624_),
    .B(_06626_),
    .Y(_06627_));
 sg13g2_inv_1 _15764_ (.Y(_06628_),
    .A(_06626_));
 sg13g2_nor2_1 _15765_ (.A(_06623_),
    .B(_06628_),
    .Y(_06629_));
 sg13g2_nor2_1 _15766_ (.A(_06627_),
    .B(_06629_),
    .Y(_06630_));
 sg13g2_a221oi_1 _15767_ (.B2(_06630_),
    .C1(_06629_),
    .B1(_06621_),
    .A1(_06578_),
    .Y(_06631_),
    .A2(_06579_));
 sg13g2_a21oi_1 _15768_ (.A1(_06575_),
    .A2(_06577_),
    .Y(_06632_),
    .B1(_06631_));
 sg13g2_xnor2_1 _15769_ (.Y(_06633_),
    .A(_06498_),
    .B(_06491_));
 sg13g2_inv_1 _15770_ (.Y(_06634_),
    .A(_06633_));
 sg13g2_nor2_1 _15771_ (.A(_06562_),
    .B(_06512_),
    .Y(_06635_));
 sg13g2_xor2_1 _15772_ (.B(_06561_),
    .A(_06635_),
    .X(_06636_));
 sg13g2_buf_1 _15773_ (.A(_06636_),
    .X(_06637_));
 sg13g2_xnor2_1 _15774_ (.Y(_06638_),
    .A(_06634_),
    .B(_06637_));
 sg13g2_inv_1 _15775_ (.Y(_06639_),
    .A(_06637_));
 sg13g2_nor2_1 _15776_ (.A(_06634_),
    .B(_06639_),
    .Y(_06640_));
 sg13g2_a21oi_1 _15777_ (.A1(_06632_),
    .A2(_06638_),
    .Y(_06641_),
    .B1(_06640_));
 sg13g2_inv_1 _15778_ (.Y(_06642_),
    .A(_06641_));
 sg13g2_inv_1 _15779_ (.Y(_06643_),
    .A(_06497_));
 sg13g2_a21oi_1 _15780_ (.A1(_06492_),
    .A2(_06643_),
    .Y(_06644_),
    .B1(_06495_));
 sg13g2_xnor2_1 _15781_ (.Y(_06645_),
    .A(_06493_),
    .B(_06644_));
 sg13g2_nor2_1 _15782_ (.A(_06645_),
    .B(net75),
    .Y(_06646_));
 sg13g2_inv_1 _15783_ (.Y(_06647_),
    .A(_06645_));
 sg13g2_nor2_1 _15784_ (.A(_06647_),
    .B(net74),
    .Y(_06648_));
 sg13g2_nor2_1 _15785_ (.A(_06646_),
    .B(_06648_),
    .Y(_06649_));
 sg13g2_a21oi_1 _15786_ (.A1(_06642_),
    .A2(_06649_),
    .Y(_06650_),
    .B1(_06648_));
 sg13g2_xnor2_1 _15787_ (.Y(_06651_),
    .A(_06573_),
    .B(_06650_));
 sg13g2_nand2_1 _15788_ (.Y(_06652_),
    .A(net135),
    .B(_00196_));
 sg13g2_o21ai_1 _15789_ (.B1(_06652_),
    .Y(_00249_),
    .A1(_06651_),
    .A2(net60));
 sg13g2_xnor2_1 _15790_ (.Y(_06653_),
    .A(_05642_),
    .B(_05168_));
 sg13g2_inv_1 _15791_ (.Y(_06654_),
    .A(_06653_));
 sg13g2_nand2_1 _15792_ (.Y(_06655_),
    .A(_06458_),
    .B(_06493_));
 sg13g2_a21oi_1 _15793_ (.A1(_06458_),
    .A2(_06501_),
    .Y(_06656_),
    .B1(_06455_));
 sg13g2_o21ai_1 _15794_ (.B1(_06656_),
    .Y(_06657_),
    .A1(_06655_),
    .A2(_06644_));
 sg13g2_xnor2_1 _15795_ (.Y(_06658_),
    .A(_06654_),
    .B(_06657_));
 sg13g2_nor2_1 _15796_ (.A(_06658_),
    .B(net75),
    .Y(_06659_));
 sg13g2_inv_1 _15797_ (.Y(_06660_),
    .A(_06658_));
 sg13g2_nor2_1 _15798_ (.A(_06660_),
    .B(net74),
    .Y(_06661_));
 sg13g2_nor2_1 _15799_ (.A(_06659_),
    .B(_06661_),
    .Y(_06662_));
 sg13g2_inv_1 _15800_ (.Y(_06663_),
    .A(_06572_));
 sg13g2_o21ai_1 _15801_ (.B1(_06663_),
    .Y(_06664_),
    .A1(_06568_),
    .A2(_06650_));
 sg13g2_xor2_1 _15802_ (.B(_06664_),
    .A(_06662_),
    .X(_06665_));
 sg13g2_nand2_1 _15803_ (.Y(_06666_),
    .A(net135),
    .B(_00197_));
 sg13g2_o21ai_1 _15804_ (.B1(_06666_),
    .Y(_00250_),
    .A1(_06665_),
    .A2(net60));
 sg13g2_inv_1 _15805_ (.Y(_06667_),
    .A(_05693_));
 sg13g2_xnor2_1 _15806_ (.Y(_06668_),
    .A(_05693_),
    .B(_05168_));
 sg13g2_inv_1 _15807_ (.Y(_06669_),
    .A(_06668_));
 sg13g2_nand3_1 _15808_ (.B(_06458_),
    .C(_06653_),
    .A(_06503_),
    .Y(_06670_));
 sg13g2_o21ai_1 _15809_ (.B1(_06456_),
    .Y(_06671_),
    .A1(_05598_),
    .A2(_05642_));
 sg13g2_nand2_1 _15810_ (.Y(_06672_),
    .A(_06670_),
    .B(_06671_));
 sg13g2_xnor2_1 _15811_ (.Y(_06673_),
    .A(_06669_),
    .B(_06672_));
 sg13g2_nor2_1 _15812_ (.A(_06673_),
    .B(net75),
    .Y(_06674_));
 sg13g2_inv_1 _15813_ (.Y(_06675_),
    .A(_06673_));
 sg13g2_nor2_1 _15814_ (.A(_06675_),
    .B(net74),
    .Y(_06676_));
 sg13g2_nor2_1 _15815_ (.A(_06674_),
    .B(_06676_),
    .Y(_06677_));
 sg13g2_nor2b_1 _15816_ (.A(_06650_),
    .B_N(_06573_),
    .Y(_06678_));
 sg13g2_a221oi_1 _15817_ (.B2(_06662_),
    .C1(_06661_),
    .B1(_06678_),
    .A1(net75),
    .Y(_06679_),
    .A2(_06504_));
 sg13g2_xnor2_1 _15818_ (.Y(_06680_),
    .A(_06677_),
    .B(_06679_));
 sg13g2_nand2_1 _15819_ (.Y(_06681_),
    .A(net64),
    .B(_06680_));
 sg13g2_o21ai_1 _15820_ (.B1(_06681_),
    .Y(_00251_),
    .A1(_06667_),
    .A2(net154));
 sg13g2_xnor2_1 _15821_ (.Y(_06682_),
    .A(_05729_),
    .B(_05168_));
 sg13g2_inv_1 _15822_ (.Y(_06683_),
    .A(_06682_));
 sg13g2_nand3_1 _15823_ (.B(_06653_),
    .C(_06668_),
    .A(_06657_),
    .Y(_06684_));
 sg13g2_o21ai_1 _15824_ (.B1(_06456_),
    .Y(_06685_),
    .A1(net202),
    .A2(_05693_));
 sg13g2_nand2_1 _15825_ (.Y(_06686_),
    .A(_06684_),
    .B(_06685_));
 sg13g2_xnor2_1 _15826_ (.Y(_06687_),
    .A(_06683_),
    .B(_06686_));
 sg13g2_inv_1 _15827_ (.Y(_06688_),
    .A(_06687_));
 sg13g2_xnor2_1 _15828_ (.Y(_06689_),
    .A(_06688_),
    .B(net75));
 sg13g2_nand2_1 _15829_ (.Y(_06690_),
    .A(_06664_),
    .B(_06662_));
 sg13g2_nor2_1 _15830_ (.A(_06661_),
    .B(_06676_),
    .Y(_06691_));
 sg13g2_o21ai_1 _15831_ (.B1(_06691_),
    .Y(_06692_),
    .A1(_06674_),
    .A2(_06690_));
 sg13g2_xor2_1 _15832_ (.B(_06692_),
    .A(_06689_),
    .X(_06693_));
 sg13g2_nand2_1 _15833_ (.Y(_06694_),
    .A(net135),
    .B(_00198_));
 sg13g2_o21ai_1 _15834_ (.B1(_06694_),
    .Y(_00252_),
    .A1(_06693_),
    .A2(net60));
 sg13g2_inv_1 _15835_ (.Y(_06695_),
    .A(_05772_));
 sg13g2_xnor2_1 _15836_ (.Y(_06696_),
    .A(_05772_),
    .B(_05168_));
 sg13g2_nand2_1 _15837_ (.Y(_06697_),
    .A(_06668_),
    .B(_06682_));
 sg13g2_inv_1 _15838_ (.Y(_06698_),
    .A(net200));
 sg13g2_a21oi_1 _15839_ (.A1(_06667_),
    .A2(_06698_),
    .Y(_06699_),
    .B1(net204));
 sg13g2_nor2_1 _15840_ (.A(_06671_),
    .B(_06697_),
    .Y(_06700_));
 sg13g2_nor2_1 _15841_ (.A(_06699_),
    .B(_06700_),
    .Y(_06701_));
 sg13g2_o21ai_1 _15842_ (.B1(_06701_),
    .Y(_06702_),
    .A1(_06697_),
    .A2(_06670_));
 sg13g2_xnor2_1 _15843_ (.Y(_06703_),
    .A(_06696_),
    .B(_06702_));
 sg13g2_xnor2_1 _15844_ (.Y(_06704_),
    .A(_06703_),
    .B(_06567_));
 sg13g2_inv_1 _15845_ (.Y(_06705_),
    .A(_06704_));
 sg13g2_nand3b_1 _15846_ (.B(_06677_),
    .C(_06689_),
    .Y(_06706_),
    .A_N(_06679_));
 sg13g2_nor2_1 _15847_ (.A(_06688_),
    .B(_06571_),
    .Y(_06707_));
 sg13g2_inv_1 _15848_ (.Y(_06708_),
    .A(_06707_));
 sg13g2_nand3b_1 _15849_ (.B(_06706_),
    .C(_06708_),
    .Y(_06709_),
    .A_N(_06676_));
 sg13g2_xnor2_1 _15850_ (.Y(_06710_),
    .A(_06705_),
    .B(_06709_));
 sg13g2_nand2_1 _15851_ (.Y(_06711_),
    .A(net64),
    .B(_06710_));
 sg13g2_o21ai_1 _15852_ (.B1(_06711_),
    .Y(_00253_),
    .A1(_06695_),
    .A2(net154));
 sg13g2_nand2_1 _15853_ (.Y(_06712_),
    .A(_06682_),
    .B(_06696_));
 sg13g2_inv_1 _15854_ (.Y(_06713_),
    .A(_06712_));
 sg13g2_inv_1 _15855_ (.Y(_06714_),
    .A(_06685_));
 sg13g2_a21oi_1 _15856_ (.A1(_06698_),
    .A2(_06695_),
    .Y(_06715_),
    .B1(net204));
 sg13g2_a21oi_1 _15857_ (.A1(_06713_),
    .A2(_06714_),
    .Y(_06716_),
    .B1(_06715_));
 sg13g2_o21ai_1 _15858_ (.B1(_06716_),
    .Y(_06717_),
    .A1(_06712_),
    .A2(_06684_));
 sg13g2_xor2_1 _15859_ (.B(net204),
    .A(_05807_),
    .X(_06718_));
 sg13g2_nand2b_1 _15860_ (.Y(_06719_),
    .B(_06718_),
    .A_N(_06717_));
 sg13g2_nand2b_1 _15861_ (.Y(_06720_),
    .B(_06717_),
    .A_N(_06718_));
 sg13g2_nand2_1 _15862_ (.Y(_06721_),
    .A(_06719_),
    .B(_06720_));
 sg13g2_buf_1 _15863_ (.A(_06721_),
    .X(_06722_));
 sg13g2_inv_1 _15864_ (.Y(_06723_),
    .A(net77));
 sg13g2_xnor2_1 _15865_ (.Y(_06724_),
    .A(_06723_),
    .B(_06567_));
 sg13g2_a21oi_1 _15866_ (.A1(_06688_),
    .A2(_06703_),
    .Y(_06725_),
    .B1(_06571_));
 sg13g2_nand3_1 _15867_ (.B(_06689_),
    .C(_06704_),
    .A(_06692_),
    .Y(_06726_));
 sg13g2_nor2b_1 _15868_ (.A(_06725_),
    .B_N(_06726_),
    .Y(_06727_));
 sg13g2_or2_1 _15869_ (.X(_06728_),
    .B(_06727_),
    .A(_06724_));
 sg13g2_nand2_1 _15870_ (.Y(_06729_),
    .A(_06727_),
    .B(_06724_));
 sg13g2_nand2_1 _15871_ (.Y(_06730_),
    .A(_06728_),
    .B(_06729_));
 sg13g2_buf_1 _15872_ (.A(_06730_),
    .X(_06731_));
 sg13g2_nand2_1 _15873_ (.Y(_06732_),
    .A(net135),
    .B(_05807_));
 sg13g2_o21ai_1 _15874_ (.B1(_06732_),
    .Y(_00254_),
    .A1(_06731_),
    .A2(net60));
 sg13g2_xnor2_1 _15875_ (.Y(_06733_),
    .A(_06588_),
    .B(_06587_));
 sg13g2_xnor2_1 _15876_ (.Y(_06734_),
    .A(_06590_),
    .B(_06733_));
 sg13g2_nand2_1 _15877_ (.Y(_06735_),
    .A(net135),
    .B(_00199_));
 sg13g2_o21ai_1 _15878_ (.B1(_06735_),
    .Y(_00255_),
    .A1(_06734_),
    .A2(net60));
 sg13g2_xnor2_1 _15879_ (.Y(_06736_),
    .A(_06592_),
    .B(_06600_));
 sg13g2_nand2_1 _15880_ (.Y(_06737_),
    .A(_06394_),
    .B(_00200_));
 sg13g2_o21ai_1 _15881_ (.B1(_06737_),
    .Y(_00256_),
    .A1(_06736_),
    .A2(_06452_));
 sg13g2_nand2_1 _15882_ (.Y(_06738_),
    .A(_06608_),
    .B(_06605_));
 sg13g2_xor2_1 _15883_ (.B(_06602_),
    .A(_06738_),
    .X(_06739_));
 sg13g2_nand2_1 _15884_ (.Y(_06740_),
    .A(_06394_),
    .B(_00201_));
 sg13g2_o21ai_1 _15885_ (.B1(_06740_),
    .Y(_00257_),
    .A1(_06739_),
    .A2(net60));
 sg13g2_nand2b_1 _15886_ (.Y(_06741_),
    .B(_06618_),
    .A_N(_06619_));
 sg13g2_xnor2_1 _15887_ (.Y(_06742_),
    .A(_06741_),
    .B(_06609_));
 sg13g2_buf_1 _15888_ (.A(_06229_),
    .X(_06743_));
 sg13g2_nand2_1 _15889_ (.Y(_06744_),
    .A(net134),
    .B(_00202_));
 sg13g2_o21ai_1 _15890_ (.B1(_06744_),
    .Y(_00258_),
    .A1(_06742_),
    .A2(net60));
 sg13g2_nand2_1 _15891_ (.Y(_06745_),
    .A(_06584_),
    .B(_06582_));
 sg13g2_nor2b_1 _15892_ (.A(_06585_),
    .B_N(_06745_),
    .Y(_06746_));
 sg13g2_nand3b_1 _15893_ (.B(_06606_),
    .C(_06608_),
    .Y(_06747_),
    .A_N(_06619_));
 sg13g2_and2_1 _15894_ (.A(_06747_),
    .B(_06618_),
    .X(_06748_));
 sg13g2_xor2_1 _15895_ (.B(_06748_),
    .A(_06746_),
    .X(_06749_));
 sg13g2_nand2_1 _15896_ (.Y(_06750_),
    .A(_06743_),
    .B(_00203_));
 sg13g2_o21ai_1 _15897_ (.B1(_06750_),
    .Y(_00259_),
    .A1(_06749_),
    .A2(net60));
 sg13g2_xor2_1 _15898_ (.B(_06621_),
    .A(_06630_),
    .X(_06751_));
 sg13g2_nand2_1 _15899_ (.Y(_06752_),
    .A(_06345_),
    .B(_06751_));
 sg13g2_o21ai_1 _15900_ (.B1(_06752_),
    .Y(_00260_),
    .A1(_06482_),
    .A2(_06343_));
 sg13g2_buf_1 _15901_ (.A(net67),
    .X(_06753_));
 sg13g2_xnor2_1 _15902_ (.Y(_06754_),
    .A(_06579_),
    .B(_06575_));
 sg13g2_nand2_1 _15903_ (.Y(_06755_),
    .A(_06748_),
    .B(_06746_));
 sg13g2_nor2b_1 _15904_ (.A(_06629_),
    .B_N(_06745_),
    .Y(_06756_));
 sg13g2_a21oi_1 _15905_ (.A1(_06755_),
    .A2(_06756_),
    .Y(_06757_),
    .B1(_06627_));
 sg13g2_xor2_1 _15906_ (.B(_06757_),
    .A(_06754_),
    .X(_06758_));
 sg13g2_nand2_1 _15907_ (.Y(_06759_),
    .A(net63),
    .B(_06758_));
 sg13g2_o21ai_1 _15908_ (.B1(_06759_),
    .Y(_00261_),
    .A1(_06460_),
    .A2(_06343_));
 sg13g2_xor2_1 _15909_ (.B(_06632_),
    .A(_06638_),
    .X(_06760_));
 sg13g2_buf_1 _15910_ (.A(_06227_),
    .X(_06761_));
 sg13g2_nand2_1 _15911_ (.Y(_06762_),
    .A(net134),
    .B(_00204_));
 sg13g2_o21ai_1 _15912_ (.B1(_06762_),
    .Y(_00262_),
    .A1(_06760_),
    .A2(net59));
 sg13g2_buf_1 _15913_ (.A(_06342_),
    .X(_06763_));
 sg13g2_xnor2_1 _15914_ (.Y(_06764_),
    .A(_06649_),
    .B(_06641_));
 sg13g2_nand2_1 _15915_ (.Y(_06765_),
    .A(net63),
    .B(_06764_));
 sg13g2_o21ai_1 _15916_ (.B1(_06765_),
    .Y(_00263_),
    .A1(_06500_),
    .A2(net153));
 sg13g2_xnor2_1 _15917_ (.Y(_06766_),
    .A(net217),
    .B(_06420_));
 sg13g2_xor2_1 _15918_ (.B(_06751_),
    .A(_06766_),
    .X(_06767_));
 sg13g2_nand2_1 _15919_ (.Y(_06768_),
    .A(net134),
    .B(net217));
 sg13g2_o21ai_1 _15920_ (.B1(_06768_),
    .Y(_00264_),
    .A1(_06767_),
    .A2(net59));
 sg13g2_xnor2_1 _15921_ (.Y(_06769_),
    .A(_06615_),
    .B(net68));
 sg13g2_inv_1 _15922_ (.Y(_06770_),
    .A(_06769_));
 sg13g2_inv_1 _15923_ (.Y(_06771_),
    .A(net68));
 sg13g2_xnor2_1 _15924_ (.Y(_06772_),
    .A(_06603_),
    .B(net68));
 sg13g2_inv_1 _15925_ (.Y(_06773_),
    .A(_06772_));
 sg13g2_xnor2_1 _15926_ (.Y(_06774_),
    .A(_06599_),
    .B(_06710_));
 sg13g2_inv_1 _15927_ (.Y(_06775_),
    .A(_06450_));
 sg13g2_nor2b_1 _15928_ (.A(_06775_),
    .B_N(_06680_),
    .Y(_06776_));
 sg13g2_nor2_1 _15929_ (.A(_06450_),
    .B(_06680_),
    .Y(_06777_));
 sg13g2_nor2_1 _15930_ (.A(_06436_),
    .B(_06438_),
    .Y(_06778_));
 sg13g2_xnor2_1 _15931_ (.Y(_06779_),
    .A(_06778_),
    .B(_06431_));
 sg13g2_xor2_1 _15932_ (.B(_06426_),
    .A(_06429_),
    .X(_06780_));
 sg13g2_nand2_1 _15933_ (.Y(_06781_),
    .A(_06764_),
    .B(_06780_));
 sg13g2_xor2_1 _15934_ (.B(_06423_),
    .A(_06424_),
    .X(_06782_));
 sg13g2_xor2_1 _15935_ (.B(_06760_),
    .A(_06782_),
    .X(_06783_));
 sg13g2_xor2_1 _15936_ (.B(_06418_),
    .A(_06421_),
    .X(_06784_));
 sg13g2_nor2b_1 _15937_ (.A(_06766_),
    .B_N(_06751_),
    .Y(_06785_));
 sg13g2_inv_1 _15938_ (.Y(_06786_),
    .A(_06785_));
 sg13g2_xor2_1 _15939_ (.B(_06758_),
    .A(_06784_),
    .X(_06787_));
 sg13g2_inv_1 _15940_ (.Y(_06788_),
    .A(_06787_));
 sg13g2_nor2_1 _15941_ (.A(_06786_),
    .B(_06788_),
    .Y(_06789_));
 sg13g2_a21o_1 _15942_ (.A2(_06784_),
    .A1(_06758_),
    .B1(_06789_),
    .X(_06790_));
 sg13g2_nand2_1 _15943_ (.Y(_06791_),
    .A(_06783_),
    .B(_06790_));
 sg13g2_nand2_1 _15944_ (.Y(_06792_),
    .A(_06760_),
    .B(_06782_));
 sg13g2_nand2_1 _15945_ (.Y(_06793_),
    .A(_06791_),
    .B(_06792_));
 sg13g2_or2_1 _15946_ (.X(_06794_),
    .B(_06764_),
    .A(_06780_));
 sg13g2_nand3_1 _15947_ (.B(_06781_),
    .C(_06794_),
    .A(_06793_),
    .Y(_06795_));
 sg13g2_buf_1 _15948_ (.A(_06795_),
    .X(_06796_));
 sg13g2_xor2_1 _15949_ (.B(_06651_),
    .A(_06779_),
    .X(_06797_));
 sg13g2_inv_1 _15950_ (.Y(_06798_),
    .A(_06797_));
 sg13g2_a21oi_1 _15951_ (.A1(_06781_),
    .A2(_06796_),
    .Y(_06799_),
    .B1(_06798_));
 sg13g2_a21o_1 _15952_ (.A2(_06779_),
    .A1(_06651_),
    .B1(_06799_),
    .X(_06800_));
 sg13g2_nand2b_1 _15953_ (.Y(_06801_),
    .B(_06445_),
    .A_N(_06447_));
 sg13g2_xor2_1 _15954_ (.B(_06439_),
    .A(_06801_),
    .X(_06802_));
 sg13g2_inv_1 _15955_ (.Y(_06803_),
    .A(_06802_));
 sg13g2_xnor2_1 _15956_ (.Y(_06804_),
    .A(_06803_),
    .B(_06665_));
 sg13g2_nor2b_1 _15957_ (.A(_06803_),
    .B_N(_06665_),
    .Y(_06805_));
 sg13g2_a21oi_1 _15958_ (.A1(_06800_),
    .A2(_06804_),
    .Y(_06806_),
    .B1(_06805_));
 sg13g2_nor2_1 _15959_ (.A(_06777_),
    .B(_06806_),
    .Y(_06807_));
 sg13g2_nor2_1 _15960_ (.A(_06776_),
    .B(_06807_),
    .Y(_06808_));
 sg13g2_nand2_1 _15961_ (.Y(_06809_),
    .A(_06693_),
    .B(_06587_));
 sg13g2_nor2_1 _15962_ (.A(_06587_),
    .B(_06693_),
    .Y(_06810_));
 sg13g2_a21oi_1 _15963_ (.A1(_06808_),
    .A2(_06809_),
    .Y(_06811_),
    .B1(_06810_));
 sg13g2_inv_1 _15964_ (.Y(_06812_),
    .A(_06811_));
 sg13g2_nor2_1 _15965_ (.A(_06774_),
    .B(_06812_),
    .Y(_06813_));
 sg13g2_a21oi_1 _15966_ (.A1(_06599_),
    .A2(_06710_),
    .Y(_06814_),
    .B1(_06813_));
 sg13g2_nor2_1 _15967_ (.A(_06773_),
    .B(_06814_),
    .Y(_06815_));
 sg13g2_a21oi_1 _15968_ (.A1(_06603_),
    .A2(_06771_),
    .Y(_06816_),
    .B1(_06815_));
 sg13g2_nor2_1 _15969_ (.A(_06770_),
    .B(_06816_),
    .Y(_06817_));
 sg13g2_buf_1 _15970_ (.A(_06225_),
    .X(_06818_));
 sg13g2_nand2_1 _15971_ (.Y(_06819_),
    .A(_06816_),
    .B(_06770_));
 sg13g2_nand3b_1 _15972_ (.B(net66),
    .C(_06819_),
    .Y(_06820_),
    .A_N(_06817_));
 sg13g2_o21ai_1 _15973_ (.B1(_06820_),
    .Y(_00265_),
    .A1(_06516_),
    .A2(net153));
 sg13g2_xnor2_1 _15974_ (.Y(_06821_),
    .A(_06584_),
    .B(net68));
 sg13g2_a21oi_1 _15975_ (.A1(_06615_),
    .A2(_06771_),
    .Y(_06822_),
    .B1(_06817_));
 sg13g2_nor2_1 _15976_ (.A(_06821_),
    .B(_06822_),
    .Y(_06823_));
 sg13g2_nand2_1 _15977_ (.Y(_06824_),
    .A(_06822_),
    .B(_06821_));
 sg13g2_nand3b_1 _15978_ (.B(_06818_),
    .C(_06824_),
    .Y(_06825_),
    .A_N(_06823_));
 sg13g2_o21ai_1 _15979_ (.B1(_06825_),
    .Y(_00266_),
    .A1(_06548_),
    .A2(net153));
 sg13g2_nor2_1 _15980_ (.A(_06584_),
    .B(net68),
    .Y(_06826_));
 sg13g2_nor2_1 _15981_ (.A(_06826_),
    .B(_06823_),
    .Y(_06827_));
 sg13g2_inv_1 _15982_ (.Y(_06828_),
    .A(_06827_));
 sg13g2_nor2_1 _15983_ (.A(_06626_),
    .B(net68),
    .Y(_06829_));
 sg13g2_nor2_1 _15984_ (.A(_06628_),
    .B(_06771_),
    .Y(_06830_));
 sg13g2_nor2_1 _15985_ (.A(_06829_),
    .B(_06830_),
    .Y(_06831_));
 sg13g2_buf_1 _15986_ (.A(_06226_),
    .X(_06832_));
 sg13g2_a21oi_1 _15987_ (.A1(_06828_),
    .A2(_06831_),
    .Y(_06833_),
    .B1(net62));
 sg13g2_o21ai_1 _15988_ (.B1(_06833_),
    .Y(_06834_),
    .A1(_06828_),
    .A2(_06831_));
 sg13g2_o21ai_1 _15989_ (.B1(_06834_),
    .Y(_00267_),
    .A1(_06555_),
    .A2(_06763_));
 sg13g2_xnor2_1 _15990_ (.Y(_06835_),
    .A(_06575_),
    .B(net68));
 sg13g2_inv_1 _15991_ (.Y(_06836_),
    .A(_06829_));
 sg13g2_o21ai_1 _15992_ (.B1(_06836_),
    .Y(_06837_),
    .A1(_06830_),
    .A2(_06827_));
 sg13g2_inv_1 _15993_ (.Y(_06838_),
    .A(_06835_));
 sg13g2_inv_1 _15994_ (.Y(_06839_),
    .A(_06837_));
 sg13g2_nor2_1 _15995_ (.A(_06838_),
    .B(_06839_),
    .Y(_06840_));
 sg13g2_nor2_1 _15996_ (.A(net62),
    .B(_06840_),
    .Y(_06841_));
 sg13g2_o21ai_1 _15997_ (.B1(_06841_),
    .Y(_06842_),
    .A1(_06835_),
    .A2(_06837_));
 sg13g2_o21ai_1 _15998_ (.B1(_06842_),
    .Y(_00268_),
    .A1(_06514_),
    .A2(_06763_));
 sg13g2_inv_1 _15999_ (.Y(_06843_),
    .A(_06508_));
 sg13g2_a21oi_1 _16000_ (.A1(_06575_),
    .A2(_06771_),
    .Y(_06844_),
    .B1(_06840_));
 sg13g2_inv_1 _16001_ (.Y(_06845_),
    .A(_06844_));
 sg13g2_nor2_1 _16002_ (.A(_06637_),
    .B(net68),
    .Y(_06846_));
 sg13g2_nor2_1 _16003_ (.A(_06639_),
    .B(_06771_),
    .Y(_06847_));
 sg13g2_nor2_1 _16004_ (.A(_06846_),
    .B(_06847_),
    .Y(_06848_));
 sg13g2_a21oi_1 _16005_ (.A1(_06845_),
    .A2(_06848_),
    .Y(_06849_),
    .B1(_06226_));
 sg13g2_o21ai_1 _16006_ (.B1(_06849_),
    .Y(_06850_),
    .A1(_06845_),
    .A2(_06848_));
 sg13g2_o21ai_1 _16007_ (.B1(_06850_),
    .Y(_00269_),
    .A1(_06843_),
    .A2(net153));
 sg13g2_xnor2_1 _16008_ (.Y(_06851_),
    .A(_06723_),
    .B(_06727_));
 sg13g2_inv_1 _16009_ (.Y(_06852_),
    .A(_06847_));
 sg13g2_a21oi_1 _16010_ (.A1(_06845_),
    .A2(_06852_),
    .Y(_06853_),
    .B1(_06846_));
 sg13g2_a21oi_1 _16011_ (.A1(_06853_),
    .A2(_06851_),
    .Y(_06854_),
    .B1(_06226_));
 sg13g2_o21ai_1 _16012_ (.B1(_06854_),
    .Y(_06855_),
    .A1(_06851_),
    .A2(_06853_));
 sg13g2_o21ai_1 _16013_ (.B1(_06855_),
    .Y(_00270_),
    .A1(net184),
    .A2(net153));
 sg13g2_nand2_1 _16014_ (.Y(_06856_),
    .A(_06788_),
    .B(_06786_));
 sg13g2_nand3b_1 _16015_ (.B(_06818_),
    .C(_06856_),
    .Y(_06857_),
    .A_N(_06789_));
 sg13g2_o21ai_1 _16016_ (.B1(_06857_),
    .Y(_00271_),
    .A1(_06416_),
    .A2(net153));
 sg13g2_xnor2_1 _16017_ (.Y(_06858_),
    .A(_06790_),
    .B(_06783_));
 sg13g2_nand2_1 _16018_ (.Y(_06859_),
    .A(net134),
    .B(_06412_));
 sg13g2_o21ai_1 _16019_ (.B1(_06859_),
    .Y(_00272_),
    .A1(_06858_),
    .A2(net59));
 sg13g2_a21oi_1 _16020_ (.A1(_06794_),
    .A2(_06781_),
    .Y(_06860_),
    .B1(_06793_));
 sg13g2_nand2b_1 _16021_ (.Y(_06861_),
    .B(_06796_),
    .A_N(_06860_));
 sg13g2_nand2_1 _16022_ (.Y(_06862_),
    .A(net134),
    .B(_06427_));
 sg13g2_o21ai_1 _16023_ (.B1(_06862_),
    .Y(_00273_),
    .A1(_06861_),
    .A2(net59));
 sg13g2_nand3_1 _16024_ (.B(_06781_),
    .C(_06796_),
    .A(_06798_),
    .Y(_06863_));
 sg13g2_nand2b_1 _16025_ (.Y(_06864_),
    .B(_06863_),
    .A_N(_06799_));
 sg13g2_nand2_1 _16026_ (.Y(_06865_),
    .A(net134),
    .B(_06433_));
 sg13g2_o21ai_1 _16027_ (.B1(_06865_),
    .Y(_00274_),
    .A1(_06864_),
    .A2(net59));
 sg13g2_xnor2_1 _16028_ (.Y(_06866_),
    .A(_06804_),
    .B(_06800_));
 sg13g2_nand2_1 _16029_ (.Y(_06867_),
    .A(net134),
    .B(_06441_));
 sg13g2_o21ai_1 _16030_ (.B1(_06867_),
    .Y(_00275_),
    .A1(_06866_),
    .A2(net59));
 sg13g2_buf_1 _16031_ (.A(_06832_),
    .X(_06868_));
 sg13g2_nor2_1 _16032_ (.A(_06777_),
    .B(_06776_),
    .Y(_06869_));
 sg13g2_xor2_1 _16033_ (.B(_06806_),
    .A(_06869_),
    .X(_06870_));
 sg13g2_nand2_1 _16034_ (.Y(_06871_),
    .A(net134),
    .B(_06405_));
 sg13g2_o21ai_1 _16035_ (.B1(_06871_),
    .Y(_00276_),
    .A1(_06868_),
    .A2(_06870_));
 sg13g2_nor2b_1 _16036_ (.A(_06810_),
    .B_N(_06809_),
    .Y(_06872_));
 sg13g2_o21ai_1 _16037_ (.B1(_06872_),
    .Y(_06873_),
    .A1(_06776_),
    .A2(_06807_));
 sg13g2_nand2b_1 _16038_ (.Y(_06874_),
    .B(_06808_),
    .A_N(_06872_));
 sg13g2_nand3_1 _16039_ (.B(_06874_),
    .C(net67),
    .A(_06873_),
    .Y(_06875_));
 sg13g2_o21ai_1 _16040_ (.B1(_06875_),
    .Y(_00277_),
    .A1(_06527_),
    .A2(net153));
 sg13g2_nand2_1 _16041_ (.Y(_06876_),
    .A(_06812_),
    .B(_06774_));
 sg13g2_nand3b_1 _16042_ (.B(_06344_),
    .C(_06876_),
    .Y(_06877_),
    .A_N(_06813_));
 sg13g2_o21ai_1 _16043_ (.B1(_06877_),
    .Y(_00278_),
    .A1(_06535_),
    .A2(net153));
 sg13g2_buf_1 _16044_ (.A(net166),
    .X(_06878_));
 sg13g2_a21oi_1 _16045_ (.A1(_06814_),
    .A2(_06773_),
    .Y(_06879_),
    .B1(_06832_));
 sg13g2_nand2b_1 _16046_ (.Y(_06880_),
    .B(_06879_),
    .A_N(_06815_));
 sg13g2_o21ai_1 _16047_ (.B1(_06880_),
    .Y(_00279_),
    .A1(_06520_),
    .A2(_06878_));
 sg13g2_inv_1 _16048_ (.Y(_06881_),
    .A(_06211_));
 sg13g2_o21ai_1 _16049_ (.B1(_06041_),
    .Y(_06882_),
    .A1(_06036_),
    .A2(_06881_));
 sg13g2_inv_1 _16050_ (.Y(_06883_),
    .A(_06040_));
 sg13g2_a21oi_1 _16051_ (.A1(_06882_),
    .A2(_06222_),
    .Y(_06884_),
    .B1(_06883_));
 sg13g2_a21o_1 _16052_ (.A2(_06345_),
    .A1(_06042_),
    .B1(_06884_),
    .X(_00280_));
 sg13g2_inv_1 _16053_ (.Y(_06885_),
    .A(_06035_));
 sg13g2_nand2_1 _16054_ (.Y(_06886_),
    .A(net63),
    .B(_06169_));
 sg13g2_o21ai_1 _16055_ (.B1(_06886_),
    .Y(_00281_),
    .A1(_06885_),
    .A2(net152));
 sg13g2_nand2_1 _16056_ (.Y(_06887_),
    .A(net63),
    .B(_06176_));
 sg13g2_o21ai_1 _16057_ (.B1(_06887_),
    .Y(_00282_),
    .A1(_06034_),
    .A2(net152));
 sg13g2_nand2_1 _16058_ (.Y(_06888_),
    .A(net63),
    .B(_06182_));
 sg13g2_o21ai_1 _16059_ (.B1(_06888_),
    .Y(_00283_),
    .A1(_06032_),
    .A2(net152));
 sg13g2_nand2_1 _16060_ (.Y(_06889_),
    .A(net63),
    .B(_06130_));
 sg13g2_o21ai_1 _16061_ (.B1(_06889_),
    .Y(_00284_),
    .A1(_06104_),
    .A2(net152));
 sg13g2_inv_1 _16062_ (.Y(_06890_),
    .A(_00205_));
 sg13g2_nand2_1 _16063_ (.Y(_06891_),
    .A(net63),
    .B(_06125_));
 sg13g2_o21ai_1 _16064_ (.B1(_06891_),
    .Y(_00285_),
    .A1(_06890_),
    .A2(net152));
 sg13g2_buf_1 _16065_ (.A(_06030_),
    .X(_06892_));
 sg13g2_nand2_1 _16066_ (.Y(_06893_),
    .A(_06743_),
    .B(net183));
 sg13g2_o21ai_1 _16067_ (.B1(_06893_),
    .Y(_00286_),
    .A1(net76),
    .A2(net59));
 sg13g2_inv_1 _16068_ (.Y(_06894_),
    .A(net231));
 sg13g2_nor2b_1 _16069_ (.A(_06043_),
    .B_N(_06042_),
    .Y(_06895_));
 sg13g2_nor3_1 _16070_ (.A(_06044_),
    .B(_06895_),
    .C(_06223_),
    .Y(_06896_));
 sg13g2_o21ai_1 _16071_ (.B1(_06896_),
    .Y(_06897_),
    .A1(_06036_),
    .A2(_06881_));
 sg13g2_o21ai_1 _16072_ (.B1(_06897_),
    .Y(_00287_),
    .A1(_06894_),
    .A2(net152));
 sg13g2_nor2_1 _16073_ (.A(_06049_),
    .B(_06051_),
    .Y(_06898_));
 sg13g2_xor2_1 _16074_ (.B(_06045_),
    .A(_06898_),
    .X(_06899_));
 sg13g2_buf_1 _16075_ (.A(_06229_),
    .X(_06900_));
 sg13g2_buf_1 _16076_ (.A(_06047_),
    .X(_06901_));
 sg13g2_nand2_1 _16077_ (.Y(_06902_),
    .A(net133),
    .B(net190));
 sg13g2_o21ai_1 _16078_ (.B1(_06902_),
    .Y(_00288_),
    .A1(_06899_),
    .A2(net59));
 sg13g2_xor2_1 _16079_ (.B(_06052_),
    .A(_06058_),
    .X(_06903_));
 sg13g2_nand2_1 _16080_ (.Y(_06904_),
    .A(net133),
    .B(net229));
 sg13g2_o21ai_1 _16081_ (.B1(_06904_),
    .Y(_00289_),
    .A1(_06903_),
    .A2(_06761_));
 sg13g2_xnor2_1 _16082_ (.Y(_06905_),
    .A(_06140_),
    .B(_06139_));
 sg13g2_nand2_1 _16083_ (.Y(_06906_),
    .A(net133),
    .B(_06060_));
 sg13g2_o21ai_1 _16084_ (.B1(_06906_),
    .Y(_00290_),
    .A1(_06905_),
    .A2(_06761_));
 sg13g2_xnor2_1 _16085_ (.Y(_06907_),
    .A(_06070_),
    .B(_06065_));
 sg13g2_buf_1 _16086_ (.A(net62),
    .X(_06908_));
 sg13g2_nand2_1 _16087_ (.Y(_06909_),
    .A(_06900_),
    .B(_06066_));
 sg13g2_o21ai_1 _16088_ (.B1(_06909_),
    .Y(_00291_),
    .A1(_06907_),
    .A2(_06908_));
 sg13g2_nand2_1 _16089_ (.Y(_06910_),
    .A(_06900_),
    .B(_06072_));
 sg13g2_o21ai_1 _16090_ (.B1(_06910_),
    .Y(_00292_),
    .A1(_06152_),
    .A2(_06908_));
 sg13g2_nand2_1 _16091_ (.Y(_06911_),
    .A(net63),
    .B(_06149_));
 sg13g2_o21ai_1 _16092_ (.B1(_06911_),
    .Y(_00293_),
    .A1(_06079_),
    .A2(net152));
 sg13g2_nand2_1 _16093_ (.Y(_06912_),
    .A(_06753_),
    .B(_06147_));
 sg13g2_o21ai_1 _16094_ (.B1(_06912_),
    .Y(_00294_),
    .A1(_06086_),
    .A2(net152));
 sg13g2_nand2_1 _16095_ (.Y(_06913_),
    .A(_06753_),
    .B(_06133_));
 sg13g2_o21ai_1 _16096_ (.B1(_06913_),
    .Y(_00295_),
    .A1(_06165_),
    .A2(_06878_));
 sg13g2_buf_1 _16097_ (.A(\vgadonut.donut.donut_visible ),
    .X(_06914_));
 sg13g2_inv_2 _16098_ (.Y(_06915_),
    .A(_06914_));
 sg13g2_buf_1 _16099_ (.A(_06915_),
    .X(_06916_));
 sg13g2_nor2_1 _16100_ (.A(\vgadonut.donut.donuthit.hit ),
    .B(net106),
    .Y(_06917_));
 sg13g2_a21oi_1 _16101_ (.A1(_06916_),
    .A2(net106),
    .Y(_00296_),
    .B1(_06917_));
 sg13g2_buf_1 _16102_ (.A(net125),
    .X(_06918_));
 sg13g2_buf_1 _16103_ (.A(net138),
    .X(_06919_));
 sg13g2_nand2_1 _16104_ (.Y(_06920_),
    .A(net120),
    .B(\vgadonut.donut.donuthit.rx[10] ));
 sg13g2_o21ai_1 _16105_ (.B1(_06920_),
    .Y(_00298_),
    .A1(_04451_),
    .A2(net109));
 sg13g2_nand2_1 _16106_ (.Y(_06921_),
    .A(net120),
    .B(\vgadonut.donut.donuthit.rx[11] ));
 sg13g2_o21ai_1 _16107_ (.B1(_06921_),
    .Y(_00299_),
    .A1(_04494_),
    .A2(net109));
 sg13g2_inv_1 _16108_ (.Y(_06922_),
    .A(_04532_));
 sg13g2_nand2_1 _16109_ (.Y(_06923_),
    .A(net120),
    .B(\vgadonut.donut.donuthit.rx[12] ));
 sg13g2_o21ai_1 _16110_ (.B1(_06923_),
    .Y(_00300_),
    .A1(_06922_),
    .A2(net109));
 sg13g2_nand2_1 _16111_ (.Y(_06924_),
    .A(net120),
    .B(\vgadonut.donut.donuthit.rx[13] ));
 sg13g2_o21ai_1 _16112_ (.B1(_06924_),
    .Y(_00301_),
    .A1(_04572_),
    .A2(net109));
 sg13g2_nand2_1 _16113_ (.Y(_06925_),
    .A(net120),
    .B(\vgadonut.donut.donuthit.rx[14] ));
 sg13g2_o21ai_1 _16114_ (.B1(_06925_),
    .Y(_00302_),
    .A1(_04601_),
    .A2(net109));
 sg13g2_nand2_1 _16115_ (.Y(_06926_),
    .A(net120),
    .B(\vgadonut.donut.donuthit.rx[15] ));
 sg13g2_o21ai_1 _16116_ (.B1(_06926_),
    .Y(_00303_),
    .A1(_04704_),
    .A2(net109));
 sg13g2_buf_1 _16117_ (.A(_04305_),
    .X(_06927_));
 sg13g2_nand2_1 _16118_ (.Y(_06928_),
    .A(net119),
    .B(\vgadonut.donut.donuthit.rx[5] ));
 sg13g2_o21ai_1 _16119_ (.B1(_06928_),
    .Y(_00304_),
    .A1(_04196_),
    .A2(net109));
 sg13g2_nand2_1 _16120_ (.Y(_06929_),
    .A(net119),
    .B(\vgadonut.donut.donuthit.rx[6] ));
 sg13g2_o21ai_1 _16121_ (.B1(_06929_),
    .Y(_00305_),
    .A1(_04307_),
    .A2(net109));
 sg13g2_buf_1 _16122_ (.A(_04303_),
    .X(_06930_));
 sg13g2_nand2_1 _16123_ (.Y(_06931_),
    .A(net119),
    .B(\vgadonut.donut.donuthit.rx[7] ));
 sg13g2_o21ai_1 _16124_ (.B1(_06931_),
    .Y(_00306_),
    .A1(_04321_),
    .A2(_06930_));
 sg13g2_nand2_1 _16125_ (.Y(_06932_),
    .A(_06927_),
    .B(\vgadonut.donut.donuthit.rx[8] ));
 sg13g2_o21ai_1 _16126_ (.B1(_06932_),
    .Y(_00307_),
    .A1(_04371_),
    .A2(net108));
 sg13g2_nand2_1 _16127_ (.Y(_06933_),
    .A(_06927_),
    .B(\vgadonut.donut.donuthit.rx[9] ));
 sg13g2_o21ai_1 _16128_ (.B1(_06933_),
    .Y(_00308_),
    .A1(_04422_),
    .A2(_06930_));
 sg13g2_inv_1 _16129_ (.Y(_06934_),
    .A(\vgadonut.donut.donuthit.ryin[10] ));
 sg13g2_nand2_1 _16130_ (.Y(_06935_),
    .A(net119),
    .B(\vgadonut.donut.donuthit.ry[10] ));
 sg13g2_o21ai_1 _16131_ (.B1(_06935_),
    .Y(_00309_),
    .A1(_06934_),
    .A2(net108));
 sg13g2_inv_1 _16132_ (.Y(_06936_),
    .A(\vgadonut.donut.donuthit.ryin[11] ));
 sg13g2_nand2_1 _16133_ (.Y(_06937_),
    .A(net119),
    .B(\vgadonut.donut.donuthit.ry[11] ));
 sg13g2_o21ai_1 _16134_ (.B1(_06937_),
    .Y(_00310_),
    .A1(_06936_),
    .A2(net108));
 sg13g2_nand2_1 _16135_ (.Y(_06938_),
    .A(net119),
    .B(\vgadonut.donut.donuthit.ry[12] ));
 sg13g2_o21ai_1 _16136_ (.B1(_06938_),
    .Y(_00311_),
    .A1(_05093_),
    .A2(net108));
 sg13g2_nand2_1 _16137_ (.Y(_06939_),
    .A(net119),
    .B(\vgadonut.donut.donuthit.ry[13] ));
 sg13g2_o21ai_1 _16138_ (.B1(_06939_),
    .Y(_00312_),
    .A1(_05133_),
    .A2(net108));
 sg13g2_nand2_1 _16139_ (.Y(_06940_),
    .A(net119),
    .B(\vgadonut.donut.donuthit.ry[14] ));
 sg13g2_o21ai_1 _16140_ (.B1(_06940_),
    .Y(_00313_),
    .A1(_05167_),
    .A2(net108));
 sg13g2_buf_1 _16141_ (.A(net138),
    .X(_06941_));
 sg13g2_nand2_1 _16142_ (.Y(_06942_),
    .A(_06941_),
    .B(\vgadonut.donut.donuthit.ry[15] ));
 sg13g2_o21ai_1 _16143_ (.B1(_06942_),
    .Y(_00314_),
    .A1(_05222_),
    .A2(net108));
 sg13g2_nand2_1 _16144_ (.Y(_06943_),
    .A(net118),
    .B(\vgadonut.donut.donuthit.ry[5] ));
 sg13g2_o21ai_1 _16145_ (.B1(_06943_),
    .Y(_00315_),
    .A1(_04839_),
    .A2(net108));
 sg13g2_inv_1 _16146_ (.Y(_06944_),
    .A(\vgadonut.donut.donuthit.ryin[6] ));
 sg13g2_buf_1 _16147_ (.A(net137),
    .X(_06945_));
 sg13g2_nand2_1 _16148_ (.Y(_06946_),
    .A(net118),
    .B(\vgadonut.donut.donuthit.ry[6] ));
 sg13g2_o21ai_1 _16149_ (.B1(_06946_),
    .Y(_00316_),
    .A1(_06944_),
    .A2(net117));
 sg13g2_inv_1 _16150_ (.Y(_06947_),
    .A(\vgadonut.donut.donuthit.ryin[7] ));
 sg13g2_nand2_1 _16151_ (.Y(_06948_),
    .A(net118),
    .B(\vgadonut.donut.donuthit.ry[7] ));
 sg13g2_o21ai_1 _16152_ (.B1(_06948_),
    .Y(_00317_),
    .A1(_06947_),
    .A2(net117));
 sg13g2_nand2_1 _16153_ (.Y(_06949_),
    .A(net118),
    .B(\vgadonut.donut.donuthit.ry[8] ));
 sg13g2_o21ai_1 _16154_ (.B1(_06949_),
    .Y(_00318_),
    .A1(_04957_),
    .A2(net117));
 sg13g2_inv_1 _16155_ (.Y(_06950_),
    .A(\vgadonut.donut.donuthit.ryin[9] ));
 sg13g2_nand2_1 _16156_ (.Y(_06951_),
    .A(net118),
    .B(\vgadonut.donut.donuthit.ry[9] ));
 sg13g2_o21ai_1 _16157_ (.B1(_06951_),
    .Y(_00319_),
    .A1(_06950_),
    .A2(net117));
 sg13g2_nand2_1 _16158_ (.Y(_06952_),
    .A(net118),
    .B(\vgadonut.donut.donuthit.rz[10] ));
 sg13g2_o21ai_1 _16159_ (.B1(_06952_),
    .Y(_00320_),
    .A1(_05640_),
    .A2(net117));
 sg13g2_inv_1 _16160_ (.Y(_06953_),
    .A(_05691_));
 sg13g2_nand2_1 _16161_ (.Y(_06954_),
    .A(net118),
    .B(\vgadonut.donut.donuthit.rz[11] ));
 sg13g2_o21ai_1 _16162_ (.B1(_06954_),
    .Y(_00321_),
    .A1(_06953_),
    .A2(_06945_));
 sg13g2_inv_1 _16163_ (.Y(_06955_),
    .A(_05727_));
 sg13g2_nand2_1 _16164_ (.Y(_06956_),
    .A(net118),
    .B(\vgadonut.donut.donuthit.rz[12] ));
 sg13g2_o21ai_1 _16165_ (.B1(_06956_),
    .Y(_00322_),
    .A1(_06955_),
    .A2(net117));
 sg13g2_inv_1 _16166_ (.Y(_06957_),
    .A(_05770_));
 sg13g2_nand2_1 _16167_ (.Y(_06958_),
    .A(_06941_),
    .B(\vgadonut.donut.donuthit.rz[13] ));
 sg13g2_o21ai_1 _16168_ (.B1(_06958_),
    .Y(_00323_),
    .A1(_06957_),
    .A2(net117));
 sg13g2_buf_1 _16169_ (.A(_04190_),
    .X(_06959_));
 sg13g2_nand2_1 _16170_ (.Y(_06960_),
    .A(net116),
    .B(\vgadonut.donut.donuthit.rz[14] ));
 sg13g2_o21ai_1 _16171_ (.B1(_06960_),
    .Y(_00324_),
    .A1(_05805_),
    .A2(net117));
 sg13g2_nand2_1 _16172_ (.Y(_06961_),
    .A(net116),
    .B(\vgadonut.donut.donuthit.rz[15] ));
 sg13g2_o21ai_1 _16173_ (.B1(_06961_),
    .Y(_00325_),
    .A1(_05889_),
    .A2(_06945_));
 sg13g2_nand2_1 _16174_ (.Y(_06962_),
    .A(net116),
    .B(\vgadonut.donut.donuthit.rz[5] ));
 sg13g2_o21ai_1 _16175_ (.B1(_06962_),
    .Y(_00326_),
    .A1(_05415_),
    .A2(net124));
 sg13g2_nand2_1 _16176_ (.Y(_06963_),
    .A(net116),
    .B(\vgadonut.donut.donuthit.rz[6] ));
 sg13g2_o21ai_1 _16177_ (.B1(_06963_),
    .Y(_00327_),
    .A1(_05420_),
    .A2(net124));
 sg13g2_nand2_1 _16178_ (.Y(_06964_),
    .A(net116),
    .B(\vgadonut.donut.donuthit.rz[7] ));
 sg13g2_o21ai_1 _16179_ (.B1(_06964_),
    .Y(_00328_),
    .A1(_05503_),
    .A2(net124));
 sg13g2_inv_1 _16180_ (.Y(_06965_),
    .A(_05551_));
 sg13g2_nand2_1 _16181_ (.Y(_06966_),
    .A(net116),
    .B(\vgadonut.donut.donuthit.rz[8] ));
 sg13g2_o21ai_1 _16182_ (.B1(_06966_),
    .Y(_00329_),
    .A1(_06965_),
    .A2(net124));
 sg13g2_inv_1 _16183_ (.Y(_06967_),
    .A(_05595_));
 sg13g2_nand2_1 _16184_ (.Y(_06968_),
    .A(net116),
    .B(\vgadonut.donut.donuthit.rz[9] ));
 sg13g2_o21ai_1 _16185_ (.B1(_06968_),
    .Y(_00330_),
    .A1(_06967_),
    .A2(net124));
 sg13g2_inv_1 _16186_ (.Y(_06969_),
    .A(\vgadonut.donut.rx6[0] ));
 sg13g2_nand3_1 _16187_ (.B(_10128_),
    .C(_05973_),
    .A(_09800_),
    .Y(_06970_));
 sg13g2_nand3_1 _16188_ (.B(_06217_),
    .C(_06335_),
    .A(_06216_),
    .Y(_06971_));
 sg13g2_inv_1 _16189_ (.Y(_06972_),
    .A(_06213_));
 sg13g2_nor2_1 _16190_ (.A(_06971_),
    .B(_06972_),
    .Y(_06973_));
 sg13g2_nor2_1 _16191_ (.A(_10004_),
    .B(_10106_),
    .Y(_06974_));
 sg13g2_buf_2 _16192_ (.A(_06974_),
    .X(_06975_));
 sg13g2_inv_1 _16193_ (.Y(_06976_),
    .A(_06975_));
 sg13g2_nor2_1 _16194_ (.A(_06973_),
    .B(_06976_),
    .Y(_06977_));
 sg13g2_inv_1 _16195_ (.Y(_06978_),
    .A(_06977_));
 sg13g2_nand2_1 _16196_ (.Y(_06979_),
    .A(_06970_),
    .B(_06978_));
 sg13g2_buf_1 _16197_ (.A(_06979_),
    .X(_06980_));
 sg13g2_buf_1 _16198_ (.A(_06980_),
    .X(_06981_));
 sg13g2_buf_1 _16199_ (.A(_06334_),
    .X(_06982_));
 sg13g2_buf_1 _16200_ (.A(net170),
    .X(_06983_));
 sg13g2_nand2_1 _16201_ (.Y(_06984_),
    .A(\vgadonut.donut.rx6[0] ),
    .B(net230));
 sg13g2_nand2_1 _16202_ (.Y(_06985_),
    .A(_06969_),
    .B(_06883_));
 sg13g2_nand4_1 _16203_ (.B(net165),
    .C(_06984_),
    .A(net107),
    .Y(_06986_),
    .D(_06985_));
 sg13g2_o21ai_1 _16204_ (.B1(_06986_),
    .Y(_00347_),
    .A1(_06969_),
    .A2(net105));
 sg13g2_inv_1 _16205_ (.Y(_06987_),
    .A(\vgadonut.donut.donuthit.rxin[4] ));
 sg13g2_inv_1 _16206_ (.Y(_06988_),
    .A(net107));
 sg13g2_buf_1 _16207_ (.A(_06988_),
    .X(_06989_));
 sg13g2_buf_1 _16208_ (.A(_06989_),
    .X(_06990_));
 sg13g2_buf_1 _16209_ (.A(net100),
    .X(_06991_));
 sg13g2_nor2_1 _16210_ (.A(\vgadonut.donut.donuthit.rxin[4] ),
    .B(_06035_),
    .Y(_06992_));
 sg13g2_nand2_1 _16211_ (.Y(_06993_),
    .A(\vgadonut.donut.donuthit.rxin[4] ),
    .B(_06035_));
 sg13g2_nor2b_1 _16212_ (.A(_06992_),
    .B_N(_06993_),
    .Y(_06994_));
 sg13g2_nor2_1 _16213_ (.A(\vgadonut.donut.rx6[5] ),
    .B(_06066_),
    .Y(_06995_));
 sg13g2_inv_1 _16214_ (.Y(_06996_),
    .A(\vgadonut.donut.rx6[1] ));
 sg13g2_xor2_1 _16215_ (.B(net231),
    .A(\vgadonut.donut.rx6[1] ),
    .X(_06997_));
 sg13g2_nand2b_1 _16216_ (.Y(_06998_),
    .B(_06997_),
    .A_N(_06984_));
 sg13g2_o21ai_1 _16217_ (.B1(_06998_),
    .Y(_06999_),
    .A1(_06996_),
    .A2(_06894_));
 sg13g2_nor2_1 _16218_ (.A(\vgadonut.donut.rx6[2] ),
    .B(net190),
    .Y(_07000_));
 sg13g2_inv_1 _16219_ (.Y(_07001_),
    .A(_07000_));
 sg13g2_nand2_1 _16220_ (.Y(_07002_),
    .A(\vgadonut.donut.rx6[2] ),
    .B(net190));
 sg13g2_inv_1 _16221_ (.Y(_07003_),
    .A(_07002_));
 sg13g2_a21oi_1 _16222_ (.A1(_06999_),
    .A2(_07001_),
    .Y(_07004_),
    .B1(_07003_));
 sg13g2_nand2_1 _16223_ (.Y(_07005_),
    .A(\vgadonut.donut.rx6[3] ),
    .B(net229));
 sg13g2_nor2_1 _16224_ (.A(\vgadonut.donut.rx6[3] ),
    .B(net229),
    .Y(_07006_));
 sg13g2_a21oi_1 _16225_ (.A1(_07004_),
    .A2(_07005_),
    .Y(_07007_),
    .B1(_07006_));
 sg13g2_nor2_1 _16226_ (.A(\vgadonut.donut.rx6[4] ),
    .B(_06060_),
    .Y(_07008_));
 sg13g2_inv_1 _16227_ (.Y(_07009_),
    .A(_07008_));
 sg13g2_nand2_1 _16228_ (.Y(_07010_),
    .A(\vgadonut.donut.rx6[4] ),
    .B(_06060_));
 sg13g2_inv_1 _16229_ (.Y(_07011_),
    .A(_07010_));
 sg13g2_a21oi_1 _16230_ (.A1(_07007_),
    .A2(_07009_),
    .Y(_07012_),
    .B1(_07011_));
 sg13g2_nand2_1 _16231_ (.Y(_07013_),
    .A(\vgadonut.donut.rx6[5] ),
    .B(_06066_));
 sg13g2_o21ai_1 _16232_ (.B1(_07013_),
    .Y(_07014_),
    .A1(_06995_),
    .A2(_07012_));
 sg13g2_nor2_1 _16233_ (.A(\vgadonut.donut.donuthit.rxin[1] ),
    .B(_06078_),
    .Y(_07015_));
 sg13g2_nand2_1 _16234_ (.Y(_07016_),
    .A(\vgadonut.donut.donuthit.rxin[1] ),
    .B(_06078_));
 sg13g2_inv_1 _16235_ (.Y(_07017_),
    .A(_07016_));
 sg13g2_nor2_1 _16236_ (.A(_07015_),
    .B(_07017_),
    .Y(_07018_));
 sg13g2_inv_1 _16237_ (.Y(_07019_),
    .A(_07018_));
 sg13g2_nor2_1 _16238_ (.A(\vgadonut.donut.donuthit.rxin[0] ),
    .B(_06072_),
    .Y(_07020_));
 sg13g2_nand2_1 _16239_ (.Y(_07021_),
    .A(\vgadonut.donut.donuthit.rxin[0] ),
    .B(_06072_));
 sg13g2_nor2b_1 _16240_ (.A(_07020_),
    .B_N(_07021_),
    .Y(_07022_));
 sg13g2_inv_1 _16241_ (.Y(_07023_),
    .A(_07022_));
 sg13g2_nor2_1 _16242_ (.A(_07019_),
    .B(_07023_),
    .Y(_07024_));
 sg13g2_a21oi_1 _16243_ (.A1(_07021_),
    .A2(_07016_),
    .Y(_07025_),
    .B1(_07015_));
 sg13g2_a21oi_1 _16244_ (.A1(_07014_),
    .A2(_07024_),
    .Y(_07026_),
    .B1(_07025_));
 sg13g2_inv_1 _16245_ (.Y(_07027_),
    .A(_07026_));
 sg13g2_nor2_1 _16246_ (.A(\vgadonut.donut.donuthit.rxin[3] ),
    .B(_06091_),
    .Y(_07028_));
 sg13g2_nand2_1 _16247_ (.Y(_07029_),
    .A(\vgadonut.donut.donuthit.rxin[3] ),
    .B(_06091_));
 sg13g2_inv_1 _16248_ (.Y(_07030_),
    .A(_07029_));
 sg13g2_nor2_1 _16249_ (.A(_07028_),
    .B(_07030_),
    .Y(_07031_));
 sg13g2_inv_1 _16250_ (.Y(_07032_),
    .A(_07031_));
 sg13g2_buf_1 _16251_ (.A(\vgadonut.donut.donuthit.rxin[2] ),
    .X(_07033_));
 sg13g2_nor2_1 _16252_ (.A(_07033_),
    .B(_06085_),
    .Y(_07034_));
 sg13g2_nand2_1 _16253_ (.Y(_07035_),
    .A(_07033_),
    .B(_06085_));
 sg13g2_inv_1 _16254_ (.Y(_07036_),
    .A(_07035_));
 sg13g2_nor2_1 _16255_ (.A(_07034_),
    .B(_07036_),
    .Y(_07037_));
 sg13g2_nor2b_1 _16256_ (.A(_07032_),
    .B_N(_07037_),
    .Y(_07038_));
 sg13g2_a21oi_1 _16257_ (.A1(_07035_),
    .A2(_07029_),
    .Y(_07039_),
    .B1(_07028_));
 sg13g2_a21oi_1 _16258_ (.A1(_07027_),
    .A2(_07038_),
    .Y(_07040_),
    .B1(_07039_));
 sg13g2_xnor2_1 _16259_ (.Y(_07041_),
    .A(_06994_),
    .B(_07040_));
 sg13g2_buf_1 _16260_ (.A(net170),
    .X(_07042_));
 sg13g2_buf_1 _16261_ (.A(_06989_),
    .X(_07043_));
 sg13g2_a21oi_1 _16262_ (.A1(_07041_),
    .A2(net164),
    .Y(_07044_),
    .B1(net99));
 sg13g2_nand2_1 _16263_ (.Y(_07045_),
    .A(_06038_),
    .B(_04206_));
 sg13g2_buf_1 _16264_ (.A(_00135_),
    .X(_07046_));
 sg13g2_nor2_1 _16265_ (.A(_06038_),
    .B(_04206_),
    .Y(_07047_));
 sg13g2_a21oi_1 _16266_ (.A1(_07045_),
    .A2(_07046_),
    .Y(_07048_),
    .B1(_07047_));
 sg13g2_buf_1 _16267_ (.A(_00136_),
    .X(_07049_));
 sg13g2_nor2_1 _16268_ (.A(_06047_),
    .B(_04205_),
    .Y(_07050_));
 sg13g2_nand2_1 _16269_ (.Y(_07051_),
    .A(_06047_),
    .B(_04205_));
 sg13g2_nor2b_1 _16270_ (.A(_07050_),
    .B_N(_07051_),
    .Y(_07052_));
 sg13g2_xnor2_1 _16271_ (.Y(_07053_),
    .A(_07049_),
    .B(_07052_));
 sg13g2_xor2_1 _16272_ (.B(_07053_),
    .A(_07048_),
    .X(_07054_));
 sg13g2_nor2_1 _16273_ (.A(_07048_),
    .B(_07053_),
    .Y(_07055_));
 sg13g2_a21oi_1 _16274_ (.A1(_07054_),
    .A2(_07046_),
    .Y(_07056_),
    .B1(_07055_));
 sg13g2_a21oi_1 _16275_ (.A1(_07051_),
    .A2(_07049_),
    .Y(_07057_),
    .B1(_07050_));
 sg13g2_buf_1 _16276_ (.A(_00137_),
    .X(_07058_));
 sg13g2_nor2_1 _16277_ (.A(net229),
    .B(net250),
    .Y(_07059_));
 sg13g2_nand2_1 _16278_ (.Y(_07060_),
    .A(_06054_),
    .B(net250));
 sg13g2_nor2b_1 _16279_ (.A(_07059_),
    .B_N(_07060_),
    .Y(_07061_));
 sg13g2_xnor2_1 _16280_ (.Y(_07062_),
    .A(_07058_),
    .B(_07061_));
 sg13g2_xor2_1 _16281_ (.B(_07062_),
    .A(_07057_),
    .X(_07063_));
 sg13g2_xnor2_1 _16282_ (.Y(_07064_),
    .A(_07049_),
    .B(_07063_));
 sg13g2_nor2_1 _16283_ (.A(_07056_),
    .B(_07064_),
    .Y(_07065_));
 sg13g2_nor2_1 _16284_ (.A(_07057_),
    .B(_07062_),
    .Y(_07066_));
 sg13g2_a21oi_1 _16285_ (.A1(_07063_),
    .A2(_07049_),
    .Y(_07067_),
    .B1(_07066_));
 sg13g2_a21oi_1 _16286_ (.A1(_07060_),
    .A2(_07058_),
    .Y(_07068_),
    .B1(_07059_));
 sg13g2_buf_1 _16287_ (.A(_00138_),
    .X(_07069_));
 sg13g2_nor2_1 _16288_ (.A(_06060_),
    .B(net252),
    .Y(_07070_));
 sg13g2_nand2_1 _16289_ (.Y(_07071_),
    .A(_06060_),
    .B(net252));
 sg13g2_nor2b_1 _16290_ (.A(_07070_),
    .B_N(_07071_),
    .Y(_07072_));
 sg13g2_xnor2_1 _16291_ (.Y(_07073_),
    .A(_07069_),
    .B(_07072_));
 sg13g2_xor2_1 _16292_ (.B(_07073_),
    .A(_07068_),
    .X(_07074_));
 sg13g2_xnor2_1 _16293_ (.Y(_07075_),
    .A(_07058_),
    .B(_07074_));
 sg13g2_xor2_1 _16294_ (.B(_07075_),
    .A(_07067_),
    .X(_07076_));
 sg13g2_xnor2_1 _16295_ (.Y(_07077_),
    .A(_07065_),
    .B(_07076_));
 sg13g2_buf_1 _16296_ (.A(_00134_),
    .X(_07078_));
 sg13g2_inv_1 _16297_ (.Y(_07079_),
    .A(_07078_));
 sg13g2_nor2_1 _16298_ (.A(net230),
    .B(_04208_),
    .Y(_07080_));
 sg13g2_nand2_1 _16299_ (.Y(_07081_),
    .A(net230),
    .B(_04208_));
 sg13g2_nor2b_1 _16300_ (.A(_07080_),
    .B_N(_07081_),
    .Y(_07082_));
 sg13g2_xnor2_1 _16301_ (.Y(_07083_),
    .A(_07079_),
    .B(_07082_));
 sg13g2_nor2_1 _16302_ (.A(_06055_),
    .B(_07083_),
    .Y(_07084_));
 sg13g2_a21oi_1 _16303_ (.A1(_07081_),
    .A2(_07078_),
    .Y(_07085_),
    .B1(_07080_));
 sg13g2_nor2b_1 _16304_ (.A(_07047_),
    .B_N(_07045_),
    .Y(_07086_));
 sg13g2_xnor2_1 _16305_ (.Y(_07087_),
    .A(_07046_),
    .B(_07086_));
 sg13g2_xor2_1 _16306_ (.B(_07087_),
    .A(_07085_),
    .X(_07088_));
 sg13g2_xnor2_1 _16307_ (.Y(_07089_),
    .A(_07078_),
    .B(_07088_));
 sg13g2_nor2_1 _16308_ (.A(_07084_),
    .B(_07089_),
    .Y(_07090_));
 sg13g2_inv_1 _16309_ (.Y(_07091_),
    .A(_07090_));
 sg13g2_nor2_1 _16310_ (.A(_07085_),
    .B(_07087_),
    .Y(_07092_));
 sg13g2_a21oi_1 _16311_ (.A1(_07088_),
    .A2(_07078_),
    .Y(_07093_),
    .B1(_07092_));
 sg13g2_xnor2_1 _16312_ (.Y(_07094_),
    .A(_07046_),
    .B(_07054_));
 sg13g2_xnor2_1 _16313_ (.Y(_07095_),
    .A(_07093_),
    .B(_07094_));
 sg13g2_xnor2_1 _16314_ (.Y(_07096_),
    .A(_07091_),
    .B(_07095_));
 sg13g2_nor2_1 _16315_ (.A(net190),
    .B(net231),
    .Y(_07097_));
 sg13g2_nand2_1 _16316_ (.Y(_07098_),
    .A(net231),
    .B(net230));
 sg13g2_nor2_1 _16317_ (.A(net190),
    .B(_07098_),
    .Y(_07099_));
 sg13g2_inv_1 _16318_ (.Y(_07100_),
    .A(_07099_));
 sg13g2_nand2_1 _16319_ (.Y(_07101_),
    .A(net190),
    .B(net231));
 sg13g2_inv_1 _16320_ (.Y(_07102_),
    .A(_07101_));
 sg13g2_xor2_1 _16321_ (.B(net229),
    .A(net190),
    .X(_07103_));
 sg13g2_nor2_1 _16322_ (.A(_07102_),
    .B(_07103_),
    .Y(_07104_));
 sg13g2_a21oi_1 _16323_ (.A1(_06055_),
    .A2(_07102_),
    .Y(_07105_),
    .B1(_07104_));
 sg13g2_a22oi_1 _16324_ (.Y(_07106_),
    .B1(_07100_),
    .B2(_07105_),
    .A2(_07097_),
    .A1(_06883_));
 sg13g2_inv_1 _16325_ (.Y(_07107_),
    .A(_07104_));
 sg13g2_inv_1 _16326_ (.Y(_07108_),
    .A(_07083_));
 sg13g2_nand2_1 _16327_ (.Y(_07109_),
    .A(_06901_),
    .B(net229));
 sg13g2_nand2_1 _16328_ (.Y(_07110_),
    .A(_07083_),
    .B(_06055_));
 sg13g2_inv_1 _16329_ (.Y(_07111_),
    .A(_07084_));
 sg13g2_a22oi_1 _16330_ (.Y(_07112_),
    .B1(_07110_),
    .B2(_07111_),
    .A2(_06054_),
    .A1(_06901_));
 sg13g2_inv_1 _16331_ (.Y(_07113_),
    .A(_07112_));
 sg13g2_o21ai_1 _16332_ (.B1(_07113_),
    .Y(_07114_),
    .A1(_07108_),
    .A2(_07109_));
 sg13g2_xnor2_1 _16333_ (.Y(_07115_),
    .A(_07107_),
    .B(_07114_));
 sg13g2_nor2_1 _16334_ (.A(_07106_),
    .B(_07115_),
    .Y(_07116_));
 sg13g2_xnor2_1 _16335_ (.Y(_07117_),
    .A(_07084_),
    .B(_07089_));
 sg13g2_nor2_1 _16336_ (.A(_07113_),
    .B(_07117_),
    .Y(_07118_));
 sg13g2_inv_1 _16337_ (.Y(_07119_),
    .A(_07118_));
 sg13g2_nand2_1 _16338_ (.Y(_07120_),
    .A(_07117_),
    .B(_07113_));
 sg13g2_nand2_2 _16339_ (.Y(_07121_),
    .A(_07119_),
    .B(_07120_));
 sg13g2_inv_1 _16340_ (.Y(_07122_),
    .A(_07121_));
 sg13g2_nor2_1 _16341_ (.A(_07107_),
    .B(_07114_),
    .Y(_07123_));
 sg13g2_inv_1 _16342_ (.Y(_07124_),
    .A(_07123_));
 sg13g2_o21ai_1 _16343_ (.B1(_07119_),
    .Y(_07125_),
    .A1(_07124_),
    .A2(_07121_));
 sg13g2_a21oi_1 _16344_ (.A1(_07116_),
    .A2(_07122_),
    .Y(_07126_),
    .B1(_07125_));
 sg13g2_nor2_1 _16345_ (.A(_07096_),
    .B(_07126_),
    .Y(_07127_));
 sg13g2_nor2_1 _16346_ (.A(_07093_),
    .B(_07094_),
    .Y(_07128_));
 sg13g2_xnor2_1 _16347_ (.Y(_07129_),
    .A(_07056_),
    .B(_07064_));
 sg13g2_xnor2_1 _16348_ (.Y(_07130_),
    .A(_07128_),
    .B(_07129_));
 sg13g2_nor2_1 _16349_ (.A(_07091_),
    .B(_07095_),
    .Y(_07131_));
 sg13g2_inv_1 _16350_ (.Y(_07132_),
    .A(_07131_));
 sg13g2_inv_1 _16351_ (.Y(_07133_),
    .A(_07130_));
 sg13g2_nor2b_1 _16352_ (.A(_07129_),
    .B_N(_07128_),
    .Y(_07134_));
 sg13g2_inv_1 _16353_ (.Y(_07135_),
    .A(_07134_));
 sg13g2_o21ai_1 _16354_ (.B1(_07135_),
    .Y(_07136_),
    .A1(_07132_),
    .A2(_07133_));
 sg13g2_a21oi_1 _16355_ (.A1(_07127_),
    .A2(_07130_),
    .Y(_07137_),
    .B1(_07136_));
 sg13g2_nor2_1 _16356_ (.A(_07077_),
    .B(_07137_),
    .Y(_07138_));
 sg13g2_inv_1 _16357_ (.Y(_07139_),
    .A(_07138_));
 sg13g2_buf_1 _16358_ (.A(_10117_),
    .X(_07140_));
 sg13g2_nand2_1 _16359_ (.Y(_07141_),
    .A(_07137_),
    .B(_07077_));
 sg13g2_nand3_1 _16360_ (.B(net151),
    .C(_07141_),
    .A(_07139_),
    .Y(_07142_));
 sg13g2_a22oi_1 _16361_ (.Y(_00348_),
    .B1(_07044_),
    .B2(_07142_),
    .A2(net93),
    .A1(_06987_));
 sg13g2_xnor2_1 _16362_ (.Y(_07143_),
    .A(net231),
    .B(net230));
 sg13g2_a21oi_1 _16363_ (.A1(_07102_),
    .A2(_06883_),
    .Y(_07144_),
    .B1(_07097_));
 sg13g2_nand2_1 _16364_ (.Y(_07145_),
    .A(_07144_),
    .B(_07100_));
 sg13g2_inv_1 _16365_ (.Y(_07146_),
    .A(_07145_));
 sg13g2_a21oi_1 _16366_ (.A1(_00133_),
    .A2(_07143_),
    .Y(_07147_),
    .B1(_07146_));
 sg13g2_inv_1 _16367_ (.Y(_07148_),
    .A(_07147_));
 sg13g2_nand2b_1 _16368_ (.Y(_07149_),
    .B(_07144_),
    .A_N(_07105_));
 sg13g2_nor2_1 _16369_ (.A(_06055_),
    .B(_07144_),
    .Y(_07150_));
 sg13g2_inv_1 _16370_ (.Y(_07151_),
    .A(_07150_));
 sg13g2_nand2_1 _16371_ (.Y(_07152_),
    .A(_07149_),
    .B(_07151_));
 sg13g2_nor2_1 _16372_ (.A(_07152_),
    .B(_07115_),
    .Y(_07153_));
 sg13g2_o21ai_1 _16373_ (.B1(_07124_),
    .Y(_07154_),
    .A1(_07151_),
    .A2(_07115_));
 sg13g2_a21oi_1 _16374_ (.A1(_07148_),
    .A2(_07153_),
    .Y(_07155_),
    .B1(_07154_));
 sg13g2_inv_1 _16375_ (.Y(_07156_),
    .A(_07155_));
 sg13g2_nor2_1 _16376_ (.A(_07096_),
    .B(_07121_),
    .Y(_07157_));
 sg13g2_o21ai_1 _16377_ (.B1(_07132_),
    .Y(_07158_),
    .A1(_07119_),
    .A2(_07096_));
 sg13g2_a21oi_1 _16378_ (.A1(_07156_),
    .A2(_07157_),
    .Y(_07159_),
    .B1(_07158_));
 sg13g2_inv_1 _16379_ (.Y(_07160_),
    .A(_07159_));
 sg13g2_nor2_1 _16380_ (.A(_07077_),
    .B(_07133_),
    .Y(_07161_));
 sg13g2_inv_1 _16381_ (.Y(_07162_),
    .A(_07065_));
 sg13g2_inv_1 _16382_ (.Y(_07163_),
    .A(_07076_));
 sg13g2_a21oi_1 _16383_ (.A1(_07135_),
    .A2(_07162_),
    .Y(_07164_),
    .B1(_07163_));
 sg13g2_a21oi_1 _16384_ (.A1(_07160_),
    .A2(_07161_),
    .Y(_07165_),
    .B1(_07164_));
 sg13g2_inv_1 _16385_ (.Y(_07166_),
    .A(_07165_));
 sg13g2_nor2_1 _16386_ (.A(_07067_),
    .B(_07075_),
    .Y(_07167_));
 sg13g2_inv_1 _16387_ (.Y(_07168_),
    .A(_07167_));
 sg13g2_nor2_1 _16388_ (.A(_07068_),
    .B(_07073_),
    .Y(_07169_));
 sg13g2_a21oi_1 _16389_ (.A1(_07074_),
    .A2(_07058_),
    .Y(_07170_),
    .B1(_07169_));
 sg13g2_a21oi_1 _16390_ (.A1(_07071_),
    .A2(_07069_),
    .Y(_07171_),
    .B1(_07070_));
 sg13g2_buf_1 _16391_ (.A(_00139_),
    .X(_07172_));
 sg13g2_nor2_1 _16392_ (.A(_06066_),
    .B(net249),
    .Y(_07173_));
 sg13g2_nand2_1 _16393_ (.Y(_07174_),
    .A(_06066_),
    .B(net249));
 sg13g2_nor2b_1 _16394_ (.A(_07173_),
    .B_N(_07174_),
    .Y(_07175_));
 sg13g2_xnor2_1 _16395_ (.Y(_07176_),
    .A(_07172_),
    .B(_07175_));
 sg13g2_xor2_1 _16396_ (.B(_07176_),
    .A(_07171_),
    .X(_07177_));
 sg13g2_xnor2_1 _16397_ (.Y(_07178_),
    .A(_07069_),
    .B(_07177_));
 sg13g2_xnor2_1 _16398_ (.Y(_07179_),
    .A(_07170_),
    .B(_07178_));
 sg13g2_nor2_1 _16399_ (.A(_07168_),
    .B(_07179_),
    .Y(_07180_));
 sg13g2_inv_1 _16400_ (.Y(_07181_),
    .A(_07180_));
 sg13g2_nand2_1 _16401_ (.Y(_07182_),
    .A(_07179_),
    .B(_07168_));
 sg13g2_nand2_1 _16402_ (.Y(_07183_),
    .A(_07181_),
    .B(_07182_));
 sg13g2_inv_1 _16403_ (.Y(_07184_),
    .A(_07183_));
 sg13g2_buf_1 _16404_ (.A(_10106_),
    .X(_07185_));
 sg13g2_a21oi_1 _16405_ (.A1(_07166_),
    .A2(_07184_),
    .Y(_07186_),
    .B1(net163));
 sg13g2_nand2_1 _16406_ (.Y(_07187_),
    .A(_07165_),
    .B(_07183_));
 sg13g2_a21oi_1 _16407_ (.A1(_07186_),
    .A2(_07187_),
    .Y(_07188_),
    .B1(net99));
 sg13g2_nor2_1 _16408_ (.A(\vgadonut.donut.donuthit.rxin[5] ),
    .B(_06033_),
    .Y(_07189_));
 sg13g2_nand2_1 _16409_ (.Y(_07190_),
    .A(\vgadonut.donut.donuthit.rxin[5] ),
    .B(_06033_));
 sg13g2_nor2b_1 _16410_ (.A(_07189_),
    .B_N(_07190_),
    .Y(_07191_));
 sg13g2_inv_1 _16411_ (.Y(_07192_),
    .A(_07014_));
 sg13g2_o21ai_1 _16412_ (.B1(_07021_),
    .Y(_07193_),
    .A1(_07020_),
    .A2(_07192_));
 sg13g2_a221oi_1 _16413_ (.B2(_07018_),
    .C1(_07017_),
    .B1(_07193_),
    .A1(_07033_),
    .Y(_07194_),
    .A2(_06085_));
 sg13g2_nor2_1 _16414_ (.A(_07034_),
    .B(_07194_),
    .Y(_07195_));
 sg13g2_nand2_1 _16415_ (.Y(_07196_),
    .A(_07195_),
    .B(_07031_));
 sg13g2_nand2_1 _16416_ (.Y(_07197_),
    .A(_06993_),
    .B(_07029_));
 sg13g2_inv_1 _16417_ (.Y(_07198_),
    .A(_07197_));
 sg13g2_a21oi_1 _16418_ (.A1(_07196_),
    .A2(_07198_),
    .Y(_07199_),
    .B1(_06992_));
 sg13g2_buf_1 _16419_ (.A(_10117_),
    .X(_07200_));
 sg13g2_a21oi_1 _16420_ (.A1(_07199_),
    .A2(_07191_),
    .Y(_07201_),
    .B1(_07200_));
 sg13g2_o21ai_1 _16421_ (.B1(_07201_),
    .Y(_07202_),
    .A1(_07191_),
    .A2(_07199_));
 sg13g2_a22oi_1 _16422_ (.Y(_00349_),
    .B1(_07188_),
    .B2(_07202_),
    .A2(net93),
    .A1(_04196_));
 sg13g2_nor2_1 _16423_ (.A(_04222_),
    .B(_06031_),
    .Y(_07203_));
 sg13g2_nand2_1 _16424_ (.Y(_07204_),
    .A(_04222_),
    .B(_06031_));
 sg13g2_inv_1 _16425_ (.Y(_07205_),
    .A(_07204_));
 sg13g2_nor2_1 _16426_ (.A(_07203_),
    .B(_07205_),
    .Y(_07206_));
 sg13g2_inv_1 _16427_ (.Y(_07207_),
    .A(_07206_));
 sg13g2_nand2b_1 _16428_ (.Y(_07208_),
    .B(_06994_),
    .A_N(_07040_));
 sg13g2_nand2_1 _16429_ (.Y(_07209_),
    .A(_06993_),
    .B(_07190_));
 sg13g2_inv_1 _16430_ (.Y(_07210_),
    .A(_07209_));
 sg13g2_a21oi_1 _16431_ (.A1(_07208_),
    .A2(_07210_),
    .Y(_07211_),
    .B1(_07189_));
 sg13g2_xnor2_1 _16432_ (.Y(_07212_),
    .A(_07207_),
    .B(_07211_));
 sg13g2_a21oi_1 _16433_ (.A1(_07212_),
    .A2(net164),
    .Y(_07213_),
    .B1(net99));
 sg13g2_nor2_1 _16434_ (.A(_07170_),
    .B(_07178_),
    .Y(_07214_));
 sg13g2_inv_1 _16435_ (.Y(_07215_),
    .A(_07214_));
 sg13g2_nor2_1 _16436_ (.A(_07171_),
    .B(_07176_),
    .Y(_07216_));
 sg13g2_a21oi_1 _16437_ (.A1(_07177_),
    .A2(_07069_),
    .Y(_07217_),
    .B1(_07216_));
 sg13g2_a21oi_1 _16438_ (.A1(_07174_),
    .A2(_07172_),
    .Y(_07218_),
    .B1(_07173_));
 sg13g2_buf_1 _16439_ (.A(_00140_),
    .X(_07219_));
 sg13g2_nor2_1 _16440_ (.A(_06072_),
    .B(net251),
    .Y(_07220_));
 sg13g2_nand2_1 _16441_ (.Y(_07221_),
    .A(_06072_),
    .B(_04198_));
 sg13g2_nor2b_1 _16442_ (.A(_07220_),
    .B_N(_07221_),
    .Y(_07222_));
 sg13g2_xnor2_1 _16443_ (.Y(_07223_),
    .A(_07219_),
    .B(_07222_));
 sg13g2_xor2_1 _16444_ (.B(_07223_),
    .A(_07218_),
    .X(_07224_));
 sg13g2_xnor2_1 _16445_ (.Y(_07225_),
    .A(_07172_),
    .B(_07224_));
 sg13g2_xnor2_1 _16446_ (.Y(_07226_),
    .A(_07217_),
    .B(_07225_));
 sg13g2_nor2_1 _16447_ (.A(_07215_),
    .B(_07226_),
    .Y(_07227_));
 sg13g2_inv_1 _16448_ (.Y(_07228_),
    .A(_07227_));
 sg13g2_nand2_1 _16449_ (.Y(_07229_),
    .A(_07226_),
    .B(_07215_));
 sg13g2_nand2_1 _16450_ (.Y(_07230_),
    .A(_07228_),
    .B(_07229_));
 sg13g2_nor3_1 _16451_ (.A(_07162_),
    .B(_07179_),
    .C(_07163_),
    .Y(_07231_));
 sg13g2_nor2_1 _16452_ (.A(_07180_),
    .B(_07231_),
    .Y(_07232_));
 sg13g2_o21ai_1 _16453_ (.B1(_07232_),
    .Y(_07233_),
    .A1(_07183_),
    .A2(_07139_));
 sg13g2_inv_1 _16454_ (.Y(_07234_),
    .A(_07233_));
 sg13g2_buf_1 _16455_ (.A(_10106_),
    .X(_07235_));
 sg13g2_buf_1 _16456_ (.A(net162),
    .X(_07236_));
 sg13g2_a21oi_1 _16457_ (.A1(_07234_),
    .A2(_07230_),
    .Y(_07237_),
    .B1(net149));
 sg13g2_o21ai_1 _16458_ (.B1(_07237_),
    .Y(_07238_),
    .A1(_07230_),
    .A2(_07234_));
 sg13g2_a22oi_1 _16459_ (.Y(_00350_),
    .B1(_07213_),
    .B2(_07238_),
    .A2(net93),
    .A1(_04307_));
 sg13g2_nor2_1 _16460_ (.A(_07180_),
    .B(_07227_),
    .Y(_07239_));
 sg13g2_nand2_1 _16461_ (.Y(_07240_),
    .A(_07166_),
    .B(_07184_));
 sg13g2_a22oi_1 _16462_ (.Y(_07241_),
    .B1(_07239_),
    .B2(_07240_),
    .A2(_07226_),
    .A1(_07215_));
 sg13g2_nor2_1 _16463_ (.A(_07217_),
    .B(_07225_),
    .Y(_07242_));
 sg13g2_inv_1 _16464_ (.Y(_07243_),
    .A(_07242_));
 sg13g2_nor2_1 _16465_ (.A(_07218_),
    .B(_07223_),
    .Y(_07244_));
 sg13g2_a21oi_1 _16466_ (.A1(_07224_),
    .A2(_07172_),
    .Y(_07245_),
    .B1(_07244_));
 sg13g2_a21oi_1 _16467_ (.A1(_07221_),
    .A2(_07219_),
    .Y(_07246_),
    .B1(_07220_));
 sg13g2_buf_1 _16468_ (.A(_00141_),
    .X(_07247_));
 sg13g2_nor2_1 _16469_ (.A(_06078_),
    .B(net248),
    .Y(_07248_));
 sg13g2_nand2_1 _16470_ (.Y(_07249_),
    .A(_06078_),
    .B(_04223_));
 sg13g2_nor2b_1 _16471_ (.A(_07248_),
    .B_N(_07249_),
    .Y(_07250_));
 sg13g2_xnor2_1 _16472_ (.Y(_07251_),
    .A(_07247_),
    .B(_07250_));
 sg13g2_xor2_1 _16473_ (.B(_07251_),
    .A(_07246_),
    .X(_07252_));
 sg13g2_xnor2_1 _16474_ (.Y(_07253_),
    .A(_07219_),
    .B(_07252_));
 sg13g2_xnor2_1 _16475_ (.Y(_07254_),
    .A(_07245_),
    .B(_07253_));
 sg13g2_nor2_1 _16476_ (.A(_07243_),
    .B(_07254_),
    .Y(_07255_));
 sg13g2_inv_1 _16477_ (.Y(_07256_),
    .A(_07255_));
 sg13g2_nand2_1 _16478_ (.Y(_07257_),
    .A(_07254_),
    .B(_07243_));
 sg13g2_nand2_1 _16479_ (.Y(_07258_),
    .A(_07256_),
    .B(_07257_));
 sg13g2_nand2b_1 _16480_ (.Y(_07259_),
    .B(_07258_),
    .A_N(_07241_));
 sg13g2_nand2b_1 _16481_ (.Y(_07260_),
    .B(_07241_),
    .A_N(_07258_));
 sg13g2_nand3_1 _16482_ (.B(net151),
    .C(_07260_),
    .A(_07259_),
    .Y(_07261_));
 sg13g2_nor2_1 _16483_ (.A(_04310_),
    .B(_06102_),
    .Y(_07262_));
 sg13g2_nand2_1 _16484_ (.Y(_07263_),
    .A(_04310_),
    .B(_06102_));
 sg13g2_inv_1 _16485_ (.Y(_07264_),
    .A(_07263_));
 sg13g2_nor2_1 _16486_ (.A(_07262_),
    .B(_07264_),
    .Y(_07265_));
 sg13g2_inv_1 _16487_ (.Y(_07266_),
    .A(_07265_));
 sg13g2_nand2_1 _16488_ (.Y(_07267_),
    .A(_07190_),
    .B(_07204_));
 sg13g2_a21oi_1 _16489_ (.A1(_07199_),
    .A2(_07191_),
    .Y(_07268_),
    .B1(_07267_));
 sg13g2_nor2_1 _16490_ (.A(_07203_),
    .B(_07268_),
    .Y(_07269_));
 sg13g2_xnor2_1 _16491_ (.Y(_07270_),
    .A(_07266_),
    .B(_07269_));
 sg13g2_buf_1 _16492_ (.A(_06989_),
    .X(_07271_));
 sg13g2_a21oi_1 _16493_ (.A1(_07270_),
    .A2(net165),
    .Y(_07272_),
    .B1(net98));
 sg13g2_a22oi_1 _16494_ (.Y(_00351_),
    .B1(_07261_),
    .B2(_07272_),
    .A2(net93),
    .A1(_04321_));
 sg13g2_buf_1 _16495_ (.A(_10117_),
    .X(_07273_));
 sg13g2_nor2_1 _16496_ (.A(_04370_),
    .B(net228),
    .Y(_07274_));
 sg13g2_nand2_1 _16497_ (.Y(_07275_),
    .A(_04370_),
    .B(net228));
 sg13g2_nor2b_1 _16498_ (.A(_07274_),
    .B_N(_07275_),
    .Y(_07276_));
 sg13g2_inv_1 _16499_ (.Y(_07277_),
    .A(_07276_));
 sg13g2_nor2_1 _16500_ (.A(_07207_),
    .B(_07266_),
    .Y(_07278_));
 sg13g2_a221oi_1 _16501_ (.B2(_07278_),
    .C1(_07264_),
    .B1(_07211_),
    .A1(_07205_),
    .Y(_07279_),
    .A2(_07265_));
 sg13g2_nor2_1 _16502_ (.A(_07277_),
    .B(_07279_),
    .Y(_07280_));
 sg13g2_nor2_1 _16503_ (.A(_07273_),
    .B(_07280_),
    .Y(_07281_));
 sg13g2_nand2_1 _16504_ (.Y(_07282_),
    .A(_07279_),
    .B(_07277_));
 sg13g2_a21oi_1 _16505_ (.A1(_07281_),
    .A2(_07282_),
    .Y(_07283_),
    .B1(net99));
 sg13g2_or2_1 _16506_ (.X(_07284_),
    .B(_07253_),
    .A(_07245_));
 sg13g2_nor2_1 _16507_ (.A(_07246_),
    .B(_07251_),
    .Y(_07285_));
 sg13g2_a21oi_1 _16508_ (.A1(_07252_),
    .A2(_07219_),
    .Y(_07286_),
    .B1(_07285_));
 sg13g2_a21oi_1 _16509_ (.A1(_07249_),
    .A2(_07247_),
    .Y(_07287_),
    .B1(_07248_));
 sg13g2_buf_1 _16510_ (.A(_00142_),
    .X(_07288_));
 sg13g2_nor2_1 _16511_ (.A(_06085_),
    .B(net213),
    .Y(_07289_));
 sg13g2_nand2_1 _16512_ (.Y(_07290_),
    .A(_06085_),
    .B(net213));
 sg13g2_nor2b_1 _16513_ (.A(_07289_),
    .B_N(_07290_),
    .Y(_07291_));
 sg13g2_xnor2_1 _16514_ (.Y(_07292_),
    .A(_07288_),
    .B(_07291_));
 sg13g2_xor2_1 _16515_ (.B(_07292_),
    .A(_07287_),
    .X(_07293_));
 sg13g2_xnor2_1 _16516_ (.Y(_07294_),
    .A(_07247_),
    .B(_07293_));
 sg13g2_xnor2_1 _16517_ (.Y(_07295_),
    .A(_07286_),
    .B(_07294_));
 sg13g2_nor2_1 _16518_ (.A(_07284_),
    .B(_07295_),
    .Y(_07296_));
 sg13g2_nand2_1 _16519_ (.Y(_07297_),
    .A(_07295_),
    .B(_07284_));
 sg13g2_nand2b_1 _16520_ (.Y(_07298_),
    .B(_07297_),
    .A_N(_07296_));
 sg13g2_nand2_1 _16521_ (.Y(_07299_),
    .A(_07228_),
    .B(_07256_));
 sg13g2_nor2_1 _16522_ (.A(_07230_),
    .B(_07258_),
    .Y(_07300_));
 sg13g2_a22oi_1 _16523_ (.Y(_07301_),
    .B1(_07300_),
    .B2(_07233_),
    .A2(_07299_),
    .A1(_07257_));
 sg13g2_nor2_1 _16524_ (.A(_07298_),
    .B(_07301_),
    .Y(_07302_));
 sg13g2_inv_1 _16525_ (.Y(_07303_),
    .A(_07302_));
 sg13g2_nand2_1 _16526_ (.Y(_07304_),
    .A(_07301_),
    .B(_07298_));
 sg13g2_nand3_1 _16527_ (.B(_07304_),
    .C(net151),
    .A(_07303_),
    .Y(_07305_));
 sg13g2_a22oi_1 _16528_ (.Y(_00352_),
    .B1(_07283_),
    .B2(_07305_),
    .A2(net93),
    .A1(_04371_));
 sg13g2_a21oi_1 _16529_ (.A1(_07255_),
    .A2(_07297_),
    .Y(_07306_),
    .B1(_07296_));
 sg13g2_o21ai_1 _16530_ (.B1(_07306_),
    .Y(_07307_),
    .A1(_07298_),
    .A2(_07260_));
 sg13g2_inv_1 _16531_ (.Y(_07308_),
    .A(_07307_));
 sg13g2_nor2_1 _16532_ (.A(_07286_),
    .B(_07294_),
    .Y(_07309_));
 sg13g2_inv_1 _16533_ (.Y(_07310_),
    .A(_07309_));
 sg13g2_nor2_1 _16534_ (.A(_07287_),
    .B(_07292_),
    .Y(_07311_));
 sg13g2_a21oi_1 _16535_ (.A1(_07293_),
    .A2(_07247_),
    .Y(_07312_),
    .B1(_07311_));
 sg13g2_a21oi_1 _16536_ (.A1(_07290_),
    .A2(_07288_),
    .Y(_07313_),
    .B1(_07289_));
 sg13g2_buf_1 _16537_ (.A(_00143_),
    .X(_07314_));
 sg13g2_nor2_1 _16538_ (.A(_06091_),
    .B(net212),
    .Y(_07315_));
 sg13g2_nand2_1 _16539_ (.Y(_07316_),
    .A(_06091_),
    .B(net212));
 sg13g2_nor2b_1 _16540_ (.A(_07315_),
    .B_N(_07316_),
    .Y(_07317_));
 sg13g2_xnor2_1 _16541_ (.Y(_07318_),
    .A(_07314_),
    .B(_07317_));
 sg13g2_xor2_1 _16542_ (.B(_07318_),
    .A(_07313_),
    .X(_07319_));
 sg13g2_xnor2_1 _16543_ (.Y(_07320_),
    .A(_07288_),
    .B(_07319_));
 sg13g2_xnor2_1 _16544_ (.Y(_07321_),
    .A(_07312_),
    .B(_07320_));
 sg13g2_nor2_1 _16545_ (.A(_07310_),
    .B(_07321_),
    .Y(_07322_));
 sg13g2_nand2_1 _16546_ (.Y(_07323_),
    .A(_07321_),
    .B(_07310_));
 sg13g2_nand2b_1 _16547_ (.Y(_07324_),
    .B(_07323_),
    .A_N(_07322_));
 sg13g2_a21oi_1 _16548_ (.A1(_07308_),
    .A2(_07324_),
    .Y(_07325_),
    .B1(_07185_));
 sg13g2_nor2_1 _16549_ (.A(_07324_),
    .B(_07308_),
    .Y(_07326_));
 sg13g2_inv_1 _16550_ (.Y(_07327_),
    .A(_07326_));
 sg13g2_a21oi_1 _16551_ (.A1(_07325_),
    .A2(_07327_),
    .Y(_07328_),
    .B1(net99));
 sg13g2_nor2_1 _16552_ (.A(_04412_),
    .B(net197),
    .Y(_07329_));
 sg13g2_inv_1 _16553_ (.Y(_07330_),
    .A(_07329_));
 sg13g2_nand2_1 _16554_ (.Y(_07331_),
    .A(_04412_),
    .B(net197));
 sg13g2_nand2_1 _16555_ (.Y(_07332_),
    .A(_07330_),
    .B(_07331_));
 sg13g2_a221oi_1 _16556_ (.B2(_07265_),
    .C1(_07264_),
    .B1(_07269_),
    .A1(_04370_),
    .Y(_07333_),
    .A2(net228));
 sg13g2_or3_1 _16557_ (.A(_07274_),
    .B(_07332_),
    .C(_07333_),
    .X(_07334_));
 sg13g2_buf_1 _16558_ (.A(net162),
    .X(_07335_));
 sg13g2_o21ai_1 _16559_ (.B1(_07332_),
    .Y(_07336_),
    .A1(_07274_),
    .A2(_07333_));
 sg13g2_nand3_1 _16560_ (.B(_07335_),
    .C(_07336_),
    .A(_07334_),
    .Y(_07337_));
 sg13g2_a22oi_1 _16561_ (.Y(_00353_),
    .B1(_07328_),
    .B2(_07337_),
    .A2(_06991_),
    .A1(_04422_));
 sg13g2_xor2_1 _16562_ (.B(_04450_),
    .A(net197),
    .X(_07338_));
 sg13g2_inv_1 _16563_ (.Y(_07339_),
    .A(_07338_));
 sg13g2_nand2_1 _16564_ (.Y(_07340_),
    .A(_07275_),
    .B(_07331_));
 sg13g2_o21ai_1 _16565_ (.B1(_07330_),
    .Y(_07341_),
    .A1(_07340_),
    .A2(_07280_));
 sg13g2_nor2_1 _16566_ (.A(_07339_),
    .B(_07341_),
    .Y(_07342_));
 sg13g2_nor2_1 _16567_ (.A(net148),
    .B(_07342_),
    .Y(_07343_));
 sg13g2_nand2_1 _16568_ (.Y(_07344_),
    .A(_07341_),
    .B(_07339_));
 sg13g2_a21oi_1 _16569_ (.A1(_07343_),
    .A2(_07344_),
    .Y(_07345_),
    .B1(_07043_));
 sg13g2_a21oi_1 _16570_ (.A1(_07296_),
    .A2(_07323_),
    .Y(_07346_),
    .B1(_07322_));
 sg13g2_o21ai_1 _16571_ (.B1(_07346_),
    .Y(_07347_),
    .A1(_07324_),
    .A2(_07303_));
 sg13g2_nor2_1 _16572_ (.A(_07312_),
    .B(_07320_),
    .Y(_07348_));
 sg13g2_inv_1 _16573_ (.Y(_07349_),
    .A(_07348_));
 sg13g2_nor2_1 _16574_ (.A(_07313_),
    .B(_07318_),
    .Y(_07350_));
 sg13g2_a21oi_1 _16575_ (.A1(_07319_),
    .A2(_07288_),
    .Y(_07351_),
    .B1(_07350_));
 sg13g2_a21oi_1 _16576_ (.A1(_07316_),
    .A2(_07314_),
    .Y(_07352_),
    .B1(_07315_));
 sg13g2_nor2_1 _16577_ (.A(_06035_),
    .B(net211),
    .Y(_07353_));
 sg13g2_nand2_1 _16578_ (.Y(_07354_),
    .A(_06035_),
    .B(net211));
 sg13g2_nor2b_1 _16579_ (.A(_07353_),
    .B_N(_07354_),
    .Y(_07355_));
 sg13g2_xnor2_1 _16580_ (.Y(_07356_),
    .A(_06111_),
    .B(_07355_));
 sg13g2_xor2_1 _16581_ (.B(_07356_),
    .A(_07352_),
    .X(_07357_));
 sg13g2_xnor2_1 _16582_ (.Y(_07358_),
    .A(_07314_),
    .B(_07357_));
 sg13g2_xnor2_1 _16583_ (.Y(_07359_),
    .A(_07351_),
    .B(_07358_));
 sg13g2_nor2_1 _16584_ (.A(_07349_),
    .B(_07359_),
    .Y(_07360_));
 sg13g2_inv_1 _16585_ (.Y(_07361_),
    .A(_07360_));
 sg13g2_nand2_1 _16586_ (.Y(_07362_),
    .A(_07359_),
    .B(_07349_));
 sg13g2_nand2_1 _16587_ (.Y(_07363_),
    .A(_07361_),
    .B(_07362_));
 sg13g2_nand2b_1 _16588_ (.Y(_07364_),
    .B(_07363_),
    .A_N(_07347_));
 sg13g2_nand2b_1 _16589_ (.Y(_07365_),
    .B(_07347_),
    .A_N(_07363_));
 sg13g2_nand3_1 _16590_ (.B(net151),
    .C(_07365_),
    .A(_07364_),
    .Y(_07366_));
 sg13g2_a22oi_1 _16591_ (.Y(_00354_),
    .B1(_07345_),
    .B2(_07366_),
    .A2(_06991_),
    .A1(_04451_));
 sg13g2_buf_1 _16592_ (.A(net100),
    .X(_07367_));
 sg13g2_a21oi_1 _16593_ (.A1(_07322_),
    .A2(_07362_),
    .Y(_07368_),
    .B1(_07360_));
 sg13g2_o21ai_1 _16594_ (.B1(_07368_),
    .Y(_07369_),
    .A1(_07363_),
    .A2(_07327_));
 sg13g2_inv_1 _16595_ (.Y(_07370_),
    .A(_07369_));
 sg13g2_nor2_1 _16596_ (.A(_07351_),
    .B(_07358_),
    .Y(_07371_));
 sg13g2_inv_1 _16597_ (.Y(_07372_),
    .A(_07371_));
 sg13g2_a21oi_1 _16598_ (.A1(_07354_),
    .A2(_06111_),
    .Y(_07373_),
    .B1(_07353_));
 sg13g2_inv_2 _16599_ (.Y(_07374_),
    .A(_00144_));
 sg13g2_xnor2_1 _16600_ (.Y(_07375_),
    .A(_06033_),
    .B(net247));
 sg13g2_xnor2_1 _16601_ (.Y(_07376_),
    .A(_07374_),
    .B(_07375_));
 sg13g2_xnor2_1 _16602_ (.Y(_07377_),
    .A(_07373_),
    .B(_07376_));
 sg13g2_xnor2_1 _16603_ (.Y(_07378_),
    .A(_06108_),
    .B(_07377_));
 sg13g2_nor2_1 _16604_ (.A(_07352_),
    .B(_07356_),
    .Y(_07379_));
 sg13g2_a21oi_1 _16605_ (.A1(_07357_),
    .A2(_07314_),
    .Y(_07380_),
    .B1(_07379_));
 sg13g2_xnor2_1 _16606_ (.Y(_07381_),
    .A(_07378_),
    .B(_07380_));
 sg13g2_nor2_1 _16607_ (.A(_07372_),
    .B(_07381_),
    .Y(_07382_));
 sg13g2_nand2_1 _16608_ (.Y(_07383_),
    .A(_07381_),
    .B(_07372_));
 sg13g2_nand2b_1 _16609_ (.Y(_07384_),
    .B(_07383_),
    .A_N(_07382_));
 sg13g2_a21oi_1 _16610_ (.A1(_07370_),
    .A2(_07384_),
    .Y(_07385_),
    .B1(_07185_));
 sg13g2_nor2_1 _16611_ (.A(_07384_),
    .B(_07370_),
    .Y(_07386_));
 sg13g2_inv_1 _16612_ (.Y(_07387_),
    .A(_07386_));
 sg13g2_a21oi_1 _16613_ (.A1(_07385_),
    .A2(_07387_),
    .Y(_07388_),
    .B1(_07043_));
 sg13g2_o21ai_1 _16614_ (.B1(net183),
    .Y(_07389_),
    .A1(_04412_),
    .A2(_04450_));
 sg13g2_o21ai_1 _16615_ (.B1(_07389_),
    .Y(_07390_),
    .A1(_07339_),
    .A2(_07334_));
 sg13g2_buf_1 _16616_ (.A(_07390_),
    .X(_07391_));
 sg13g2_xor2_1 _16617_ (.B(_04493_),
    .A(net183),
    .X(_07392_));
 sg13g2_a21oi_1 _16618_ (.A1(_07391_),
    .A2(_07392_),
    .Y(_07393_),
    .B1(_07273_));
 sg13g2_o21ai_1 _16619_ (.B1(_07393_),
    .Y(_07394_),
    .A1(_07391_),
    .A2(_07392_));
 sg13g2_a22oi_1 _16620_ (.Y(_00355_),
    .B1(_07388_),
    .B2(_07394_),
    .A2(net92),
    .A1(_04494_));
 sg13g2_xor2_1 _16621_ (.B(_04532_),
    .A(net197),
    .X(_07395_));
 sg13g2_inv_1 _16622_ (.Y(_07396_),
    .A(_07395_));
 sg13g2_nand2_1 _16623_ (.Y(_07397_),
    .A(_07342_),
    .B(_07392_));
 sg13g2_o21ai_1 _16624_ (.B1(net183),
    .Y(_07398_),
    .A1(_04450_),
    .A2(_04493_));
 sg13g2_nand2_1 _16625_ (.Y(_07399_),
    .A(_07397_),
    .B(_07398_));
 sg13g2_xnor2_1 _16626_ (.Y(_07400_),
    .A(_07396_),
    .B(_07399_));
 sg13g2_buf_1 _16627_ (.A(_06989_),
    .X(_07401_));
 sg13g2_a21oi_1 _16628_ (.A1(_07400_),
    .A2(_07042_),
    .Y(_07402_),
    .B1(net97));
 sg13g2_o21ai_1 _16629_ (.B1(_07383_),
    .Y(_07403_),
    .A1(_07382_),
    .A2(_07360_));
 sg13g2_o21ai_1 _16630_ (.B1(_07403_),
    .Y(_07404_),
    .A1(_07384_),
    .A2(_07365_));
 sg13g2_nor2_1 _16631_ (.A(_07378_),
    .B(_07380_),
    .Y(_07405_));
 sg13g2_inv_1 _16632_ (.Y(_07406_),
    .A(_07405_));
 sg13g2_nand2_1 _16633_ (.Y(_07407_),
    .A(_06034_),
    .B(_06067_));
 sg13g2_a21oi_1 _16634_ (.A1(_06033_),
    .A2(net247),
    .Y(_07408_),
    .B1(_07374_));
 sg13g2_a21oi_1 _16635_ (.A1(_07374_),
    .A2(_07407_),
    .Y(_07409_),
    .B1(_07408_));
 sg13g2_xnor2_1 _16636_ (.Y(_07410_),
    .A(_06031_),
    .B(net210));
 sg13g2_xnor2_1 _16637_ (.Y(_07411_),
    .A(_06029_),
    .B(_07410_));
 sg13g2_xnor2_1 _16638_ (.Y(_07412_),
    .A(_07409_),
    .B(_07411_));
 sg13g2_nor2_1 _16639_ (.A(_07373_),
    .B(_07376_),
    .Y(_07413_));
 sg13g2_nor2_1 _16640_ (.A(net228),
    .B(_07377_),
    .Y(_07414_));
 sg13g2_nor2_1 _16641_ (.A(_07413_),
    .B(_07414_),
    .Y(_07415_));
 sg13g2_xnor2_1 _16642_ (.Y(_07416_),
    .A(_07412_),
    .B(_07415_));
 sg13g2_inv_1 _16643_ (.Y(_07417_),
    .A(_07416_));
 sg13g2_nor2_1 _16644_ (.A(_07406_),
    .B(_07417_),
    .Y(_07418_));
 sg13g2_inv_1 _16645_ (.Y(_07419_),
    .A(_07418_));
 sg13g2_nand2_1 _16646_ (.Y(_07420_),
    .A(_07417_),
    .B(_07406_));
 sg13g2_nand2_1 _16647_ (.Y(_07421_),
    .A(_07419_),
    .B(_07420_));
 sg13g2_nand2b_1 _16648_ (.Y(_07422_),
    .B(_07421_),
    .A_N(_07404_));
 sg13g2_nand2b_1 _16649_ (.Y(_07423_),
    .B(_07404_),
    .A_N(_07421_));
 sg13g2_nand3_1 _16650_ (.B(_07140_),
    .C(_07423_),
    .A(_07422_),
    .Y(_07424_));
 sg13g2_a22oi_1 _16651_ (.Y(_00356_),
    .B1(_07402_),
    .B2(_07424_),
    .A2(net92),
    .A1(_06922_));
 sg13g2_a21oi_1 _16652_ (.A1(_07382_),
    .A2(_07420_),
    .Y(_07425_),
    .B1(_07418_));
 sg13g2_o21ai_1 _16653_ (.B1(_07425_),
    .Y(_07426_),
    .A1(_07421_),
    .A2(_07387_));
 sg13g2_inv_1 _16654_ (.Y(_07427_),
    .A(_07426_));
 sg13g2_nand2b_1 _16655_ (.Y(_07428_),
    .B(_07407_),
    .A_N(_07408_));
 sg13g2_nand2_1 _16656_ (.Y(_07429_),
    .A(_07410_),
    .B(net197));
 sg13g2_o21ai_1 _16657_ (.B1(_07429_),
    .Y(_07430_),
    .A1(_07410_),
    .A2(_07428_));
 sg13g2_nor2_1 _16658_ (.A(_06102_),
    .B(net209),
    .Y(_07431_));
 sg13g2_inv_1 _16659_ (.Y(_07432_),
    .A(_07431_));
 sg13g2_nand2_1 _16660_ (.Y(_07433_),
    .A(_06102_),
    .B(net209));
 sg13g2_nand2_1 _16661_ (.Y(_07434_),
    .A(_07432_),
    .B(_07433_));
 sg13g2_xnor2_1 _16662_ (.Y(_07435_),
    .A(_06029_),
    .B(_07434_));
 sg13g2_nor2_1 _16663_ (.A(_06031_),
    .B(_04496_),
    .Y(_07436_));
 sg13g2_a21oi_1 _16664_ (.A1(_06031_),
    .A2(net210),
    .Y(_07437_),
    .B1(_07374_));
 sg13g2_nor2_1 _16665_ (.A(_07436_),
    .B(_07437_),
    .Y(_07438_));
 sg13g2_a21oi_1 _16666_ (.A1(_07438_),
    .A2(_07374_),
    .Y(_07439_),
    .B1(_07437_));
 sg13g2_xnor2_1 _16667_ (.Y(_07440_),
    .A(_07435_),
    .B(_07439_));
 sg13g2_xor2_1 _16668_ (.B(_07440_),
    .A(_07430_),
    .X(_07441_));
 sg13g2_nor2b_1 _16669_ (.A(_07415_),
    .B_N(_07412_),
    .Y(_07442_));
 sg13g2_inv_1 _16670_ (.Y(_07443_),
    .A(_07442_));
 sg13g2_nor2_1 _16671_ (.A(_07441_),
    .B(_07443_),
    .Y(_07444_));
 sg13g2_nand2_1 _16672_ (.Y(_07445_),
    .A(_07443_),
    .B(_07441_));
 sg13g2_inv_1 _16673_ (.Y(_07446_),
    .A(_07445_));
 sg13g2_nor2_1 _16674_ (.A(_07444_),
    .B(_07446_),
    .Y(_07447_));
 sg13g2_inv_1 _16675_ (.Y(_07448_),
    .A(_07447_));
 sg13g2_a21oi_1 _16676_ (.A1(_07427_),
    .A2(_07448_),
    .Y(_07449_),
    .B1(net147));
 sg13g2_nor2_1 _16677_ (.A(_07448_),
    .B(_07427_),
    .Y(_07450_));
 sg13g2_inv_1 _16678_ (.Y(_07451_),
    .A(_07450_));
 sg13g2_nand2_1 _16679_ (.Y(_07452_),
    .A(_07449_),
    .B(_07451_));
 sg13g2_xor2_1 _16680_ (.B(_04571_),
    .A(_06030_),
    .X(_07453_));
 sg13g2_inv_1 _16681_ (.Y(_07454_),
    .A(_07453_));
 sg13g2_nand2_1 _16682_ (.Y(_07455_),
    .A(_07392_),
    .B(_07395_));
 sg13g2_inv_1 _16683_ (.Y(_07456_),
    .A(_07391_));
 sg13g2_o21ai_1 _16684_ (.B1(net183),
    .Y(_07457_),
    .A1(_04493_),
    .A2(_04532_));
 sg13g2_o21ai_1 _16685_ (.B1(_07457_),
    .Y(_07458_),
    .A1(_07455_),
    .A2(_07456_));
 sg13g2_xnor2_1 _16686_ (.Y(_07459_),
    .A(_07454_),
    .B(_07458_));
 sg13g2_a21oi_1 _16687_ (.A1(_07459_),
    .A2(_06983_),
    .Y(_07460_),
    .B1(_07271_));
 sg13g2_a22oi_1 _16688_ (.Y(_00357_),
    .B1(_07452_),
    .B2(_07460_),
    .A2(net92),
    .A1(_04572_));
 sg13g2_nand2b_1 _16689_ (.Y(_07461_),
    .B(_06984_),
    .A_N(_06997_));
 sg13g2_nand4_1 _16690_ (.B(net165),
    .C(_06998_),
    .A(net107),
    .Y(_07462_),
    .D(_07461_));
 sg13g2_o21ai_1 _16691_ (.B1(_07462_),
    .Y(_00358_),
    .A1(_06996_),
    .A2(net105));
 sg13g2_xor2_1 _16692_ (.B(\vgadonut.donut.donuthit.rxin[14] ),
    .A(net183),
    .X(_07463_));
 sg13g2_inv_1 _16693_ (.Y(_07464_),
    .A(_07397_));
 sg13g2_nor2_1 _16694_ (.A(_07396_),
    .B(_07454_),
    .Y(_07465_));
 sg13g2_inv_1 _16695_ (.Y(_07466_),
    .A(_07465_));
 sg13g2_o21ai_1 _16696_ (.B1(_06892_),
    .Y(_07467_),
    .A1(_04532_),
    .A2(_04571_));
 sg13g2_o21ai_1 _16697_ (.B1(_07467_),
    .Y(_07468_),
    .A1(_07398_),
    .A2(_07466_));
 sg13g2_a21oi_1 _16698_ (.A1(_07464_),
    .A2(_07465_),
    .Y(_07469_),
    .B1(_07468_));
 sg13g2_xnor2_1 _16699_ (.Y(_07470_),
    .A(_07463_),
    .B(_07469_));
 sg13g2_a21oi_1 _16700_ (.A1(_07470_),
    .A2(_07042_),
    .Y(_07471_),
    .B1(net97));
 sg13g2_nor3_1 _16701_ (.A(_07436_),
    .B(_07437_),
    .C(_07434_),
    .Y(_07472_));
 sg13g2_a21oi_1 _16702_ (.A1(net197),
    .A2(_07434_),
    .Y(_07473_),
    .B1(_07472_));
 sg13g2_a21oi_1 _16703_ (.A1(_06102_),
    .A2(net209),
    .Y(_07474_),
    .B1(_07374_));
 sg13g2_a21oi_1 _16704_ (.A1(_07374_),
    .A2(_07432_),
    .Y(_07475_),
    .B1(_07474_));
 sg13g2_nor2_1 _16705_ (.A(net228),
    .B(net246),
    .Y(_07476_));
 sg13g2_nand2_1 _16706_ (.Y(_07477_),
    .A(net228),
    .B(net246));
 sg13g2_nand2b_1 _16707_ (.Y(_07478_),
    .B(_07477_),
    .A_N(_07476_));
 sg13g2_xnor2_1 _16708_ (.Y(_07479_),
    .A(net197),
    .B(_07478_));
 sg13g2_xnor2_1 _16709_ (.Y(_07480_),
    .A(_07475_),
    .B(_07479_));
 sg13g2_xnor2_1 _16710_ (.Y(_07481_),
    .A(_07473_),
    .B(_07480_));
 sg13g2_nor2b_1 _16711_ (.A(_07430_),
    .B_N(_07440_),
    .Y(_07482_));
 sg13g2_inv_1 _16712_ (.Y(_07483_),
    .A(_07482_));
 sg13g2_nor2_1 _16713_ (.A(_07481_),
    .B(_07483_),
    .Y(_07484_));
 sg13g2_nand2_1 _16714_ (.Y(_07485_),
    .A(_07483_),
    .B(_07481_));
 sg13g2_inv_1 _16715_ (.Y(_07486_),
    .A(_07485_));
 sg13g2_nor2_1 _16716_ (.A(_07484_),
    .B(_07486_),
    .Y(_07487_));
 sg13g2_nor2_1 _16717_ (.A(_07444_),
    .B(_07418_),
    .Y(_07488_));
 sg13g2_a21oi_1 _16718_ (.A1(_07423_),
    .A2(_07488_),
    .Y(_07489_),
    .B1(_07446_));
 sg13g2_a21oi_1 _16719_ (.A1(_07489_),
    .A2(_07487_),
    .Y(_07490_),
    .B1(_07236_));
 sg13g2_o21ai_1 _16720_ (.B1(_07490_),
    .Y(_07491_),
    .A1(_07487_),
    .A2(_07489_));
 sg13g2_a22oi_1 _16721_ (.Y(_00359_),
    .B1(_07471_),
    .B2(_07491_),
    .A2(_07367_),
    .A1(_04601_));
 sg13g2_xnor2_1 _16722_ (.Y(_07492_),
    .A(net183),
    .B(_04660_));
 sg13g2_nand2_1 _16723_ (.Y(_07493_),
    .A(_07453_),
    .B(_07463_));
 sg13g2_nor2_1 _16724_ (.A(_07455_),
    .B(_07493_),
    .Y(_07494_));
 sg13g2_o21ai_1 _16725_ (.B1(_06892_),
    .Y(_07495_),
    .A1(_04571_),
    .A2(\vgadonut.donut.donuthit.rxin[14] ));
 sg13g2_o21ai_1 _16726_ (.B1(_07495_),
    .Y(_07496_),
    .A1(_07457_),
    .A2(_07493_));
 sg13g2_a21oi_1 _16727_ (.A1(_07391_),
    .A2(_07494_),
    .Y(_07497_),
    .B1(_07496_));
 sg13g2_xor2_1 _16728_ (.B(_07497_),
    .A(_07492_),
    .X(_07498_));
 sg13g2_buf_1 _16729_ (.A(net170),
    .X(_07499_));
 sg13g2_a21oi_1 _16730_ (.A1(_07498_),
    .A2(_07499_),
    .Y(_07500_),
    .B1(net97));
 sg13g2_nor2_1 _16731_ (.A(_07484_),
    .B(_07444_),
    .Y(_07501_));
 sg13g2_a21oi_1 _16732_ (.A1(_07451_),
    .A2(_07501_),
    .Y(_07502_),
    .B1(_07486_));
 sg13g2_nand2_1 _16733_ (.Y(_07503_),
    .A(_07480_),
    .B(_07473_));
 sg13g2_a21oi_1 _16734_ (.A1(_07477_),
    .A2(_00144_),
    .Y(_07504_),
    .B1(_07476_));
 sg13g2_xnor2_1 _16735_ (.Y(_07505_),
    .A(_06116_),
    .B(_07504_));
 sg13g2_nor3_1 _16736_ (.A(_07431_),
    .B(_07474_),
    .C(_07478_),
    .Y(_07506_));
 sg13g2_a21oi_1 _16737_ (.A1(net183),
    .A2(_07478_),
    .Y(_07507_),
    .B1(_07506_));
 sg13g2_xnor2_1 _16738_ (.Y(_07508_),
    .A(_07505_),
    .B(_07507_));
 sg13g2_xor2_1 _16739_ (.B(_07508_),
    .A(_07503_),
    .X(_07509_));
 sg13g2_nand2b_1 _16740_ (.Y(_07510_),
    .B(_07509_),
    .A_N(_07502_));
 sg13g2_nand2b_1 _16741_ (.Y(_07511_),
    .B(_07502_),
    .A_N(_07509_));
 sg13g2_nand3_1 _16742_ (.B(_07140_),
    .C(_07511_),
    .A(_07510_),
    .Y(_07512_));
 sg13g2_a22oi_1 _16743_ (.Y(_00360_),
    .B1(_07500_),
    .B2(_07512_),
    .A2(net92),
    .A1(_04704_));
 sg13g2_nor2_1 _16744_ (.A(_07000_),
    .B(_07003_),
    .Y(_07513_));
 sg13g2_o21ai_1 _16745_ (.B1(net162),
    .Y(_07514_),
    .A1(_07513_),
    .A2(_06999_));
 sg13g2_a21oi_1 _16746_ (.A1(_06999_),
    .A2(_07513_),
    .Y(_07515_),
    .B1(_07514_));
 sg13g2_a21oi_1 _16747_ (.A1(net230),
    .A2(net150),
    .Y(_07516_),
    .B1(_07515_));
 sg13g2_buf_1 _16748_ (.A(_06980_),
    .X(_07517_));
 sg13g2_nor2_1 _16749_ (.A(\vgadonut.donut.rx6[2] ),
    .B(net104),
    .Y(_07518_));
 sg13g2_a21oi_1 _16750_ (.A1(_06981_),
    .A2(_07516_),
    .Y(_00361_),
    .B1(_07518_));
 sg13g2_nand2b_1 _16751_ (.Y(_07519_),
    .B(_07005_),
    .A_N(_07006_));
 sg13g2_xor2_1 _16752_ (.B(_07004_),
    .A(_07519_),
    .X(_07520_));
 sg13g2_buf_1 _16753_ (.A(_06982_),
    .X(_07521_));
 sg13g2_buf_1 _16754_ (.A(net162),
    .X(_07522_));
 sg13g2_nor2_1 _16755_ (.A(_06894_),
    .B(net146),
    .Y(_07523_));
 sg13g2_a21oi_1 _16756_ (.A1(_07520_),
    .A2(net160),
    .Y(_07524_),
    .B1(_07523_));
 sg13g2_nor2_1 _16757_ (.A(\vgadonut.donut.rx6[3] ),
    .B(net104),
    .Y(_07525_));
 sg13g2_a21oi_1 _16758_ (.A1(_07524_),
    .A2(_06981_),
    .Y(_00362_),
    .B1(_07525_));
 sg13g2_inv_1 _16759_ (.Y(_07526_),
    .A(\vgadonut.donut.rx6[4] ));
 sg13g2_nand2_1 _16760_ (.Y(_07527_),
    .A(_07009_),
    .B(_07010_));
 sg13g2_xnor2_1 _16761_ (.Y(_07528_),
    .A(_07527_),
    .B(_07007_));
 sg13g2_xnor2_1 _16762_ (.Y(_07529_),
    .A(net190),
    .B(net230));
 sg13g2_a21oi_1 _16763_ (.A1(net148),
    .A2(_07529_),
    .Y(_07530_),
    .B1(net100));
 sg13g2_o21ai_1 _16764_ (.B1(_07530_),
    .Y(_07531_),
    .A1(net150),
    .A2(_07528_));
 sg13g2_o21ai_1 _16765_ (.B1(_07531_),
    .Y(_00363_),
    .A1(_07526_),
    .A2(_07517_));
 sg13g2_buf_1 _16766_ (.A(net100),
    .X(_07532_));
 sg13g2_inv_1 _16767_ (.Y(_07533_),
    .A(net170));
 sg13g2_xnor2_1 _16768_ (.Y(_07534_),
    .A(_07148_),
    .B(_07152_));
 sg13g2_nand2b_1 _16769_ (.Y(_07535_),
    .B(_07013_),
    .A_N(_06995_));
 sg13g2_or2_1 _16770_ (.X(_07536_),
    .B(_07012_),
    .A(_07535_));
 sg13g2_a21oi_1 _16771_ (.A1(_07012_),
    .A2(_07535_),
    .Y(_07537_),
    .B1(_10117_));
 sg13g2_a22oi_1 _16772_ (.Y(_07538_),
    .B1(_07536_),
    .B2(_07537_),
    .A2(_07534_),
    .A1(_07533_));
 sg13g2_nand2_1 _16773_ (.Y(_07539_),
    .A(net98),
    .B(\vgadonut.donut.rx6[5] ));
 sg13g2_o21ai_1 _16774_ (.B1(_07539_),
    .Y(_00364_),
    .A1(net91),
    .A2(_07538_));
 sg13g2_inv_1 _16775_ (.Y(_07540_),
    .A(\vgadonut.donut.donuthit.rxin[0] ));
 sg13g2_nand2_1 _16776_ (.Y(_07541_),
    .A(_07115_),
    .B(_07106_));
 sg13g2_nand3b_1 _16777_ (.B(_07200_),
    .C(_07541_),
    .Y(_07542_),
    .A_N(_07116_));
 sg13g2_xnor2_1 _16778_ (.Y(_07543_),
    .A(_07023_),
    .B(_07014_));
 sg13g2_a21oi_1 _16779_ (.A1(_07543_),
    .A2(_06983_),
    .Y(_07544_),
    .B1(_07271_));
 sg13g2_a22oi_1 _16780_ (.Y(_00365_),
    .B1(_07542_),
    .B2(_07544_),
    .A2(net92),
    .A1(_07540_));
 sg13g2_inv_1 _16781_ (.Y(_07545_),
    .A(\vgadonut.donut.donuthit.rxin[1] ));
 sg13g2_xnor2_1 _16782_ (.Y(_07546_),
    .A(_07019_),
    .B(_07193_));
 sg13g2_a21oi_1 _16783_ (.A1(_07546_),
    .A2(net161),
    .Y(_07547_),
    .B1(_07401_));
 sg13g2_a21oi_1 _16784_ (.A1(_07155_),
    .A2(_07121_),
    .Y(_07548_),
    .B1(_07236_));
 sg13g2_o21ai_1 _16785_ (.B1(_07548_),
    .Y(_07549_),
    .A1(_07121_),
    .A2(_07155_));
 sg13g2_a22oi_1 _16786_ (.Y(_00366_),
    .B1(_07547_),
    .B2(_07549_),
    .A2(net92),
    .A1(_07545_));
 sg13g2_inv_1 _16787_ (.Y(_07550_),
    .A(_07033_));
 sg13g2_xnor2_1 _16788_ (.Y(_07551_),
    .A(_07037_),
    .B(_07026_));
 sg13g2_a21oi_1 _16789_ (.A1(_07551_),
    .A2(_07499_),
    .Y(_07552_),
    .B1(_07401_));
 sg13g2_a21oi_1 _16790_ (.A1(_07126_),
    .A2(_07096_),
    .Y(_07553_),
    .B1(_07335_));
 sg13g2_nand2b_1 _16791_ (.Y(_07554_),
    .B(_07553_),
    .A_N(_07127_));
 sg13g2_a22oi_1 _16792_ (.Y(_00367_),
    .B1(_07552_),
    .B2(_07554_),
    .A2(_07367_),
    .A1(_07550_));
 sg13g2_o21ai_1 _16793_ (.B1(_07032_),
    .Y(_07555_),
    .A1(_07034_),
    .A2(_07194_));
 sg13g2_nand3_1 _16794_ (.B(_07235_),
    .C(_07196_),
    .A(_07555_),
    .Y(_07556_));
 sg13g2_a21oi_1 _16795_ (.A1(_07160_),
    .A2(_07130_),
    .Y(_07557_),
    .B1(_07235_));
 sg13g2_o21ai_1 _16796_ (.B1(_07557_),
    .Y(_07558_),
    .A1(_07130_),
    .A2(_07160_));
 sg13g2_a21oi_1 _16797_ (.A1(_07556_),
    .A2(_07558_),
    .Y(_07559_),
    .B1(_06990_));
 sg13g2_a21o_1 _16798_ (.A2(net98),
    .A1(\vgadonut.donut.donuthit.rxin[3] ),
    .B1(_07559_),
    .X(_00368_));
 sg13g2_inv_1 _16799_ (.Y(_07560_),
    .A(\vgadonut.donut.ry6[0] ));
 sg13g2_inv_1 _16800_ (.Y(_07561_),
    .A(\vgadonut.donut.ycA[0] ));
 sg13g2_buf_2 _16801_ (.A(\vgadonut.donut.sAsB[0] ),
    .X(_07562_));
 sg13g2_nand2_1 _16802_ (.Y(_07563_),
    .A(\vgadonut.donut.ry6[0] ),
    .B(_07562_));
 sg13g2_inv_1 _16803_ (.Y(_07564_),
    .A(_07562_));
 sg13g2_nand2_1 _16804_ (.Y(_07565_),
    .A(_07560_),
    .B(_07564_));
 sg13g2_nand3_1 _16805_ (.B(_07563_),
    .C(_07565_),
    .A(_06334_),
    .Y(_07566_));
 sg13g2_o21ai_1 _16806_ (.B1(_07566_),
    .Y(_07567_),
    .A1(_07561_),
    .A2(net170));
 sg13g2_nand2_1 _16807_ (.Y(_07568_),
    .A(net104),
    .B(_07567_));
 sg13g2_o21ai_1 _16808_ (.B1(_07568_),
    .Y(_00369_),
    .A1(_07560_),
    .A2(net104));
 sg13g2_buf_1 _16809_ (.A(\vgadonut.donut.sAsB[4] ),
    .X(_07569_));
 sg13g2_buf_1 _16810_ (.A(\vgadonut.donut.sAsB[2] ),
    .X(_07570_));
 sg13g2_buf_1 _16811_ (.A(\vgadonut.donut.sAsB[3] ),
    .X(_07571_));
 sg13g2_buf_1 _16812_ (.A(\vgadonut.donut.sAsB[1] ),
    .X(_07572_));
 sg13g2_nor2_1 _16813_ (.A(_07562_),
    .B(_07572_),
    .Y(_07573_));
 sg13g2_inv_1 _16814_ (.Y(_07574_),
    .A(_07573_));
 sg13g2_nor3_1 _16815_ (.A(_07570_),
    .B(_07571_),
    .C(_07574_),
    .Y(_07575_));
 sg13g2_inv_1 _16816_ (.Y(_07576_),
    .A(_07575_));
 sg13g2_nor3_1 _16817_ (.A(_07569_),
    .B(_06420_),
    .C(_07576_),
    .Y(_07577_));
 sg13g2_xnor2_1 _16818_ (.Y(_07578_),
    .A(_06417_),
    .B(_07577_));
 sg13g2_buf_2 _16819_ (.A(_07578_),
    .X(_07579_));
 sg13g2_inv_1 _16820_ (.Y(_07580_),
    .A(_07579_));
 sg13g2_buf_1 _16821_ (.A(\vgadonut.donut.ycA[7] ),
    .X(_07581_));
 sg13g2_inv_1 _16822_ (.Y(_07582_),
    .A(_07581_));
 sg13g2_nand2_1 _16823_ (.Y(_07583_),
    .A(_07562_),
    .B(_07572_));
 sg13g2_nand2_1 _16824_ (.Y(_07584_),
    .A(_07574_),
    .B(_07583_));
 sg13g2_buf_2 _16825_ (.A(_07584_),
    .X(_07585_));
 sg13g2_xnor2_1 _16826_ (.Y(_07586_),
    .A(_07581_),
    .B(_04824_));
 sg13g2_nand2_1 _16827_ (.Y(_07587_),
    .A(_07585_),
    .B(_07586_));
 sg13g2_o21ai_1 _16828_ (.B1(_07587_),
    .Y(_07588_),
    .A1(_07582_),
    .A2(_04824_));
 sg13g2_buf_1 _16829_ (.A(\vgadonut.donut.ycA[8] ),
    .X(_07589_));
 sg13g2_xnor2_1 _16830_ (.Y(_07590_),
    .A(_07589_),
    .B(_04823_));
 sg13g2_xnor2_1 _16831_ (.Y(_07591_),
    .A(_07570_),
    .B(_07573_));
 sg13g2_buf_1 _16832_ (.A(_07591_),
    .X(_07592_));
 sg13g2_xor2_1 _16833_ (.B(_07592_),
    .A(_07590_),
    .X(_07593_));
 sg13g2_xnor2_1 _16834_ (.Y(_07594_),
    .A(_07588_),
    .B(_07593_));
 sg13g2_nor2b_1 _16835_ (.A(_07593_),
    .B_N(_07588_),
    .Y(_07595_));
 sg13g2_a21oi_1 _16836_ (.A1(_07580_),
    .A2(_07594_),
    .Y(_07596_),
    .B1(_07595_));
 sg13g2_inv_1 _16837_ (.Y(_07597_),
    .A(_07589_));
 sg13g2_inv_1 _16838_ (.Y(_07598_),
    .A(_07592_));
 sg13g2_nand2_1 _16839_ (.Y(_07599_),
    .A(_07598_),
    .B(_07590_));
 sg13g2_o21ai_1 _16840_ (.B1(_07599_),
    .Y(_07600_),
    .A1(_07597_),
    .A2(_04823_));
 sg13g2_buf_1 _16841_ (.A(\vgadonut.donut.ycA[9] ),
    .X(_07601_));
 sg13g2_xnor2_1 _16842_ (.Y(_07602_),
    .A(_07601_),
    .B(_04820_));
 sg13g2_inv_1 _16843_ (.Y(_07603_),
    .A(_00121_));
 sg13g2_nor3_1 _16844_ (.A(_07572_),
    .B(_07570_),
    .C(_07603_),
    .Y(_07604_));
 sg13g2_xnor2_1 _16845_ (.Y(_07605_),
    .A(_07571_),
    .B(_07604_));
 sg13g2_buf_1 _16846_ (.A(_07605_),
    .X(_07606_));
 sg13g2_xor2_1 _16847_ (.B(_07606_),
    .A(_07602_),
    .X(_07607_));
 sg13g2_xor2_1 _16848_ (.B(_07607_),
    .A(_07600_),
    .X(_07608_));
 sg13g2_inv_1 _16849_ (.Y(_07609_),
    .A(_07604_));
 sg13g2_nor3_1 _16850_ (.A(_07571_),
    .B(_07569_),
    .C(_07609_),
    .Y(_07610_));
 sg13g2_inv_1 _16851_ (.Y(_07611_),
    .A(_07610_));
 sg13g2_nor3_2 _16852_ (.A(_06420_),
    .B(_06417_),
    .C(_07611_),
    .Y(_07612_));
 sg13g2_xnor2_1 _16853_ (.Y(_07613_),
    .A(_06414_),
    .B(_07612_));
 sg13g2_buf_2 _16854_ (.A(_07613_),
    .X(_07614_));
 sg13g2_xnor2_1 _16855_ (.Y(_07615_),
    .A(_07608_),
    .B(_07614_));
 sg13g2_nor2_1 _16856_ (.A(_07596_),
    .B(_07615_),
    .Y(_07616_));
 sg13g2_xnor2_1 _16857_ (.Y(_07617_),
    .A(_07596_),
    .B(_07615_));
 sg13g2_nor2_1 _16858_ (.A(_07579_),
    .B(_07617_),
    .Y(_07618_));
 sg13g2_nor2_1 _16859_ (.A(_07616_),
    .B(_07618_),
    .Y(_07619_));
 sg13g2_nor2b_1 _16860_ (.A(_07607_),
    .B_N(_07600_),
    .Y(_07620_));
 sg13g2_nor2_1 _16861_ (.A(_07608_),
    .B(_07614_),
    .Y(_07621_));
 sg13g2_nor2_1 _16862_ (.A(_07620_),
    .B(_07621_),
    .Y(_07622_));
 sg13g2_inv_1 _16863_ (.Y(_07623_),
    .A(_07606_));
 sg13g2_inv_1 _16864_ (.Y(_07624_),
    .A(_07601_));
 sg13g2_nor2_1 _16865_ (.A(_04820_),
    .B(_07624_),
    .Y(_07625_));
 sg13g2_a21oi_1 _16866_ (.A1(_07623_),
    .A2(_07602_),
    .Y(_07626_),
    .B1(_07625_));
 sg13g2_buf_1 _16867_ (.A(\vgadonut.donut.ycA[10] ),
    .X(_07627_));
 sg13g2_xnor2_1 _16868_ (.Y(_07628_),
    .A(_07627_),
    .B(_04815_));
 sg13g2_xnor2_1 _16869_ (.Y(_07629_),
    .A(_07569_),
    .B(_07575_));
 sg13g2_buf_2 _16870_ (.A(_07629_),
    .X(_07630_));
 sg13g2_xor2_1 _16871_ (.B(_07630_),
    .A(_07628_),
    .X(_07631_));
 sg13g2_xnor2_1 _16872_ (.Y(_07632_),
    .A(_07626_),
    .B(_07631_));
 sg13g2_inv_1 _16873_ (.Y(_07633_),
    .A(_07577_));
 sg13g2_nor3_1 _16874_ (.A(_06417_),
    .B(_06414_),
    .C(_07633_),
    .Y(_07634_));
 sg13g2_xnor2_1 _16875_ (.Y(_07635_),
    .A(_06428_),
    .B(_07634_));
 sg13g2_buf_2 _16876_ (.A(_07635_),
    .X(_07636_));
 sg13g2_xnor2_1 _16877_ (.Y(_07637_),
    .A(_07632_),
    .B(_07636_));
 sg13g2_xnor2_1 _16878_ (.Y(_07638_),
    .A(_07622_),
    .B(_07637_));
 sg13g2_xnor2_1 _16879_ (.Y(_07639_),
    .A(_07614_),
    .B(_07638_));
 sg13g2_xnor2_1 _16880_ (.Y(_07640_),
    .A(_07619_),
    .B(_07639_));
 sg13g2_xnor2_1 _16881_ (.Y(_07641_),
    .A(_07586_),
    .B(_07585_));
 sg13g2_buf_1 _16882_ (.A(\vgadonut.donut.ycA[6] ),
    .X(_07642_));
 sg13g2_inv_1 _16883_ (.Y(_07643_),
    .A(_07642_));
 sg13g2_xnor2_1 _16884_ (.Y(_07644_),
    .A(_07642_),
    .B(_04826_));
 sg13g2_nand2_1 _16885_ (.Y(_07645_),
    .A(_07644_),
    .B(_00121_));
 sg13g2_o21ai_1 _16886_ (.B1(_07645_),
    .Y(_07646_),
    .A1(_07643_),
    .A2(_04826_));
 sg13g2_xnor2_1 _16887_ (.Y(_07647_),
    .A(_07641_),
    .B(_07646_));
 sg13g2_xnor2_1 _16888_ (.Y(_07648_),
    .A(_06420_),
    .B(_07610_));
 sg13g2_buf_2 _16889_ (.A(_07648_),
    .X(_07649_));
 sg13g2_inv_1 _16890_ (.Y(_07650_),
    .A(_07649_));
 sg13g2_nor2b_1 _16891_ (.A(_07641_),
    .B_N(_07646_),
    .Y(_07651_));
 sg13g2_a21oi_1 _16892_ (.A1(_07647_),
    .A2(_07650_),
    .Y(_07652_),
    .B1(_07651_));
 sg13g2_xor2_1 _16893_ (.B(_07579_),
    .A(_07594_),
    .X(_07653_));
 sg13g2_nor2_1 _16894_ (.A(_07652_),
    .B(_07653_),
    .Y(_07654_));
 sg13g2_xnor2_1 _16895_ (.Y(_07655_),
    .A(_07652_),
    .B(_07653_));
 sg13g2_nor2_1 _16896_ (.A(_07649_),
    .B(_07655_),
    .Y(_07656_));
 sg13g2_nor2_1 _16897_ (.A(_07654_),
    .B(_07656_),
    .Y(_07657_));
 sg13g2_xnor2_1 _16898_ (.Y(_07658_),
    .A(_07579_),
    .B(_07617_));
 sg13g2_nor2_1 _16899_ (.A(_07657_),
    .B(_07658_),
    .Y(_07659_));
 sg13g2_inv_1 _16900_ (.Y(_07660_),
    .A(_07659_));
 sg13g2_nand2_1 _16901_ (.Y(_07661_),
    .A(_07658_),
    .B(_07657_));
 sg13g2_nand2_1 _16902_ (.Y(_07662_),
    .A(_07660_),
    .B(_07661_));
 sg13g2_buf_2 _16903_ (.A(\vgadonut.donut.ycA[4] ),
    .X(_07663_));
 sg13g2_inv_1 _16904_ (.Y(_07664_),
    .A(_07663_));
 sg13g2_xnor2_1 _16905_ (.Y(_07665_),
    .A(_07664_),
    .B(_07592_));
 sg13g2_inv_1 _16906_ (.Y(_07666_),
    .A(_00122_));
 sg13g2_a21oi_1 _16907_ (.A1(_07665_),
    .A2(_07666_),
    .Y(_07667_),
    .B1(_07585_));
 sg13g2_nand2_1 _16908_ (.Y(_07668_),
    .A(_07592_),
    .B(_07663_));
 sg13g2_buf_1 _16909_ (.A(\vgadonut.donut.ycA[5] ),
    .X(_07669_));
 sg13g2_inv_1 _16910_ (.Y(_07670_),
    .A(_07669_));
 sg13g2_xnor2_1 _16911_ (.Y(_07671_),
    .A(_07670_),
    .B(_07606_));
 sg13g2_xnor2_1 _16912_ (.Y(_07672_),
    .A(_07668_),
    .B(_07671_));
 sg13g2_nor2b_1 _16913_ (.A(_07667_),
    .B_N(_07672_),
    .Y(_07673_));
 sg13g2_inv_1 _16914_ (.Y(_07674_),
    .A(_07673_));
 sg13g2_a21oi_1 _16915_ (.A1(_07574_),
    .A2(_07583_),
    .Y(_07675_),
    .B1(_07666_));
 sg13g2_nor2_1 _16916_ (.A(_00122_),
    .B(_07585_),
    .Y(_07676_));
 sg13g2_o21ai_1 _16917_ (.B1(_07562_),
    .Y(_07677_),
    .A1(_07675_),
    .A2(_07676_));
 sg13g2_xnor2_1 _16918_ (.Y(_07678_),
    .A(_07676_),
    .B(_07665_));
 sg13g2_nand2b_1 _16919_ (.Y(_07679_),
    .B(_07678_),
    .A_N(_07677_));
 sg13g2_buf_2 _16920_ (.A(\vgadonut.donut.ycA[2] ),
    .X(_07680_));
 sg13g2_buf_1 _16921_ (.A(\vgadonut.donut.ycA[3] ),
    .X(_07681_));
 sg13g2_xnor2_1 _16922_ (.Y(_07682_),
    .A(_07572_),
    .B(_07681_));
 sg13g2_inv_1 _16923_ (.Y(_07683_),
    .A(_07682_));
 sg13g2_nor3_1 _16924_ (.A(_07564_),
    .B(_07680_),
    .C(_07683_),
    .Y(_07684_));
 sg13g2_inv_1 _16925_ (.Y(_07685_),
    .A(_07684_));
 sg13g2_nor2b_1 _16926_ (.A(_07678_),
    .B_N(_07677_),
    .Y(_07686_));
 sg13g2_a21oi_1 _16927_ (.A1(_07679_),
    .A2(_07685_),
    .Y(_07687_),
    .B1(_07686_));
 sg13g2_nor2b_1 _16928_ (.A(_07672_),
    .B_N(_07667_),
    .Y(_07688_));
 sg13g2_a21oi_1 _16929_ (.A1(_07674_),
    .A2(_07687_),
    .Y(_07689_),
    .B1(_07688_));
 sg13g2_nand2_1 _16930_ (.Y(_07690_),
    .A(_07606_),
    .B(_07669_));
 sg13g2_xnor2_1 _16931_ (.Y(_07691_),
    .A(_07603_),
    .B(_07644_));
 sg13g2_inv_1 _16932_ (.Y(_07692_),
    .A(_07691_));
 sg13g2_xnor2_1 _16933_ (.Y(_07693_),
    .A(_07692_),
    .B(_07630_));
 sg13g2_xnor2_1 _16934_ (.Y(_07694_),
    .A(_07690_),
    .B(_07693_));
 sg13g2_inv_1 _16935_ (.Y(_07695_),
    .A(_07694_));
 sg13g2_a21oi_1 _16936_ (.A1(_07671_),
    .A2(_07663_),
    .Y(_07696_),
    .B1(_07598_));
 sg13g2_nand2_1 _16937_ (.Y(_07697_),
    .A(_07695_),
    .B(_07696_));
 sg13g2_nor2_1 _16938_ (.A(_07696_),
    .B(_07695_),
    .Y(_07698_));
 sg13g2_a21oi_1 _16939_ (.A1(_07689_),
    .A2(_07697_),
    .Y(_07699_),
    .B1(_07698_));
 sg13g2_inv_1 _16940_ (.Y(_07700_),
    .A(_07699_));
 sg13g2_a21oi_1 _16941_ (.A1(_07693_),
    .A2(_07669_),
    .Y(_07701_),
    .B1(_07623_));
 sg13g2_nand2_1 _16942_ (.Y(_07702_),
    .A(_07630_),
    .B(_07691_));
 sg13g2_xor2_1 _16943_ (.B(_07647_),
    .A(_07649_),
    .X(_07703_));
 sg13g2_xnor2_1 _16944_ (.Y(_07704_),
    .A(_07702_),
    .B(_07703_));
 sg13g2_nor2_1 _16945_ (.A(_07701_),
    .B(_07704_),
    .Y(_07705_));
 sg13g2_inv_1 _16946_ (.Y(_07706_),
    .A(_07705_));
 sg13g2_nand2_1 _16947_ (.Y(_07707_),
    .A(_07704_),
    .B(_07701_));
 sg13g2_nand2_1 _16948_ (.Y(_07708_),
    .A(_07706_),
    .B(_07707_));
 sg13g2_xnor2_1 _16949_ (.Y(_07709_),
    .A(_07649_),
    .B(_07655_));
 sg13g2_o21ai_1 _16950_ (.B1(_07630_),
    .Y(_07710_),
    .A1(_07692_),
    .A2(_07703_));
 sg13g2_nor2b_1 _16951_ (.A(_07709_),
    .B_N(_07710_),
    .Y(_07711_));
 sg13g2_inv_1 _16952_ (.Y(_07712_),
    .A(_07711_));
 sg13g2_nand2b_1 _16953_ (.Y(_07713_),
    .B(_07709_),
    .A_N(_07710_));
 sg13g2_nand2_1 _16954_ (.Y(_07714_),
    .A(_07712_),
    .B(_07713_));
 sg13g2_nor2_1 _16955_ (.A(_07708_),
    .B(_07714_),
    .Y(_07715_));
 sg13g2_o21ai_1 _16956_ (.B1(_07712_),
    .Y(_07716_),
    .A1(_07706_),
    .A2(_07714_));
 sg13g2_a21oi_1 _16957_ (.A1(_07700_),
    .A2(_07715_),
    .Y(_07717_),
    .B1(_07716_));
 sg13g2_inv_1 _16958_ (.Y(_07718_),
    .A(_07717_));
 sg13g2_nand2b_1 _16959_ (.Y(_07719_),
    .B(_07718_),
    .A_N(_07662_));
 sg13g2_nand2_1 _16960_ (.Y(_07720_),
    .A(_07719_),
    .B(_07660_));
 sg13g2_xnor2_1 _16961_ (.Y(_07721_),
    .A(_07640_),
    .B(_07720_));
 sg13g2_inv_1 _16962_ (.Y(_07722_),
    .A(_06414_));
 sg13g2_inv_1 _16963_ (.Y(_07723_),
    .A(_06428_));
 sg13g2_nand3_1 _16964_ (.B(_07722_),
    .C(_07723_),
    .A(_07612_),
    .Y(_07724_));
 sg13g2_xnor2_1 _16965_ (.Y(_07725_),
    .A(_06434_),
    .B(_07724_));
 sg13g2_inv_2 _16966_ (.Y(_07726_),
    .A(_07725_));
 sg13g2_nor2_1 _16967_ (.A(\vgadonut.donut.donuthit.ryin[3] ),
    .B(_07726_),
    .Y(_07727_));
 sg13g2_nor2_1 _16968_ (.A(\vgadonut.donut.ry6[4] ),
    .B(_07630_),
    .Y(_07728_));
 sg13g2_inv_1 _16969_ (.Y(_07729_),
    .A(\vgadonut.donut.ry6[3] ));
 sg13g2_nor2_1 _16970_ (.A(_07729_),
    .B(_07623_),
    .Y(_07730_));
 sg13g2_nor2_1 _16971_ (.A(\vgadonut.donut.ry6[2] ),
    .B(_07592_),
    .Y(_07731_));
 sg13g2_xnor2_1 _16972_ (.Y(_07732_),
    .A(\vgadonut.donut.ry6[1] ),
    .B(_07585_));
 sg13g2_inv_1 _16973_ (.Y(_07733_),
    .A(_07563_));
 sg13g2_nor2b_1 _16974_ (.A(_07585_),
    .B_N(\vgadonut.donut.ry6[1] ),
    .Y(_07734_));
 sg13g2_a21oi_1 _16975_ (.A1(_07732_),
    .A2(_07733_),
    .Y(_07735_),
    .B1(_07734_));
 sg13g2_inv_1 _16976_ (.Y(_07736_),
    .A(\vgadonut.donut.ry6[2] ));
 sg13g2_nor2_1 _16977_ (.A(_07736_),
    .B(_07598_),
    .Y(_07737_));
 sg13g2_inv_1 _16978_ (.Y(_07738_),
    .A(_07737_));
 sg13g2_o21ai_1 _16979_ (.B1(_07738_),
    .Y(_07739_),
    .A1(_07731_),
    .A2(_07735_));
 sg13g2_nor2_1 _16980_ (.A(\vgadonut.donut.ry6[3] ),
    .B(_07606_),
    .Y(_07740_));
 sg13g2_inv_1 _16981_ (.Y(_07741_),
    .A(_07740_));
 sg13g2_o21ai_1 _16982_ (.B1(_07741_),
    .Y(_07742_),
    .A1(_07730_),
    .A2(_07739_));
 sg13g2_inv_1 _16983_ (.Y(_07743_),
    .A(\vgadonut.donut.ry6[4] ));
 sg13g2_inv_1 _16984_ (.Y(_07744_),
    .A(_07630_));
 sg13g2_nor2_1 _16985_ (.A(_07743_),
    .B(_07744_),
    .Y(_07745_));
 sg13g2_inv_1 _16986_ (.Y(_07746_),
    .A(_07745_));
 sg13g2_o21ai_1 _16987_ (.B1(_07746_),
    .Y(_07747_),
    .A1(_07728_),
    .A2(_07742_));
 sg13g2_nor2_1 _16988_ (.A(\vgadonut.donut.ry6[5] ),
    .B(_07649_),
    .Y(_07748_));
 sg13g2_inv_1 _16989_ (.Y(_07749_),
    .A(_07748_));
 sg13g2_inv_1 _16990_ (.Y(_07750_),
    .A(\vgadonut.donut.ry6[5] ));
 sg13g2_nor2_1 _16991_ (.A(_07750_),
    .B(_07650_),
    .Y(_07751_));
 sg13g2_a21oi_1 _16992_ (.A1(_07747_),
    .A2(_07749_),
    .Y(_07752_),
    .B1(_07751_));
 sg13g2_nor2_1 _16993_ (.A(\vgadonut.donut.donuthit.ryin[0] ),
    .B(_07579_),
    .Y(_07753_));
 sg13g2_inv_1 _16994_ (.Y(_07754_),
    .A(\vgadonut.donut.donuthit.ryin[0] ));
 sg13g2_nor2_1 _16995_ (.A(_07754_),
    .B(_07580_),
    .Y(_07755_));
 sg13g2_nor2_1 _16996_ (.A(_07753_),
    .B(_07755_),
    .Y(_07756_));
 sg13g2_nand2b_1 _16997_ (.Y(_07757_),
    .B(_07756_),
    .A_N(_07752_));
 sg13g2_inv_1 _16998_ (.Y(_07758_),
    .A(\vgadonut.donut.donuthit.ryin[1] ));
 sg13g2_inv_1 _16999_ (.Y(_07759_),
    .A(_07614_));
 sg13g2_nor2_1 _17000_ (.A(_07758_),
    .B(_07759_),
    .Y(_07760_));
 sg13g2_nor2_1 _17001_ (.A(_07755_),
    .B(_07760_),
    .Y(_07761_));
 sg13g2_nor2_1 _17002_ (.A(\vgadonut.donut.donuthit.ryin[1] ),
    .B(_07614_),
    .Y(_07762_));
 sg13g2_a21oi_1 _17003_ (.A1(_07757_),
    .A2(_07761_),
    .Y(_07763_),
    .B1(_07762_));
 sg13g2_nor2_1 _17004_ (.A(\vgadonut.donut.donuthit.ryin[2] ),
    .B(_07636_),
    .Y(_07764_));
 sg13g2_inv_1 _17005_ (.Y(_07765_),
    .A(\vgadonut.donut.donuthit.ryin[2] ));
 sg13g2_inv_1 _17006_ (.Y(_07766_),
    .A(_07636_));
 sg13g2_nor2_1 _17007_ (.A(_07765_),
    .B(_07766_),
    .Y(_07767_));
 sg13g2_nor2_1 _17008_ (.A(_07764_),
    .B(_07767_),
    .Y(_07768_));
 sg13g2_a221oi_1 _17009_ (.B2(_07768_),
    .C1(_07767_),
    .B1(_07763_),
    .A1(\vgadonut.donut.donuthit.ryin[3] ),
    .Y(_07769_),
    .A2(_07726_));
 sg13g2_nor2_1 _17010_ (.A(_07727_),
    .B(_07769_),
    .Y(_07770_));
 sg13g2_nand3_1 _17011_ (.B(_07723_),
    .C(_06435_),
    .A(_07634_),
    .Y(_07771_));
 sg13g2_buf_1 _17012_ (.A(_07771_),
    .X(_07772_));
 sg13g2_xnor2_1 _17013_ (.Y(_07773_),
    .A(_06443_),
    .B(_07772_));
 sg13g2_buf_2 _17014_ (.A(_07773_),
    .X(_07774_));
 sg13g2_nor2_1 _17015_ (.A(\vgadonut.donut.donuthit.ryin[4] ),
    .B(_07774_),
    .Y(_07775_));
 sg13g2_inv_1 _17016_ (.Y(_07776_),
    .A(_07774_));
 sg13g2_nor2b_1 _17017_ (.A(_07776_),
    .B_N(\vgadonut.donut.donuthit.ryin[4] ),
    .Y(_07777_));
 sg13g2_nor2_1 _17018_ (.A(_07775_),
    .B(_07777_),
    .Y(_07778_));
 sg13g2_nand2_1 _17019_ (.Y(_07779_),
    .A(_07770_),
    .B(_07778_));
 sg13g2_nor2_1 _17020_ (.A(_07778_),
    .B(_07770_),
    .Y(_07780_));
 sg13g2_nor2_1 _17021_ (.A(net148),
    .B(_07780_),
    .Y(_07781_));
 sg13g2_a22oi_1 _17022_ (.Y(_07782_),
    .B1(_07779_),
    .B2(_07781_),
    .A2(_07721_),
    .A1(_07533_));
 sg13g2_nand2_1 _17023_ (.Y(_07783_),
    .A(net98),
    .B(\vgadonut.donut.donuthit.ryin[4] ));
 sg13g2_o21ai_1 _17024_ (.B1(_07783_),
    .Y(_00370_),
    .A1(net91),
    .A2(_07782_));
 sg13g2_nor2_1 _17025_ (.A(_07626_),
    .B(_07631_),
    .Y(_07784_));
 sg13g2_nor2_1 _17026_ (.A(_07632_),
    .B(_07636_),
    .Y(_07785_));
 sg13g2_nor2_1 _17027_ (.A(_07784_),
    .B(_07785_),
    .Y(_07786_));
 sg13g2_inv_1 _17028_ (.Y(_07787_),
    .A(_07627_));
 sg13g2_nand2_1 _17029_ (.Y(_07788_),
    .A(_07744_),
    .B(_07628_));
 sg13g2_o21ai_1 _17030_ (.B1(_07788_),
    .Y(_07789_),
    .A1(_07787_),
    .A2(_04815_));
 sg13g2_buf_1 _17031_ (.A(\vgadonut.donut.ycA[11] ),
    .X(_07790_));
 sg13g2_xnor2_1 _17032_ (.Y(_07791_),
    .A(_07790_),
    .B(net243));
 sg13g2_xor2_1 _17033_ (.B(_07649_),
    .A(_07791_),
    .X(_07792_));
 sg13g2_xor2_1 _17034_ (.B(_07792_),
    .A(_07789_),
    .X(_07793_));
 sg13g2_xnor2_1 _17035_ (.Y(_07794_),
    .A(_07726_),
    .B(_07793_));
 sg13g2_xnor2_1 _17036_ (.Y(_07795_),
    .A(_07786_),
    .B(_07794_));
 sg13g2_xnor2_1 _17037_ (.Y(_07796_),
    .A(_07636_),
    .B(_07795_));
 sg13g2_nor2_1 _17038_ (.A(_07622_),
    .B(_07637_),
    .Y(_07797_));
 sg13g2_nor2_1 _17039_ (.A(_07614_),
    .B(_07638_),
    .Y(_07798_));
 sg13g2_nor2_1 _17040_ (.A(_07797_),
    .B(_07798_),
    .Y(_07799_));
 sg13g2_xnor2_1 _17041_ (.Y(_07800_),
    .A(_07796_),
    .B(_07799_));
 sg13g2_nor2_1 _17042_ (.A(_07662_),
    .B(_07640_),
    .Y(_07801_));
 sg13g2_nor2_1 _17043_ (.A(_07619_),
    .B(_07639_),
    .Y(_07802_));
 sg13g2_inv_1 _17044_ (.Y(_07803_),
    .A(_07802_));
 sg13g2_o21ai_1 _17045_ (.B1(_07803_),
    .Y(_07804_),
    .A1(_07660_),
    .A2(_07640_));
 sg13g2_a21oi_1 _17046_ (.A1(_07718_),
    .A2(_07801_),
    .Y(_07805_),
    .B1(_07804_));
 sg13g2_a21oi_1 _17047_ (.A1(_07805_),
    .A2(_07800_),
    .Y(_07806_),
    .B1(net146));
 sg13g2_o21ai_1 _17048_ (.B1(_07806_),
    .Y(_07807_),
    .A1(_07800_),
    .A2(_07805_));
 sg13g2_nor2_1 _17049_ (.A(_06434_),
    .B(_06442_),
    .Y(_07808_));
 sg13g2_nor2b_1 _17050_ (.A(_07724_),
    .B_N(_07808_),
    .Y(_07809_));
 sg13g2_xnor2_1 _17051_ (.Y(_07810_),
    .A(_06406_),
    .B(_07809_));
 sg13g2_buf_2 _17052_ (.A(_07810_),
    .X(_07811_));
 sg13g2_xnor2_1 _17053_ (.Y(_07812_),
    .A(_04839_),
    .B(_07811_));
 sg13g2_nand2b_1 _17054_ (.Y(_07813_),
    .B(_07779_),
    .A_N(_07777_));
 sg13g2_xor2_1 _17055_ (.B(_07813_),
    .A(_07812_),
    .X(_07814_));
 sg13g2_a21oi_1 _17056_ (.A1(_07814_),
    .A2(net165),
    .Y(_07815_),
    .B1(net98));
 sg13g2_a22oi_1 _17057_ (.Y(_00371_),
    .B1(_07807_),
    .B2(_07815_),
    .A2(net92),
    .A1(_04839_));
 sg13g2_nor2_1 _17058_ (.A(_07786_),
    .B(_07794_),
    .Y(_07816_));
 sg13g2_nor2_1 _17059_ (.A(_07636_),
    .B(_07795_),
    .Y(_07817_));
 sg13g2_nor2_1 _17060_ (.A(_07816_),
    .B(_07817_),
    .Y(_07818_));
 sg13g2_nor2b_1 _17061_ (.A(_07792_),
    .B_N(_07789_),
    .Y(_07819_));
 sg13g2_nor2_1 _17062_ (.A(_07726_),
    .B(_07793_),
    .Y(_07820_));
 sg13g2_nor2_1 _17063_ (.A(_07819_),
    .B(_07820_),
    .Y(_07821_));
 sg13g2_inv_1 _17064_ (.Y(_07822_),
    .A(_07790_));
 sg13g2_nor2_1 _17065_ (.A(net243),
    .B(_07822_),
    .Y(_07823_));
 sg13g2_a21oi_1 _17066_ (.A1(_07650_),
    .A2(_07791_),
    .Y(_07824_),
    .B1(_07823_));
 sg13g2_buf_1 _17067_ (.A(\vgadonut.donut.ycA[12] ),
    .X(_07825_));
 sg13g2_xnor2_1 _17068_ (.Y(_07826_),
    .A(_07825_),
    .B(_04816_));
 sg13g2_inv_1 _17069_ (.Y(_07827_),
    .A(_07826_));
 sg13g2_xnor2_1 _17070_ (.Y(_07828_),
    .A(_07827_),
    .B(_07579_));
 sg13g2_xnor2_1 _17071_ (.Y(_07829_),
    .A(_07824_),
    .B(_07828_));
 sg13g2_xnor2_1 _17072_ (.Y(_07830_),
    .A(_07774_),
    .B(_07829_));
 sg13g2_xnor2_1 _17073_ (.Y(_07831_),
    .A(_07821_),
    .B(_07830_));
 sg13g2_xnor2_1 _17074_ (.Y(_07832_),
    .A(_07726_),
    .B(_07831_));
 sg13g2_nor2_1 _17075_ (.A(_07818_),
    .B(_07832_),
    .Y(_07833_));
 sg13g2_inv_1 _17076_ (.Y(_07834_),
    .A(_07833_));
 sg13g2_nand2_1 _17077_ (.Y(_07835_),
    .A(_07832_),
    .B(_07818_));
 sg13g2_nand2_1 _17078_ (.Y(_07836_),
    .A(_07834_),
    .B(_07835_));
 sg13g2_nor2_1 _17079_ (.A(_07799_),
    .B(_07796_),
    .Y(_07837_));
 sg13g2_nor2_1 _17080_ (.A(_07802_),
    .B(_07837_),
    .Y(_07838_));
 sg13g2_nand2b_1 _17081_ (.Y(_07839_),
    .B(_07720_),
    .A_N(_07640_));
 sg13g2_a22oi_1 _17082_ (.Y(_07840_),
    .B1(_07838_),
    .B2(_07839_),
    .A2(_07796_),
    .A1(_07799_));
 sg13g2_xnor2_1 _17083_ (.Y(_07841_),
    .A(_07836_),
    .B(_07840_));
 sg13g2_nand3b_1 _17084_ (.B(_06443_),
    .C(_06407_),
    .Y(_07842_),
    .A_N(_07772_));
 sg13g2_xnor2_1 _17085_ (.Y(_07843_),
    .A(_06529_),
    .B(_07842_));
 sg13g2_buf_2 _17086_ (.A(_07843_),
    .X(_07844_));
 sg13g2_xnor2_1 _17087_ (.Y(_07845_),
    .A(_06944_),
    .B(_07844_));
 sg13g2_inv_1 _17088_ (.Y(_07846_),
    .A(_07845_));
 sg13g2_inv_1 _17089_ (.Y(_07847_),
    .A(_00123_));
 sg13g2_a22oi_1 _17090_ (.Y(_07848_),
    .B1(_07812_),
    .B2(_07813_),
    .A2(_07811_),
    .A1(_07847_));
 sg13g2_nor2_1 _17091_ (.A(_07846_),
    .B(_07848_),
    .Y(_07849_));
 sg13g2_inv_1 _17092_ (.Y(_07850_),
    .A(_07849_));
 sg13g2_a21oi_1 _17093_ (.A1(_07848_),
    .A2(_07846_),
    .Y(_07851_),
    .B1(_10117_));
 sg13g2_a22oi_1 _17094_ (.Y(_07852_),
    .B1(_07850_),
    .B2(_07851_),
    .A2(_07841_),
    .A1(_07533_));
 sg13g2_nand2_1 _17095_ (.Y(_07853_),
    .A(net98),
    .B(\vgadonut.donut.donuthit.ryin[6] ));
 sg13g2_o21ai_1 _17096_ (.B1(_07853_),
    .Y(_00372_),
    .A1(net91),
    .A2(_07852_));
 sg13g2_nor2_1 _17097_ (.A(_07824_),
    .B(_07828_),
    .Y(_07854_));
 sg13g2_nor2_1 _17098_ (.A(_07774_),
    .B(_07829_),
    .Y(_07855_));
 sg13g2_nor2_1 _17099_ (.A(_07854_),
    .B(_07855_),
    .Y(_07856_));
 sg13g2_inv_1 _17100_ (.Y(_07857_),
    .A(_07825_));
 sg13g2_nor2_1 _17101_ (.A(net244),
    .B(_07857_),
    .Y(_07858_));
 sg13g2_a21oi_1 _17102_ (.A1(_07580_),
    .A2(_07826_),
    .Y(_07859_),
    .B1(_07858_));
 sg13g2_buf_1 _17103_ (.A(\vgadonut.donut.ycA[13] ),
    .X(_07860_));
 sg13g2_xnor2_1 _17104_ (.Y(_07861_),
    .A(_07860_),
    .B(_04842_));
 sg13g2_xor2_1 _17105_ (.B(_07614_),
    .A(_07861_),
    .X(_07862_));
 sg13g2_xnor2_1 _17106_ (.Y(_07863_),
    .A(_07859_),
    .B(_07862_));
 sg13g2_xnor2_1 _17107_ (.Y(_07864_),
    .A(_07811_),
    .B(_07863_));
 sg13g2_xnor2_1 _17108_ (.Y(_07865_),
    .A(_07856_),
    .B(_07864_));
 sg13g2_xnor2_1 _17109_ (.Y(_07866_),
    .A(_07774_),
    .B(_07865_));
 sg13g2_nor2_1 _17110_ (.A(_07821_),
    .B(_07830_),
    .Y(_07867_));
 sg13g2_nor2_1 _17111_ (.A(_07726_),
    .B(_07831_),
    .Y(_07868_));
 sg13g2_nor2_1 _17112_ (.A(_07867_),
    .B(_07868_),
    .Y(_07869_));
 sg13g2_xnor2_1 _17113_ (.Y(_07870_),
    .A(_07866_),
    .B(_07869_));
 sg13g2_nor2_1 _17114_ (.A(_07837_),
    .B(_07833_),
    .Y(_07871_));
 sg13g2_o21ai_1 _17115_ (.B1(_07871_),
    .Y(_07872_),
    .A1(_07800_),
    .A2(_07805_));
 sg13g2_nand2_1 _17116_ (.Y(_07873_),
    .A(_07872_),
    .B(_07835_));
 sg13g2_a21oi_1 _17117_ (.A1(_07873_),
    .A2(_07870_),
    .Y(_07874_),
    .B1(net146));
 sg13g2_o21ai_1 _17118_ (.B1(_07874_),
    .Y(_07875_),
    .A1(_07870_),
    .A2(_07873_));
 sg13g2_nand3_1 _17119_ (.B(_06407_),
    .C(_06529_),
    .A(_07809_),
    .Y(_07876_));
 sg13g2_xnor2_1 _17120_ (.Y(_07877_),
    .A(_06533_),
    .B(_07876_));
 sg13g2_buf_2 _17121_ (.A(_07877_),
    .X(_07878_));
 sg13g2_xnor2_1 _17122_ (.Y(_07879_),
    .A(\vgadonut.donut.donuthit.ryin[7] ),
    .B(_07878_));
 sg13g2_inv_1 _17123_ (.Y(_07880_),
    .A(_07844_));
 sg13g2_nor2_1 _17124_ (.A(_00124_),
    .B(_07880_),
    .Y(_07881_));
 sg13g2_nor2_1 _17125_ (.A(_07881_),
    .B(_07849_),
    .Y(_07882_));
 sg13g2_xnor2_1 _17126_ (.Y(_07883_),
    .A(_07879_),
    .B(_07882_));
 sg13g2_a21oi_1 _17127_ (.A1(_07883_),
    .A2(net165),
    .Y(_07884_),
    .B1(net98));
 sg13g2_a22oi_1 _17128_ (.Y(_00373_),
    .B1(_07875_),
    .B2(_07884_),
    .A2(net92),
    .A1(_06947_));
 sg13g2_buf_1 _17129_ (.A(net100),
    .X(_07885_));
 sg13g2_nor2_1 _17130_ (.A(_07856_),
    .B(_07864_),
    .Y(_07886_));
 sg13g2_nor2_1 _17131_ (.A(_07774_),
    .B(_07865_),
    .Y(_07887_));
 sg13g2_nor2_1 _17132_ (.A(_07886_),
    .B(_07887_),
    .Y(_07888_));
 sg13g2_nor2_1 _17133_ (.A(_07859_),
    .B(_07862_),
    .Y(_07889_));
 sg13g2_nor2_1 _17134_ (.A(_07811_),
    .B(_07863_),
    .Y(_07890_));
 sg13g2_nor2_1 _17135_ (.A(_07889_),
    .B(_07890_),
    .Y(_07891_));
 sg13g2_inv_1 _17136_ (.Y(_07892_),
    .A(_07860_));
 sg13g2_nand2_1 _17137_ (.Y(_07893_),
    .A(_07759_),
    .B(_07861_));
 sg13g2_o21ai_1 _17138_ (.B1(_07893_),
    .Y(_07894_),
    .A1(_07892_),
    .A2(_04842_));
 sg13g2_buf_2 _17139_ (.A(\vgadonut.donut.ycA[14] ),
    .X(_07895_));
 sg13g2_xnor2_1 _17140_ (.Y(_07896_),
    .A(_07895_),
    .B(_04944_));
 sg13g2_xor2_1 _17141_ (.B(_07636_),
    .A(_07896_),
    .X(_07897_));
 sg13g2_xor2_1 _17142_ (.B(_07897_),
    .A(_07894_),
    .X(_07898_));
 sg13g2_xnor2_1 _17143_ (.Y(_07899_),
    .A(_07844_),
    .B(_07898_));
 sg13g2_xnor2_1 _17144_ (.Y(_07900_),
    .A(_07891_),
    .B(_07899_));
 sg13g2_xnor2_1 _17145_ (.Y(_07901_),
    .A(_07811_),
    .B(_07900_));
 sg13g2_xnor2_1 _17146_ (.Y(_07902_),
    .A(_07888_),
    .B(_07901_));
 sg13g2_nor2_1 _17147_ (.A(_07836_),
    .B(_07870_),
    .Y(_07903_));
 sg13g2_nand2b_1 _17148_ (.Y(_07904_),
    .B(_07833_),
    .A_N(_07870_));
 sg13g2_o21ai_1 _17149_ (.B1(_07904_),
    .Y(_07905_),
    .A1(_07869_),
    .A2(_07866_));
 sg13g2_a21oi_1 _17150_ (.A1(_07840_),
    .A2(_07903_),
    .Y(_07906_),
    .B1(_07905_));
 sg13g2_nor2_1 _17151_ (.A(_07902_),
    .B(_07906_),
    .Y(_07907_));
 sg13g2_nand2_1 _17152_ (.Y(_07908_),
    .A(_07906_),
    .B(_07902_));
 sg13g2_nand3b_1 _17153_ (.B(net150),
    .C(_07908_),
    .Y(_07909_),
    .A_N(_07907_));
 sg13g2_inv_1 _17154_ (.Y(_07910_),
    .A(_07882_));
 sg13g2_nor2_1 _17155_ (.A(_00125_),
    .B(_07878_),
    .Y(_07911_));
 sg13g2_a21oi_1 _17156_ (.A1(_07910_),
    .A2(_07879_),
    .Y(_07912_),
    .B1(_07911_));
 sg13g2_nor2_1 _17157_ (.A(_06406_),
    .B(_06525_),
    .Y(_07913_));
 sg13g2_nand3_1 _17158_ (.B(_06443_),
    .C(_06538_),
    .A(_07913_),
    .Y(_07914_));
 sg13g2_nor2_1 _17159_ (.A(_07914_),
    .B(_07772_),
    .Y(_07915_));
 sg13g2_xnor2_1 _17160_ (.Y(_07916_),
    .A(_06541_),
    .B(_07915_));
 sg13g2_buf_2 _17161_ (.A(_07916_),
    .X(_07917_));
 sg13g2_xnor2_1 _17162_ (.Y(_07918_),
    .A(_04957_),
    .B(_07917_));
 sg13g2_a21oi_1 _17163_ (.A1(_07912_),
    .A2(_07918_),
    .Y(_07919_),
    .B1(net148));
 sg13g2_or2_1 _17164_ (.X(_07920_),
    .B(_07912_),
    .A(_07918_));
 sg13g2_a21oi_1 _17165_ (.A1(_07919_),
    .A2(_07920_),
    .Y(_07921_),
    .B1(net98));
 sg13g2_a22oi_1 _17166_ (.Y(_00374_),
    .B1(_07909_),
    .B2(_07921_),
    .A2(net90),
    .A1(_04957_));
 sg13g2_nor2_1 _17167_ (.A(_07891_),
    .B(_07899_),
    .Y(_07922_));
 sg13g2_nor2_1 _17168_ (.A(_07811_),
    .B(_07900_),
    .Y(_07923_));
 sg13g2_nor2_1 _17169_ (.A(_07922_),
    .B(_07923_),
    .Y(_07924_));
 sg13g2_nor2b_1 _17170_ (.A(_07897_),
    .B_N(_07894_),
    .Y(_07925_));
 sg13g2_nor2_1 _17171_ (.A(_07844_),
    .B(_07898_),
    .Y(_07926_));
 sg13g2_nor2_1 _17172_ (.A(_07925_),
    .B(_07926_),
    .Y(_07927_));
 sg13g2_buf_2 _17173_ (.A(\vgadonut.donut.ycA[15] ),
    .X(_07928_));
 sg13g2_xnor2_1 _17174_ (.Y(_07929_),
    .A(_07928_),
    .B(_04959_));
 sg13g2_xnor2_1 _17175_ (.Y(_07930_),
    .A(_07929_),
    .B(_07725_));
 sg13g2_inv_1 _17176_ (.Y(_07931_),
    .A(_07895_));
 sg13g2_nand2_1 _17177_ (.Y(_07932_),
    .A(_07766_),
    .B(_07896_));
 sg13g2_o21ai_1 _17178_ (.B1(_07932_),
    .Y(_07933_),
    .A1(_07931_),
    .A2(_04944_));
 sg13g2_xor2_1 _17179_ (.B(_07933_),
    .A(_07930_),
    .X(_07934_));
 sg13g2_xor2_1 _17180_ (.B(_07934_),
    .A(_07878_),
    .X(_07935_));
 sg13g2_xnor2_1 _17181_ (.Y(_07936_),
    .A(_07927_),
    .B(_07935_));
 sg13g2_xnor2_1 _17182_ (.Y(_07937_),
    .A(_07844_),
    .B(_07936_));
 sg13g2_nor2_1 _17183_ (.A(_07924_),
    .B(_07937_),
    .Y(_07938_));
 sg13g2_inv_1 _17184_ (.Y(_07939_),
    .A(_07938_));
 sg13g2_nand2_1 _17185_ (.Y(_07940_),
    .A(_07937_),
    .B(_07924_));
 sg13g2_nand2_1 _17186_ (.Y(_07941_),
    .A(_07939_),
    .B(_07940_));
 sg13g2_nor2_1 _17187_ (.A(_07888_),
    .B(_07901_),
    .Y(_07942_));
 sg13g2_nor2_1 _17188_ (.A(_07942_),
    .B(_07907_),
    .Y(_07943_));
 sg13g2_a21oi_1 _17189_ (.A1(_07943_),
    .A2(_07941_),
    .Y(_07944_),
    .B1(net146));
 sg13g2_o21ai_1 _17190_ (.B1(_07944_),
    .Y(_07945_),
    .A1(_07941_),
    .A2(_07943_));
 sg13g2_nor2_1 _17191_ (.A(_06414_),
    .B(_06428_),
    .Y(_07946_));
 sg13g2_nor4_1 _17192_ (.A(_06406_),
    .B(_06525_),
    .C(_06533_),
    .D(_06518_),
    .Y(_07947_));
 sg13g2_nand4_1 _17193_ (.B(_07946_),
    .C(_07808_),
    .A(_07612_),
    .Y(_07948_),
    .D(_07947_));
 sg13g2_nand2b_1 _17194_ (.Y(_07949_),
    .B(_06517_),
    .A_N(_07948_));
 sg13g2_nand2_1 _17195_ (.Y(_07950_),
    .A(_07948_),
    .B(net191));
 sg13g2_nand2_1 _17196_ (.Y(_07951_),
    .A(_07949_),
    .B(_07950_));
 sg13g2_buf_2 _17197_ (.A(_07951_),
    .X(_07952_));
 sg13g2_xnor2_1 _17198_ (.Y(_07953_),
    .A(\vgadonut.donut.donuthit.ryin[9] ),
    .B(_07952_));
 sg13g2_o21ai_1 _17199_ (.B1(_07920_),
    .Y(_07954_),
    .A1(_00126_),
    .A2(_07917_));
 sg13g2_xor2_1 _17200_ (.B(_07954_),
    .A(_07953_),
    .X(_07955_));
 sg13g2_buf_1 _17201_ (.A(_06989_),
    .X(_07956_));
 sg13g2_a21oi_1 _17202_ (.A1(_07955_),
    .A2(net165),
    .Y(_07957_),
    .B1(net96));
 sg13g2_a22oi_1 _17203_ (.Y(_00375_),
    .B1(_07945_),
    .B2(_07957_),
    .A2(net90),
    .A1(_06950_));
 sg13g2_nor2b_1 _17204_ (.A(_07930_),
    .B_N(_07933_),
    .Y(_07958_));
 sg13g2_nor2b_1 _17205_ (.A(_07934_),
    .B_N(_07878_),
    .Y(_07959_));
 sg13g2_nor2_1 _17206_ (.A(_07958_),
    .B(_07959_),
    .Y(_07960_));
 sg13g2_inv_1 _17207_ (.Y(_07961_),
    .A(_07928_));
 sg13g2_nor2_1 _17208_ (.A(_04959_),
    .B(_07961_),
    .Y(_07962_));
 sg13g2_a21oi_1 _17209_ (.A1(_07725_),
    .A2(_07929_),
    .Y(_07963_),
    .B1(_07962_));
 sg13g2_buf_2 _17210_ (.A(\vgadonut.donut.ycA[16] ),
    .X(_07964_));
 sg13g2_xnor2_1 _17211_ (.Y(_07965_),
    .A(_07964_),
    .B(_04990_));
 sg13g2_inv_1 _17212_ (.Y(_07966_),
    .A(_07965_));
 sg13g2_xnor2_1 _17213_ (.Y(_07967_),
    .A(_07966_),
    .B(_07774_));
 sg13g2_nor2_1 _17214_ (.A(_07963_),
    .B(_07967_),
    .Y(_07968_));
 sg13g2_nand2_1 _17215_ (.Y(_07969_),
    .A(_07967_),
    .B(_07963_));
 sg13g2_nor2b_1 _17216_ (.A(_07968_),
    .B_N(_07969_),
    .Y(_07970_));
 sg13g2_xnor2_1 _17217_ (.Y(_07971_),
    .A(_07917_),
    .B(_07970_));
 sg13g2_xnor2_1 _17218_ (.Y(_07972_),
    .A(_07960_),
    .B(_07971_));
 sg13g2_xor2_1 _17219_ (.B(_07972_),
    .A(_07878_),
    .X(_07973_));
 sg13g2_nor2_1 _17220_ (.A(_07927_),
    .B(_07935_),
    .Y(_07974_));
 sg13g2_nor2_1 _17221_ (.A(_07844_),
    .B(_07936_),
    .Y(_07975_));
 sg13g2_nor2_1 _17222_ (.A(_07974_),
    .B(_07975_),
    .Y(_07976_));
 sg13g2_xnor2_1 _17223_ (.Y(_07977_),
    .A(_07973_),
    .B(_07976_));
 sg13g2_inv_1 _17224_ (.Y(_07978_),
    .A(_07943_));
 sg13g2_a21oi_1 _17225_ (.A1(_07978_),
    .A2(_07940_),
    .Y(_07979_),
    .B1(_07938_));
 sg13g2_nor2_1 _17226_ (.A(_07977_),
    .B(_07979_),
    .Y(_07980_));
 sg13g2_nand2_1 _17227_ (.Y(_07981_),
    .A(_07979_),
    .B(_07977_));
 sg13g2_nand3b_1 _17228_ (.B(net150),
    .C(_07981_),
    .Y(_07982_),
    .A_N(_07980_));
 sg13g2_xnor2_1 _17229_ (.Y(_07983_),
    .A(_06934_),
    .B(_07952_));
 sg13g2_inv_1 _17230_ (.Y(_07984_),
    .A(_07983_));
 sg13g2_nor2_1 _17231_ (.A(_00127_),
    .B(_07952_),
    .Y(_07985_));
 sg13g2_nand2_1 _17232_ (.Y(_07986_),
    .A(_07954_),
    .B(_07953_));
 sg13g2_nand2b_1 _17233_ (.Y(_07987_),
    .B(_07986_),
    .A_N(_07985_));
 sg13g2_nor2_1 _17234_ (.A(_07984_),
    .B(_07987_),
    .Y(_07988_));
 sg13g2_nor2_1 _17235_ (.A(net148),
    .B(_07988_),
    .Y(_07989_));
 sg13g2_nand2_1 _17236_ (.Y(_07990_),
    .A(_07987_),
    .B(_07984_));
 sg13g2_a21oi_1 _17237_ (.A1(_07989_),
    .A2(_07990_),
    .Y(_07991_),
    .B1(net96));
 sg13g2_a22oi_1 _17238_ (.Y(_00376_),
    .B1(_07982_),
    .B2(_07991_),
    .A2(net90),
    .A1(_06934_));
 sg13g2_nand2_1 _17239_ (.Y(_07992_),
    .A(_07971_),
    .B(_07960_));
 sg13g2_nor2_1 _17240_ (.A(_07960_),
    .B(_07971_),
    .Y(_07993_));
 sg13g2_a21oi_1 _17241_ (.A1(_07992_),
    .A2(_07878_),
    .Y(_07994_),
    .B1(_07993_));
 sg13g2_a21oi_2 _17242_ (.B1(_07968_),
    .Y(_07995_),
    .A2(_07917_),
    .A1(_07969_));
 sg13g2_inv_2 _17243_ (.Y(_07996_),
    .A(_07952_));
 sg13g2_buf_2 _17244_ (.A(\vgadonut.donut.ycA[17] ),
    .X(_07997_));
 sg13g2_xnor2_1 _17245_ (.Y(_07998_),
    .A(_07997_),
    .B(_05025_));
 sg13g2_inv_1 _17246_ (.Y(_07999_),
    .A(_07998_));
 sg13g2_xnor2_1 _17247_ (.Y(_08000_),
    .A(_07999_),
    .B(_07811_));
 sg13g2_inv_1 _17248_ (.Y(_08001_),
    .A(_07964_));
 sg13g2_nor2_1 _17249_ (.A(_04990_),
    .B(_08001_),
    .Y(_08002_));
 sg13g2_a21oi_1 _17250_ (.A1(_07776_),
    .A2(_07965_),
    .Y(_08003_),
    .B1(_08002_));
 sg13g2_xnor2_1 _17251_ (.Y(_08004_),
    .A(_08000_),
    .B(_08003_));
 sg13g2_xnor2_1 _17252_ (.Y(_08005_),
    .A(_07996_),
    .B(_08004_));
 sg13g2_xnor2_1 _17253_ (.Y(_08006_),
    .A(_07995_),
    .B(_08005_));
 sg13g2_xor2_1 _17254_ (.B(_08006_),
    .A(_07917_),
    .X(_08007_));
 sg13g2_nor2_1 _17255_ (.A(_07994_),
    .B(_08007_),
    .Y(_08008_));
 sg13g2_inv_1 _17256_ (.Y(_08009_),
    .A(_08008_));
 sg13g2_nand2_1 _17257_ (.Y(_08010_),
    .A(_08007_),
    .B(_07994_));
 sg13g2_nand2_1 _17258_ (.Y(_08011_),
    .A(_08009_),
    .B(_08010_));
 sg13g2_nor2_1 _17259_ (.A(_07941_),
    .B(_07977_),
    .Y(_08012_));
 sg13g2_nor2_1 _17260_ (.A(_07976_),
    .B(_07973_),
    .Y(_08013_));
 sg13g2_inv_1 _17261_ (.Y(_08014_),
    .A(_08013_));
 sg13g2_o21ai_1 _17262_ (.B1(_08014_),
    .Y(_08015_),
    .A1(_07939_),
    .A2(_07977_));
 sg13g2_a21oi_1 _17263_ (.A1(_07978_),
    .A2(_08012_),
    .Y(_08016_),
    .B1(_08015_));
 sg13g2_a21oi_1 _17264_ (.A1(_08016_),
    .A2(_08011_),
    .Y(_08017_),
    .B1(net146));
 sg13g2_o21ai_1 _17265_ (.B1(_08017_),
    .Y(_08018_),
    .A1(_08011_),
    .A2(_08016_));
 sg13g2_xnor2_1 _17266_ (.Y(_08019_),
    .A(_06936_),
    .B(_07952_));
 sg13g2_nor2_1 _17267_ (.A(_00128_),
    .B(_07952_),
    .Y(_08020_));
 sg13g2_a21oi_1 _17268_ (.A1(_07985_),
    .A2(_06934_),
    .Y(_08021_),
    .B1(_08020_));
 sg13g2_o21ai_1 _17269_ (.B1(_08021_),
    .Y(_08022_),
    .A1(_07983_),
    .A2(_07986_));
 sg13g2_xnor2_1 _17270_ (.Y(_08023_),
    .A(_08019_),
    .B(_08022_));
 sg13g2_a21oi_1 _17271_ (.A1(_08023_),
    .A2(net165),
    .Y(_08024_),
    .B1(net96));
 sg13g2_a22oi_1 _17272_ (.Y(_00377_),
    .B1(_08018_),
    .B2(_08024_),
    .A2(net90),
    .A1(_06936_));
 sg13g2_nor2_1 _17273_ (.A(_08000_),
    .B(_08003_),
    .Y(_08025_));
 sg13g2_nor2_1 _17274_ (.A(_07996_),
    .B(_08004_),
    .Y(_08026_));
 sg13g2_nor2_1 _17275_ (.A(_08025_),
    .B(_08026_),
    .Y(_08027_));
 sg13g2_nor2_1 _17276_ (.A(_07999_),
    .B(_07811_),
    .Y(_08028_));
 sg13g2_a21oi_1 _17277_ (.A1(_07997_),
    .A2(_06485_),
    .Y(_08029_),
    .B1(_08028_));
 sg13g2_buf_1 _17278_ (.A(\vgadonut.donut.ycA[18] ),
    .X(_08030_));
 sg13g2_xnor2_1 _17279_ (.Y(_08031_),
    .A(_08030_),
    .B(_05062_));
 sg13g2_inv_1 _17280_ (.Y(_08032_),
    .A(_08031_));
 sg13g2_xnor2_1 _17281_ (.Y(_08033_),
    .A(_08032_),
    .B(_07844_));
 sg13g2_nor2_1 _17282_ (.A(_08029_),
    .B(_08033_),
    .Y(_08034_));
 sg13g2_inv_1 _17283_ (.Y(_08035_),
    .A(_08034_));
 sg13g2_nand2_1 _17284_ (.Y(_08036_),
    .A(_08033_),
    .B(_08029_));
 sg13g2_nand2_1 _17285_ (.Y(_08037_),
    .A(_08035_),
    .B(_08036_));
 sg13g2_xnor2_1 _17286_ (.Y(_08038_),
    .A(_08027_),
    .B(_08037_));
 sg13g2_nand2_1 _17287_ (.Y(_08039_),
    .A(_08005_),
    .B(_07995_));
 sg13g2_nor2_1 _17288_ (.A(_07995_),
    .B(_08005_),
    .Y(_08040_));
 sg13g2_a21oi_1 _17289_ (.A1(_08039_),
    .A2(_07917_),
    .Y(_08041_),
    .B1(_08040_));
 sg13g2_nor2_1 _17290_ (.A(_08038_),
    .B(_08041_),
    .Y(_08042_));
 sg13g2_nand2_1 _17291_ (.Y(_08043_),
    .A(_08041_),
    .B(_08038_));
 sg13g2_nand2b_1 _17292_ (.Y(_08044_),
    .B(_08043_),
    .A_N(_08042_));
 sg13g2_nand2_1 _17293_ (.Y(_08045_),
    .A(_08014_),
    .B(_08009_));
 sg13g2_o21ai_1 _17294_ (.B1(_08010_),
    .Y(_08046_),
    .A1(_08045_),
    .A2(_07980_));
 sg13g2_a21oi_1 _17295_ (.A1(_08046_),
    .A2(_08044_),
    .Y(_08047_),
    .B1(_07522_));
 sg13g2_o21ai_1 _17296_ (.B1(_08047_),
    .Y(_08048_),
    .A1(_08044_),
    .A2(_08046_));
 sg13g2_buf_1 _17297_ (.A(_07952_),
    .X(_08049_));
 sg13g2_xnor2_1 _17298_ (.Y(_08050_),
    .A(_05093_),
    .B(net115));
 sg13g2_inv_1 _17299_ (.Y(_08051_),
    .A(_00129_));
 sg13g2_a22oi_1 _17300_ (.Y(_08052_),
    .B1(_06936_),
    .B2(_08020_),
    .A2(_08051_),
    .A1(_07996_));
 sg13g2_o21ai_1 _17301_ (.B1(_08052_),
    .Y(_08053_),
    .A1(_08019_),
    .A2(_07990_));
 sg13g2_xnor2_1 _17302_ (.Y(_08054_),
    .A(_08050_),
    .B(_08053_));
 sg13g2_a21oi_1 _17303_ (.A1(_08054_),
    .A2(net165),
    .Y(_08055_),
    .B1(net96));
 sg13g2_a22oi_1 _17304_ (.Y(_00378_),
    .B1(_08048_),
    .B2(_08055_),
    .A2(net90),
    .A1(_05093_));
 sg13g2_buf_1 _17305_ (.A(\vgadonut.donut.ycA[19] ),
    .X(_08056_));
 sg13g2_xnor2_1 _17306_ (.Y(_08057_),
    .A(_08056_),
    .B(_05095_));
 sg13g2_xnor2_1 _17307_ (.Y(_08058_),
    .A(_08057_),
    .B(_07878_));
 sg13g2_inv_1 _17308_ (.Y(_08059_),
    .A(_08030_));
 sg13g2_nor2_1 _17309_ (.A(_05062_),
    .B(_08059_),
    .Y(_08060_));
 sg13g2_a21oi_1 _17310_ (.A1(_07880_),
    .A2(_08031_),
    .Y(_08061_),
    .B1(_08060_));
 sg13g2_nor2_1 _17311_ (.A(_08058_),
    .B(_08061_),
    .Y(_08062_));
 sg13g2_inv_1 _17312_ (.Y(_08063_),
    .A(_08062_));
 sg13g2_nand2_1 _17313_ (.Y(_08064_),
    .A(_08061_),
    .B(_08058_));
 sg13g2_nand2_1 _17314_ (.Y(_08065_),
    .A(_08063_),
    .B(_08064_));
 sg13g2_a21oi_1 _17315_ (.A1(_08036_),
    .A2(net115),
    .Y(_08066_),
    .B1(_08034_));
 sg13g2_xnor2_1 _17316_ (.Y(_08067_),
    .A(_08065_),
    .B(_08066_));
 sg13g2_mux2_1 _17317_ (.A0(_08027_),
    .A1(_07996_),
    .S(_08037_),
    .X(_08068_));
 sg13g2_nor2_1 _17318_ (.A(_08067_),
    .B(_08068_),
    .Y(_08069_));
 sg13g2_nand2_1 _17319_ (.Y(_08070_),
    .A(_08068_),
    .B(_08067_));
 sg13g2_nor2b_1 _17320_ (.A(_08069_),
    .B_N(_08070_),
    .Y(_08071_));
 sg13g2_nor2_1 _17321_ (.A(_08011_),
    .B(_08016_),
    .Y(_08072_));
 sg13g2_nor3_1 _17322_ (.A(_08008_),
    .B(_08042_),
    .C(_08072_),
    .Y(_08073_));
 sg13g2_nor2b_1 _17323_ (.A(_08073_),
    .B_N(_08043_),
    .Y(_08074_));
 sg13g2_a21oi_1 _17324_ (.A1(_08074_),
    .A2(_08071_),
    .Y(_08075_),
    .B1(_07522_));
 sg13g2_o21ai_1 _17325_ (.B1(_08075_),
    .Y(_08076_),
    .A1(_08071_),
    .A2(_08074_));
 sg13g2_xnor2_1 _17326_ (.Y(_08077_),
    .A(\vgadonut.donut.donuthit.ryin[13] ),
    .B(net115));
 sg13g2_nand2b_1 _17327_ (.Y(_08078_),
    .B(_08053_),
    .A_N(_08050_));
 sg13g2_o21ai_1 _17328_ (.B1(_08078_),
    .Y(_08079_),
    .A1(_00130_),
    .A2(net115));
 sg13g2_xor2_1 _17329_ (.B(_08079_),
    .A(_08077_),
    .X(_08080_));
 sg13g2_a21oi_1 _17330_ (.A1(_08080_),
    .A2(net147),
    .Y(_08081_),
    .B1(_07956_));
 sg13g2_a22oi_1 _17331_ (.Y(_00379_),
    .B1(_08076_),
    .B2(_08081_),
    .A2(_07885_),
    .A1(_05133_));
 sg13g2_xnor2_1 _17332_ (.Y(_08082_),
    .A(_07563_),
    .B(_07732_));
 sg13g2_buf_1 _17333_ (.A(\vgadonut.donut.ycA[1] ),
    .X(_08083_));
 sg13g2_nor2b_1 _17334_ (.A(net163),
    .B_N(_08083_),
    .Y(_08084_));
 sg13g2_a21oi_1 _17335_ (.A1(_08082_),
    .A2(net160),
    .Y(_08085_),
    .B1(_08084_));
 sg13g2_nor2_1 _17336_ (.A(\vgadonut.donut.ry6[1] ),
    .B(net104),
    .Y(_08086_));
 sg13g2_a21oi_1 _17337_ (.A1(net105),
    .A2(_08085_),
    .Y(_00380_),
    .B1(_08086_));
 sg13g2_buf_1 _17338_ (.A(\vgadonut.donut.ycA[20] ),
    .X(_08087_));
 sg13g2_xnor2_1 _17339_ (.Y(_08088_),
    .A(_08087_),
    .B(_05135_));
 sg13g2_xor2_1 _17340_ (.B(_07917_),
    .A(_08088_),
    .X(_08089_));
 sg13g2_inv_1 _17341_ (.Y(_08090_),
    .A(_08056_));
 sg13g2_nand2_1 _17342_ (.Y(_08091_),
    .A(_07878_),
    .B(_08057_));
 sg13g2_o21ai_1 _17343_ (.B1(_08091_),
    .Y(_08092_),
    .A1(_08090_),
    .A2(_05095_));
 sg13g2_xnor2_1 _17344_ (.Y(_08093_),
    .A(_08089_),
    .B(_08092_));
 sg13g2_a21oi_1 _17345_ (.A1(_08064_),
    .A2(net115),
    .Y(_08094_),
    .B1(_08062_));
 sg13g2_xnor2_1 _17346_ (.Y(_08095_),
    .A(_08093_),
    .B(_08094_));
 sg13g2_mux2_1 _17347_ (.A0(_08066_),
    .A1(_07996_),
    .S(_08065_),
    .X(_08096_));
 sg13g2_xor2_1 _17348_ (.B(_08096_),
    .A(_08095_),
    .X(_08097_));
 sg13g2_inv_1 _17349_ (.Y(_08098_),
    .A(_08097_));
 sg13g2_o21ai_1 _17350_ (.B1(_08070_),
    .Y(_08099_),
    .A1(_08069_),
    .A2(_08074_));
 sg13g2_nor2_1 _17351_ (.A(_08098_),
    .B(_08099_),
    .Y(_08100_));
 sg13g2_a21oi_1 _17352_ (.A1(_08099_),
    .A2(_08098_),
    .Y(_08101_),
    .B1(net147));
 sg13g2_nand2b_1 _17353_ (.Y(_08102_),
    .B(_08101_),
    .A_N(_08100_));
 sg13g2_xnor2_1 _17354_ (.Y(_08103_),
    .A(_05167_),
    .B(net115));
 sg13g2_nand2_1 _17355_ (.Y(_08104_),
    .A(_08079_),
    .B(_08077_));
 sg13g2_o21ai_1 _17356_ (.B1(_08104_),
    .Y(_08105_),
    .A1(_00131_),
    .A2(net115));
 sg13g2_xnor2_1 _17357_ (.Y(_08106_),
    .A(_08103_),
    .B(_08105_));
 sg13g2_a21oi_1 _17358_ (.A1(_08106_),
    .A2(net164),
    .Y(_08107_),
    .B1(_07956_));
 sg13g2_a22oi_1 _17359_ (.Y(_00381_),
    .B1(_08102_),
    .B2(_08107_),
    .A2(_07885_),
    .A1(_05167_));
 sg13g2_mux2_1 _17360_ (.A0(_08094_),
    .A1(_07996_),
    .S(_08093_),
    .X(_08108_));
 sg13g2_xnor2_1 _17361_ (.Y(_08109_),
    .A(\vgadonut.donut.ycA[21] ),
    .B(_05169_));
 sg13g2_xor2_1 _17362_ (.B(net115),
    .A(_08109_),
    .X(_08110_));
 sg13g2_inv_1 _17363_ (.Y(_08111_),
    .A(_08087_));
 sg13g2_nor2_1 _17364_ (.A(_05135_),
    .B(_08111_),
    .Y(_08112_));
 sg13g2_a21oi_1 _17365_ (.A1(_07917_),
    .A2(_08088_),
    .Y(_08113_),
    .B1(_08112_));
 sg13g2_xor2_1 _17366_ (.B(_08113_),
    .A(_08110_),
    .X(_08114_));
 sg13g2_nand2_1 _17367_ (.Y(_08115_),
    .A(_08092_),
    .B(_08089_));
 sg13g2_o21ai_1 _17368_ (.B1(_08115_),
    .Y(_08116_),
    .A1(_07996_),
    .A2(_08093_));
 sg13g2_xor2_1 _17369_ (.B(_08116_),
    .A(_08114_),
    .X(_08117_));
 sg13g2_xnor2_1 _17370_ (.Y(_08118_),
    .A(_08108_),
    .B(_08117_));
 sg13g2_nor2_1 _17371_ (.A(_08095_),
    .B(_08096_),
    .Y(_08119_));
 sg13g2_nor2_1 _17372_ (.A(_08119_),
    .B(_08100_),
    .Y(_08120_));
 sg13g2_or2_1 _17373_ (.X(_08121_),
    .B(_08120_),
    .A(_08118_));
 sg13g2_a21oi_1 _17374_ (.A1(_08120_),
    .A2(_08118_),
    .Y(_08122_),
    .B1(net162));
 sg13g2_nor2_1 _17375_ (.A(_00132_),
    .B(_08049_),
    .Y(_08123_));
 sg13g2_a221oi_1 _17376_ (.B2(_05167_),
    .C1(_08123_),
    .B1(_08105_),
    .A1(_08049_),
    .Y(_08124_),
    .A2(_08104_));
 sg13g2_xnor2_1 _17377_ (.Y(_08125_),
    .A(_05222_),
    .B(_08124_));
 sg13g2_buf_1 _17378_ (.A(_06989_),
    .X(_08126_));
 sg13g2_a221oi_1 _17379_ (.B2(_06982_),
    .C1(net95),
    .B1(_08125_),
    .A1(_08121_),
    .Y(_08127_),
    .A2(_08122_));
 sg13g2_a21oi_1 _17380_ (.A1(_05222_),
    .A2(net93),
    .Y(_00382_),
    .B1(_08127_));
 sg13g2_nor2_1 _17381_ (.A(_07731_),
    .B(_07737_),
    .Y(_08128_));
 sg13g2_xnor2_1 _17382_ (.Y(_08129_),
    .A(_08128_),
    .B(_07735_));
 sg13g2_xnor2_1 _17383_ (.Y(_08130_),
    .A(_07562_),
    .B(_07680_));
 sg13g2_nor2_1 _17384_ (.A(_08130_),
    .B(net146),
    .Y(_08131_));
 sg13g2_a21oi_1 _17385_ (.A1(_08129_),
    .A2(net160),
    .Y(_08132_),
    .B1(_08131_));
 sg13g2_nor2_1 _17386_ (.A(\vgadonut.donut.ry6[2] ),
    .B(net107),
    .Y(_08133_));
 sg13g2_a21oi_1 _17387_ (.A1(_08132_),
    .A2(net105),
    .Y(_00383_),
    .B1(_08133_));
 sg13g2_nor2_1 _17388_ (.A(_07740_),
    .B(_07730_),
    .Y(_08134_));
 sg13g2_o21ai_1 _17389_ (.B1(net163),
    .Y(_08135_),
    .A1(_08134_),
    .A2(_07739_));
 sg13g2_a21o_1 _17390_ (.A2(_08134_),
    .A1(_07739_),
    .B1(_08135_),
    .X(_08136_));
 sg13g2_inv_1 _17391_ (.Y(_08137_),
    .A(_07680_));
 sg13g2_a21oi_1 _17392_ (.A1(_07562_),
    .A2(_08137_),
    .Y(_08138_),
    .B1(_07682_));
 sg13g2_nor2_1 _17393_ (.A(_08138_),
    .B(_07684_),
    .Y(_08139_));
 sg13g2_inv_1 _17394_ (.Y(_08140_),
    .A(_08139_));
 sg13g2_a21oi_1 _17395_ (.A1(net151),
    .A2(_08140_),
    .Y(_08141_),
    .B1(net96));
 sg13g2_a22oi_1 _17396_ (.Y(_00384_),
    .B1(_08136_),
    .B2(_08141_),
    .A2(net90),
    .A1(_07729_));
 sg13g2_nand2b_1 _17397_ (.Y(_08142_),
    .B(_07679_),
    .A_N(_07686_));
 sg13g2_nand2b_1 _17398_ (.Y(_08143_),
    .B(_07685_),
    .A_N(_08142_));
 sg13g2_a21oi_1 _17399_ (.A1(_08142_),
    .A2(_07684_),
    .Y(_08144_),
    .B1(net162));
 sg13g2_nor2_1 _17400_ (.A(_07728_),
    .B(_07745_),
    .Y(_08145_));
 sg13g2_xnor2_1 _17401_ (.Y(_08146_),
    .A(_08145_),
    .B(_07742_));
 sg13g2_a221oi_1 _17402_ (.B2(net170),
    .C1(net95),
    .B1(_08146_),
    .A1(_08143_),
    .Y(_08147_),
    .A2(_08144_));
 sg13g2_a21oi_1 _17403_ (.A1(_07743_),
    .A2(net93),
    .Y(_00385_),
    .B1(_08147_));
 sg13g2_nor3_1 _17404_ (.A(_07688_),
    .B(_07673_),
    .C(_07687_),
    .Y(_08148_));
 sg13g2_o21ai_1 _17405_ (.B1(_07687_),
    .Y(_08149_),
    .A1(_07688_),
    .A2(_07673_));
 sg13g2_nand3b_1 _17406_ (.B(net150),
    .C(_08149_),
    .Y(_08150_),
    .A_N(_08148_));
 sg13g2_nor2_1 _17407_ (.A(_07748_),
    .B(_07751_),
    .Y(_08151_));
 sg13g2_xor2_1 _17408_ (.B(_07747_),
    .A(_08151_),
    .X(_08152_));
 sg13g2_a21oi_1 _17409_ (.A1(_08152_),
    .A2(net164),
    .Y(_08153_),
    .B1(net96));
 sg13g2_a22oi_1 _17410_ (.Y(_00386_),
    .B1(_08150_),
    .B2(_08153_),
    .A2(net90),
    .A1(_07750_));
 sg13g2_xnor2_1 _17411_ (.Y(_08154_),
    .A(_07756_),
    .B(_07752_));
 sg13g2_nand2b_1 _17412_ (.Y(_08155_),
    .B(_07697_),
    .A_N(_07698_));
 sg13g2_a21oi_1 _17413_ (.A1(_08155_),
    .A2(_07689_),
    .Y(_08156_),
    .B1(_10106_));
 sg13g2_o21ai_1 _17414_ (.B1(_08156_),
    .Y(_08157_),
    .A1(_07689_),
    .A2(_08155_));
 sg13g2_nor2b_1 _17415_ (.A(net100),
    .B_N(_08157_),
    .Y(_08158_));
 sg13g2_o21ai_1 _17416_ (.B1(_08158_),
    .Y(_08159_),
    .A1(net150),
    .A2(_08154_));
 sg13g2_o21ai_1 _17417_ (.B1(_08159_),
    .Y(_00387_),
    .A1(_07754_),
    .A2(_07517_));
 sg13g2_a21oi_1 _17418_ (.A1(_07699_),
    .A2(_07708_),
    .Y(_08160_),
    .B1(net163));
 sg13g2_nand2b_1 _17419_ (.Y(_08161_),
    .B(_07700_),
    .A_N(_07708_));
 sg13g2_a21oi_1 _17420_ (.A1(_08160_),
    .A2(_08161_),
    .Y(_08162_),
    .B1(net97));
 sg13g2_nor2_1 _17421_ (.A(_07762_),
    .B(_07760_),
    .Y(_08163_));
 sg13g2_inv_1 _17422_ (.Y(_08164_),
    .A(_07755_));
 sg13g2_o21ai_1 _17423_ (.B1(_08164_),
    .Y(_08165_),
    .A1(_07753_),
    .A2(_07752_));
 sg13g2_a21oi_1 _17424_ (.A1(_08165_),
    .A2(_08163_),
    .Y(_08166_),
    .B1(net148));
 sg13g2_o21ai_1 _17425_ (.B1(_08166_),
    .Y(_08167_),
    .A1(_08163_),
    .A2(_08165_));
 sg13g2_a22oi_1 _17426_ (.Y(_00388_),
    .B1(_08162_),
    .B2(_08167_),
    .A2(net90),
    .A1(_07758_));
 sg13g2_buf_1 _17427_ (.A(net100),
    .X(_08168_));
 sg13g2_a21oi_1 _17428_ (.A1(_07700_),
    .A2(_07707_),
    .Y(_08169_),
    .B1(_07705_));
 sg13g2_nor2_1 _17429_ (.A(_07714_),
    .B(_08169_),
    .Y(_08170_));
 sg13g2_nand2_1 _17430_ (.Y(_08171_),
    .A(_08169_),
    .B(_07714_));
 sg13g2_nand3b_1 _17431_ (.B(net150),
    .C(_08171_),
    .Y(_08172_),
    .A_N(_08170_));
 sg13g2_inv_1 _17432_ (.Y(_08173_),
    .A(_07768_));
 sg13g2_xnor2_1 _17433_ (.Y(_08174_),
    .A(_08173_),
    .B(_07763_));
 sg13g2_a21oi_1 _17434_ (.A1(_08174_),
    .A2(net164),
    .Y(_08175_),
    .B1(net96));
 sg13g2_a22oi_1 _17435_ (.Y(_00389_),
    .B1(_08172_),
    .B2(_08175_),
    .A2(net89),
    .A1(_07765_));
 sg13g2_inv_1 _17436_ (.Y(_08176_),
    .A(\vgadonut.donut.donuthit.ryin[3] ));
 sg13g2_nand2_1 _17437_ (.Y(_08177_),
    .A(_07717_),
    .B(_07662_));
 sg13g2_nand3_1 _17438_ (.B(net151),
    .C(_08177_),
    .A(_07719_),
    .Y(_08178_));
 sg13g2_nor2_1 _17439_ (.A(_08176_),
    .B(_07725_),
    .Y(_08179_));
 sg13g2_nor2_1 _17440_ (.A(_08179_),
    .B(_07727_),
    .Y(_08180_));
 sg13g2_a221oi_1 _17441_ (.B2(_08163_),
    .C1(_07760_),
    .B1(_08165_),
    .A1(\vgadonut.donut.donuthit.ryin[2] ),
    .Y(_08181_),
    .A2(_07636_));
 sg13g2_nor2_1 _17442_ (.A(_07764_),
    .B(_08181_),
    .Y(_08182_));
 sg13g2_xor2_1 _17443_ (.B(_08182_),
    .A(_08180_),
    .X(_08183_));
 sg13g2_a21oi_1 _17444_ (.A1(_08183_),
    .A2(net164),
    .Y(_08184_),
    .B1(net96));
 sg13g2_a22oi_1 _17445_ (.Y(_00390_),
    .B1(_08178_),
    .B2(_08184_),
    .A2(net89),
    .A1(_08176_));
 sg13g2_inv_1 _17446_ (.Y(_08185_),
    .A(\vgadonut.donut.rz6[0] ));
 sg13g2_inv_1 _17447_ (.Y(_08186_),
    .A(\vgadonut.donut.ysA[0] ));
 sg13g2_nand2_1 _17448_ (.Y(_08187_),
    .A(\vgadonut.donut.rz6[0] ),
    .B(net217));
 sg13g2_nand2b_1 _17449_ (.Y(_08188_),
    .B(_08185_),
    .A_N(net217));
 sg13g2_nand3_1 _17450_ (.B(_08187_),
    .C(_08188_),
    .A(_06334_),
    .Y(_08189_));
 sg13g2_o21ai_1 _17451_ (.B1(_08189_),
    .Y(_08190_),
    .A1(_08186_),
    .A2(net170));
 sg13g2_nand2_1 _17452_ (.Y(_08191_),
    .A(net104),
    .B(_08190_));
 sg13g2_o21ai_1 _17453_ (.B1(_08191_),
    .Y(_00391_),
    .A1(_08185_),
    .A2(net104));
 sg13g2_inv_1 _17454_ (.Y(_08192_),
    .A(\vgadonut.donut.donuthit.rzin[4] ));
 sg13g2_nor2_1 _17455_ (.A(\vgadonut.donut.donuthit.rzin[4] ),
    .B(_06515_),
    .Y(_08193_));
 sg13g2_nand2_1 _17456_ (.Y(_08194_),
    .A(\vgadonut.donut.donuthit.rzin[4] ),
    .B(_06515_));
 sg13g2_nor2b_1 _17457_ (.A(_08193_),
    .B_N(_08194_),
    .Y(_08195_));
 sg13g2_nand2_1 _17458_ (.Y(_08196_),
    .A(\vgadonut.donut.donuthit.rzin[2] ),
    .B(_06534_));
 sg13g2_inv_1 _17459_ (.Y(_08197_),
    .A(_08196_));
 sg13g2_nor2_1 _17460_ (.A(\vgadonut.donut.donuthit.rzin[3] ),
    .B(_06519_),
    .Y(_08198_));
 sg13g2_nand2_1 _17461_ (.Y(_08199_),
    .A(\vgadonut.donut.donuthit.rzin[3] ),
    .B(_06519_));
 sg13g2_inv_1 _17462_ (.Y(_08200_),
    .A(_08199_));
 sg13g2_nor2_1 _17463_ (.A(_08198_),
    .B(_08200_),
    .Y(_08201_));
 sg13g2_nor2_1 _17464_ (.A(\vgadonut.donut.rz6[5] ),
    .B(_06441_),
    .Y(_08202_));
 sg13g2_xor2_1 _17465_ (.B(_06415_),
    .A(\vgadonut.donut.rz6[1] ),
    .X(_08203_));
 sg13g2_inv_1 _17466_ (.Y(_08204_),
    .A(_08203_));
 sg13g2_nand2_1 _17467_ (.Y(_08205_),
    .A(\vgadonut.donut.rz6[1] ),
    .B(_06415_));
 sg13g2_o21ai_1 _17468_ (.B1(_08205_),
    .Y(_08206_),
    .A1(_08187_),
    .A2(_08204_));
 sg13g2_nor2_1 _17469_ (.A(\vgadonut.donut.rz6[2] ),
    .B(_06412_),
    .Y(_08207_));
 sg13g2_inv_1 _17470_ (.Y(_08208_),
    .A(_08207_));
 sg13g2_nand2_1 _17471_ (.Y(_08209_),
    .A(\vgadonut.donut.rz6[2] ),
    .B(_06412_));
 sg13g2_inv_1 _17472_ (.Y(_08210_),
    .A(_08209_));
 sg13g2_a21oi_1 _17473_ (.A1(_08206_),
    .A2(_08208_),
    .Y(_08211_),
    .B1(_08210_));
 sg13g2_nand2_1 _17474_ (.Y(_08212_),
    .A(\vgadonut.donut.rz6[3] ),
    .B(_06427_));
 sg13g2_nor2_1 _17475_ (.A(\vgadonut.donut.rz6[3] ),
    .B(_06427_),
    .Y(_08213_));
 sg13g2_a21oi_1 _17476_ (.A1(_08211_),
    .A2(_08212_),
    .Y(_08214_),
    .B1(_08213_));
 sg13g2_nor2_1 _17477_ (.A(\vgadonut.donut.rz6[4] ),
    .B(_06433_),
    .Y(_08215_));
 sg13g2_inv_1 _17478_ (.Y(_08216_),
    .A(_08215_));
 sg13g2_nand2_1 _17479_ (.Y(_08217_),
    .A(\vgadonut.donut.rz6[4] ),
    .B(_06433_));
 sg13g2_inv_1 _17480_ (.Y(_08218_),
    .A(_08217_));
 sg13g2_a21oi_1 _17481_ (.A1(_08214_),
    .A2(_08216_),
    .Y(_08219_),
    .B1(_08218_));
 sg13g2_nand2_1 _17482_ (.Y(_08220_),
    .A(\vgadonut.donut.rz6[5] ),
    .B(_06441_));
 sg13g2_o21ai_1 _17483_ (.B1(_08220_),
    .Y(_08221_),
    .A1(_08202_),
    .A2(_08219_));
 sg13g2_nor2_1 _17484_ (.A(\vgadonut.donut.donuthit.rzin[0] ),
    .B(_06405_),
    .Y(_08222_));
 sg13g2_nand2_1 _17485_ (.Y(_08223_),
    .A(\vgadonut.donut.donuthit.rzin[0] ),
    .B(_06405_));
 sg13g2_inv_1 _17486_ (.Y(_08224_),
    .A(_08223_));
 sg13g2_nor2_1 _17487_ (.A(_08222_),
    .B(_08224_),
    .Y(_08225_));
 sg13g2_inv_1 _17488_ (.Y(_08226_),
    .A(_08225_));
 sg13g2_nor2_1 _17489_ (.A(\vgadonut.donut.donuthit.rzin[1] ),
    .B(_06526_),
    .Y(_08227_));
 sg13g2_nand2_1 _17490_ (.Y(_08228_),
    .A(\vgadonut.donut.donuthit.rzin[1] ),
    .B(_06526_));
 sg13g2_inv_1 _17491_ (.Y(_08229_),
    .A(_08228_));
 sg13g2_nor2_1 _17492_ (.A(_08227_),
    .B(_08229_),
    .Y(_08230_));
 sg13g2_inv_1 _17493_ (.Y(_08231_),
    .A(_08230_));
 sg13g2_nor2_1 _17494_ (.A(_08226_),
    .B(_08231_),
    .Y(_08232_));
 sg13g2_a21oi_1 _17495_ (.A1(_08223_),
    .A2(_08228_),
    .Y(_08233_),
    .B1(_08227_));
 sg13g2_a21oi_1 _17496_ (.A1(_08221_),
    .A2(_08232_),
    .Y(_08234_),
    .B1(_08233_));
 sg13g2_inv_1 _17497_ (.Y(_08235_),
    .A(_08234_));
 sg13g2_nor2_1 _17498_ (.A(\vgadonut.donut.donuthit.rzin[2] ),
    .B(_06534_),
    .Y(_08236_));
 sg13g2_nor2_1 _17499_ (.A(_08236_),
    .B(_08197_),
    .Y(_08237_));
 sg13g2_inv_1 _17500_ (.Y(_08238_),
    .A(_08237_));
 sg13g2_inv_1 _17501_ (.Y(_08239_),
    .A(_08201_));
 sg13g2_nor2_1 _17502_ (.A(_08238_),
    .B(_08239_),
    .Y(_08240_));
 sg13g2_a221oi_1 _17503_ (.B2(_08240_),
    .C1(_08200_),
    .B1(_08235_),
    .A1(_08197_),
    .Y(_08241_),
    .A2(_08201_));
 sg13g2_xnor2_1 _17504_ (.Y(_08242_),
    .A(_08195_),
    .B(_08241_));
 sg13g2_a21oi_1 _17505_ (.A1(_08242_),
    .A2(net161),
    .Y(_08243_),
    .B1(net97));
 sg13g2_inv_1 _17506_ (.Y(_08244_),
    .A(_00109_));
 sg13g2_buf_1 _17507_ (.A(\vgadonut.donut.ysA[7] ),
    .X(_08245_));
 sg13g2_xnor2_1 _17508_ (.Y(_08246_),
    .A(_08245_),
    .B(_05396_));
 sg13g2_nand2_1 _17509_ (.Y(_08247_),
    .A(_08245_),
    .B(_05396_));
 sg13g2_o21ai_1 _17510_ (.B1(_08247_),
    .Y(_08248_),
    .A1(_08244_),
    .A2(_08246_));
 sg13g2_buf_1 _17511_ (.A(\vgadonut.donut.ysA[8] ),
    .X(_08249_));
 sg13g2_inv_1 _17512_ (.Y(_08250_),
    .A(_08249_));
 sg13g2_nand2_1 _17513_ (.Y(_08251_),
    .A(_08250_),
    .B(_05405_));
 sg13g2_nand2_1 _17514_ (.Y(_08252_),
    .A(_08249_),
    .B(_05390_));
 sg13g2_buf_2 _17515_ (.A(_00110_),
    .X(_08253_));
 sg13g2_a21oi_1 _17516_ (.A1(_08251_),
    .A2(_08252_),
    .Y(_08254_),
    .B1(_08253_));
 sg13g2_nand3_1 _17517_ (.B(_08253_),
    .C(_08252_),
    .A(_08251_),
    .Y(_08255_));
 sg13g2_nand2b_1 _17518_ (.Y(_08256_),
    .B(_08255_),
    .A_N(_08254_));
 sg13g2_xnor2_1 _17519_ (.Y(_08257_),
    .A(_08248_),
    .B(_08256_));
 sg13g2_buf_2 _17520_ (.A(_00111_),
    .X(_08258_));
 sg13g2_nor2b_1 _17521_ (.A(_08256_),
    .B_N(_08248_),
    .Y(_08259_));
 sg13g2_a21oi_1 _17522_ (.A1(_08257_),
    .A2(_08258_),
    .Y(_08260_),
    .B1(_08259_));
 sg13g2_buf_2 _17523_ (.A(_00112_),
    .X(_08261_));
 sg13g2_nand2_1 _17524_ (.Y(_08262_),
    .A(_08255_),
    .B(_08252_));
 sg13g2_buf_1 _17525_ (.A(\vgadonut.donut.ysA[9] ),
    .X(_08263_));
 sg13g2_inv_1 _17526_ (.Y(_08264_),
    .A(_08263_));
 sg13g2_nand2_1 _17527_ (.Y(_08265_),
    .A(_08264_),
    .B(_05401_));
 sg13g2_nand2_1 _17528_ (.Y(_08266_),
    .A(_08263_),
    .B(_05380_));
 sg13g2_a21oi_1 _17529_ (.A1(_08265_),
    .A2(_08266_),
    .Y(_08267_),
    .B1(_08258_));
 sg13g2_nand3_1 _17530_ (.B(_08258_),
    .C(_08266_),
    .A(_08265_),
    .Y(_08268_));
 sg13g2_nand2b_1 _17531_ (.Y(_08269_),
    .B(_08268_),
    .A_N(_08267_));
 sg13g2_xnor2_1 _17532_ (.Y(_08270_),
    .A(_08262_),
    .B(_08269_));
 sg13g2_xnor2_1 _17533_ (.Y(_08271_),
    .A(_08261_),
    .B(_08270_));
 sg13g2_nor2_1 _17534_ (.A(_08260_),
    .B(_08271_),
    .Y(_08272_));
 sg13g2_inv_2 _17535_ (.Y(_08273_),
    .A(_00107_));
 sg13g2_xnor2_1 _17536_ (.Y(_08274_),
    .A(_08260_),
    .B(_08271_));
 sg13g2_nor2_1 _17537_ (.A(_08273_),
    .B(_08274_),
    .Y(_08275_));
 sg13g2_nor2_1 _17538_ (.A(_08272_),
    .B(_08275_),
    .Y(_08276_));
 sg13g2_nor2b_1 _17539_ (.A(_08269_),
    .B_N(_08262_),
    .Y(_08277_));
 sg13g2_a21oi_1 _17540_ (.A1(_08270_),
    .A2(_08261_),
    .Y(_08278_),
    .B1(_08277_));
 sg13g2_buf_2 _17541_ (.A(_00113_),
    .X(_08279_));
 sg13g2_nand2_1 _17542_ (.Y(_08280_),
    .A(_08268_),
    .B(_08266_));
 sg13g2_buf_1 _17543_ (.A(\vgadonut.donut.ysA[10] ),
    .X(_08281_));
 sg13g2_inv_1 _17544_ (.Y(_08282_),
    .A(_08281_));
 sg13g2_nand2_1 _17545_ (.Y(_08283_),
    .A(_08282_),
    .B(_06464_));
 sg13g2_nand2_1 _17546_ (.Y(_08284_),
    .A(_08281_),
    .B(net236));
 sg13g2_a21oi_1 _17547_ (.A1(_08283_),
    .A2(_08284_),
    .Y(_08285_),
    .B1(_08261_));
 sg13g2_nand3_1 _17548_ (.B(_08261_),
    .C(_08284_),
    .A(_08283_),
    .Y(_08286_));
 sg13g2_nand2b_1 _17549_ (.Y(_08287_),
    .B(_08286_),
    .A_N(_08285_));
 sg13g2_xnor2_1 _17550_ (.Y(_08288_),
    .A(_08280_),
    .B(_08287_));
 sg13g2_xnor2_1 _17551_ (.Y(_08289_),
    .A(_08279_),
    .B(_08288_));
 sg13g2_xnor2_1 _17552_ (.Y(_08290_),
    .A(_08278_),
    .B(_08289_));
 sg13g2_xnor2_1 _17553_ (.Y(_08291_),
    .A(_08244_),
    .B(_08290_));
 sg13g2_nor2_1 _17554_ (.A(_08276_),
    .B(_08291_),
    .Y(_08292_));
 sg13g2_inv_1 _17555_ (.Y(_08293_),
    .A(_08292_));
 sg13g2_nand2_1 _17556_ (.Y(_08294_),
    .A(_08291_),
    .B(_08276_));
 sg13g2_nand2_1 _17557_ (.Y(_08295_),
    .A(_08293_),
    .B(_08294_));
 sg13g2_inv_1 _17558_ (.Y(_08296_),
    .A(_00097_));
 sg13g2_xnor2_1 _17559_ (.Y(_08297_),
    .A(_08244_),
    .B(_08246_));
 sg13g2_buf_1 _17560_ (.A(\vgadonut.donut.ysA[6] ),
    .X(_08298_));
 sg13g2_xnor2_1 _17561_ (.Y(_08299_),
    .A(_08298_),
    .B(_05403_));
 sg13g2_nand2_1 _17562_ (.Y(_08300_),
    .A(_08298_),
    .B(_05403_));
 sg13g2_o21ai_1 _17563_ (.B1(_08300_),
    .Y(_08301_),
    .A1(_08273_),
    .A2(_08299_));
 sg13g2_xnor2_1 _17564_ (.Y(_08302_),
    .A(_08297_),
    .B(_08301_));
 sg13g2_xnor2_1 _17565_ (.Y(_08303_),
    .A(_08253_),
    .B(_08302_));
 sg13g2_xnor2_1 _17566_ (.Y(_08304_),
    .A(_08273_),
    .B(_08299_));
 sg13g2_buf_1 _17567_ (.A(\vgadonut.donut.ysA[5] ),
    .X(_08305_));
 sg13g2_inv_1 _17568_ (.Y(_08306_),
    .A(_08305_));
 sg13g2_xnor2_1 _17569_ (.Y(_08307_),
    .A(_06412_),
    .B(_08305_));
 sg13g2_nand2_1 _17570_ (.Y(_08308_),
    .A(_08307_),
    .B(_00107_));
 sg13g2_o21ai_1 _17571_ (.B1(_08308_),
    .Y(_08309_),
    .A1(_06412_),
    .A2(_08306_));
 sg13g2_xnor2_1 _17572_ (.Y(_08310_),
    .A(_08304_),
    .B(_08309_));
 sg13g2_nor2b_1 _17573_ (.A(_08304_),
    .B_N(_08309_),
    .Y(_08311_));
 sg13g2_a21oi_1 _17574_ (.A1(_08310_),
    .A2(_00109_),
    .Y(_08312_),
    .B1(_08311_));
 sg13g2_xnor2_1 _17575_ (.Y(_08313_),
    .A(_08303_),
    .B(_08312_));
 sg13g2_xnor2_1 _17576_ (.Y(_08314_),
    .A(_08296_),
    .B(_08313_));
 sg13g2_xnor2_1 _17577_ (.Y(_08315_),
    .A(_00109_),
    .B(_08310_));
 sg13g2_xnor2_1 _17578_ (.Y(_08316_),
    .A(_08273_),
    .B(_08307_));
 sg13g2_buf_2 _17579_ (.A(\vgadonut.donut.ysA[4] ),
    .X(_08317_));
 sg13g2_inv_1 _17580_ (.Y(_08318_),
    .A(_08317_));
 sg13g2_xnor2_1 _17581_ (.Y(_08319_),
    .A(_06415_),
    .B(_08317_));
 sg13g2_nand2_1 _17582_ (.Y(_08320_),
    .A(_08319_),
    .B(_00105_));
 sg13g2_o21ai_1 _17583_ (.B1(_08320_),
    .Y(_08321_),
    .A1(_06415_),
    .A2(_08318_));
 sg13g2_or2_1 _17584_ (.X(_08322_),
    .B(_08321_),
    .A(_08316_));
 sg13g2_nor2b_1 _17585_ (.A(_08315_),
    .B_N(_08322_),
    .Y(_08323_));
 sg13g2_xor2_1 _17586_ (.B(_08315_),
    .A(_08322_),
    .X(_08324_));
 sg13g2_nor2b_1 _17587_ (.A(_08324_),
    .B_N(_00108_),
    .Y(_08325_));
 sg13g2_nor2_1 _17588_ (.A(_08323_),
    .B(_08325_),
    .Y(_08326_));
 sg13g2_nor2_1 _17589_ (.A(_08314_),
    .B(_08326_),
    .Y(_08327_));
 sg13g2_inv_1 _17590_ (.Y(_08328_),
    .A(_00105_));
 sg13g2_xnor2_1 _17591_ (.Y(_08329_),
    .A(_08328_),
    .B(_08319_));
 sg13g2_buf_1 _17592_ (.A(\vgadonut.donut.ysA[3] ),
    .X(_08330_));
 sg13g2_inv_1 _17593_ (.Y(_08331_),
    .A(_08330_));
 sg13g2_xnor2_1 _17594_ (.Y(_08332_),
    .A(net217),
    .B(_08330_));
 sg13g2_nand2_1 _17595_ (.Y(_08333_),
    .A(_08332_),
    .B(_00097_));
 sg13g2_o21ai_1 _17596_ (.B1(_08333_),
    .Y(_08334_),
    .A1(_06419_),
    .A2(_08331_));
 sg13g2_nor2_1 _17597_ (.A(_08329_),
    .B(_08334_),
    .Y(_08335_));
 sg13g2_xnor2_1 _17598_ (.Y(_08336_),
    .A(_08316_),
    .B(_08321_));
 sg13g2_nor2b_1 _17599_ (.A(_08335_),
    .B_N(_08336_),
    .Y(_08337_));
 sg13g2_inv_1 _17600_ (.Y(_08338_),
    .A(_08337_));
 sg13g2_xor2_1 _17601_ (.B(_08324_),
    .A(_00108_),
    .X(_08339_));
 sg13g2_nor2_1 _17602_ (.A(_08338_),
    .B(_08339_),
    .Y(_08340_));
 sg13g2_buf_1 _17603_ (.A(\vgadonut.donut.ysA[2] ),
    .X(_08341_));
 sg13g2_nand2b_1 _17604_ (.Y(_08342_),
    .B(net217),
    .A_N(_08341_));
 sg13g2_xnor2_1 _17605_ (.Y(_08343_),
    .A(_00097_),
    .B(_08332_));
 sg13g2_nor2b_1 _17606_ (.A(_08342_),
    .B_N(_08343_),
    .Y(_08344_));
 sg13g2_inv_1 _17607_ (.Y(_08345_),
    .A(_08344_));
 sg13g2_xnor2_1 _17608_ (.Y(_08346_),
    .A(_08329_),
    .B(_08334_));
 sg13g2_nor2_1 _17609_ (.A(_08345_),
    .B(_08346_),
    .Y(_08347_));
 sg13g2_xor2_1 _17610_ (.B(_08336_),
    .A(_08335_),
    .X(_08348_));
 sg13g2_nor2_1 _17611_ (.A(_08347_),
    .B(_08348_),
    .Y(_08349_));
 sg13g2_inv_1 _17612_ (.Y(_08350_),
    .A(_08349_));
 sg13g2_xnor2_1 _17613_ (.Y(_08351_),
    .A(_08338_),
    .B(_08339_));
 sg13g2_nor2_1 _17614_ (.A(_08350_),
    .B(_08351_),
    .Y(_08352_));
 sg13g2_nor2_1 _17615_ (.A(_08340_),
    .B(_08352_),
    .Y(_08353_));
 sg13g2_inv_1 _17616_ (.Y(_08354_),
    .A(_08353_));
 sg13g2_nand2_1 _17617_ (.Y(_08355_),
    .A(_08326_),
    .B(_08314_));
 sg13g2_o21ai_1 _17618_ (.B1(_08355_),
    .Y(_08356_),
    .A1(_08327_),
    .A2(_08354_));
 sg13g2_inv_1 _17619_ (.Y(_08357_),
    .A(_08356_));
 sg13g2_nor2b_1 _17620_ (.A(_08297_),
    .B_N(_08301_),
    .Y(_08358_));
 sg13g2_a21oi_1 _17621_ (.A1(_08302_),
    .A2(_08253_),
    .Y(_08359_),
    .B1(_08358_));
 sg13g2_xnor2_1 _17622_ (.Y(_08360_),
    .A(_08258_),
    .B(_08257_));
 sg13g2_nor2_1 _17623_ (.A(_08359_),
    .B(_08360_),
    .Y(_08361_));
 sg13g2_xnor2_1 _17624_ (.Y(_08362_),
    .A(_08359_),
    .B(_08360_));
 sg13g2_nor2_1 _17625_ (.A(_08328_),
    .B(_08362_),
    .Y(_08363_));
 sg13g2_nor2_1 _17626_ (.A(_08361_),
    .B(_08363_),
    .Y(_08364_));
 sg13g2_xnor2_1 _17627_ (.Y(_08365_),
    .A(_08273_),
    .B(_08274_));
 sg13g2_xnor2_1 _17628_ (.Y(_08366_),
    .A(_08364_),
    .B(_08365_));
 sg13g2_nor2_1 _17629_ (.A(_08303_),
    .B(_08312_),
    .Y(_08367_));
 sg13g2_nor2_1 _17630_ (.A(_08296_),
    .B(_08313_),
    .Y(_08368_));
 sg13g2_nor2_1 _17631_ (.A(_08367_),
    .B(_08368_),
    .Y(_08369_));
 sg13g2_xnor2_1 _17632_ (.Y(_08370_),
    .A(_08328_),
    .B(_08362_));
 sg13g2_nor2_1 _17633_ (.A(_08369_),
    .B(_08370_),
    .Y(_08371_));
 sg13g2_inv_1 _17634_ (.Y(_08372_),
    .A(_08371_));
 sg13g2_nand2_1 _17635_ (.Y(_08373_),
    .A(_08370_),
    .B(_08369_));
 sg13g2_nand2_1 _17636_ (.Y(_08374_),
    .A(_08372_),
    .B(_08373_));
 sg13g2_nor2_1 _17637_ (.A(_08366_),
    .B(_08374_),
    .Y(_08375_));
 sg13g2_nand2b_1 _17638_ (.Y(_08376_),
    .B(_08371_),
    .A_N(_08366_));
 sg13g2_o21ai_1 _17639_ (.B1(_08376_),
    .Y(_08377_),
    .A1(_08364_),
    .A2(_08365_));
 sg13g2_a21oi_1 _17640_ (.A1(_08357_),
    .A2(_08375_),
    .Y(_08378_),
    .B1(_08377_));
 sg13g2_a21oi_1 _17641_ (.A1(_08378_),
    .A2(_08295_),
    .Y(_08379_),
    .B1(net149));
 sg13g2_o21ai_1 _17642_ (.B1(_08379_),
    .Y(_08380_),
    .A1(_08295_),
    .A2(_08378_));
 sg13g2_a22oi_1 _17643_ (.Y(_00392_),
    .B1(_08243_),
    .B2(_08380_),
    .A2(net89),
    .A1(_08192_));
 sg13g2_nor2_1 _17644_ (.A(\vgadonut.donut.donuthit.rzin[5] ),
    .B(_06546_),
    .Y(_08381_));
 sg13g2_nand2_1 _17645_ (.Y(_08382_),
    .A(\vgadonut.donut.donuthit.rzin[5] ),
    .B(_06546_));
 sg13g2_inv_1 _17646_ (.Y(_08383_),
    .A(_08382_));
 sg13g2_nor2_1 _17647_ (.A(_08381_),
    .B(_08383_),
    .Y(_08384_));
 sg13g2_inv_1 _17648_ (.Y(_08385_),
    .A(_08384_));
 sg13g2_inv_1 _17649_ (.Y(_08386_),
    .A(_08222_));
 sg13g2_a21oi_1 _17650_ (.A1(_08221_),
    .A2(_08386_),
    .Y(_08387_),
    .B1(_08224_));
 sg13g2_inv_1 _17651_ (.Y(_08388_),
    .A(_08387_));
 sg13g2_nor2_1 _17652_ (.A(_08238_),
    .B(_08231_),
    .Y(_08389_));
 sg13g2_a21oi_1 _17653_ (.A1(_08196_),
    .A2(_08228_),
    .Y(_08390_),
    .B1(_08236_));
 sg13g2_a21oi_1 _17654_ (.A1(_08388_),
    .A2(_08389_),
    .Y(_08391_),
    .B1(_08390_));
 sg13g2_nand2b_1 _17655_ (.Y(_08392_),
    .B(_08201_),
    .A_N(_08391_));
 sg13g2_nand2_1 _17656_ (.Y(_08393_),
    .A(_08194_),
    .B(_08199_));
 sg13g2_inv_1 _17657_ (.Y(_08394_),
    .A(_08393_));
 sg13g2_a21oi_1 _17658_ (.A1(_08392_),
    .A2(_08394_),
    .Y(_08395_),
    .B1(_08193_));
 sg13g2_xnor2_1 _17659_ (.Y(_08396_),
    .A(_08385_),
    .B(_08395_));
 sg13g2_a21oi_1 _17660_ (.A1(_08396_),
    .A2(net161),
    .Y(_08397_),
    .B1(net97));
 sg13g2_nor2_1 _17661_ (.A(_08278_),
    .B(_08289_),
    .Y(_08398_));
 sg13g2_nor2_1 _17662_ (.A(_08244_),
    .B(_08290_),
    .Y(_08399_));
 sg13g2_nor2_1 _17663_ (.A(_08398_),
    .B(_08399_),
    .Y(_08400_));
 sg13g2_nor2b_1 _17664_ (.A(_08287_),
    .B_N(_08280_),
    .Y(_08401_));
 sg13g2_a21oi_2 _17665_ (.B1(_08401_),
    .Y(_08402_),
    .A2(_08279_),
    .A1(_08288_));
 sg13g2_buf_2 _17666_ (.A(_00114_),
    .X(_08403_));
 sg13g2_nand2_1 _17667_ (.Y(_08404_),
    .A(_08286_),
    .B(_08284_));
 sg13g2_buf_1 _17668_ (.A(\vgadonut.donut.ysA[11] ),
    .X(_08405_));
 sg13g2_inv_1 _17669_ (.Y(_08406_),
    .A(_08405_));
 sg13g2_nand2_1 _17670_ (.Y(_08407_),
    .A(_08406_),
    .B(_06462_));
 sg13g2_nand2_1 _17671_ (.Y(_08408_),
    .A(_08405_),
    .B(net237));
 sg13g2_a21oi_1 _17672_ (.A1(_08407_),
    .A2(_08408_),
    .Y(_08409_),
    .B1(_08279_));
 sg13g2_nand3_1 _17673_ (.B(_08279_),
    .C(_08408_),
    .A(_08407_),
    .Y(_08410_));
 sg13g2_nand2b_1 _17674_ (.Y(_08411_),
    .B(_08410_),
    .A_N(_08409_));
 sg13g2_xnor2_1 _17675_ (.Y(_08412_),
    .A(_08404_),
    .B(_08411_));
 sg13g2_xnor2_1 _17676_ (.Y(_08413_),
    .A(_08403_),
    .B(_08412_));
 sg13g2_xnor2_1 _17677_ (.Y(_08414_),
    .A(_08402_),
    .B(_08413_));
 sg13g2_xor2_1 _17678_ (.B(_08414_),
    .A(_08253_),
    .X(_08415_));
 sg13g2_xnor2_1 _17679_ (.Y(_08416_),
    .A(_08400_),
    .B(_08415_));
 sg13g2_inv_1 _17680_ (.Y(_08417_),
    .A(_08378_));
 sg13g2_a21oi_1 _17681_ (.A1(_08417_),
    .A2(_08294_),
    .Y(_08418_),
    .B1(_08292_));
 sg13g2_a21oi_1 _17682_ (.A1(_08418_),
    .A2(_08416_),
    .Y(_08419_),
    .B1(net149));
 sg13g2_o21ai_1 _17683_ (.B1(_08419_),
    .Y(_08420_),
    .A1(_08416_),
    .A2(_08418_));
 sg13g2_a22oi_1 _17684_ (.Y(_00393_),
    .B1(_08397_),
    .B2(_08420_),
    .A2(net89),
    .A1(_05415_));
 sg13g2_nand2_1 _17685_ (.Y(_08421_),
    .A(_08413_),
    .B(_08402_));
 sg13g2_nor2_1 _17686_ (.A(_08402_),
    .B(_08413_),
    .Y(_08422_));
 sg13g2_a21oi_1 _17687_ (.A1(_08421_),
    .A2(_08253_),
    .Y(_08423_),
    .B1(_08422_));
 sg13g2_nor2b_1 _17688_ (.A(_08411_),
    .B_N(_08404_),
    .Y(_08424_));
 sg13g2_a21oi_2 _17689_ (.B1(_08424_),
    .Y(_08425_),
    .A2(_08403_),
    .A1(_08412_));
 sg13g2_buf_2 _17690_ (.A(_00115_),
    .X(_08426_));
 sg13g2_nand2_1 _17691_ (.Y(_08427_),
    .A(_08410_),
    .B(_08408_));
 sg13g2_buf_1 _17692_ (.A(\vgadonut.donut.ysA[12] ),
    .X(_08428_));
 sg13g2_inv_1 _17693_ (.Y(_08429_),
    .A(_08428_));
 sg13g2_nand2_1 _17694_ (.Y(_08430_),
    .A(_08429_),
    .B(_06482_));
 sg13g2_nand2_1 _17695_ (.Y(_08431_),
    .A(_08428_),
    .B(_05385_));
 sg13g2_a21oi_1 _17696_ (.A1(_08430_),
    .A2(_08431_),
    .Y(_08432_),
    .B1(_08403_));
 sg13g2_nand3_1 _17697_ (.B(_08403_),
    .C(_08431_),
    .A(_08430_),
    .Y(_08433_));
 sg13g2_nand2b_1 _17698_ (.Y(_08434_),
    .B(_08433_),
    .A_N(_08432_));
 sg13g2_xnor2_1 _17699_ (.Y(_08435_),
    .A(_08427_),
    .B(_08434_));
 sg13g2_xnor2_1 _17700_ (.Y(_08436_),
    .A(_08426_),
    .B(_08435_));
 sg13g2_xnor2_1 _17701_ (.Y(_08437_),
    .A(_08425_),
    .B(_08436_));
 sg13g2_xor2_1 _17702_ (.B(_08437_),
    .A(_08258_),
    .X(_08438_));
 sg13g2_nor2_1 _17703_ (.A(_08423_),
    .B(_08438_),
    .Y(_08439_));
 sg13g2_inv_1 _17704_ (.Y(_08440_),
    .A(_08439_));
 sg13g2_nand2_1 _17705_ (.Y(_08441_),
    .A(_08438_),
    .B(_08423_));
 sg13g2_nand2_1 _17706_ (.Y(_08442_),
    .A(_08440_),
    .B(_08441_));
 sg13g2_nor2_1 _17707_ (.A(_08416_),
    .B(_08295_),
    .Y(_08443_));
 sg13g2_nand2b_1 _17708_ (.Y(_08444_),
    .B(_08292_),
    .A_N(_08416_));
 sg13g2_o21ai_1 _17709_ (.B1(_08444_),
    .Y(_08445_),
    .A1(_08400_),
    .A2(_08415_));
 sg13g2_a21oi_1 _17710_ (.A1(_08417_),
    .A2(_08443_),
    .Y(_08446_),
    .B1(_08445_));
 sg13g2_a21oi_1 _17711_ (.A1(_08446_),
    .A2(_08442_),
    .Y(_08447_),
    .B1(net163));
 sg13g2_o21ai_1 _17712_ (.B1(_08447_),
    .Y(_08448_),
    .A1(_08442_),
    .A2(_08446_));
 sg13g2_nor2_1 _17713_ (.A(\vgadonut.donut.donuthit.rzin[6] ),
    .B(_06552_),
    .Y(_08449_));
 sg13g2_nand2_1 _17714_ (.Y(_08450_),
    .A(\vgadonut.donut.donuthit.rzin[6] ),
    .B(_06552_));
 sg13g2_inv_1 _17715_ (.Y(_08451_),
    .A(_08450_));
 sg13g2_nor2_1 _17716_ (.A(_08449_),
    .B(_08451_),
    .Y(_08452_));
 sg13g2_inv_1 _17717_ (.Y(_08453_),
    .A(_08452_));
 sg13g2_nand2b_1 _17718_ (.Y(_08454_),
    .B(_08195_),
    .A_N(_08241_));
 sg13g2_nand3_1 _17719_ (.B(_08194_),
    .C(_08382_),
    .A(_08454_),
    .Y(_08455_));
 sg13g2_nor2b_1 _17720_ (.A(_08381_),
    .B_N(_08455_),
    .Y(_08456_));
 sg13g2_xnor2_1 _17721_ (.Y(_08457_),
    .A(_08453_),
    .B(_08456_));
 sg13g2_a21oi_1 _17722_ (.A1(_08457_),
    .A2(net164),
    .Y(_08458_),
    .B1(net99));
 sg13g2_a22oi_1 _17723_ (.Y(_00394_),
    .B1(_08448_),
    .B2(_08458_),
    .A2(net89),
    .A1(_05420_));
 sg13g2_nor2_1 _17724_ (.A(_05502_),
    .B(_06513_),
    .Y(_08459_));
 sg13g2_nand2_1 _17725_ (.Y(_08460_),
    .A(_05502_),
    .B(_06513_));
 sg13g2_inv_1 _17726_ (.Y(_08461_),
    .A(_08460_));
 sg13g2_nor2_1 _17727_ (.A(_08459_),
    .B(_08461_),
    .Y(_08462_));
 sg13g2_nor2_1 _17728_ (.A(_08385_),
    .B(_08453_),
    .Y(_08463_));
 sg13g2_a221oi_1 _17729_ (.B2(_08463_),
    .C1(_08451_),
    .B1(_08395_),
    .A1(_08383_),
    .Y(_08464_),
    .A2(_08452_));
 sg13g2_xnor2_1 _17730_ (.Y(_08465_),
    .A(_08462_),
    .B(_08464_));
 sg13g2_a21oi_1 _17731_ (.A1(_08465_),
    .A2(net161),
    .Y(_08466_),
    .B1(net97));
 sg13g2_nand2_1 _17732_ (.Y(_08467_),
    .A(_08436_),
    .B(_08425_));
 sg13g2_nor2_1 _17733_ (.A(_08425_),
    .B(_08436_),
    .Y(_08468_));
 sg13g2_a21oi_2 _17734_ (.B1(_08468_),
    .Y(_08469_),
    .A2(_08258_),
    .A1(_08467_));
 sg13g2_nor2b_1 _17735_ (.A(_08434_),
    .B_N(_08427_),
    .Y(_08470_));
 sg13g2_a21oi_2 _17736_ (.B1(_08470_),
    .Y(_08471_),
    .A2(_08426_),
    .A1(_08435_));
 sg13g2_buf_2 _17737_ (.A(_00116_),
    .X(_08472_));
 sg13g2_nand2_1 _17738_ (.Y(_08473_),
    .A(_08433_),
    .B(_08431_));
 sg13g2_buf_1 _17739_ (.A(\vgadonut.donut.ysA[13] ),
    .X(_08474_));
 sg13g2_inv_1 _17740_ (.Y(_08475_),
    .A(_08474_));
 sg13g2_nand2_1 _17741_ (.Y(_08476_),
    .A(_08475_),
    .B(_06460_));
 sg13g2_nand2_1 _17742_ (.Y(_08477_),
    .A(_08474_),
    .B(_05421_));
 sg13g2_a21oi_1 _17743_ (.A1(_08476_),
    .A2(_08477_),
    .Y(_08478_),
    .B1(_08426_));
 sg13g2_nand3_1 _17744_ (.B(_08426_),
    .C(_08477_),
    .A(_08476_),
    .Y(_08479_));
 sg13g2_nand2b_1 _17745_ (.Y(_08480_),
    .B(_08479_),
    .A_N(_08478_));
 sg13g2_xnor2_1 _17746_ (.Y(_08481_),
    .A(_08473_),
    .B(_08480_));
 sg13g2_xnor2_1 _17747_ (.Y(_08482_),
    .A(_08472_),
    .B(_08481_));
 sg13g2_xnor2_1 _17748_ (.Y(_08483_),
    .A(_08471_),
    .B(_08482_));
 sg13g2_xor2_1 _17749_ (.B(_08483_),
    .A(_08261_),
    .X(_08484_));
 sg13g2_xnor2_1 _17750_ (.Y(_08485_),
    .A(_08469_),
    .B(_08484_));
 sg13g2_inv_1 _17751_ (.Y(_08486_),
    .A(_08446_));
 sg13g2_a21oi_1 _17752_ (.A1(_08486_),
    .A2(_08441_),
    .Y(_08487_),
    .B1(_08439_));
 sg13g2_a21oi_1 _17753_ (.A1(_08487_),
    .A2(_08485_),
    .Y(_08488_),
    .B1(net149));
 sg13g2_o21ai_1 _17754_ (.B1(_08488_),
    .Y(_08489_),
    .A1(_08485_),
    .A2(_08487_));
 sg13g2_a22oi_1 _17755_ (.Y(_00395_),
    .B1(_08466_),
    .B2(_08489_),
    .A2(net89),
    .A1(_05503_));
 sg13g2_inv_1 _17756_ (.Y(_08490_),
    .A(_08487_));
 sg13g2_nand2_1 _17757_ (.Y(_08491_),
    .A(_08484_),
    .B(_08469_));
 sg13g2_nor2_1 _17758_ (.A(_08469_),
    .B(_08484_),
    .Y(_08492_));
 sg13g2_a21oi_1 _17759_ (.A1(_08490_),
    .A2(_08491_),
    .Y(_08493_),
    .B1(_08492_));
 sg13g2_nand2_1 _17760_ (.Y(_08494_),
    .A(_08482_),
    .B(_08471_));
 sg13g2_nor2_1 _17761_ (.A(_08471_),
    .B(_08482_),
    .Y(_08495_));
 sg13g2_a21oi_2 _17762_ (.B1(_08495_),
    .Y(_08496_),
    .A2(_08261_),
    .A1(_08494_));
 sg13g2_nor2b_1 _17763_ (.A(_08480_),
    .B_N(_08473_),
    .Y(_08497_));
 sg13g2_a21oi_2 _17764_ (.B1(_08497_),
    .Y(_08498_),
    .A2(_08472_),
    .A1(_08481_));
 sg13g2_buf_2 _17765_ (.A(_00117_),
    .X(_08499_));
 sg13g2_nand2_1 _17766_ (.Y(_08500_),
    .A(_08479_),
    .B(_08477_));
 sg13g2_buf_1 _17767_ (.A(\vgadonut.donut.ysA[14] ),
    .X(_08501_));
 sg13g2_inv_1 _17768_ (.Y(_08502_),
    .A(_08501_));
 sg13g2_nand2_1 _17769_ (.Y(_08503_),
    .A(_08502_),
    .B(_06494_));
 sg13g2_nand2_1 _17770_ (.Y(_08504_),
    .A(_08501_),
    .B(net233));
 sg13g2_a21oi_1 _17771_ (.A1(_08503_),
    .A2(_08504_),
    .Y(_08505_),
    .B1(_08472_));
 sg13g2_nand3_1 _17772_ (.B(_08472_),
    .C(_08504_),
    .A(_08503_),
    .Y(_08506_));
 sg13g2_nand2b_1 _17773_ (.Y(_08507_),
    .B(_08506_),
    .A_N(_08505_));
 sg13g2_xnor2_1 _17774_ (.Y(_08508_),
    .A(_08500_),
    .B(_08507_));
 sg13g2_xnor2_1 _17775_ (.Y(_08509_),
    .A(_08499_),
    .B(_08508_));
 sg13g2_xnor2_1 _17776_ (.Y(_08510_),
    .A(_08498_),
    .B(_08509_));
 sg13g2_xor2_1 _17777_ (.B(_08510_),
    .A(_08279_),
    .X(_08511_));
 sg13g2_xnor2_1 _17778_ (.Y(_08512_),
    .A(_08496_),
    .B(_08511_));
 sg13g2_a21oi_1 _17779_ (.A1(_08493_),
    .A2(_08512_),
    .Y(_08513_),
    .B1(net147));
 sg13g2_nor2_1 _17780_ (.A(_08512_),
    .B(_08493_),
    .Y(_08514_));
 sg13g2_inv_1 _17781_ (.Y(_08515_),
    .A(_08514_));
 sg13g2_nand2_1 _17782_ (.Y(_08516_),
    .A(_08513_),
    .B(_08515_));
 sg13g2_xor2_1 _17783_ (.B(_06508_),
    .A(_05551_),
    .X(_08517_));
 sg13g2_a221oi_1 _17784_ (.B2(_08452_),
    .C1(_08451_),
    .B1(_08456_),
    .A1(_05502_),
    .Y(_08518_),
    .A2(_06513_));
 sg13g2_nor2_1 _17785_ (.A(_08459_),
    .B(_08518_),
    .Y(_08519_));
 sg13g2_xor2_1 _17786_ (.B(_08519_),
    .A(_08517_),
    .X(_08520_));
 sg13g2_a21oi_1 _17787_ (.A1(_08520_),
    .A2(net164),
    .Y(_08521_),
    .B1(net99));
 sg13g2_a22oi_1 _17788_ (.Y(_00396_),
    .B1(_08516_),
    .B2(_08521_),
    .A2(net89),
    .A1(_06965_));
 sg13g2_nand2_1 _17789_ (.Y(_08522_),
    .A(_06967_),
    .B(net184));
 sg13g2_nand2_1 _17790_ (.Y(_08523_),
    .A(_05595_),
    .B(_06505_));
 sg13g2_nand2_1 _17791_ (.Y(_08524_),
    .A(_08522_),
    .B(_08523_));
 sg13g2_nand2_1 _17792_ (.Y(_08525_),
    .A(_08462_),
    .B(_08517_));
 sg13g2_nand2_1 _17793_ (.Y(_08526_),
    .A(_05551_),
    .B(_06508_));
 sg13g2_inv_1 _17794_ (.Y(_08527_),
    .A(_08526_));
 sg13g2_a21oi_1 _17795_ (.A1(_08517_),
    .A2(_08461_),
    .Y(_08528_),
    .B1(_08527_));
 sg13g2_o21ai_1 _17796_ (.B1(_08528_),
    .Y(_08529_),
    .A1(_08525_),
    .A2(_08464_));
 sg13g2_xnor2_1 _17797_ (.Y(_08530_),
    .A(_08524_),
    .B(_08529_));
 sg13g2_a21oi_1 _17798_ (.A1(_08530_),
    .A2(net161),
    .Y(_08531_),
    .B1(net97));
 sg13g2_nand2_1 _17799_ (.Y(_08532_),
    .A(_08509_),
    .B(_08498_));
 sg13g2_nor2_1 _17800_ (.A(_08498_),
    .B(_08509_),
    .Y(_08533_));
 sg13g2_a21oi_1 _17801_ (.A1(_08532_),
    .A2(_08279_),
    .Y(_08534_),
    .B1(_08533_));
 sg13g2_nor2b_1 _17802_ (.A(_08507_),
    .B_N(_08500_),
    .Y(_08535_));
 sg13g2_a21oi_2 _17803_ (.B1(_08535_),
    .Y(_08536_),
    .A2(_08499_),
    .A1(_08508_));
 sg13g2_buf_2 _17804_ (.A(_00118_),
    .X(_08537_));
 sg13g2_nand2_1 _17805_ (.Y(_08538_),
    .A(_08506_),
    .B(_08504_));
 sg13g2_buf_1 _17806_ (.A(\vgadonut.donut.ysA[15] ),
    .X(_08539_));
 sg13g2_inv_1 _17807_ (.Y(_08540_),
    .A(_08539_));
 sg13g2_nand2_1 _17808_ (.Y(_08541_),
    .A(_08540_),
    .B(_06500_));
 sg13g2_nand2_1 _17809_ (.Y(_08542_),
    .A(_08539_),
    .B(net232));
 sg13g2_a21oi_1 _17810_ (.A1(_08541_),
    .A2(_08542_),
    .Y(_08543_),
    .B1(_08499_));
 sg13g2_nand3_1 _17811_ (.B(_08499_),
    .C(_08542_),
    .A(_08541_),
    .Y(_08544_));
 sg13g2_nand2b_1 _17812_ (.Y(_08545_),
    .B(_08544_),
    .A_N(_08543_));
 sg13g2_xnor2_1 _17813_ (.Y(_08546_),
    .A(_08538_),
    .B(_08545_));
 sg13g2_xnor2_1 _17814_ (.Y(_08547_),
    .A(_08537_),
    .B(_08546_));
 sg13g2_xnor2_1 _17815_ (.Y(_08548_),
    .A(_08536_),
    .B(_08547_));
 sg13g2_xor2_1 _17816_ (.B(_08548_),
    .A(_08403_),
    .X(_08549_));
 sg13g2_nor2_1 _17817_ (.A(_08534_),
    .B(_08549_),
    .Y(_08550_));
 sg13g2_nand2_1 _17818_ (.Y(_08551_),
    .A(_08549_),
    .B(_08534_));
 sg13g2_nand2b_1 _17819_ (.Y(_08552_),
    .B(_08551_),
    .A_N(_08550_));
 sg13g2_nor2_1 _17820_ (.A(_08496_),
    .B(_08511_),
    .Y(_08553_));
 sg13g2_a21oi_1 _17821_ (.A1(_08496_),
    .A2(_08511_),
    .Y(_08554_),
    .B1(_08493_));
 sg13g2_nor2_1 _17822_ (.A(_08553_),
    .B(_08554_),
    .Y(_08555_));
 sg13g2_a21oi_1 _17823_ (.A1(_08555_),
    .A2(_08552_),
    .Y(_08556_),
    .B1(net149));
 sg13g2_o21ai_1 _17824_ (.B1(_08556_),
    .Y(_08557_),
    .A1(_08552_),
    .A2(_08555_));
 sg13g2_a22oi_1 _17825_ (.Y(_00397_),
    .B1(_08531_),
    .B2(_08557_),
    .A2(net89),
    .A1(_06967_));
 sg13g2_a21oi_1 _17826_ (.A1(_08553_),
    .A2(_08551_),
    .Y(_08558_),
    .B1(_08550_));
 sg13g2_o21ai_1 _17827_ (.B1(_08558_),
    .Y(_08559_),
    .A1(_08552_),
    .A2(_08515_));
 sg13g2_inv_1 _17828_ (.Y(_08560_),
    .A(_08559_));
 sg13g2_nand2_1 _17829_ (.Y(_08561_),
    .A(_08547_),
    .B(_08536_));
 sg13g2_nor2_1 _17830_ (.A(_08536_),
    .B(_08547_),
    .Y(_08562_));
 sg13g2_a21oi_1 _17831_ (.A1(_08561_),
    .A2(_08403_),
    .Y(_08563_),
    .B1(_08562_));
 sg13g2_nor2b_1 _17832_ (.A(_08545_),
    .B_N(_08538_),
    .Y(_08564_));
 sg13g2_a21oi_2 _17833_ (.B1(_08564_),
    .Y(_08565_),
    .A2(_08537_),
    .A1(_08546_));
 sg13g2_buf_2 _17834_ (.A(_00119_),
    .X(_08566_));
 sg13g2_nand2_1 _17835_ (.Y(_08567_),
    .A(_08544_),
    .B(_08542_));
 sg13g2_buf_1 _17836_ (.A(\vgadonut.donut.ysA[16] ),
    .X(_08568_));
 sg13g2_inv_1 _17837_ (.Y(_08569_),
    .A(_08568_));
 sg13g2_nand2_1 _17838_ (.Y(_08570_),
    .A(_08569_),
    .B(_06454_));
 sg13g2_nand2_1 _17839_ (.Y(_08571_),
    .A(_08568_),
    .B(net203));
 sg13g2_a21oi_1 _17840_ (.A1(_08570_),
    .A2(_08571_),
    .Y(_08572_),
    .B1(_08537_));
 sg13g2_nand3_1 _17841_ (.B(_08537_),
    .C(_08571_),
    .A(_08570_),
    .Y(_08573_));
 sg13g2_nand2b_1 _17842_ (.Y(_08574_),
    .B(_08573_),
    .A_N(_08572_));
 sg13g2_xnor2_1 _17843_ (.Y(_08575_),
    .A(_08567_),
    .B(_08574_));
 sg13g2_xnor2_1 _17844_ (.Y(_08576_),
    .A(_08566_),
    .B(_08575_));
 sg13g2_xnor2_1 _17845_ (.Y(_08577_),
    .A(_08565_),
    .B(_08576_));
 sg13g2_xor2_1 _17846_ (.B(_08577_),
    .A(_08426_),
    .X(_08578_));
 sg13g2_nor2_1 _17847_ (.A(_08563_),
    .B(_08578_),
    .Y(_08579_));
 sg13g2_nand2_1 _17848_ (.Y(_08580_),
    .A(_08578_),
    .B(_08563_));
 sg13g2_nand2b_1 _17849_ (.Y(_08581_),
    .B(_08580_),
    .A_N(_08579_));
 sg13g2_a21oi_1 _17850_ (.A1(_08560_),
    .A2(_08581_),
    .Y(_08582_),
    .B1(net147));
 sg13g2_nor2_1 _17851_ (.A(_08581_),
    .B(_08560_),
    .Y(_08583_));
 sg13g2_inv_1 _17852_ (.Y(_08584_),
    .A(_08583_));
 sg13g2_nand2_1 _17853_ (.Y(_08585_),
    .A(_08582_),
    .B(_08584_));
 sg13g2_buf_1 _17854_ (.A(_06505_),
    .X(_08586_));
 sg13g2_xor2_1 _17855_ (.B(_05639_),
    .A(net189),
    .X(_08587_));
 sg13g2_inv_1 _17856_ (.Y(_08588_),
    .A(_08587_));
 sg13g2_nand2_1 _17857_ (.Y(_08589_),
    .A(_08526_),
    .B(_08523_));
 sg13g2_nand2_1 _17858_ (.Y(_08590_),
    .A(_08519_),
    .B(_08517_));
 sg13g2_inv_1 _17859_ (.Y(_08591_),
    .A(_08590_));
 sg13g2_o21ai_1 _17860_ (.B1(_08522_),
    .Y(_08592_),
    .A1(_08589_),
    .A2(_08591_));
 sg13g2_nor2_1 _17861_ (.A(_08588_),
    .B(_08592_),
    .Y(_08593_));
 sg13g2_nor2_1 _17862_ (.A(net148),
    .B(_08593_),
    .Y(_08594_));
 sg13g2_nand2_1 _17863_ (.Y(_08595_),
    .A(_08592_),
    .B(_08588_));
 sg13g2_a21oi_1 _17864_ (.A1(_08594_),
    .A2(_08595_),
    .Y(_08596_),
    .B1(net99));
 sg13g2_a22oi_1 _17865_ (.Y(_00398_),
    .B1(_08585_),
    .B2(_08596_),
    .A2(_08168_),
    .A1(_05640_));
 sg13g2_xor2_1 _17866_ (.B(_05691_),
    .A(_06505_),
    .X(_08597_));
 sg13g2_inv_1 _17867_ (.Y(_08598_),
    .A(_08597_));
 sg13g2_nand4_1 _17868_ (.B(_08523_),
    .C(_08522_),
    .A(_08529_),
    .Y(_08599_),
    .D(_08587_));
 sg13g2_o21ai_1 _17869_ (.B1(net189),
    .Y(_08600_),
    .A1(_05595_),
    .A2(_05639_));
 sg13g2_nand2_1 _17870_ (.Y(_08601_),
    .A(_08599_),
    .B(_08600_));
 sg13g2_xnor2_1 _17871_ (.Y(_08602_),
    .A(_08598_),
    .B(_08601_));
 sg13g2_a21oi_1 _17872_ (.A1(_08602_),
    .A2(net161),
    .Y(_08603_),
    .B1(net95));
 sg13g2_nand2_1 _17873_ (.Y(_08604_),
    .A(_08576_),
    .B(_08565_));
 sg13g2_nor2_1 _17874_ (.A(_08565_),
    .B(_08576_),
    .Y(_08605_));
 sg13g2_a21oi_1 _17875_ (.A1(_08604_),
    .A2(_08426_),
    .Y(_08606_),
    .B1(_08605_));
 sg13g2_nor2b_1 _17876_ (.A(_08574_),
    .B_N(_08567_),
    .Y(_08607_));
 sg13g2_a21oi_2 _17877_ (.B1(_08607_),
    .Y(_08608_),
    .A2(_08566_),
    .A1(_08575_));
 sg13g2_buf_1 _17878_ (.A(_00120_),
    .X(_08609_));
 sg13g2_nand2_1 _17879_ (.Y(_08610_),
    .A(_08573_),
    .B(_08571_));
 sg13g2_buf_1 _17880_ (.A(\vgadonut.donut.ysA[17] ),
    .X(_08611_));
 sg13g2_inv_1 _17881_ (.Y(_08612_),
    .A(_08611_));
 sg13g2_nand2b_1 _17882_ (.Y(_08613_),
    .B(_08612_),
    .A_N(_05643_));
 sg13g2_nand2_1 _17883_ (.Y(_08614_),
    .A(_08611_),
    .B(_05643_));
 sg13g2_a21oi_1 _17884_ (.A1(_08613_),
    .A2(_08614_),
    .Y(_08615_),
    .B1(_08566_));
 sg13g2_nand3_1 _17885_ (.B(_08566_),
    .C(_08614_),
    .A(_08613_),
    .Y(_08616_));
 sg13g2_nand2b_1 _17886_ (.Y(_08617_),
    .B(_08616_),
    .A_N(_08615_));
 sg13g2_xnor2_1 _17887_ (.Y(_08618_),
    .A(_08610_),
    .B(_08617_));
 sg13g2_xnor2_1 _17888_ (.Y(_08619_),
    .A(_08609_),
    .B(_08618_));
 sg13g2_xnor2_1 _17889_ (.Y(_08620_),
    .A(_08608_),
    .B(_08619_));
 sg13g2_xor2_1 _17890_ (.B(_08620_),
    .A(_08472_),
    .X(_08621_));
 sg13g2_nor2_1 _17891_ (.A(_08606_),
    .B(_08621_),
    .Y(_08622_));
 sg13g2_nand2_1 _17892_ (.Y(_08623_),
    .A(_08621_),
    .B(_08606_));
 sg13g2_nand2b_1 _17893_ (.Y(_08624_),
    .B(_08623_),
    .A_N(_08622_));
 sg13g2_a21oi_1 _17894_ (.A1(_08559_),
    .A2(_08580_),
    .Y(_08625_),
    .B1(_08579_));
 sg13g2_a21oi_1 _17895_ (.A1(_08625_),
    .A2(_08624_),
    .Y(_08626_),
    .B1(net149));
 sg13g2_o21ai_1 _17896_ (.B1(_08626_),
    .Y(_08627_),
    .A1(_08624_),
    .A2(_08625_));
 sg13g2_a22oi_1 _17897_ (.Y(_00399_),
    .B1(_08603_),
    .B2(_08627_),
    .A2(_08168_),
    .A1(_06953_));
 sg13g2_xor2_1 _17898_ (.B(_05727_),
    .A(_06505_),
    .X(_08628_));
 sg13g2_o21ai_1 _17899_ (.B1(_08586_),
    .Y(_08629_),
    .A1(_05639_),
    .A2(_05691_));
 sg13g2_inv_1 _17900_ (.Y(_08630_),
    .A(_08629_));
 sg13g2_nand2_1 _17901_ (.Y(_08631_),
    .A(_08593_),
    .B(_08597_));
 sg13g2_inv_1 _17902_ (.Y(_08632_),
    .A(_08631_));
 sg13g2_nor2_1 _17903_ (.A(_08630_),
    .B(_08632_),
    .Y(_08633_));
 sg13g2_xnor2_1 _17904_ (.Y(_08634_),
    .A(_08628_),
    .B(_08633_));
 sg13g2_a21oi_1 _17905_ (.A1(_08634_),
    .A2(net161),
    .Y(_08635_),
    .B1(net95));
 sg13g2_nand2_1 _17906_ (.Y(_08636_),
    .A(_08619_),
    .B(_08608_));
 sg13g2_nor2_1 _17907_ (.A(_08608_),
    .B(_08619_),
    .Y(_08637_));
 sg13g2_a21oi_1 _17908_ (.A1(_08636_),
    .A2(_08472_),
    .Y(_08638_),
    .B1(_08637_));
 sg13g2_inv_1 _17909_ (.Y(_08639_),
    .A(_08499_));
 sg13g2_inv_2 _17910_ (.Y(_08640_),
    .A(_08609_));
 sg13g2_nand2_1 _17911_ (.Y(_08641_),
    .A(_08616_),
    .B(_08614_));
 sg13g2_buf_2 _17912_ (.A(\vgadonut.donut.ysA[18] ),
    .X(_08642_));
 sg13g2_xnor2_1 _17913_ (.Y(_08643_),
    .A(_08642_),
    .B(net201));
 sg13g2_xnor2_1 _17914_ (.Y(_08644_),
    .A(net184),
    .B(_08643_));
 sg13g2_xnor2_1 _17915_ (.Y(_08645_),
    .A(_08641_),
    .B(_08644_));
 sg13g2_xnor2_1 _17916_ (.Y(_08646_),
    .A(_08640_),
    .B(_08645_));
 sg13g2_nor2b_1 _17917_ (.A(_08617_),
    .B_N(_08610_),
    .Y(_08647_));
 sg13g2_a21oi_1 _17918_ (.A1(_08618_),
    .A2(_08609_),
    .Y(_08648_),
    .B1(_08647_));
 sg13g2_xnor2_1 _17919_ (.Y(_08649_),
    .A(_08646_),
    .B(_08648_));
 sg13g2_xnor2_1 _17920_ (.Y(_08650_),
    .A(_08639_),
    .B(_08649_));
 sg13g2_nor2_1 _17921_ (.A(_08638_),
    .B(_08650_),
    .Y(_08651_));
 sg13g2_nand2_1 _17922_ (.Y(_08652_),
    .A(_08650_),
    .B(_08638_));
 sg13g2_nor2b_1 _17923_ (.A(_08651_),
    .B_N(_08652_),
    .Y(_08653_));
 sg13g2_a21oi_1 _17924_ (.A1(_08623_),
    .A2(_08579_),
    .Y(_08654_),
    .B1(_08622_));
 sg13g2_o21ai_1 _17925_ (.B1(_08654_),
    .Y(_08655_),
    .A1(_08624_),
    .A2(_08584_));
 sg13g2_a21oi_1 _17926_ (.A1(_08655_),
    .A2(_08653_),
    .Y(_08656_),
    .B1(net149));
 sg13g2_o21ai_1 _17927_ (.B1(_08656_),
    .Y(_08657_),
    .A1(_08653_),
    .A2(_08655_));
 sg13g2_a22oi_1 _17928_ (.Y(_00400_),
    .B1(_08635_),
    .B2(_08657_),
    .A2(net91),
    .A1(_06955_));
 sg13g2_xor2_1 _17929_ (.B(_05770_),
    .A(net189),
    .X(_08658_));
 sg13g2_inv_1 _17930_ (.Y(_08659_),
    .A(_08658_));
 sg13g2_inv_1 _17931_ (.Y(_08660_),
    .A(_08628_));
 sg13g2_nor2_1 _17932_ (.A(_08598_),
    .B(_08660_),
    .Y(_08661_));
 sg13g2_inv_1 _17933_ (.Y(_08662_),
    .A(_08661_));
 sg13g2_nor2_1 _17934_ (.A(_08600_),
    .B(_08662_),
    .Y(_08663_));
 sg13g2_nand2_1 _17935_ (.Y(_08664_),
    .A(net189),
    .B(_05691_));
 sg13g2_inv_1 _17936_ (.Y(_08665_),
    .A(_08664_));
 sg13g2_nand2_1 _17937_ (.Y(_08666_),
    .A(net189),
    .B(_05727_));
 sg13g2_inv_1 _17938_ (.Y(_08667_),
    .A(_08666_));
 sg13g2_nor2_1 _17939_ (.A(_08665_),
    .B(_08667_),
    .Y(_08668_));
 sg13g2_nor2b_1 _17940_ (.A(_08663_),
    .B_N(_08668_),
    .Y(_08669_));
 sg13g2_o21ai_1 _17941_ (.B1(_08669_),
    .Y(_08670_),
    .A1(_08662_),
    .A2(_08599_));
 sg13g2_xnor2_1 _17942_ (.Y(_08671_),
    .A(_08659_),
    .B(_08670_));
 sg13g2_a21oi_1 _17943_ (.A1(_08671_),
    .A2(net161),
    .Y(_08672_),
    .B1(net95));
 sg13g2_a21oi_1 _17944_ (.A1(_08655_),
    .A2(_08652_),
    .Y(_08673_),
    .B1(_08651_));
 sg13g2_inv_1 _17945_ (.Y(_08674_),
    .A(_08673_));
 sg13g2_nand2_1 _17946_ (.Y(_08675_),
    .A(_08643_),
    .B(_06505_));
 sg13g2_o21ai_1 _17947_ (.B1(_08675_),
    .Y(_08676_),
    .A1(_08643_),
    .A2(_08641_));
 sg13g2_nand2_1 _17948_ (.Y(_08677_),
    .A(_08642_),
    .B(_05694_));
 sg13g2_inv_1 _17949_ (.Y(_08678_),
    .A(_08642_));
 sg13g2_a21oi_1 _17950_ (.A1(_08678_),
    .A2(_06667_),
    .Y(_08679_),
    .B1(_08640_));
 sg13g2_a21oi_1 _17951_ (.A1(_08640_),
    .A2(_08677_),
    .Y(_08680_),
    .B1(_08679_));
 sg13g2_buf_2 _17952_ (.A(\vgadonut.donut.ysA[19] ),
    .X(_08681_));
 sg13g2_nor2_1 _17953_ (.A(_08681_),
    .B(_05730_),
    .Y(_08682_));
 sg13g2_nand2_1 _17954_ (.Y(_08683_),
    .A(_08681_),
    .B(_05730_));
 sg13g2_inv_1 _17955_ (.Y(_08684_),
    .A(_08683_));
 sg13g2_nor2_1 _17956_ (.A(_08682_),
    .B(_08684_),
    .Y(_08685_));
 sg13g2_xnor2_1 _17957_ (.Y(_08686_),
    .A(net184),
    .B(_08685_));
 sg13g2_xnor2_1 _17958_ (.Y(_08687_),
    .A(_08680_),
    .B(_08686_));
 sg13g2_xor2_1 _17959_ (.B(_08687_),
    .A(_08676_),
    .X(_08688_));
 sg13g2_xnor2_1 _17960_ (.Y(_08689_),
    .A(_08537_),
    .B(_08688_));
 sg13g2_inv_1 _17961_ (.Y(_08690_),
    .A(_08689_));
 sg13g2_nor2_1 _17962_ (.A(_08646_),
    .B(_08648_),
    .Y(_08691_));
 sg13g2_nor2_1 _17963_ (.A(_08639_),
    .B(_08649_),
    .Y(_08692_));
 sg13g2_nor2_1 _17964_ (.A(_08691_),
    .B(_08692_),
    .Y(_08693_));
 sg13g2_nor2_1 _17965_ (.A(_08690_),
    .B(_08693_),
    .Y(_08694_));
 sg13g2_nand2_1 _17966_ (.Y(_08695_),
    .A(_08693_),
    .B(_08690_));
 sg13g2_nor2b_1 _17967_ (.A(_08694_),
    .B_N(_08695_),
    .Y(_08696_));
 sg13g2_nand2_1 _17968_ (.Y(_08697_),
    .A(_08674_),
    .B(_08696_));
 sg13g2_nand2b_1 _17969_ (.Y(_08698_),
    .B(_08673_),
    .A_N(_08696_));
 sg13g2_nand3_1 _17970_ (.B(net151),
    .C(_08698_),
    .A(_08697_),
    .Y(_08699_));
 sg13g2_a22oi_1 _17971_ (.Y(_00401_),
    .B1(_08672_),
    .B2(_08699_),
    .A2(net91),
    .A1(_06957_));
 sg13g2_xnor2_1 _17972_ (.Y(_08700_),
    .A(_08187_),
    .B(_08203_));
 sg13g2_buf_1 _17973_ (.A(\vgadonut.donut.ysA[1] ),
    .X(_08701_));
 sg13g2_nor2b_1 _17974_ (.A(net170),
    .B_N(_08701_),
    .Y(_08702_));
 sg13g2_a21oi_1 _17975_ (.A1(net160),
    .A2(_08700_),
    .Y(_08703_),
    .B1(_08702_));
 sg13g2_nor2_1 _17976_ (.A(\vgadonut.donut.rz6[1] ),
    .B(net107),
    .Y(_08704_));
 sg13g2_a21oi_1 _17977_ (.A1(net105),
    .A2(_08703_),
    .Y(_00402_),
    .B1(_08704_));
 sg13g2_xor2_1 _17978_ (.B(\vgadonut.donut.donuthit.rzin[14] ),
    .A(net189),
    .X(_08705_));
 sg13g2_nor2_1 _17979_ (.A(_08660_),
    .B(_08659_),
    .Y(_08706_));
 sg13g2_a21oi_1 _17980_ (.A1(_08706_),
    .A2(_08630_),
    .Y(_08707_),
    .B1(_08667_));
 sg13g2_o21ai_1 _17981_ (.B1(_08707_),
    .Y(_08708_),
    .A1(net184),
    .A2(_06957_));
 sg13g2_a21oi_1 _17982_ (.A1(_08632_),
    .A2(_08706_),
    .Y(_08709_),
    .B1(_08708_));
 sg13g2_xnor2_1 _17983_ (.Y(_08710_),
    .A(_08705_),
    .B(_08709_));
 sg13g2_a21oi_1 _17984_ (.A1(_08710_),
    .A2(_07521_),
    .Y(_08711_),
    .B1(_08126_));
 sg13g2_inv_1 _17985_ (.Y(_08712_),
    .A(_08566_));
 sg13g2_nor2b_1 _17986_ (.A(_08679_),
    .B_N(_08677_),
    .Y(_08713_));
 sg13g2_nor2_1 _17987_ (.A(net184),
    .B(_08685_),
    .Y(_08714_));
 sg13g2_a21oi_1 _17988_ (.A1(_08713_),
    .A2(_08685_),
    .Y(_08715_),
    .B1(_08714_));
 sg13g2_nor2_1 _17989_ (.A(_08640_),
    .B(_08682_),
    .Y(_08716_));
 sg13g2_a21oi_1 _17990_ (.A1(_08640_),
    .A2(_08683_),
    .Y(_08717_),
    .B1(_08716_));
 sg13g2_buf_1 _17991_ (.A(\vgadonut.donut.ysA[20] ),
    .X(_08718_));
 sg13g2_nor2_1 _17992_ (.A(_08718_),
    .B(net199),
    .Y(_08719_));
 sg13g2_nand2_1 _17993_ (.Y(_08720_),
    .A(_08718_),
    .B(net199));
 sg13g2_nor2b_1 _17994_ (.A(_08719_),
    .B_N(_08720_),
    .Y(_08721_));
 sg13g2_xnor2_1 _17995_ (.Y(_08722_),
    .A(net184),
    .B(_08721_));
 sg13g2_xnor2_1 _17996_ (.Y(_08723_),
    .A(_08717_),
    .B(_08722_));
 sg13g2_xnor2_1 _17997_ (.Y(_08724_),
    .A(_08715_),
    .B(_08723_));
 sg13g2_xnor2_1 _17998_ (.Y(_08725_),
    .A(_08712_),
    .B(_08724_));
 sg13g2_inv_1 _17999_ (.Y(_08726_),
    .A(_08537_));
 sg13g2_nand2b_1 _18000_ (.Y(_08727_),
    .B(_08687_),
    .A_N(_08676_));
 sg13g2_o21ai_1 _18001_ (.B1(_08727_),
    .Y(_08728_),
    .A1(_08726_),
    .A2(_08688_));
 sg13g2_inv_1 _18002_ (.Y(_08729_),
    .A(_08728_));
 sg13g2_nor2_1 _18003_ (.A(_08725_),
    .B(_08729_),
    .Y(_08730_));
 sg13g2_nand2_1 _18004_ (.Y(_08731_),
    .A(_08729_),
    .B(_08725_));
 sg13g2_nor2b_1 _18005_ (.A(_08730_),
    .B_N(_08731_),
    .Y(_08732_));
 sg13g2_a21oi_1 _18006_ (.A1(_08674_),
    .A2(_08695_),
    .Y(_08733_),
    .B1(_08694_));
 sg13g2_inv_1 _18007_ (.Y(_08734_),
    .A(_08733_));
 sg13g2_a21oi_1 _18008_ (.A1(_08734_),
    .A2(_08732_),
    .Y(_08735_),
    .B1(net149));
 sg13g2_o21ai_1 _18009_ (.B1(_08735_),
    .Y(_08736_),
    .A1(_08732_),
    .A2(_08734_));
 sg13g2_a22oi_1 _18010_ (.Y(_00403_),
    .B1(_08711_),
    .B2(_08736_),
    .A2(_07532_),
    .A1(_05805_));
 sg13g2_xnor2_1 _18011_ (.Y(_08737_),
    .A(net189),
    .B(_05861_));
 sg13g2_nand2_1 _18012_ (.Y(_08738_),
    .A(_08658_),
    .B(_08705_));
 sg13g2_nor2_1 _18013_ (.A(_08738_),
    .B(_08662_),
    .Y(_08739_));
 sg13g2_o21ai_1 _18014_ (.B1(net189),
    .Y(_08740_),
    .A1(_05770_),
    .A2(\vgadonut.donut.donuthit.rzin[14] ));
 sg13g2_o21ai_1 _18015_ (.B1(_08740_),
    .Y(_08741_),
    .A1(_08668_),
    .A2(_08738_));
 sg13g2_a21oi_1 _18016_ (.A1(_08601_),
    .A2(_08739_),
    .Y(_08742_),
    .B1(_08741_));
 sg13g2_xor2_1 _18017_ (.B(_08742_),
    .A(_08737_),
    .X(_08743_));
 sg13g2_a21oi_1 _18018_ (.A1(_08743_),
    .A2(_07521_),
    .Y(_08744_),
    .B1(_08126_));
 sg13g2_a21oi_1 _18019_ (.A1(_08734_),
    .A2(_08731_),
    .Y(_08745_),
    .B1(_08730_));
 sg13g2_nor2_1 _18020_ (.A(_08684_),
    .B(_08716_),
    .Y(_08746_));
 sg13g2_nor2_1 _18021_ (.A(_06507_),
    .B(_08721_),
    .Y(_08747_));
 sg13g2_a21oi_1 _18022_ (.A1(_08746_),
    .A2(_08721_),
    .Y(_08748_),
    .B1(_08747_));
 sg13g2_o21ai_1 _18023_ (.B1(_08720_),
    .Y(_08749_),
    .A1(_08640_),
    .A2(_08719_));
 sg13g2_xnor2_1 _18024_ (.Y(_08750_),
    .A(\vgadonut.donut.ysA[21] ),
    .B(_05807_));
 sg13g2_xnor2_1 _18025_ (.Y(_08751_),
    .A(_08586_),
    .B(_08750_));
 sg13g2_xnor2_1 _18026_ (.Y(_08752_),
    .A(_08749_),
    .B(_08751_));
 sg13g2_xnor2_1 _18027_ (.Y(_08753_),
    .A(_08748_),
    .B(_08752_));
 sg13g2_nor2_1 _18028_ (.A(_08712_),
    .B(_08724_),
    .Y(_08754_));
 sg13g2_a21oi_1 _18029_ (.A1(_08715_),
    .A2(_08723_),
    .Y(_08755_),
    .B1(_08754_));
 sg13g2_xnor2_1 _18030_ (.Y(_08756_),
    .A(_08753_),
    .B(_08755_));
 sg13g2_o21ai_1 _18031_ (.B1(net148),
    .Y(_08757_),
    .A1(_08756_),
    .A2(_08745_));
 sg13g2_a21o_1 _18032_ (.A2(_08756_),
    .A1(_08745_),
    .B1(_08757_),
    .X(_08758_));
 sg13g2_a22oi_1 _18033_ (.Y(_00404_),
    .B1(_08744_),
    .B2(_08758_),
    .A2(_07532_),
    .A1(_05889_));
 sg13g2_xor2_1 _18034_ (.B(_08341_),
    .A(net217),
    .X(_08759_));
 sg13g2_nor2_1 _18035_ (.A(_08207_),
    .B(_08210_),
    .Y(_08760_));
 sg13g2_o21ai_1 _18036_ (.B1(net162),
    .Y(_08761_),
    .A1(_08760_),
    .A2(_08206_));
 sg13g2_a21oi_1 _18037_ (.A1(_08206_),
    .A2(_08760_),
    .Y(_08762_),
    .B1(_08761_));
 sg13g2_a21oi_1 _18038_ (.A1(net150),
    .A2(_08759_),
    .Y(_08763_),
    .B1(_08762_));
 sg13g2_nor2_1 _18039_ (.A(\vgadonut.donut.rz6[2] ),
    .B(net107),
    .Y(_08764_));
 sg13g2_a21oi_1 _18040_ (.A1(net105),
    .A2(_08763_),
    .Y(_00405_),
    .B1(_08764_));
 sg13g2_nor2b_1 _18041_ (.A(_08213_),
    .B_N(_08212_),
    .Y(_08765_));
 sg13g2_xnor2_1 _18042_ (.Y(_08766_),
    .A(_08765_),
    .B(_08211_));
 sg13g2_nand2b_1 _18043_ (.Y(_08767_),
    .B(_08342_),
    .A_N(_08343_));
 sg13g2_a21oi_1 _18044_ (.A1(_08345_),
    .A2(_08767_),
    .Y(_08768_),
    .B1(net163));
 sg13g2_a21oi_1 _18045_ (.A1(_08766_),
    .A2(net160),
    .Y(_08769_),
    .B1(_08768_));
 sg13g2_nor2_1 _18046_ (.A(\vgadonut.donut.rz6[3] ),
    .B(net107),
    .Y(_08770_));
 sg13g2_a21oi_1 _18047_ (.A1(_08769_),
    .A2(net105),
    .Y(_00406_),
    .B1(_08770_));
 sg13g2_nand2_1 _18048_ (.Y(_08771_),
    .A(_08216_),
    .B(_08217_));
 sg13g2_xnor2_1 _18049_ (.Y(_08772_),
    .A(_08771_),
    .B(_08214_));
 sg13g2_xnor2_1 _18050_ (.Y(_08773_),
    .A(_08344_),
    .B(_08346_));
 sg13g2_nor2_1 _18051_ (.A(net163),
    .B(_08773_),
    .Y(_08774_));
 sg13g2_a21oi_1 _18052_ (.A1(_08772_),
    .A2(net160),
    .Y(_08775_),
    .B1(_08774_));
 sg13g2_nor2_1 _18053_ (.A(\vgadonut.donut.rz6[4] ),
    .B(net107),
    .Y(_08776_));
 sg13g2_a21oi_1 _18054_ (.A1(_08775_),
    .A2(net105),
    .Y(_00407_),
    .B1(_08776_));
 sg13g2_inv_1 _18055_ (.Y(_08777_),
    .A(\vgadonut.donut.rz6[5] ));
 sg13g2_nand2_1 _18056_ (.Y(_08778_),
    .A(_08347_),
    .B(_08336_));
 sg13g2_nor2_1 _18057_ (.A(net162),
    .B(_08349_),
    .Y(_08779_));
 sg13g2_nor2b_1 _18058_ (.A(_08202_),
    .B_N(_08220_),
    .Y(_08780_));
 sg13g2_xnor2_1 _18059_ (.Y(_08781_),
    .A(_08780_),
    .B(_08219_));
 sg13g2_a221oi_1 _18060_ (.B2(net147),
    .C1(net100),
    .B1(_08781_),
    .A1(_08778_),
    .Y(_08782_),
    .A2(_08779_));
 sg13g2_a21oi_1 _18061_ (.A1(_08777_),
    .A2(net93),
    .Y(_00408_),
    .B1(_08782_));
 sg13g2_inv_1 _18062_ (.Y(_08783_),
    .A(\vgadonut.donut.donuthit.rzin[0] ));
 sg13g2_xnor2_1 _18063_ (.Y(_08784_),
    .A(_08226_),
    .B(_08221_));
 sg13g2_a21oi_1 _18064_ (.A1(_08784_),
    .A2(net160),
    .Y(_08785_),
    .B1(net95));
 sg13g2_nand2_1 _18065_ (.Y(_08786_),
    .A(_08351_),
    .B(_08350_));
 sg13g2_nand3b_1 _18066_ (.B(net151),
    .C(_08786_),
    .Y(_08787_),
    .A_N(_08352_));
 sg13g2_a22oi_1 _18067_ (.Y(_00409_),
    .B1(_08785_),
    .B2(_08787_),
    .A2(net91),
    .A1(_08783_));
 sg13g2_inv_1 _18068_ (.Y(_08788_),
    .A(\vgadonut.donut.donuthit.rzin[1] ));
 sg13g2_xnor2_1 _18069_ (.Y(_08789_),
    .A(_08230_),
    .B(_08387_));
 sg13g2_a21oi_1 _18070_ (.A1(_08789_),
    .A2(net147),
    .Y(_08790_),
    .B1(net95));
 sg13g2_nand2b_1 _18071_ (.Y(_08791_),
    .B(_08355_),
    .A_N(_08327_));
 sg13g2_a21oi_1 _18072_ (.A1(_08353_),
    .A2(_08791_),
    .Y(_08792_),
    .B1(net146));
 sg13g2_o21ai_1 _18073_ (.B1(_08792_),
    .Y(_08793_),
    .A1(_08353_),
    .A2(_08791_));
 sg13g2_a22oi_1 _18074_ (.Y(_00410_),
    .B1(_08790_),
    .B2(_08793_),
    .A2(net91),
    .A1(_08788_));
 sg13g2_inv_1 _18075_ (.Y(_08794_),
    .A(\vgadonut.donut.donuthit.rzin[2] ));
 sg13g2_xnor2_1 _18076_ (.Y(_08795_),
    .A(_08237_),
    .B(_08234_));
 sg13g2_a21oi_1 _18077_ (.A1(_08795_),
    .A2(net160),
    .Y(_08796_),
    .B1(net95));
 sg13g2_a21oi_1 _18078_ (.A1(_08356_),
    .A2(_08374_),
    .Y(_08797_),
    .B1(net146));
 sg13g2_o21ai_1 _18079_ (.B1(_08797_),
    .Y(_08798_),
    .A1(_08356_),
    .A2(_08374_));
 sg13g2_a22oi_1 _18080_ (.Y(_00411_),
    .B1(_08796_),
    .B2(_08798_),
    .A2(net91),
    .A1(_08794_));
 sg13g2_inv_1 _18081_ (.Y(_08799_),
    .A(\vgadonut.donut.donuthit.rzin[3] ));
 sg13g2_a21oi_1 _18082_ (.A1(_08357_),
    .A2(_08373_),
    .Y(_08800_),
    .B1(_08371_));
 sg13g2_xor2_1 _18083_ (.B(_08800_),
    .A(_08366_),
    .X(_08801_));
 sg13g2_xnor2_1 _18084_ (.Y(_08802_),
    .A(_08239_),
    .B(_08391_));
 sg13g2_a21oi_1 _18085_ (.A1(_08802_),
    .A2(net163),
    .Y(_08803_),
    .B1(_06989_));
 sg13g2_o21ai_1 _18086_ (.B1(_08803_),
    .Y(_08804_),
    .A1(net147),
    .A2(_08801_));
 sg13g2_o21ai_1 _18087_ (.B1(_08804_),
    .Y(_00412_),
    .A1(_08799_),
    .A2(net104));
 sg13g2_inv_1 _18088_ (.Y(_08805_),
    .A(\vgadonut.donut.sA[0] ));
 sg13g2_xnor2_1 _18089_ (.Y(_08806_),
    .A(_08805_),
    .B(_06393_));
 sg13g2_nand2_1 _18090_ (.Y(_08807_),
    .A(net133),
    .B(_00206_));
 sg13g2_o21ai_1 _18091_ (.B1(_08807_),
    .Y(_00413_),
    .A1(_08806_),
    .A2(net57));
 sg13g2_inv_1 _18092_ (.Y(_08808_),
    .A(_06382_));
 sg13g2_nor2_1 _18093_ (.A(_06288_),
    .B(_08808_),
    .Y(_08809_));
 sg13g2_inv_1 _18094_ (.Y(_08810_),
    .A(_08809_));
 sg13g2_nand2_1 _18095_ (.Y(_08811_),
    .A(_08808_),
    .B(_06288_));
 sg13g2_nand2_1 _18096_ (.Y(_08812_),
    .A(_08810_),
    .B(_08811_));
 sg13g2_nor2_1 _18097_ (.A(net193),
    .B(_06369_),
    .Y(_08813_));
 sg13g2_nand2_1 _18098_ (.Y(_08814_),
    .A(_06369_),
    .B(net193));
 sg13g2_inv_1 _18099_ (.Y(_08815_),
    .A(_08814_));
 sg13g2_nor2_2 _18100_ (.A(_08813_),
    .B(_08815_),
    .Y(_08816_));
 sg13g2_nor2_1 _18101_ (.A(_06255_),
    .B(_06357_),
    .Y(_08817_));
 sg13g2_nor2_1 _18102_ (.A(net223),
    .B(_06358_),
    .Y(_08818_));
 sg13g2_nor2_1 _18103_ (.A(_08817_),
    .B(_08818_),
    .Y(_08819_));
 sg13g2_nand2_1 _18104_ (.Y(_08820_),
    .A(_08816_),
    .B(_08819_));
 sg13g2_buf_1 _18105_ (.A(\vgadonut.donut.sA[4] ),
    .X(_08821_));
 sg13g2_nor2_1 _18106_ (.A(net215),
    .B(_06402_),
    .Y(_08822_));
 sg13g2_inv_1 _18107_ (.Y(_08823_),
    .A(net215));
 sg13g2_nor2b_1 _18108_ (.A(_08823_),
    .B_N(_06402_),
    .Y(_08824_));
 sg13g2_buf_1 _18109_ (.A(_08824_),
    .X(_08825_));
 sg13g2_nor2_1 _18110_ (.A(_08822_),
    .B(_08825_),
    .Y(_08826_));
 sg13g2_inv_1 _18111_ (.Y(_08827_),
    .A(_08826_));
 sg13g2_nor2_1 _18112_ (.A(net198),
    .B(_06305_),
    .Y(_08828_));
 sg13g2_nand2_1 _18113_ (.Y(_08829_),
    .A(_06305_),
    .B(net198));
 sg13g2_inv_1 _18114_ (.Y(_08830_),
    .A(_08829_));
 sg13g2_nor2_2 _18115_ (.A(_08828_),
    .B(_08830_),
    .Y(_08831_));
 sg13g2_inv_1 _18116_ (.Y(_08832_),
    .A(_08831_));
 sg13g2_inv_1 _18117_ (.Y(_08833_),
    .A(_06328_));
 sg13g2_nor2_1 _18118_ (.A(_06263_),
    .B(_08833_),
    .Y(_08834_));
 sg13g2_nand2_1 _18119_ (.Y(_08835_),
    .A(_08833_),
    .B(_06263_));
 sg13g2_nand2b_1 _18120_ (.Y(_08836_),
    .B(_08835_),
    .A_N(_08834_));
 sg13g2_nor2_1 _18121_ (.A(net195),
    .B(_06350_),
    .Y(_08837_));
 sg13g2_nand2_1 _18122_ (.Y(_08838_),
    .A(_06350_),
    .B(net195));
 sg13g2_inv_1 _18123_ (.Y(_08839_),
    .A(_08838_));
 sg13g2_nor3_1 _18124_ (.A(_08836_),
    .B(_08837_),
    .C(_08839_),
    .Y(_08840_));
 sg13g2_inv_1 _18125_ (.Y(_08841_),
    .A(_08840_));
 sg13g2_nor3_1 _18126_ (.A(_08827_),
    .B(_08832_),
    .C(_08841_),
    .Y(_08842_));
 sg13g2_buf_1 _18127_ (.A(\vgadonut.donut.sA[1] ),
    .X(_08843_));
 sg13g2_inv_1 _18128_ (.Y(_08844_),
    .A(_08843_));
 sg13g2_xnor2_1 _18129_ (.Y(_08845_),
    .A(_08844_),
    .B(_06396_));
 sg13g2_nor2b_1 _18130_ (.A(_08805_),
    .B_N(_06393_),
    .Y(_08846_));
 sg13g2_nor2b_1 _18131_ (.A(_08844_),
    .B_N(_06396_),
    .Y(_08847_));
 sg13g2_a21oi_1 _18132_ (.A1(_08845_),
    .A2(_08846_),
    .Y(_08848_),
    .B1(_08847_));
 sg13g2_inv_1 _18133_ (.Y(_08849_),
    .A(_08848_));
 sg13g2_inv_1 _18134_ (.Y(_08850_),
    .A(_06398_));
 sg13g2_buf_1 _18135_ (.A(\vgadonut.donut.sA[2] ),
    .X(_08851_));
 sg13g2_inv_1 _18136_ (.Y(_08852_),
    .A(_08851_));
 sg13g2_nand2_1 _18137_ (.Y(_08853_),
    .A(_08850_),
    .B(_08852_));
 sg13g2_nor2_1 _18138_ (.A(_08852_),
    .B(_08850_),
    .Y(_08854_));
 sg13g2_a21oi_2 _18139_ (.B1(_08854_),
    .Y(_08855_),
    .A2(_08853_),
    .A1(_08849_));
 sg13g2_buf_2 _18140_ (.A(\vgadonut.donut.sA[3] ),
    .X(_08856_));
 sg13g2_nand2_1 _18141_ (.Y(_08857_),
    .A(_06400_),
    .B(_08856_));
 sg13g2_nor2_1 _18142_ (.A(_08856_),
    .B(_06400_),
    .Y(_08858_));
 sg13g2_a21oi_1 _18143_ (.A1(_08855_),
    .A2(_08857_),
    .Y(_08859_),
    .B1(_08858_));
 sg13g2_a21oi_1 _18144_ (.A1(_08831_),
    .A2(_08825_),
    .Y(_08860_),
    .B1(_08830_));
 sg13g2_nor2_1 _18145_ (.A(_08837_),
    .B(_08839_),
    .Y(_08861_));
 sg13g2_a21oi_1 _18146_ (.A1(_08861_),
    .A2(_08834_),
    .Y(_08862_),
    .B1(_08839_));
 sg13g2_o21ai_1 _18147_ (.B1(_08862_),
    .Y(_08863_),
    .A1(_08860_),
    .A2(_08841_));
 sg13g2_a21oi_1 _18148_ (.A1(_08842_),
    .A2(_08859_),
    .Y(_08864_),
    .B1(_08863_));
 sg13g2_a21oi_1 _18149_ (.A1(_08816_),
    .A2(_08817_),
    .Y(_08865_),
    .B1(_08815_));
 sg13g2_o21ai_1 _18150_ (.B1(_08865_),
    .Y(_08866_),
    .A1(_08820_),
    .A2(_08864_));
 sg13g2_xnor2_1 _18151_ (.Y(_08867_),
    .A(_08812_),
    .B(_08866_));
 sg13g2_nand2_1 _18152_ (.Y(_08868_),
    .A(net133),
    .B(_00207_));
 sg13g2_o21ai_1 _18153_ (.B1(_08868_),
    .Y(_00414_),
    .A1(_08867_),
    .A2(net57));
 sg13g2_nor2_1 _18154_ (.A(_06295_),
    .B(_08808_),
    .Y(_08869_));
 sg13g2_inv_1 _18155_ (.Y(_08870_),
    .A(_08869_));
 sg13g2_nor2_1 _18156_ (.A(_06291_),
    .B(_06382_),
    .Y(_08871_));
 sg13g2_inv_1 _18157_ (.Y(_08872_),
    .A(_08871_));
 sg13g2_nand2_1 _18158_ (.Y(_08873_),
    .A(_08870_),
    .B(_08872_));
 sg13g2_nor2_1 _18159_ (.A(_08809_),
    .B(_08815_),
    .Y(_08874_));
 sg13g2_inv_1 _18160_ (.Y(_08875_),
    .A(_08857_));
 sg13g2_a21o_1 _18161_ (.A2(_08875_),
    .A1(_08826_),
    .B1(_08825_),
    .X(_08876_));
 sg13g2_inv_1 _18162_ (.Y(_08877_),
    .A(_08876_));
 sg13g2_nor2_1 _18163_ (.A(_08858_),
    .B(_08875_),
    .Y(_08878_));
 sg13g2_inv_1 _18164_ (.Y(_08879_),
    .A(_08855_));
 sg13g2_nand3_1 _18165_ (.B(_08826_),
    .C(_08879_),
    .A(_08878_),
    .Y(_08880_));
 sg13g2_nand2_1 _18166_ (.Y(_08881_),
    .A(_08877_),
    .B(_08880_));
 sg13g2_a221oi_1 _18167_ (.B2(_08831_),
    .C1(_08830_),
    .B1(_08881_),
    .A1(net194),
    .Y(_08882_),
    .A2(_06328_));
 sg13g2_nor2b_1 _18168_ (.A(_08882_),
    .B_N(_08835_),
    .Y(_08883_));
 sg13g2_nand2_1 _18169_ (.Y(_08884_),
    .A(_08883_),
    .B(_08861_));
 sg13g2_nor2_1 _18170_ (.A(_08817_),
    .B(_08839_),
    .Y(_08885_));
 sg13g2_a21oi_1 _18171_ (.A1(_08884_),
    .A2(_08885_),
    .Y(_08886_),
    .B1(_08818_));
 sg13g2_nand2_1 _18172_ (.Y(_08887_),
    .A(_08886_),
    .B(_08816_));
 sg13g2_a22oi_1 _18173_ (.Y(_08888_),
    .B1(_08874_),
    .B2(_08887_),
    .A2(_08808_),
    .A1(_06288_));
 sg13g2_xnor2_1 _18174_ (.Y(_08889_),
    .A(_08873_),
    .B(_08888_));
 sg13g2_nand2_1 _18175_ (.Y(_08890_),
    .A(net133),
    .B(_00208_));
 sg13g2_o21ai_1 _18176_ (.B1(_08890_),
    .Y(_00415_),
    .A1(_08889_),
    .A2(net57));
 sg13g2_xnor2_1 _18177_ (.Y(_08891_),
    .A(_06249_),
    .B(_06382_));
 sg13g2_nand4_1 _18178_ (.B(_08811_),
    .C(_08810_),
    .A(_08866_),
    .Y(_08892_),
    .D(_08872_));
 sg13g2_nand3_1 _18179_ (.B(_08810_),
    .C(_08870_),
    .A(_08892_),
    .Y(_08893_));
 sg13g2_xnor2_1 _18180_ (.Y(_08894_),
    .A(_08891_),
    .B(_08893_));
 sg13g2_nand2_1 _18181_ (.Y(_08895_),
    .A(net133),
    .B(net224));
 sg13g2_o21ai_1 _18182_ (.B1(_08895_),
    .Y(_00416_),
    .A1(_08894_),
    .A2(net57));
 sg13g2_inv_1 _18183_ (.Y(_08896_),
    .A(net226));
 sg13g2_xnor2_1 _18184_ (.Y(_08897_),
    .A(_08896_),
    .B(_06382_));
 sg13g2_nor2_1 _18185_ (.A(_06249_),
    .B(_08808_),
    .Y(_08898_));
 sg13g2_a21oi_1 _18186_ (.A1(_08888_),
    .A2(_08891_),
    .Y(_08899_),
    .B1(_08898_));
 sg13g2_o21ai_1 _18187_ (.B1(_08870_),
    .Y(_08900_),
    .A1(_08871_),
    .A2(_08899_));
 sg13g2_xor2_1 _18188_ (.B(_08900_),
    .A(_08897_),
    .X(_08901_));
 sg13g2_nand2_1 _18189_ (.Y(_08902_),
    .A(net133),
    .B(_00209_));
 sg13g2_o21ai_1 _18190_ (.B1(_08902_),
    .Y(_00417_),
    .A1(_08901_),
    .A2(net57));
 sg13g2_nor2_1 _18191_ (.A(net196),
    .B(_06382_),
    .Y(_08903_));
 sg13g2_nand2_1 _18192_ (.Y(_08904_),
    .A(_06382_),
    .B(net196));
 sg13g2_nand2b_1 _18193_ (.Y(_08905_),
    .B(_08904_),
    .A_N(_08903_));
 sg13g2_nor2_1 _18194_ (.A(_08896_),
    .B(_08808_),
    .Y(_08906_));
 sg13g2_a21oi_1 _18195_ (.A1(_08900_),
    .A2(_08897_),
    .Y(_08907_),
    .B1(_08906_));
 sg13g2_xnor2_1 _18196_ (.Y(_08908_),
    .A(_08905_),
    .B(_08907_));
 sg13g2_buf_1 _18197_ (.A(_06229_),
    .X(_08909_));
 sg13g2_nand2_1 _18198_ (.Y(_08910_),
    .A(_08909_),
    .B(net196));
 sg13g2_o21ai_1 _18199_ (.B1(_08910_),
    .Y(_00418_),
    .A1(_08908_),
    .A2(net57));
 sg13g2_buf_1 _18200_ (.A(_06371_),
    .X(_08911_));
 sg13g2_buf_1 _18201_ (.A(net188),
    .X(_08912_));
 sg13g2_xnor2_1 _18202_ (.Y(_08913_),
    .A(_08912_),
    .B(_06378_));
 sg13g2_o21ai_1 _18203_ (.B1(_08904_),
    .Y(_08914_),
    .A1(_08903_),
    .A2(_08907_));
 sg13g2_xnor2_1 _18204_ (.Y(_08915_),
    .A(_08913_),
    .B(_08914_));
 sg13g2_buf_1 _18205_ (.A(net192),
    .X(_08916_));
 sg13g2_buf_1 _18206_ (.A(net180),
    .X(_08917_));
 sg13g2_nand2_1 _18207_ (.Y(_08918_),
    .A(_08909_),
    .B(net177));
 sg13g2_o21ai_1 _18208_ (.B1(_08918_),
    .Y(_00419_),
    .A1(_08915_),
    .A2(net57));
 sg13g2_xor2_1 _18209_ (.B(_08845_),
    .A(_08846_),
    .X(_08919_));
 sg13g2_nand2_1 _18210_ (.Y(_08920_),
    .A(net132),
    .B(_00210_));
 sg13g2_o21ai_1 _18211_ (.B1(_08920_),
    .Y(_00420_),
    .A1(_08919_),
    .A2(net57));
 sg13g2_nor2b_1 _18212_ (.A(_08854_),
    .B_N(_08853_),
    .Y(_08921_));
 sg13g2_xnor2_1 _18213_ (.Y(_08922_),
    .A(_08848_),
    .B(_08921_));
 sg13g2_buf_1 _18214_ (.A(net62),
    .X(_08923_));
 sg13g2_nand2_1 _18215_ (.Y(_08924_),
    .A(net132),
    .B(_00211_));
 sg13g2_o21ai_1 _18216_ (.B1(_08924_),
    .Y(_00421_),
    .A1(_08922_),
    .A2(net56));
 sg13g2_xnor2_1 _18217_ (.Y(_08925_),
    .A(_08855_),
    .B(_08878_));
 sg13g2_nand2_1 _18218_ (.Y(_08926_),
    .A(net132),
    .B(_00212_));
 sg13g2_o21ai_1 _18219_ (.B1(_08926_),
    .Y(_00422_),
    .A1(_08925_),
    .A2(net56));
 sg13g2_xnor2_1 _18220_ (.Y(_08927_),
    .A(_08827_),
    .B(_08859_));
 sg13g2_nand2_1 _18221_ (.Y(_08928_),
    .A(net132),
    .B(_00213_));
 sg13g2_o21ai_1 _18222_ (.B1(_08928_),
    .Y(_00423_),
    .A1(_08927_),
    .A2(net56));
 sg13g2_xor2_1 _18223_ (.B(_08881_),
    .A(_08831_),
    .X(_08929_));
 sg13g2_nand2_1 _18224_ (.Y(_08930_),
    .A(net132),
    .B(_00214_));
 sg13g2_o21ai_1 _18225_ (.B1(_08930_),
    .Y(_00424_),
    .A1(_08929_),
    .A2(net56));
 sg13g2_a221oi_1 _18226_ (.B2(_06305_),
    .C1(_08825_),
    .B1(net198),
    .A1(_08859_),
    .Y(_08931_),
    .A2(_08826_));
 sg13g2_nor2_1 _18227_ (.A(_08828_),
    .B(_08931_),
    .Y(_08932_));
 sg13g2_xor2_1 _18228_ (.B(_08932_),
    .A(_08836_),
    .X(_08933_));
 sg13g2_nand2_1 _18229_ (.Y(_08934_),
    .A(net132),
    .B(net194));
 sg13g2_o21ai_1 _18230_ (.B1(_08934_),
    .Y(_00425_),
    .A1(_08933_),
    .A2(net56));
 sg13g2_xnor2_1 _18231_ (.Y(_08935_),
    .A(_08861_),
    .B(_08883_));
 sg13g2_nand2_1 _18232_ (.Y(_08936_),
    .A(net132),
    .B(net195));
 sg13g2_o21ai_1 _18233_ (.B1(_08936_),
    .Y(_00426_),
    .A1(_08935_),
    .A2(net56));
 sg13g2_xnor2_1 _18234_ (.Y(_08937_),
    .A(_08819_),
    .B(_08864_));
 sg13g2_nand2_1 _18235_ (.Y(_08938_),
    .A(net132),
    .B(_00215_));
 sg13g2_o21ai_1 _18236_ (.B1(_08938_),
    .Y(_00427_),
    .A1(_08937_),
    .A2(_08923_));
 sg13g2_xnor2_1 _18237_ (.Y(_08939_),
    .A(_08816_),
    .B(_08886_));
 sg13g2_buf_1 _18238_ (.A(_06229_),
    .X(_08940_));
 sg13g2_nand2_1 _18239_ (.Y(_08941_),
    .A(_08940_),
    .B(net193));
 sg13g2_o21ai_1 _18240_ (.B1(_08941_),
    .Y(_00428_),
    .A1(_08939_),
    .A2(_08923_));
 sg13g2_inv_1 _18241_ (.Y(_08942_),
    .A(_06417_));
 sg13g2_nor2_1 _18242_ (.A(_08942_),
    .B(_06584_),
    .Y(_08943_));
 sg13g2_nand2_1 _18243_ (.Y(_08944_),
    .A(_06584_),
    .B(_08942_));
 sg13g2_nand2b_1 _18244_ (.Y(_08945_),
    .B(_08944_),
    .A_N(_08943_));
 sg13g2_inv_1 _18245_ (.Y(_08946_),
    .A(_07569_));
 sg13g2_inv_1 _18246_ (.Y(_08947_),
    .A(_06603_));
 sg13g2_nor2_1 _18247_ (.A(_08946_),
    .B(_08947_),
    .Y(_08948_));
 sg13g2_inv_1 _18248_ (.Y(_08949_),
    .A(_07571_));
 sg13g2_inv_1 _18249_ (.Y(_08950_),
    .A(_06599_));
 sg13g2_inv_1 _18250_ (.Y(_08951_),
    .A(_07570_));
 sg13g2_inv_1 _18251_ (.Y(_08952_),
    .A(_06587_));
 sg13g2_inv_1 _18252_ (.Y(_08953_),
    .A(_07572_));
 sg13g2_xnor2_1 _18253_ (.Y(_08954_),
    .A(_08953_),
    .B(_06450_));
 sg13g2_nor2_1 _18254_ (.A(_07564_),
    .B(_06803_),
    .Y(_08955_));
 sg13g2_nand2_1 _18255_ (.Y(_08956_),
    .A(_08954_),
    .B(_08955_));
 sg13g2_o21ai_1 _18256_ (.B1(_08956_),
    .Y(_08957_),
    .A1(_08953_),
    .A2(_06775_));
 sg13g2_xnor2_1 _18257_ (.Y(_08958_),
    .A(_08951_),
    .B(_06587_));
 sg13g2_nand2_1 _18258_ (.Y(_08959_),
    .A(_08957_),
    .B(_08958_));
 sg13g2_o21ai_1 _18259_ (.B1(_08959_),
    .Y(_08960_),
    .A1(_08951_),
    .A2(_08952_));
 sg13g2_xnor2_1 _18260_ (.Y(_08961_),
    .A(_08949_),
    .B(_06599_));
 sg13g2_nand2_1 _18261_ (.Y(_08962_),
    .A(_08960_),
    .B(_08961_));
 sg13g2_o21ai_1 _18262_ (.B1(_08962_),
    .Y(_08963_),
    .A1(_08949_),
    .A2(_08950_));
 sg13g2_nand2_1 _18263_ (.Y(_08964_),
    .A(_08947_),
    .B(_08946_));
 sg13g2_o21ai_1 _18264_ (.B1(_08964_),
    .Y(_08965_),
    .A1(_08948_),
    .A2(_08963_));
 sg13g2_inv_1 _18265_ (.Y(_08966_),
    .A(_06420_));
 sg13g2_nor2_1 _18266_ (.A(_08966_),
    .B(_06614_),
    .Y(_08967_));
 sg13g2_inv_1 _18267_ (.Y(_08968_),
    .A(_08967_));
 sg13g2_nor2_1 _18268_ (.A(_06420_),
    .B(_06615_),
    .Y(_08969_));
 sg13g2_a21oi_1 _18269_ (.A1(_08965_),
    .A2(_08968_),
    .Y(_08970_),
    .B1(_08969_));
 sg13g2_xor2_1 _18270_ (.B(_08970_),
    .A(_08945_),
    .X(_08971_));
 sg13g2_xnor2_1 _18271_ (.Y(_08972_),
    .A(_06581_),
    .B(_08971_));
 sg13g2_xnor2_1 _18272_ (.Y(_08973_),
    .A(_04826_),
    .B(_08972_));
 sg13g2_nand2_1 _18273_ (.Y(_08974_),
    .A(net131),
    .B(_00216_));
 sg13g2_o21ai_1 _18274_ (.B1(_08974_),
    .Y(_00429_),
    .A1(_08973_),
    .A2(net56));
 sg13g2_nor2_1 _18275_ (.A(_06442_),
    .B(_06570_),
    .Y(_08975_));
 sg13g2_nor2_1 _18276_ (.A(_06435_),
    .B(_06637_),
    .Y(_08976_));
 sg13g2_o21ai_1 _18277_ (.B1(_08944_),
    .Y(_08977_),
    .A1(_08943_),
    .A2(_08970_));
 sg13g2_inv_1 _18278_ (.Y(_08978_),
    .A(_08977_));
 sg13g2_nor2_1 _18279_ (.A(_06414_),
    .B(_06628_),
    .Y(_08979_));
 sg13g2_inv_1 _18280_ (.Y(_08980_),
    .A(_08979_));
 sg13g2_nor2_1 _18281_ (.A(_07722_),
    .B(_06626_),
    .Y(_08981_));
 sg13g2_a21oi_1 _18282_ (.A1(_08978_),
    .A2(_08980_),
    .Y(_08982_),
    .B1(_08981_));
 sg13g2_inv_1 _18283_ (.Y(_08983_),
    .A(_08982_));
 sg13g2_nor2_1 _18284_ (.A(_06428_),
    .B(_06575_),
    .Y(_08984_));
 sg13g2_inv_1 _18285_ (.Y(_08985_),
    .A(_08984_));
 sg13g2_nor2_1 _18286_ (.A(_07723_),
    .B(_06578_),
    .Y(_08986_));
 sg13g2_a21oi_1 _18287_ (.A1(_08983_),
    .A2(_08985_),
    .Y(_08987_),
    .B1(_08986_));
 sg13g2_xnor2_1 _18288_ (.Y(_08988_),
    .A(_06434_),
    .B(_06637_));
 sg13g2_nor2b_1 _18289_ (.A(_08987_),
    .B_N(_08988_),
    .Y(_08989_));
 sg13g2_nor2_1 _18290_ (.A(_08976_),
    .B(_08989_),
    .Y(_08990_));
 sg13g2_nand2_1 _18291_ (.Y(_08991_),
    .A(_06570_),
    .B(_06442_));
 sg13g2_o21ai_1 _18292_ (.B1(_08991_),
    .Y(_08992_),
    .A1(_08975_),
    .A2(_08990_));
 sg13g2_xnor2_1 _18293_ (.Y(_08993_),
    .A(_06525_),
    .B(_06566_));
 sg13g2_xnor2_1 _18294_ (.Y(_08994_),
    .A(_06406_),
    .B(_06566_));
 sg13g2_nand3_1 _18295_ (.B(_08993_),
    .C(_08994_),
    .A(_08992_),
    .Y(_08995_));
 sg13g2_xnor2_1 _18296_ (.Y(_08996_),
    .A(_06518_),
    .B(net75));
 sg13g2_xnor2_1 _18297_ (.Y(_08997_),
    .A(_06533_),
    .B(_06566_));
 sg13g2_nand3b_1 _18298_ (.B(_08996_),
    .C(_08997_),
    .Y(_08998_),
    .A_N(_08995_));
 sg13g2_nand3_1 _18299_ (.B(net74),
    .C(_07947_),
    .A(_08998_),
    .Y(_08999_));
 sg13g2_o21ai_1 _18300_ (.B1(_08999_),
    .Y(_09000_),
    .A1(net74),
    .A2(_08998_));
 sg13g2_xnor2_1 _18301_ (.Y(_09001_),
    .A(net191),
    .B(_09000_));
 sg13g2_buf_1 _18302_ (.A(_09001_),
    .X(_09002_));
 sg13g2_xnor2_1 _18303_ (.Y(_09003_),
    .A(net207),
    .B(_06703_));
 sg13g2_inv_1 _18304_ (.Y(_09004_),
    .A(_04958_));
 sg13g2_nor2_1 _18305_ (.A(_09004_),
    .B(_06703_),
    .Y(_09005_));
 sg13g2_a21oi_1 _18306_ (.A1(_09002_),
    .A2(_09003_),
    .Y(_09006_),
    .B1(_09005_));
 sg13g2_xnor2_1 _18307_ (.Y(_09007_),
    .A(net240),
    .B(_06721_));
 sg13g2_xnor2_1 _18308_ (.Y(_09008_),
    .A(_09007_),
    .B(_09002_));
 sg13g2_nor2_1 _18309_ (.A(_09006_),
    .B(_09008_),
    .Y(_09009_));
 sg13g2_inv_1 _18310_ (.Y(_09010_),
    .A(_09009_));
 sg13g2_nand2_1 _18311_ (.Y(_09011_),
    .A(_09008_),
    .B(_09006_));
 sg13g2_nand2_1 _18312_ (.Y(_09012_),
    .A(_09010_),
    .B(_09011_));
 sg13g2_nand2_1 _18313_ (.Y(_09013_),
    .A(_08997_),
    .B(_08993_));
 sg13g2_nand2b_1 _18314_ (.Y(_09014_),
    .B(_08991_),
    .A_N(_08975_));
 sg13g2_nor2_1 _18315_ (.A(_09014_),
    .B(_08990_),
    .Y(_09015_));
 sg13g2_nand2_1 _18316_ (.Y(_09016_),
    .A(_09015_),
    .B(_08994_));
 sg13g2_nand2_1 _18317_ (.Y(_09017_),
    .A(net74),
    .B(_07914_));
 sg13g2_o21ai_1 _18318_ (.B1(_09017_),
    .Y(_09018_),
    .A1(_09013_),
    .A2(_09016_));
 sg13g2_xnor2_1 _18319_ (.Y(_09019_),
    .A(_08996_),
    .B(_09018_));
 sg13g2_inv_1 _18320_ (.Y(_09020_),
    .A(net241));
 sg13g2_xnor2_1 _18321_ (.Y(_09021_),
    .A(_09020_),
    .B(_06687_));
 sg13g2_nor2_1 _18322_ (.A(_09020_),
    .B(_06688_),
    .Y(_09022_));
 sg13g2_a21oi_1 _18323_ (.A1(_09019_),
    .A2(_09021_),
    .Y(_09023_),
    .B1(_09022_));
 sg13g2_xnor2_1 _18324_ (.Y(_09024_),
    .A(_09003_),
    .B(_09002_));
 sg13g2_nor2_1 _18325_ (.A(_09023_),
    .B(_09024_),
    .Y(_09025_));
 sg13g2_o21ai_1 _18326_ (.B1(_08995_),
    .Y(_09026_),
    .A1(net75),
    .A2(_07913_));
 sg13g2_xnor2_1 _18327_ (.Y(_09027_),
    .A(_08997_),
    .B(_09026_));
 sg13g2_inv_1 _18328_ (.Y(_09028_),
    .A(net242));
 sg13g2_xnor2_1 _18329_ (.Y(_09029_),
    .A(_09028_),
    .B(_06673_));
 sg13g2_nor2_1 _18330_ (.A(_09028_),
    .B(_06675_),
    .Y(_09030_));
 sg13g2_a21oi_1 _18331_ (.A1(_09027_),
    .A2(_09029_),
    .Y(_09031_),
    .B1(_09030_));
 sg13g2_xnor2_1 _18332_ (.Y(_09032_),
    .A(_09021_),
    .B(_09019_));
 sg13g2_xnor2_1 _18333_ (.Y(_09033_),
    .A(_09032_),
    .B(_09031_));
 sg13g2_inv_1 _18334_ (.Y(_09034_),
    .A(net244));
 sg13g2_o21ai_1 _18335_ (.B1(net74),
    .Y(_09035_),
    .A1(_06442_),
    .A2(_06406_));
 sg13g2_nand2_1 _18336_ (.Y(_09036_),
    .A(_09016_),
    .B(_09035_));
 sg13g2_xnor2_1 _18337_ (.Y(_09037_),
    .A(_08993_),
    .B(_09036_));
 sg13g2_xnor2_1 _18338_ (.Y(_09038_),
    .A(_09034_),
    .B(_06658_));
 sg13g2_nand2_1 _18339_ (.Y(_09039_),
    .A(_09037_),
    .B(_09038_));
 sg13g2_o21ai_1 _18340_ (.B1(_09039_),
    .Y(_09040_),
    .A1(_09034_),
    .A2(_06660_));
 sg13g2_buf_1 _18341_ (.A(_09040_),
    .X(_09041_));
 sg13g2_xor2_1 _18342_ (.B(_09027_),
    .A(_09029_),
    .X(_09042_));
 sg13g2_nor2_1 _18343_ (.A(_09041_),
    .B(_09042_),
    .Y(_09043_));
 sg13g2_xor2_1 _18344_ (.B(_08990_),
    .A(_09014_),
    .X(_09044_));
 sg13g2_inv_1 _18345_ (.Y(_09045_),
    .A(_09044_));
 sg13g2_inv_1 _18346_ (.Y(_09046_),
    .A(_04815_));
 sg13g2_xnor2_1 _18347_ (.Y(_09047_),
    .A(_09046_),
    .B(_06645_));
 sg13g2_nor2_1 _18348_ (.A(_09046_),
    .B(_06647_),
    .Y(_09048_));
 sg13g2_a21oi_2 _18349_ (.B1(_09048_),
    .Y(_09049_),
    .A2(_09047_),
    .A1(_09045_));
 sg13g2_inv_1 _18350_ (.Y(_09050_),
    .A(net243));
 sg13g2_xnor2_1 _18351_ (.Y(_09051_),
    .A(_09050_),
    .B(_06504_));
 sg13g2_xor2_1 _18352_ (.B(_08992_),
    .A(_08994_),
    .X(_09052_));
 sg13g2_xor2_1 _18353_ (.B(_09052_),
    .A(_09051_),
    .X(_09053_));
 sg13g2_inv_1 _18354_ (.Y(_09054_),
    .A(_04823_));
 sg13g2_nand2b_1 _18355_ (.Y(_09055_),
    .B(_08985_),
    .A_N(_08986_));
 sg13g2_xor2_1 _18356_ (.B(_08982_),
    .A(_09055_),
    .X(_09056_));
 sg13g2_inv_1 _18357_ (.Y(_09057_),
    .A(_09056_));
 sg13g2_xnor2_1 _18358_ (.Y(_09058_),
    .A(_04823_),
    .B(_06577_));
 sg13g2_nand2_1 _18359_ (.Y(_09059_),
    .A(_09057_),
    .B(_09058_));
 sg13g2_o21ai_1 _18360_ (.B1(_09059_),
    .Y(_09060_),
    .A1(_09054_),
    .A2(_06577_));
 sg13g2_inv_1 _18361_ (.Y(_09061_),
    .A(_04820_));
 sg13g2_xnor2_1 _18362_ (.Y(_09062_),
    .A(_09061_),
    .B(_06633_));
 sg13g2_xnor2_1 _18363_ (.Y(_09063_),
    .A(_08988_),
    .B(_08987_));
 sg13g2_xor2_1 _18364_ (.B(_09063_),
    .A(_09062_),
    .X(_09064_));
 sg13g2_xnor2_1 _18365_ (.Y(_09065_),
    .A(_09060_),
    .B(_09064_));
 sg13g2_xor2_1 _18366_ (.B(_09056_),
    .A(_09058_),
    .X(_09066_));
 sg13g2_inv_1 _18367_ (.Y(_09067_),
    .A(_04824_));
 sg13g2_nor2_1 _18368_ (.A(_08981_),
    .B(_08979_),
    .Y(_09068_));
 sg13g2_xor2_1 _18369_ (.B(_08977_),
    .A(_09068_),
    .X(_09069_));
 sg13g2_xnor2_1 _18370_ (.Y(_09070_),
    .A(_04824_),
    .B(_06623_));
 sg13g2_nand2_1 _18371_ (.Y(_09071_),
    .A(_09069_),
    .B(_09070_));
 sg13g2_o21ai_1 _18372_ (.B1(_09071_),
    .Y(_09072_),
    .A1(_09067_),
    .A2(_06623_));
 sg13g2_nor2b_1 _18373_ (.A(_09066_),
    .B_N(_09072_),
    .Y(_09073_));
 sg13g2_nor2b_1 _18374_ (.A(_09064_),
    .B_N(_09060_),
    .Y(_09074_));
 sg13g2_a21oi_1 _18375_ (.A1(_09065_),
    .A2(_09073_),
    .Y(_09075_),
    .B1(_09074_));
 sg13g2_xnor2_1 _18376_ (.Y(_09076_),
    .A(_09070_),
    .B(_09069_));
 sg13g2_nand2b_1 _18377_ (.Y(_09077_),
    .B(_06581_),
    .A_N(_08971_));
 sg13g2_nor2b_1 _18378_ (.A(_09076_),
    .B_N(_09077_),
    .Y(_09078_));
 sg13g2_xnor2_1 _18379_ (.Y(_09079_),
    .A(_09077_),
    .B(_09076_));
 sg13g2_nor2b_1 _18380_ (.A(_08972_),
    .B_N(_04826_),
    .Y(_09080_));
 sg13g2_nand2_1 _18381_ (.Y(_09081_),
    .A(_09079_),
    .B(_09080_));
 sg13g2_inv_1 _18382_ (.Y(_09082_),
    .A(_09081_));
 sg13g2_nor2_1 _18383_ (.A(_09078_),
    .B(_09082_),
    .Y(_09083_));
 sg13g2_inv_1 _18384_ (.Y(_09084_),
    .A(_09083_));
 sg13g2_xnor2_1 _18385_ (.Y(_09085_),
    .A(_09072_),
    .B(_09066_));
 sg13g2_nand3_1 _18386_ (.B(_09084_),
    .C(_09085_),
    .A(_09065_),
    .Y(_09086_));
 sg13g2_nand2_1 _18387_ (.Y(_09087_),
    .A(_09075_),
    .B(_09086_));
 sg13g2_inv_1 _18388_ (.Y(_09088_),
    .A(_09063_));
 sg13g2_nor2_1 _18389_ (.A(_09061_),
    .B(_06634_),
    .Y(_09089_));
 sg13g2_a21oi_1 _18390_ (.A1(_09088_),
    .A2(_09062_),
    .Y(_09090_),
    .B1(_09089_));
 sg13g2_xor2_1 _18391_ (.B(_09044_),
    .A(_09047_),
    .X(_09091_));
 sg13g2_nor2_1 _18392_ (.A(_09090_),
    .B(_09091_),
    .Y(_09092_));
 sg13g2_nand2_1 _18393_ (.Y(_09093_),
    .A(_09091_),
    .B(_09090_));
 sg13g2_nor2b_1 _18394_ (.A(_09092_),
    .B_N(_09093_),
    .Y(_09094_));
 sg13g2_nand2_1 _18395_ (.Y(_09095_),
    .A(_09087_),
    .B(_09094_));
 sg13g2_nor2_1 _18396_ (.A(_09049_),
    .B(_09053_),
    .Y(_09096_));
 sg13g2_nor2_1 _18397_ (.A(_09092_),
    .B(_09096_),
    .Y(_09097_));
 sg13g2_a22oi_1 _18398_ (.Y(_09098_),
    .B1(_09095_),
    .B2(_09097_),
    .A2(_09053_),
    .A1(_09049_));
 sg13g2_xnor2_1 _18399_ (.Y(_09099_),
    .A(_09038_),
    .B(_09037_));
 sg13g2_inv_1 _18400_ (.Y(_09100_),
    .A(_09052_));
 sg13g2_nor2_1 _18401_ (.A(_09050_),
    .B(_06569_),
    .Y(_09101_));
 sg13g2_a21oi_1 _18402_ (.A1(_09100_),
    .A2(_09051_),
    .Y(_09102_),
    .B1(_09101_));
 sg13g2_nand2_1 _18403_ (.Y(_09103_),
    .A(_09099_),
    .B(_09102_));
 sg13g2_nor2_1 _18404_ (.A(_09102_),
    .B(_09099_),
    .Y(_09104_));
 sg13g2_a221oi_1 _18405_ (.B2(_09103_),
    .C1(_09104_),
    .B1(_09098_),
    .A1(_09041_),
    .Y(_09105_),
    .A2(_09042_));
 sg13g2_nor2_1 _18406_ (.A(_09043_),
    .B(_09105_),
    .Y(_09106_));
 sg13g2_nand2b_1 _18407_ (.Y(_09107_),
    .B(_09106_),
    .A_N(_09033_));
 sg13g2_o21ai_1 _18408_ (.B1(_09107_),
    .Y(_09108_),
    .A1(_09031_),
    .A2(_09032_));
 sg13g2_buf_1 _18409_ (.A(_09108_),
    .X(_09109_));
 sg13g2_nand2_1 _18410_ (.Y(_09110_),
    .A(_09024_),
    .B(_09023_));
 sg13g2_o21ai_1 _18411_ (.B1(_09110_),
    .Y(_09111_),
    .A1(_09025_),
    .A2(_09109_));
 sg13g2_xor2_1 _18412_ (.B(_09111_),
    .A(_09012_),
    .X(_09112_));
 sg13g2_nand2_1 _18413_ (.Y(_09113_),
    .A(net131),
    .B(_00217_));
 sg13g2_o21ai_1 _18414_ (.B1(_09113_),
    .Y(_00430_),
    .A1(net65),
    .A2(_09112_));
 sg13g2_xnor2_1 _18415_ (.Y(_09114_),
    .A(net239),
    .B(net77));
 sg13g2_buf_1 _18416_ (.A(_09002_),
    .X(_09115_));
 sg13g2_xnor2_1 _18417_ (.Y(_09116_),
    .A(_09114_),
    .B(net69));
 sg13g2_nand2_1 _18418_ (.Y(_09117_),
    .A(net69),
    .B(_09007_));
 sg13g2_o21ai_1 _18419_ (.B1(_09117_),
    .Y(_09118_),
    .A1(_06478_),
    .A2(net77));
 sg13g2_inv_1 _18420_ (.Y(_09119_),
    .A(_09118_));
 sg13g2_nor2_1 _18421_ (.A(_09116_),
    .B(_09119_),
    .Y(_09120_));
 sg13g2_inv_1 _18422_ (.Y(_09121_),
    .A(_09120_));
 sg13g2_nand2_1 _18423_ (.Y(_09122_),
    .A(_09119_),
    .B(_09116_));
 sg13g2_nand2_1 _18424_ (.Y(_09123_),
    .A(_09121_),
    .B(_09122_));
 sg13g2_nor2_1 _18425_ (.A(_09025_),
    .B(_09009_),
    .Y(_09124_));
 sg13g2_nor2b_1 _18426_ (.A(_09025_),
    .B_N(_09110_),
    .Y(_09125_));
 sg13g2_nand2_1 _18427_ (.Y(_09126_),
    .A(_09109_),
    .B(_09125_));
 sg13g2_a22oi_1 _18428_ (.Y(_09127_),
    .B1(_09124_),
    .B2(_09126_),
    .A2(_09008_),
    .A1(_09006_));
 sg13g2_xnor2_1 _18429_ (.Y(_09128_),
    .A(_09123_),
    .B(_09127_));
 sg13g2_nand2_1 _18430_ (.Y(_09129_),
    .A(net131),
    .B(_00218_));
 sg13g2_o21ai_1 _18431_ (.B1(_09129_),
    .Y(_00431_),
    .A1(net65),
    .A2(_09128_));
 sg13g2_buf_1 _18432_ (.A(net166),
    .X(_09130_));
 sg13g2_xnor2_1 _18433_ (.Y(_09131_),
    .A(net238),
    .B(_06722_));
 sg13g2_xnor2_1 _18434_ (.Y(_09132_),
    .A(_09131_),
    .B(net69));
 sg13g2_nand2_1 _18435_ (.Y(_09133_),
    .A(net69),
    .B(_09114_));
 sg13g2_o21ai_1 _18436_ (.B1(_09133_),
    .Y(_09134_),
    .A1(_06485_),
    .A2(net77));
 sg13g2_xor2_1 _18437_ (.B(_09134_),
    .A(_09132_),
    .X(_09135_));
 sg13g2_nor2_1 _18438_ (.A(_09012_),
    .B(_09111_),
    .Y(_09136_));
 sg13g2_nor3_1 _18439_ (.A(_09009_),
    .B(_09120_),
    .C(_09136_),
    .Y(_09137_));
 sg13g2_nor2b_1 _18440_ (.A(_09137_),
    .B_N(_09122_),
    .Y(_09138_));
 sg13g2_xnor2_1 _18441_ (.Y(_09139_),
    .A(_09135_),
    .B(_09138_));
 sg13g2_nand2_1 _18442_ (.Y(_09140_),
    .A(_09139_),
    .B(net66));
 sg13g2_o21ai_1 _18443_ (.B1(_09140_),
    .Y(_00432_),
    .A1(_06488_),
    .A2(net145));
 sg13g2_xnor2_1 _18444_ (.Y(_09141_),
    .A(net206),
    .B(net77));
 sg13g2_xor2_1 _18445_ (.B(net69),
    .A(_09141_),
    .X(_09142_));
 sg13g2_nand2_1 _18446_ (.Y(_09143_),
    .A(net69),
    .B(_09131_));
 sg13g2_o21ai_1 _18447_ (.B1(_09143_),
    .Y(_09144_),
    .A1(_06488_),
    .A2(net77));
 sg13g2_buf_1 _18448_ (.A(_09144_),
    .X(_09145_));
 sg13g2_or2_1 _18449_ (.X(_09146_),
    .B(_09145_),
    .A(_09142_));
 sg13g2_nand2_1 _18450_ (.Y(_09147_),
    .A(_09145_),
    .B(_09142_));
 sg13g2_nand2_1 _18451_ (.Y(_09148_),
    .A(_09146_),
    .B(_09147_));
 sg13g2_inv_1 _18452_ (.Y(_09149_),
    .A(_09134_));
 sg13g2_nor2_1 _18453_ (.A(_09132_),
    .B(_09149_),
    .Y(_09150_));
 sg13g2_nor2_1 _18454_ (.A(_09120_),
    .B(_09150_),
    .Y(_09151_));
 sg13g2_inv_1 _18455_ (.Y(_09152_),
    .A(_09123_));
 sg13g2_nand2_1 _18456_ (.Y(_09153_),
    .A(_09127_),
    .B(_09152_));
 sg13g2_a22oi_1 _18457_ (.Y(_09154_),
    .B1(_09151_),
    .B2(_09153_),
    .A2(_09132_),
    .A1(_09149_));
 sg13g2_xnor2_1 _18458_ (.Y(_09155_),
    .A(_09148_),
    .B(_09154_));
 sg13g2_nand2_1 _18459_ (.Y(_09156_),
    .A(_08940_),
    .B(_00219_));
 sg13g2_o21ai_1 _18460_ (.B1(_09156_),
    .Y(_00433_),
    .A1(net65),
    .A2(_09155_));
 sg13g2_xnor2_1 _18461_ (.Y(_09157_),
    .A(net205),
    .B(net77));
 sg13g2_xnor2_1 _18462_ (.Y(_09158_),
    .A(_09157_),
    .B(net69));
 sg13g2_inv_1 _18463_ (.Y(_09159_),
    .A(_09158_));
 sg13g2_nand2_1 _18464_ (.Y(_09160_),
    .A(net69),
    .B(_09141_));
 sg13g2_o21ai_1 _18465_ (.B1(_09160_),
    .Y(_09161_),
    .A1(_06496_),
    .A2(net77));
 sg13g2_buf_1 _18466_ (.A(_09161_),
    .X(_09162_));
 sg13g2_xnor2_1 _18467_ (.Y(_09163_),
    .A(_09159_),
    .B(_09162_));
 sg13g2_inv_1 _18468_ (.Y(_09164_),
    .A(_09135_));
 sg13g2_a221oi_1 _18469_ (.B2(_09164_),
    .C1(_09150_),
    .B1(_09138_),
    .A1(_09145_),
    .Y(_09165_),
    .A2(_09142_));
 sg13g2_nor2b_1 _18470_ (.A(_09165_),
    .B_N(_09146_),
    .Y(_09166_));
 sg13g2_xor2_1 _18471_ (.B(_09166_),
    .A(_09163_),
    .X(_09167_));
 sg13g2_nand2_1 _18472_ (.Y(_09168_),
    .A(net131),
    .B(net205));
 sg13g2_o21ai_1 _18473_ (.B1(_09168_),
    .Y(_00434_),
    .A1(net65),
    .A2(_09167_));
 sg13g2_nand2b_1 _18474_ (.Y(_09169_),
    .B(_09154_),
    .A_N(_09148_));
 sg13g2_a22oi_1 _18475_ (.Y(_09170_),
    .B1(_09162_),
    .B2(_09159_),
    .A2(_09142_),
    .A1(_09145_));
 sg13g2_nor2_1 _18476_ (.A(_09159_),
    .B(_09162_),
    .Y(_09171_));
 sg13g2_a21oi_1 _18477_ (.A1(_09169_),
    .A2(_09170_),
    .Y(_09172_),
    .B1(_09171_));
 sg13g2_inv_1 _18478_ (.Y(_09173_),
    .A(_05134_));
 sg13g2_o21ai_1 _18479_ (.B1(_09115_),
    .Y(_09174_),
    .A1(_09173_),
    .A2(_06723_));
 sg13g2_o21ai_1 _18480_ (.B1(_09174_),
    .Y(_09175_),
    .A1(net205),
    .A2(_06722_));
 sg13g2_xnor2_1 _18481_ (.Y(_09176_),
    .A(net204),
    .B(_09175_));
 sg13g2_nand2b_1 _18482_ (.Y(_09177_),
    .B(_09176_),
    .A_N(_09172_));
 sg13g2_nand2b_1 _18483_ (.Y(_09178_),
    .B(_09172_),
    .A_N(_09176_));
 sg13g2_nand2_1 _18484_ (.Y(_09179_),
    .A(_09177_),
    .B(_09178_));
 sg13g2_buf_1 _18485_ (.A(_09179_),
    .X(_09180_));
 sg13g2_nand2_1 _18486_ (.Y(_09181_),
    .A(net131),
    .B(net204));
 sg13g2_o21ai_1 _18487_ (.B1(_09181_),
    .Y(_00435_),
    .A1(net65),
    .A2(_09180_));
 sg13g2_xor2_1 _18488_ (.B(_09079_),
    .A(_09080_),
    .X(_09182_));
 sg13g2_nand2_1 _18489_ (.Y(_09183_),
    .A(net131),
    .B(_00220_));
 sg13g2_o21ai_1 _18490_ (.B1(_09183_),
    .Y(_00436_),
    .A1(_09182_),
    .A2(net56));
 sg13g2_xnor2_1 _18491_ (.Y(_09184_),
    .A(_09083_),
    .B(_09085_));
 sg13g2_buf_1 _18492_ (.A(net62),
    .X(_09185_));
 sg13g2_nand2_1 _18493_ (.Y(_09186_),
    .A(net131),
    .B(_00221_));
 sg13g2_o21ai_1 _18494_ (.B1(_09186_),
    .Y(_00437_),
    .A1(_09184_),
    .A2(net55));
 sg13g2_a21oi_1 _18495_ (.A1(_09084_),
    .A2(_09085_),
    .Y(_09187_),
    .B1(_09073_));
 sg13g2_xnor2_1 _18496_ (.Y(_09188_),
    .A(_09065_),
    .B(_09187_));
 sg13g2_nand2_1 _18497_ (.Y(_09189_),
    .A(net131),
    .B(_00222_));
 sg13g2_o21ai_1 _18498_ (.B1(_09189_),
    .Y(_00438_),
    .A1(_09188_),
    .A2(net55));
 sg13g2_xor2_1 _18499_ (.B(_09087_),
    .A(_09094_),
    .X(_09190_));
 sg13g2_buf_1 _18500_ (.A(_06229_),
    .X(_09191_));
 sg13g2_nand2_1 _18501_ (.Y(_09192_),
    .A(net130),
    .B(_00223_));
 sg13g2_o21ai_1 _18502_ (.B1(_09192_),
    .Y(_00439_),
    .A1(_09190_),
    .A2(net55));
 sg13g2_xor2_1 _18503_ (.B(_09053_),
    .A(_09049_),
    .X(_09193_));
 sg13g2_a21o_1 _18504_ (.A2(_09093_),
    .A1(_09087_),
    .B1(_09092_),
    .X(_09194_));
 sg13g2_xor2_1 _18505_ (.B(_09194_),
    .A(_09193_),
    .X(_09195_));
 sg13g2_nand2_1 _18506_ (.Y(_09196_),
    .A(net130),
    .B(_00224_));
 sg13g2_o21ai_1 _18507_ (.B1(_09196_),
    .Y(_00440_),
    .A1(_09195_),
    .A2(net55));
 sg13g2_nor2b_1 _18508_ (.A(_09104_),
    .B_N(_09103_),
    .Y(_09197_));
 sg13g2_xor2_1 _18509_ (.B(_09098_),
    .A(_09197_),
    .X(_09198_));
 sg13g2_nand2_1 _18510_ (.Y(_09199_),
    .A(net66),
    .B(_09198_));
 sg13g2_o21ai_1 _18511_ (.B1(_09199_),
    .Y(_00441_),
    .A1(_09034_),
    .A2(_09130_));
 sg13g2_xnor2_1 _18512_ (.Y(_09200_),
    .A(_09041_),
    .B(_09042_));
 sg13g2_nor2_1 _18513_ (.A(_09096_),
    .B(_09104_),
    .Y(_09201_));
 sg13g2_nand2_1 _18514_ (.Y(_09202_),
    .A(_09194_),
    .B(_09193_));
 sg13g2_a22oi_1 _18515_ (.Y(_09203_),
    .B1(_09201_),
    .B2(_09202_),
    .A2(_09099_),
    .A1(_09102_));
 sg13g2_xnor2_1 _18516_ (.Y(_09204_),
    .A(_09200_),
    .B(_09203_));
 sg13g2_nand2_1 _18517_ (.Y(_09205_),
    .A(_09204_),
    .B(net66));
 sg13g2_o21ai_1 _18518_ (.B1(_09205_),
    .Y(_00442_),
    .A1(_09028_),
    .A2(net145));
 sg13g2_xnor2_1 _18519_ (.Y(_09206_),
    .A(_09033_),
    .B(_09106_));
 sg13g2_nand2_1 _18520_ (.Y(_09207_),
    .A(net130),
    .B(_00225_));
 sg13g2_o21ai_1 _18521_ (.B1(_09207_),
    .Y(_00443_),
    .A1(net65),
    .A2(_09206_));
 sg13g2_xor2_1 _18522_ (.B(_09109_),
    .A(_09125_),
    .X(_09208_));
 sg13g2_nand2_1 _18523_ (.Y(_09209_),
    .A(_09208_),
    .B(net66));
 sg13g2_o21ai_1 _18524_ (.B1(_09209_),
    .Y(_00444_),
    .A1(_09004_),
    .A2(net145));
 sg13g2_xnor2_1 _18525_ (.Y(_09210_),
    .A(_07564_),
    .B(_06802_));
 sg13g2_xnor2_1 _18526_ (.Y(_09211_),
    .A(_09210_),
    .B(_09198_));
 sg13g2_nand2_1 _18527_ (.Y(_09212_),
    .A(net130),
    .B(_07562_));
 sg13g2_o21ai_1 _18528_ (.B1(_09212_),
    .Y(_00445_),
    .A1(_06227_),
    .A2(_09211_));
 sg13g2_xnor2_1 _18529_ (.Y(_09213_),
    .A(_09044_),
    .B(net54));
 sg13g2_inv_1 _18530_ (.Y(_09214_),
    .A(_09213_));
 sg13g2_inv_1 _18531_ (.Y(_09215_),
    .A(_09179_));
 sg13g2_xnor2_1 _18532_ (.Y(_09216_),
    .A(_09063_),
    .B(_09179_));
 sg13g2_inv_1 _18533_ (.Y(_09217_),
    .A(_09216_));
 sg13g2_nor2_1 _18534_ (.A(_09057_),
    .B(_09167_),
    .Y(_09218_));
 sg13g2_nor2b_1 _18535_ (.A(_09056_),
    .B_N(_09167_),
    .Y(_09219_));
 sg13g2_inv_1 _18536_ (.Y(_09220_),
    .A(_09139_));
 sg13g2_xnor2_1 _18537_ (.Y(_09221_),
    .A(_08961_),
    .B(_08960_));
 sg13g2_inv_1 _18538_ (.Y(_09222_),
    .A(_09208_));
 sg13g2_nor2_1 _18539_ (.A(_09221_),
    .B(_09222_),
    .Y(_09223_));
 sg13g2_xor2_1 _18540_ (.B(_09208_),
    .A(_09221_),
    .X(_09224_));
 sg13g2_xor2_1 _18541_ (.B(_08957_),
    .A(_08958_),
    .X(_09225_));
 sg13g2_xor2_1 _18542_ (.B(_09206_),
    .A(_09225_),
    .X(_09226_));
 sg13g2_inv_1 _18543_ (.Y(_09227_),
    .A(_09226_));
 sg13g2_xor2_1 _18544_ (.B(_08954_),
    .A(_08955_),
    .X(_09228_));
 sg13g2_and2_1 _18545_ (.A(_09198_),
    .B(_09210_),
    .X(_09229_));
 sg13g2_inv_1 _18546_ (.Y(_09230_),
    .A(_09229_));
 sg13g2_xnor2_1 _18547_ (.Y(_09231_),
    .A(_09228_),
    .B(_09204_));
 sg13g2_nor2_1 _18548_ (.A(_09230_),
    .B(_09231_),
    .Y(_09232_));
 sg13g2_a21o_1 _18549_ (.A2(_09228_),
    .A1(_09204_),
    .B1(_09232_),
    .X(_09233_));
 sg13g2_inv_1 _18550_ (.Y(_09234_),
    .A(_09233_));
 sg13g2_nor2_1 _18551_ (.A(_09227_),
    .B(_09234_),
    .Y(_09235_));
 sg13g2_a21o_1 _18552_ (.A2(_09225_),
    .A1(_09206_),
    .B1(_09235_),
    .X(_09236_));
 sg13g2_inv_1 _18553_ (.Y(_09237_),
    .A(_09236_));
 sg13g2_nor2_1 _18554_ (.A(_09224_),
    .B(_09237_),
    .Y(_09238_));
 sg13g2_nand2b_1 _18555_ (.Y(_09239_),
    .B(_08964_),
    .A_N(_08948_));
 sg13g2_xnor2_1 _18556_ (.Y(_09240_),
    .A(_09239_),
    .B(_08963_));
 sg13g2_xor2_1 _18557_ (.B(_09112_),
    .A(_09240_),
    .X(_09241_));
 sg13g2_o21ai_1 _18558_ (.B1(_09241_),
    .Y(_09242_),
    .A1(_09223_),
    .A2(_09238_));
 sg13g2_nand2_1 _18559_ (.Y(_09243_),
    .A(_09112_),
    .B(_09240_));
 sg13g2_nand2_1 _18560_ (.Y(_09244_),
    .A(_09242_),
    .B(_09243_));
 sg13g2_nor2_1 _18561_ (.A(_08967_),
    .B(_08969_),
    .Y(_09245_));
 sg13g2_xor2_1 _18562_ (.B(_08965_),
    .A(_09245_),
    .X(_09246_));
 sg13g2_xnor2_1 _18563_ (.Y(_09247_),
    .A(_09246_),
    .B(_09128_));
 sg13g2_nor2b_1 _18564_ (.A(_09246_),
    .B_N(_09128_),
    .Y(_09248_));
 sg13g2_a21oi_1 _18565_ (.A1(_09244_),
    .A2(_09247_),
    .Y(_09249_),
    .B1(_09248_));
 sg13g2_xnor2_1 _18566_ (.Y(_09250_),
    .A(_08971_),
    .B(_09139_));
 sg13g2_nand2b_1 _18567_ (.Y(_09251_),
    .B(_09250_),
    .A_N(_09249_));
 sg13g2_o21ai_1 _18568_ (.B1(_09251_),
    .Y(_09252_),
    .A1(_08971_),
    .A2(_09220_));
 sg13g2_buf_1 _18569_ (.A(_09252_),
    .X(_09253_));
 sg13g2_xnor2_1 _18570_ (.Y(_09254_),
    .A(_09069_),
    .B(_09155_));
 sg13g2_nor2b_1 _18571_ (.A(_09069_),
    .B_N(_09155_),
    .Y(_09255_));
 sg13g2_a21oi_1 _18572_ (.A1(_09253_),
    .A2(_09254_),
    .Y(_09256_),
    .B1(_09255_));
 sg13g2_nor2_1 _18573_ (.A(_09219_),
    .B(_09256_),
    .Y(_09257_));
 sg13g2_nor2_1 _18574_ (.A(_09218_),
    .B(_09257_),
    .Y(_09258_));
 sg13g2_nor2_1 _18575_ (.A(_09217_),
    .B(_09258_),
    .Y(_09259_));
 sg13g2_a21oi_1 _18576_ (.A1(_09063_),
    .A2(_09215_),
    .Y(_09260_),
    .B1(_09259_));
 sg13g2_nor2_1 _18577_ (.A(_09214_),
    .B(_09260_),
    .Y(_09261_));
 sg13g2_nand2_1 _18578_ (.Y(_09262_),
    .A(_09260_),
    .B(_09214_));
 sg13g2_nand3b_1 _18579_ (.B(net67),
    .C(_09262_),
    .Y(_09263_),
    .A_N(_09261_));
 sg13g2_o21ai_1 _18580_ (.B1(_09263_),
    .Y(_00446_),
    .A1(_06443_),
    .A2(net145));
 sg13g2_nor2_1 _18581_ (.A(_09100_),
    .B(net54),
    .Y(_09264_));
 sg13g2_inv_1 _18582_ (.Y(_09265_),
    .A(_09264_));
 sg13g2_nand2_1 _18583_ (.Y(_09266_),
    .A(net54),
    .B(_09100_));
 sg13g2_a21oi_1 _18584_ (.A1(_09044_),
    .A2(_09215_),
    .Y(_09267_),
    .B1(_09261_));
 sg13g2_inv_1 _18585_ (.Y(_09268_),
    .A(_09267_));
 sg13g2_a21oi_1 _18586_ (.A1(_09265_),
    .A2(_09266_),
    .Y(_09269_),
    .B1(_09268_));
 sg13g2_nand2_1 _18587_ (.Y(_09270_),
    .A(_09268_),
    .B(_09266_));
 sg13g2_o21ai_1 _18588_ (.B1(net67),
    .Y(_09271_),
    .A1(_09264_),
    .A2(_09270_));
 sg13g2_nand2_1 _18589_ (.Y(_09272_),
    .A(net130),
    .B(_06406_));
 sg13g2_o21ai_1 _18590_ (.B1(_09272_),
    .Y(_00447_),
    .A1(_09269_),
    .A2(_09271_));
 sg13g2_inv_1 _18591_ (.Y(_09273_),
    .A(_09270_));
 sg13g2_nor2_1 _18592_ (.A(_09264_),
    .B(_09273_),
    .Y(_09274_));
 sg13g2_nor2_1 _18593_ (.A(_09037_),
    .B(net54),
    .Y(_09275_));
 sg13g2_nor2b_1 _18594_ (.A(_09215_),
    .B_N(_09037_),
    .Y(_09276_));
 sg13g2_nor2_1 _18595_ (.A(_09275_),
    .B(_09276_),
    .Y(_09277_));
 sg13g2_nor2b_1 _18596_ (.A(_09274_),
    .B_N(_09277_),
    .Y(_09278_));
 sg13g2_nand2b_1 _18597_ (.Y(_09279_),
    .B(_09274_),
    .A_N(_09277_));
 sg13g2_nand3b_1 _18598_ (.B(net67),
    .C(_09279_),
    .Y(_09280_),
    .A_N(_09278_));
 sg13g2_o21ai_1 _18599_ (.B1(_09280_),
    .Y(_00448_),
    .A1(_06529_),
    .A2(_09130_));
 sg13g2_xor2_1 _18600_ (.B(net54),
    .A(_09027_),
    .X(_09281_));
 sg13g2_inv_1 _18601_ (.Y(_09282_),
    .A(_09275_));
 sg13g2_o21ai_1 _18602_ (.B1(_09282_),
    .Y(_09283_),
    .A1(_09276_),
    .A2(_09274_));
 sg13g2_and2_1 _18603_ (.A(_09283_),
    .B(_09281_),
    .X(_09284_));
 sg13g2_nor2_1 _18604_ (.A(net62),
    .B(_09284_),
    .Y(_09285_));
 sg13g2_o21ai_1 _18605_ (.B1(_09285_),
    .Y(_09286_),
    .A1(_09281_),
    .A2(_09283_));
 sg13g2_o21ai_1 _18606_ (.B1(_09286_),
    .Y(_00449_),
    .A1(_06538_),
    .A2(net145));
 sg13g2_nor2_1 _18607_ (.A(_09027_),
    .B(net54),
    .Y(_09287_));
 sg13g2_a21oi_1 _18608_ (.A1(_09278_),
    .A2(_09281_),
    .Y(_09288_),
    .B1(_09275_));
 sg13g2_nand2b_1 _18609_ (.Y(_09289_),
    .B(_09288_),
    .A_N(_09287_));
 sg13g2_xor2_1 _18610_ (.B(net54),
    .A(_09019_),
    .X(_09290_));
 sg13g2_a21oi_1 _18611_ (.A1(_09289_),
    .A2(_09290_),
    .Y(_09291_),
    .B1(_06226_));
 sg13g2_o21ai_1 _18612_ (.B1(_09291_),
    .Y(_09292_),
    .A1(_09289_),
    .A2(_09290_));
 sg13g2_o21ai_1 _18613_ (.B1(_09292_),
    .Y(_00450_),
    .A1(_06541_),
    .A2(net145));
 sg13g2_a21oi_1 _18614_ (.A1(_09284_),
    .A2(_09290_),
    .Y(_09293_),
    .B1(_09287_));
 sg13g2_o21ai_1 _18615_ (.B1(_09293_),
    .Y(_09294_),
    .A1(_09019_),
    .A2(net54));
 sg13g2_xnor2_1 _18616_ (.Y(_09295_),
    .A(_09115_),
    .B(_09180_));
 sg13g2_nand2b_1 _18617_ (.Y(_09296_),
    .B(_09295_),
    .A_N(_09294_));
 sg13g2_nand2b_1 _18618_ (.Y(_09297_),
    .B(_09294_),
    .A_N(_09295_));
 sg13g2_nand3_1 _18619_ (.B(net66),
    .C(_09297_),
    .A(_09296_),
    .Y(_09298_));
 sg13g2_o21ai_1 _18620_ (.B1(_09298_),
    .Y(_00451_),
    .A1(_06517_),
    .A2(net145));
 sg13g2_nand2_1 _18621_ (.Y(_09299_),
    .A(_09231_),
    .B(_09230_));
 sg13g2_nand3b_1 _18622_ (.B(_06344_),
    .C(_09299_),
    .Y(_09300_),
    .A_N(_09232_));
 sg13g2_o21ai_1 _18623_ (.B1(_09300_),
    .Y(_00452_),
    .A1(_08953_),
    .A2(net145));
 sg13g2_nor2_1 _18624_ (.A(net62),
    .B(_09235_),
    .Y(_09301_));
 sg13g2_o21ai_1 _18625_ (.B1(_09301_),
    .Y(_09302_),
    .A1(_09226_),
    .A2(_09233_));
 sg13g2_o21ai_1 _18626_ (.B1(_09302_),
    .Y(_00453_),
    .A1(_08951_),
    .A2(net166));
 sg13g2_a21oi_1 _18627_ (.A1(_09237_),
    .A2(_09224_),
    .Y(_09303_),
    .B1(net62));
 sg13g2_nand2b_1 _18628_ (.Y(_09304_),
    .B(_09303_),
    .A_N(_09238_));
 sg13g2_o21ai_1 _18629_ (.B1(_09304_),
    .Y(_00454_),
    .A1(_08949_),
    .A2(net166));
 sg13g2_nor3_1 _18630_ (.A(_09241_),
    .B(_09223_),
    .C(_09238_),
    .Y(_09305_));
 sg13g2_nand3b_1 _18631_ (.B(_09242_),
    .C(net67),
    .Y(_09306_),
    .A_N(_09305_));
 sg13g2_o21ai_1 _18632_ (.B1(_09306_),
    .Y(_00455_),
    .A1(_08946_),
    .A2(net166));
 sg13g2_o21ai_1 _18633_ (.B1(_06225_),
    .Y(_09307_),
    .A1(_09247_),
    .A2(_09244_));
 sg13g2_a21oi_1 _18634_ (.A1(_09247_),
    .A2(_09244_),
    .Y(_09308_),
    .B1(_09307_));
 sg13g2_a21o_1 _18635_ (.A2(net136),
    .A1(_06420_),
    .B1(_09308_),
    .X(_00456_));
 sg13g2_nand2b_1 _18636_ (.Y(_09309_),
    .B(_09249_),
    .A_N(_09250_));
 sg13g2_nand3_1 _18637_ (.B(net66),
    .C(_09309_),
    .A(_09251_),
    .Y(_09310_));
 sg13g2_o21ai_1 _18638_ (.B1(_09310_),
    .Y(_00457_),
    .A1(_08942_),
    .A2(net166));
 sg13g2_o21ai_1 _18639_ (.B1(_06225_),
    .Y(_09311_),
    .A1(_09254_),
    .A2(_09253_));
 sg13g2_a21oi_1 _18640_ (.A1(_09254_),
    .A2(_09253_),
    .Y(_09312_),
    .B1(_09311_));
 sg13g2_a21o_1 _18641_ (.A2(net136),
    .A1(_06414_),
    .B1(_09312_),
    .X(_00458_));
 sg13g2_nor2_1 _18642_ (.A(_09218_),
    .B(_09219_),
    .Y(_09313_));
 sg13g2_nand2b_1 _18643_ (.Y(_09314_),
    .B(_09313_),
    .A_N(_09256_));
 sg13g2_nand2b_1 _18644_ (.Y(_09315_),
    .B(_09256_),
    .A_N(_09313_));
 sg13g2_nand3_1 _18645_ (.B(net66),
    .C(_09315_),
    .A(_09314_),
    .Y(_09316_));
 sg13g2_o21ai_1 _18646_ (.B1(_09316_),
    .Y(_00459_),
    .A1(_07723_),
    .A2(net166));
 sg13g2_nand2_1 _18647_ (.Y(_09317_),
    .A(_09258_),
    .B(_09217_));
 sg13g2_nand3b_1 _18648_ (.B(net67),
    .C(_09317_),
    .Y(_09318_),
    .A_N(_09259_));
 sg13g2_o21ai_1 _18649_ (.B1(_09318_),
    .Y(_00460_),
    .A1(_06435_),
    .A2(net166));
 sg13g2_xnor2_1 _18650_ (.Y(_09319_),
    .A(_06151_),
    .B(_06152_));
 sg13g2_nand2_1 _18651_ (.Y(_09320_),
    .A(net130),
    .B(_04208_));
 sg13g2_o21ai_1 _18652_ (.B1(_09320_),
    .Y(_00461_),
    .A1(_09319_),
    .A2(net55));
 sg13g2_xor2_1 _18653_ (.B(_06194_),
    .A(_06195_),
    .X(_09321_));
 sg13g2_nand2_1 _18654_ (.Y(_09322_),
    .A(net130),
    .B(net211));
 sg13g2_o21ai_1 _18655_ (.B1(_09322_),
    .Y(_00462_),
    .A1(_09321_),
    .A2(net55));
 sg13g2_xnor2_1 _18656_ (.Y(_09323_),
    .A(_06198_),
    .B(_06197_));
 sg13g2_nand2_1 _18657_ (.Y(_09324_),
    .A(net130),
    .B(net247));
 sg13g2_o21ai_1 _18658_ (.B1(_09324_),
    .Y(_00463_),
    .A1(_09323_),
    .A2(net55));
 sg13g2_nand2b_1 _18659_ (.Y(_09325_),
    .B(_06199_),
    .A_N(_06201_));
 sg13g2_xnor2_1 _18660_ (.Y(_09326_),
    .A(_06122_),
    .B(_09325_));
 sg13g2_nand2_1 _18661_ (.Y(_09327_),
    .A(_09191_),
    .B(net210));
 sg13g2_o21ai_1 _18662_ (.B1(_09327_),
    .Y(_00464_),
    .A1(_09326_),
    .A2(net55));
 sg13g2_xnor2_1 _18663_ (.Y(_09328_),
    .A(_06208_),
    .B(_06205_));
 sg13g2_nand2_1 _18664_ (.Y(_09329_),
    .A(_09191_),
    .B(net209));
 sg13g2_o21ai_1 _18665_ (.B1(_09329_),
    .Y(_00465_),
    .A1(_09328_),
    .A2(_09185_));
 sg13g2_nand3_1 _18666_ (.B(_06208_),
    .C(_06122_),
    .A(_09325_),
    .Y(_09330_));
 sg13g2_o21ai_1 _18667_ (.B1(_09330_),
    .Y(_09331_),
    .A1(_06115_),
    .A2(net76));
 sg13g2_a21oi_1 _18668_ (.A1(_06208_),
    .A2(_06203_),
    .Y(_09332_),
    .B1(_09331_));
 sg13g2_xor2_1 _18669_ (.B(_09332_),
    .A(_06207_),
    .X(_09333_));
 sg13g2_buf_1 _18670_ (.A(_06223_),
    .X(_09334_));
 sg13g2_nand2_1 _18671_ (.Y(_09335_),
    .A(net140),
    .B(net246));
 sg13g2_o21ai_1 _18672_ (.B1(_09335_),
    .Y(_00466_),
    .A1(_09333_),
    .A2(_09185_));
 sg13g2_nor2_1 _18673_ (.A(_04603_),
    .B(_06222_),
    .Y(_09336_));
 sg13g2_a21oi_1 _18674_ (.A1(_06211_),
    .A2(_06222_),
    .Y(_00467_),
    .B1(_09336_));
 sg13g2_xnor2_1 _18675_ (.Y(_09337_),
    .A(_06153_),
    .B(_06150_));
 sg13g2_nand2_1 _18676_ (.Y(_09338_),
    .A(net140),
    .B(_04206_));
 sg13g2_o21ai_1 _18677_ (.B1(_09338_),
    .Y(_00468_),
    .A1(_09337_),
    .A2(net58));
 sg13g2_xnor2_1 _18678_ (.Y(_09339_),
    .A(_06156_),
    .B(_06158_));
 sg13g2_nand2_1 _18679_ (.Y(_09340_),
    .A(net140),
    .B(_04205_));
 sg13g2_o21ai_1 _18680_ (.B1(_09340_),
    .Y(_00469_),
    .A1(_09339_),
    .A2(net58));
 sg13g2_xnor2_1 _18681_ (.Y(_09341_),
    .A(_06135_),
    .B(_06159_));
 sg13g2_nand2_1 _18682_ (.Y(_09342_),
    .A(net140),
    .B(_04202_));
 sg13g2_o21ai_1 _18683_ (.B1(_09342_),
    .Y(_00470_),
    .A1(_09341_),
    .A2(_06868_));
 sg13g2_xnor2_1 _18684_ (.Y(_09343_),
    .A(_06170_),
    .B(_06161_));
 sg13g2_nand2_1 _18685_ (.Y(_09344_),
    .A(net140),
    .B(net252));
 sg13g2_o21ai_1 _18686_ (.B1(_09344_),
    .Y(_00471_),
    .A1(_09343_),
    .A2(net58));
 sg13g2_xor2_1 _18687_ (.B(_06174_),
    .A(_06177_),
    .X(_09345_));
 sg13g2_nand2_1 _18688_ (.Y(_09346_),
    .A(_09334_),
    .B(_04203_));
 sg13g2_o21ai_1 _18689_ (.B1(_09346_),
    .Y(_00472_),
    .A1(_09345_),
    .A2(net58));
 sg13g2_xor2_1 _18690_ (.B(_06180_),
    .A(_06183_),
    .X(_09347_));
 sg13g2_nand2_1 _18691_ (.Y(_09348_),
    .A(net140),
    .B(net251));
 sg13g2_o21ai_1 _18692_ (.B1(_09348_),
    .Y(_00473_),
    .A1(_09347_),
    .A2(net58));
 sg13g2_xor2_1 _18693_ (.B(_06185_),
    .A(_06131_),
    .X(_09349_));
 sg13g2_nand2_1 _18694_ (.Y(_09350_),
    .A(net140),
    .B(net248));
 sg13g2_o21ai_1 _18695_ (.B1(_09350_),
    .Y(_00474_),
    .A1(_09349_),
    .A2(net58));
 sg13g2_xnor2_1 _18696_ (.Y(_09351_),
    .A(_06128_),
    .B(_06187_));
 sg13g2_nand2_1 _18697_ (.Y(_09352_),
    .A(net140),
    .B(_04312_));
 sg13g2_o21ai_1 _18698_ (.B1(_09352_),
    .Y(_00475_),
    .A1(_09351_),
    .A2(net58));
 sg13g2_xor2_1 _18699_ (.B(_06189_),
    .A(_06191_),
    .X(_09353_));
 sg13g2_nand2_1 _18700_ (.Y(_09354_),
    .A(_09334_),
    .B(net212));
 sg13g2_o21ai_1 _18701_ (.B1(_09354_),
    .Y(_00476_),
    .A1(_09353_),
    .A2(net58));
 sg13g2_inv_2 _18702_ (.Y(_09355_),
    .A(_06973_));
 sg13g2_buf_1 _18703_ (.A(_09355_),
    .X(_09356_));
 sg13g2_nand2_1 _18704_ (.Y(_09357_),
    .A(\vgadonut.donut.ycA[0] ),
    .B(_06260_));
 sg13g2_nand2_1 _18705_ (.Y(_09358_),
    .A(net159),
    .B(_09357_));
 sg13g2_inv_1 _18706_ (.Y(_09359_),
    .A(_06260_));
 sg13g2_nor2_1 _18707_ (.A(_09359_),
    .B(_06976_),
    .Y(_09360_));
 sg13g2_inv_1 _18708_ (.Y(_09361_),
    .A(_09360_));
 sg13g2_a22oi_1 _18709_ (.Y(_00477_),
    .B1(_07561_),
    .B2(_09361_),
    .A2(_06975_),
    .A1(_09358_));
 sg13g2_nor2_1 _18710_ (.A(_10004_),
    .B(_06334_),
    .Y(_09362_));
 sg13g2_buf_1 _18711_ (.A(_09362_),
    .X(_09363_));
 sg13g2_buf_1 _18712_ (.A(_09363_),
    .X(_09364_));
 sg13g2_buf_1 _18713_ (.A(_06340_),
    .X(_09365_));
 sg13g2_nor2_1 _18714_ (.A(_06245_),
    .B(_06277_),
    .Y(_09366_));
 sg13g2_nor2_1 _18715_ (.A(_06276_),
    .B(_06301_),
    .Y(_09367_));
 sg13g2_inv_1 _18716_ (.Y(_09368_),
    .A(_09367_));
 sg13g2_nand2b_1 _18717_ (.Y(_09369_),
    .B(_09368_),
    .A_N(_09366_));
 sg13g2_nor2_1 _18718_ (.A(_06292_),
    .B(_09359_),
    .Y(_09370_));
 sg13g2_xnor2_1 _18719_ (.Y(_09371_),
    .A(_06252_),
    .B(net225));
 sg13g2_nor2b_1 _18720_ (.A(_09370_),
    .B_N(_09371_),
    .Y(_09372_));
 sg13g2_a21oi_1 _18721_ (.A1(_06253_),
    .A2(net225),
    .Y(_09373_),
    .B1(_09372_));
 sg13g2_xnor2_1 _18722_ (.Y(_09374_),
    .A(_09369_),
    .B(_09373_));
 sg13g2_nor2_1 _18723_ (.A(_07627_),
    .B(_06330_),
    .Y(_09375_));
 sg13g2_nand2_1 _18724_ (.Y(_09376_),
    .A(_07627_),
    .B(_06330_));
 sg13g2_nor2b_1 _18725_ (.A(_09375_),
    .B_N(_09376_),
    .Y(_09377_));
 sg13g2_nor2_1 _18726_ (.A(_07589_),
    .B(net227),
    .Y(_09378_));
 sg13g2_nand2_1 _18727_ (.Y(_09379_),
    .A(_07589_),
    .B(net227));
 sg13g2_nand2b_1 _18728_ (.Y(_09380_),
    .B(_09379_),
    .A_N(_09378_));
 sg13g2_nor2_1 _18729_ (.A(_07642_),
    .B(_06245_),
    .Y(_09381_));
 sg13g2_nand2_1 _18730_ (.Y(_09382_),
    .A(_07642_),
    .B(_06245_));
 sg13g2_nand2b_1 _18731_ (.Y(_09383_),
    .B(_09382_),
    .A_N(_09381_));
 sg13g2_nor2_1 _18732_ (.A(_07669_),
    .B(net225),
    .Y(_09384_));
 sg13g2_nor2_1 _18733_ (.A(_07681_),
    .B(_06284_),
    .Y(_09385_));
 sg13g2_xor2_1 _18734_ (.B(_06252_),
    .A(_08083_),
    .X(_09386_));
 sg13g2_inv_1 _18735_ (.Y(_09387_),
    .A(_09386_));
 sg13g2_nand2_1 _18736_ (.Y(_09388_),
    .A(_08083_),
    .B(_06252_));
 sg13g2_o21ai_1 _18737_ (.B1(_09388_),
    .Y(_09389_),
    .A1(_09357_),
    .A2(_09387_));
 sg13g2_nor2_1 _18738_ (.A(_07680_),
    .B(_06276_),
    .Y(_09390_));
 sg13g2_nand2_1 _18739_ (.Y(_09391_),
    .A(_07680_),
    .B(_06276_));
 sg13g2_inv_1 _18740_ (.Y(_09392_),
    .A(_09391_));
 sg13g2_nor2_1 _18741_ (.A(_09390_),
    .B(_09392_),
    .Y(_09393_));
 sg13g2_nand2_1 _18742_ (.Y(_09394_),
    .A(_07681_),
    .B(_06284_));
 sg13g2_nand2_1 _18743_ (.Y(_09395_),
    .A(_09394_),
    .B(_09391_));
 sg13g2_a21oi_1 _18744_ (.A1(_09389_),
    .A2(_09393_),
    .Y(_09396_),
    .B1(_09395_));
 sg13g2_nor2_1 _18745_ (.A(_09385_),
    .B(_09396_),
    .Y(_09397_));
 sg13g2_xor2_1 _18746_ (.B(_06292_),
    .A(_07663_),
    .X(_09398_));
 sg13g2_nand2_1 _18747_ (.Y(_09399_),
    .A(_09397_),
    .B(_09398_));
 sg13g2_nand2_1 _18748_ (.Y(_09400_),
    .A(_07669_),
    .B(net225));
 sg13g2_nand2_1 _18749_ (.Y(_09401_),
    .A(_07663_),
    .B(_06292_));
 sg13g2_nand3_1 _18750_ (.B(_09400_),
    .C(_09401_),
    .A(_09399_),
    .Y(_09402_));
 sg13g2_nor2b_1 _18751_ (.A(_09384_),
    .B_N(_09402_),
    .Y(_09403_));
 sg13g2_nand2b_1 _18752_ (.Y(_09404_),
    .B(_09403_),
    .A_N(_09383_));
 sg13g2_nand2_1 _18753_ (.Y(_09405_),
    .A(_07581_),
    .B(_06235_));
 sg13g2_nand2_1 _18754_ (.Y(_09406_),
    .A(_09382_),
    .B(_09405_));
 sg13g2_inv_1 _18755_ (.Y(_09407_),
    .A(_09406_));
 sg13g2_nor2_1 _18756_ (.A(_07581_),
    .B(_06235_),
    .Y(_09408_));
 sg13g2_a21oi_1 _18757_ (.A1(_09404_),
    .A2(_09407_),
    .Y(_09409_),
    .B1(_09408_));
 sg13g2_nand2b_1 _18758_ (.Y(_09410_),
    .B(_09409_),
    .A_N(_09380_));
 sg13g2_nand2_1 _18759_ (.Y(_09411_),
    .A(_07601_),
    .B(net220));
 sg13g2_nand2_1 _18760_ (.Y(_09412_),
    .A(_09379_),
    .B(_09411_));
 sg13g2_inv_1 _18761_ (.Y(_09413_),
    .A(_09412_));
 sg13g2_nor2_1 _18762_ (.A(_07601_),
    .B(net220),
    .Y(_09414_));
 sg13g2_a21oi_1 _18763_ (.A1(_09410_),
    .A2(_09413_),
    .Y(_09415_),
    .B1(_09414_));
 sg13g2_buf_1 _18764_ (.A(_06973_),
    .X(_09416_));
 sg13g2_a21oi_1 _18765_ (.A1(_09415_),
    .A2(_09377_),
    .Y(_09417_),
    .B1(net168));
 sg13g2_o21ai_1 _18766_ (.B1(_09417_),
    .Y(_09418_),
    .A1(_09377_),
    .A2(_09415_));
 sg13g2_o21ai_1 _18767_ (.B1(_09418_),
    .Y(_09419_),
    .A1(net169),
    .A2(_09374_));
 sg13g2_buf_1 _18768_ (.A(_09363_),
    .X(_09420_));
 sg13g2_nand2_1 _18769_ (.Y(_09421_),
    .A(_09419_),
    .B(net143));
 sg13g2_o21ai_1 _18770_ (.B1(_09421_),
    .Y(_00478_),
    .A1(_07787_),
    .A2(net144));
 sg13g2_buf_1 _18771_ (.A(_06976_),
    .X(_09422_));
 sg13g2_buf_1 _18772_ (.A(net129),
    .X(_09423_));
 sg13g2_buf_1 _18773_ (.A(_06976_),
    .X(_09424_));
 sg13g2_nor2_1 _18774_ (.A(_06284_),
    .B(_06240_),
    .Y(_09425_));
 sg13g2_inv_1 _18775_ (.Y(_09426_),
    .A(_09425_));
 sg13g2_nor2_1 _18776_ (.A(_06235_),
    .B(_06285_),
    .Y(_09427_));
 sg13g2_inv_1 _18777_ (.Y(_09428_),
    .A(_09427_));
 sg13g2_o21ai_1 _18778_ (.B1(_09368_),
    .Y(_09429_),
    .A1(_09366_),
    .A2(_09373_));
 sg13g2_a21oi_1 _18779_ (.A1(_09426_),
    .A2(_09428_),
    .Y(_09430_),
    .B1(_09429_));
 sg13g2_nand2_1 _18780_ (.Y(_09431_),
    .A(_09429_),
    .B(_09428_));
 sg13g2_nor2_1 _18781_ (.A(_09425_),
    .B(_09431_),
    .Y(_09432_));
 sg13g2_nor3_1 _18782_ (.A(net159),
    .B(_09430_),
    .C(_09432_),
    .Y(_09433_));
 sg13g2_nor2_1 _18783_ (.A(_09424_),
    .B(_09433_),
    .Y(_09434_));
 sg13g2_nor2_1 _18784_ (.A(_07790_),
    .B(net219),
    .Y(_09435_));
 sg13g2_nand2_1 _18785_ (.Y(_09436_),
    .A(_07790_),
    .B(net219));
 sg13g2_nor2b_1 _18786_ (.A(_09435_),
    .B_N(_09436_),
    .Y(_09437_));
 sg13g2_nand2_1 _18787_ (.Y(_09438_),
    .A(_09401_),
    .B(_09394_));
 sg13g2_inv_1 _18788_ (.Y(_09439_),
    .A(_09438_));
 sg13g2_inv_1 _18789_ (.Y(_09440_),
    .A(_09390_));
 sg13g2_a21oi_1 _18790_ (.A1(_09389_),
    .A2(_09440_),
    .Y(_09441_),
    .B1(_09392_));
 sg13g2_nor2b_1 _18791_ (.A(_09385_),
    .B_N(_09394_),
    .Y(_09442_));
 sg13g2_nand2b_1 _18792_ (.Y(_09443_),
    .B(_09442_),
    .A_N(_09441_));
 sg13g2_a22oi_1 _18793_ (.Y(_09444_),
    .B1(_09439_),
    .B2(_09443_),
    .A2(_06293_),
    .A1(_07664_));
 sg13g2_nor2b_1 _18794_ (.A(_09384_),
    .B_N(_09400_),
    .Y(_09445_));
 sg13g2_nand2_1 _18795_ (.Y(_09446_),
    .A(_09382_),
    .B(_09400_));
 sg13g2_a21oi_1 _18796_ (.A1(_09444_),
    .A2(_09445_),
    .Y(_09447_),
    .B1(_09446_));
 sg13g2_a21oi_1 _18797_ (.A1(_07643_),
    .A2(_06301_),
    .Y(_09448_),
    .B1(_09447_));
 sg13g2_nor2b_1 _18798_ (.A(_09408_),
    .B_N(_09405_),
    .Y(_09449_));
 sg13g2_nand2_1 _18799_ (.Y(_09450_),
    .A(_09448_),
    .B(_09449_));
 sg13g2_nand2_1 _18800_ (.Y(_09451_),
    .A(_09379_),
    .B(_09405_));
 sg13g2_inv_1 _18801_ (.Y(_09452_),
    .A(_09451_));
 sg13g2_a21oi_1 _18802_ (.A1(_09450_),
    .A2(_09452_),
    .Y(_09453_),
    .B1(_09378_));
 sg13g2_nor2b_1 _18803_ (.A(_09414_),
    .B_N(_09411_),
    .Y(_09454_));
 sg13g2_nand2_1 _18804_ (.Y(_09455_),
    .A(_09376_),
    .B(_09411_));
 sg13g2_a21oi_1 _18805_ (.A1(_09453_),
    .A2(_09454_),
    .Y(_09456_),
    .B1(_09455_));
 sg13g2_nor2_1 _18806_ (.A(_09375_),
    .B(_09456_),
    .Y(_09457_));
 sg13g2_buf_1 _18807_ (.A(net168),
    .X(_09458_));
 sg13g2_a21oi_1 _18808_ (.A1(_09457_),
    .A2(_09437_),
    .Y(_09459_),
    .B1(net158));
 sg13g2_o21ai_1 _18809_ (.B1(_09459_),
    .Y(_09460_),
    .A1(_09437_),
    .A2(_09457_));
 sg13g2_a22oi_1 _18810_ (.Y(_00479_),
    .B1(_09434_),
    .B2(_09460_),
    .A2(net114),
    .A1(_07822_));
 sg13g2_nor2_1 _18811_ (.A(_06233_),
    .B(_06293_),
    .Y(_09461_));
 sg13g2_nor2_1 _18812_ (.A(_06292_),
    .B(_06311_),
    .Y(_09462_));
 sg13g2_inv_1 _18813_ (.Y(_09463_),
    .A(_09462_));
 sg13g2_nand2b_1 _18814_ (.Y(_09464_),
    .B(_09463_),
    .A_N(_09461_));
 sg13g2_nand2_1 _18815_ (.Y(_09465_),
    .A(_09431_),
    .B(_09426_));
 sg13g2_xor2_1 _18816_ (.B(_09465_),
    .A(_09464_),
    .X(_09466_));
 sg13g2_nor2_1 _18817_ (.A(_07825_),
    .B(net218),
    .Y(_09467_));
 sg13g2_nand2_1 _18818_ (.Y(_09468_),
    .A(_07825_),
    .B(net218));
 sg13g2_nor2b_1 _18819_ (.A(_09467_),
    .B_N(_09468_),
    .Y(_09469_));
 sg13g2_nand2_1 _18820_ (.Y(_09470_),
    .A(_09376_),
    .B(_09436_));
 sg13g2_a21oi_1 _18821_ (.A1(_09415_),
    .A2(_09377_),
    .Y(_09471_),
    .B1(_09470_));
 sg13g2_nor2_1 _18822_ (.A(_09435_),
    .B(_09471_),
    .Y(_09472_));
 sg13g2_a21oi_1 _18823_ (.A1(_09472_),
    .A2(_09469_),
    .Y(_09473_),
    .B1(_09416_));
 sg13g2_o21ai_1 _18824_ (.B1(_09473_),
    .Y(_09474_),
    .A1(_09469_),
    .A2(_09472_));
 sg13g2_o21ai_1 _18825_ (.B1(_09474_),
    .Y(_09475_),
    .A1(net169),
    .A2(_09466_));
 sg13g2_nand2_1 _18826_ (.Y(_09476_),
    .A(_09475_),
    .B(net143));
 sg13g2_o21ai_1 _18827_ (.B1(_09476_),
    .Y(_00480_),
    .A1(_07857_),
    .A2(net144));
 sg13g2_nor2_1 _18828_ (.A(_06307_),
    .B(_06314_),
    .Y(_09477_));
 sg13g2_inv_1 _18829_ (.Y(_09478_),
    .A(net220));
 sg13g2_nor2_1 _18830_ (.A(_06247_),
    .B(_09478_),
    .Y(_09479_));
 sg13g2_inv_1 _18831_ (.Y(_09480_),
    .A(_09479_));
 sg13g2_nand2b_1 _18832_ (.Y(_09481_),
    .B(_09480_),
    .A_N(_09477_));
 sg13g2_inv_1 _18833_ (.Y(_09482_),
    .A(_09465_));
 sg13g2_a21oi_1 _18834_ (.A1(_09482_),
    .A2(_09463_),
    .Y(_09483_),
    .B1(_09461_));
 sg13g2_xor2_1 _18835_ (.B(_09483_),
    .A(_09481_),
    .X(_09484_));
 sg13g2_nor2_1 _18836_ (.A(_07860_),
    .B(_06371_),
    .Y(_09485_));
 sg13g2_nand2_1 _18837_ (.Y(_09486_),
    .A(_07860_),
    .B(_06371_));
 sg13g2_nor2b_1 _18838_ (.A(_09485_),
    .B_N(_09486_),
    .Y(_09487_));
 sg13g2_nand2_1 _18839_ (.Y(_09488_),
    .A(_09436_),
    .B(_09468_));
 sg13g2_a21oi_1 _18840_ (.A1(_09457_),
    .A2(_09437_),
    .Y(_09489_),
    .B1(_09488_));
 sg13g2_nor2_1 _18841_ (.A(_09467_),
    .B(_09489_),
    .Y(_09490_));
 sg13g2_inv_1 _18842_ (.Y(_09491_),
    .A(_06221_));
 sg13g2_a21oi_1 _18843_ (.A1(_09490_),
    .A2(_09487_),
    .Y(_09492_),
    .B1(_09491_));
 sg13g2_o21ai_1 _18844_ (.B1(_09492_),
    .Y(_09493_),
    .A1(_09487_),
    .A2(_09490_));
 sg13g2_o21ai_1 _18845_ (.B1(_09493_),
    .Y(_09494_),
    .A1(net169),
    .A2(_09484_));
 sg13g2_nand2_1 _18846_ (.Y(_09495_),
    .A(_09494_),
    .B(net143));
 sg13g2_o21ai_1 _18847_ (.B1(_09495_),
    .Y(_00481_),
    .A1(_07892_),
    .A2(net144));
 sg13g2_nor2_1 _18848_ (.A(_06330_),
    .B(_06301_),
    .Y(_09496_));
 sg13g2_nor2_1 _18849_ (.A(_06245_),
    .B(_06331_),
    .Y(_09497_));
 sg13g2_inv_1 _18850_ (.Y(_09498_),
    .A(_09497_));
 sg13g2_nand2b_1 _18851_ (.Y(_09499_),
    .B(_09498_),
    .A_N(_09496_));
 sg13g2_inv_1 _18852_ (.Y(_09500_),
    .A(_09483_));
 sg13g2_a21oi_1 _18853_ (.A1(_09500_),
    .A2(_09480_),
    .Y(_09501_),
    .B1(_09477_));
 sg13g2_xor2_1 _18854_ (.B(_09501_),
    .A(_09499_),
    .X(_09502_));
 sg13g2_nand2_1 _18855_ (.Y(_09503_),
    .A(_09468_),
    .B(_09486_));
 sg13g2_a21oi_1 _18856_ (.A1(_09472_),
    .A2(_09469_),
    .Y(_09504_),
    .B1(_09503_));
 sg13g2_xor2_1 _18857_ (.B(net188),
    .A(_07895_),
    .X(_09505_));
 sg13g2_inv_1 _18858_ (.Y(_09506_),
    .A(_09505_));
 sg13g2_o21ai_1 _18859_ (.B1(_09506_),
    .Y(_09507_),
    .A1(_09485_),
    .A2(_09504_));
 sg13g2_nor2_1 _18860_ (.A(_09485_),
    .B(_09504_),
    .Y(_09508_));
 sg13g2_nand2_1 _18861_ (.Y(_09509_),
    .A(_09508_),
    .B(_09505_));
 sg13g2_nand3_1 _18862_ (.B(_06221_),
    .C(_09509_),
    .A(_09507_),
    .Y(_09510_));
 sg13g2_o21ai_1 _18863_ (.B1(_09510_),
    .Y(_09511_),
    .A1(net169),
    .A2(_09502_));
 sg13g2_nand2_1 _18864_ (.Y(_09512_),
    .A(_09511_),
    .B(net143));
 sg13g2_o21ai_1 _18865_ (.B1(_09512_),
    .Y(_00482_),
    .A1(_07931_),
    .A2(net144));
 sg13g2_nor2_1 _18866_ (.A(_06352_),
    .B(_06240_),
    .Y(_09513_));
 sg13g2_nor2_1 _18867_ (.A(_06235_),
    .B(_06364_),
    .Y(_09514_));
 sg13g2_inv_1 _18868_ (.Y(_09515_),
    .A(_09514_));
 sg13g2_nand2b_1 _18869_ (.Y(_09516_),
    .B(_09515_),
    .A_N(_09513_));
 sg13g2_inv_1 _18870_ (.Y(_09517_),
    .A(_09501_));
 sg13g2_a21oi_1 _18871_ (.A1(_09517_),
    .A2(_09498_),
    .Y(_09518_),
    .B1(_09496_));
 sg13g2_xor2_1 _18872_ (.B(_09518_),
    .A(_09516_),
    .X(_09519_));
 sg13g2_nor2b_1 _18873_ (.A(_09506_),
    .B_N(_09487_),
    .Y(_09520_));
 sg13g2_o21ai_1 _18874_ (.B1(net181),
    .Y(_09521_),
    .A1(_07860_),
    .A2(_07895_));
 sg13g2_inv_1 _18875_ (.Y(_09522_),
    .A(_09521_));
 sg13g2_a21oi_1 _18876_ (.A1(_09490_),
    .A2(_09520_),
    .Y(_09523_),
    .B1(_09522_));
 sg13g2_xor2_1 _18877_ (.B(net188),
    .A(_07928_),
    .X(_09524_));
 sg13g2_inv_1 _18878_ (.Y(_09525_),
    .A(_09524_));
 sg13g2_a21oi_1 _18879_ (.A1(_09523_),
    .A2(_09525_),
    .Y(_09526_),
    .B1(_09416_));
 sg13g2_o21ai_1 _18880_ (.B1(_09526_),
    .Y(_09527_),
    .A1(_09523_),
    .A2(_09525_));
 sg13g2_o21ai_1 _18881_ (.B1(_09527_),
    .Y(_09528_),
    .A1(net169),
    .A2(_09519_));
 sg13g2_nand2_1 _18882_ (.Y(_09529_),
    .A(_09528_),
    .B(net143));
 sg13g2_o21ai_1 _18883_ (.B1(_09529_),
    .Y(_00483_),
    .A1(_07961_),
    .A2(_09364_));
 sg13g2_nor2_1 _18884_ (.A(net227),
    .B(_06361_),
    .Y(_09530_));
 sg13g2_nor2_1 _18885_ (.A(_06360_),
    .B(_06311_),
    .Y(_09531_));
 sg13g2_nor2_1 _18886_ (.A(_09530_),
    .B(_09531_),
    .Y(_09532_));
 sg13g2_inv_1 _18887_ (.Y(_09533_),
    .A(_09518_));
 sg13g2_a21oi_1 _18888_ (.A1(_09533_),
    .A2(_09515_),
    .Y(_09534_),
    .B1(_09513_));
 sg13g2_xnor2_1 _18889_ (.Y(_09535_),
    .A(_09532_),
    .B(_09534_));
 sg13g2_o21ai_1 _18890_ (.B1(net188),
    .Y(_09536_),
    .A1(_07895_),
    .A2(_07928_));
 sg13g2_o21ai_1 _18891_ (.B1(_09536_),
    .Y(_09537_),
    .A1(_09525_),
    .A2(_09509_));
 sg13g2_xor2_1 _18892_ (.B(net188),
    .A(_07964_),
    .X(_09538_));
 sg13g2_inv_1 _18893_ (.Y(_09539_),
    .A(_09538_));
 sg13g2_nand2b_1 _18894_ (.Y(_09540_),
    .B(_09539_),
    .A_N(_09537_));
 sg13g2_nand2_1 _18895_ (.Y(_09541_),
    .A(_09537_),
    .B(_09538_));
 sg13g2_nand3_1 _18896_ (.B(_06221_),
    .C(_09541_),
    .A(_09540_),
    .Y(_09542_));
 sg13g2_o21ai_1 _18897_ (.B1(_09542_),
    .Y(_09543_),
    .A1(_09365_),
    .A2(_09535_));
 sg13g2_nand2_1 _18898_ (.Y(_09544_),
    .A(_09543_),
    .B(_09420_));
 sg13g2_o21ai_1 _18899_ (.B1(_09544_),
    .Y(_00484_),
    .A1(_08001_),
    .A2(_09364_));
 sg13g2_inv_1 _18900_ (.Y(_09545_),
    .A(_07997_));
 sg13g2_buf_1 _18901_ (.A(_06221_),
    .X(_09546_));
 sg13g2_nor2_2 _18902_ (.A(net220),
    .B(_06372_),
    .Y(_09547_));
 sg13g2_nor2_1 _18903_ (.A(net188),
    .B(_09478_),
    .Y(_09548_));
 sg13g2_inv_1 _18904_ (.Y(_09549_),
    .A(_09534_));
 sg13g2_inv_1 _18905_ (.Y(_09550_),
    .A(_09530_));
 sg13g2_a21oi_1 _18906_ (.A1(_09549_),
    .A2(_09550_),
    .Y(_09551_),
    .B1(_09531_));
 sg13g2_inv_1 _18907_ (.Y(_09552_),
    .A(_09551_));
 sg13g2_nor3_1 _18908_ (.A(_09547_),
    .B(_09548_),
    .C(_09552_),
    .Y(_09553_));
 sg13g2_nor2_1 _18909_ (.A(net157),
    .B(_09553_),
    .Y(_09554_));
 sg13g2_o21ai_1 _18910_ (.B1(_09552_),
    .Y(_09555_),
    .A1(_09547_),
    .A2(_09548_));
 sg13g2_buf_1 _18911_ (.A(_06976_),
    .X(_09556_));
 sg13g2_a21oi_1 _18912_ (.A1(_09554_),
    .A2(_09555_),
    .Y(_09557_),
    .B1(net127));
 sg13g2_nor2_1 _18913_ (.A(_09525_),
    .B(_09539_),
    .Y(_09558_));
 sg13g2_nand3_1 _18914_ (.B(_09520_),
    .C(_09558_),
    .A(_09490_),
    .Y(_09559_));
 sg13g2_o21ai_1 _18915_ (.B1(net181),
    .Y(_09560_),
    .A1(_07928_),
    .A2(_07964_));
 sg13g2_inv_1 _18916_ (.Y(_09561_),
    .A(_09560_));
 sg13g2_a21oi_1 _18917_ (.A1(_09558_),
    .A2(_09522_),
    .Y(_09562_),
    .B1(_09561_));
 sg13g2_nand2_1 _18918_ (.Y(_09563_),
    .A(_09559_),
    .B(_09562_));
 sg13g2_xor2_1 _18919_ (.B(net188),
    .A(_07997_),
    .X(_09564_));
 sg13g2_o21ai_1 _18920_ (.B1(_09355_),
    .Y(_09565_),
    .A1(_09564_),
    .A2(_09563_));
 sg13g2_a21o_1 _18921_ (.A2(_09564_),
    .A1(_09563_),
    .B1(_09565_),
    .X(_09566_));
 sg13g2_a22oi_1 _18922_ (.Y(_00485_),
    .B1(_09557_),
    .B2(_09566_),
    .A2(net114),
    .A1(_09545_));
 sg13g2_nor2_1 _18923_ (.A(_06330_),
    .B(_06372_),
    .Y(_09567_));
 sg13g2_nor2_1 _18924_ (.A(net188),
    .B(_06331_),
    .Y(_09568_));
 sg13g2_nor2_1 _18925_ (.A(_09567_),
    .B(_09568_),
    .Y(_09569_));
 sg13g2_nor2_1 _18926_ (.A(_09548_),
    .B(_09552_),
    .Y(_09570_));
 sg13g2_nor3_1 _18927_ (.A(_09547_),
    .B(_09569_),
    .C(_09570_),
    .Y(_09571_));
 sg13g2_inv_1 _18928_ (.Y(_09572_),
    .A(_09570_));
 sg13g2_inv_1 _18929_ (.Y(_09573_),
    .A(_09547_));
 sg13g2_inv_1 _18930_ (.Y(_09574_),
    .A(_09569_));
 sg13g2_a21oi_1 _18931_ (.A1(_09572_),
    .A2(_09573_),
    .Y(_09575_),
    .B1(_09574_));
 sg13g2_nor3_1 _18932_ (.A(_09546_),
    .B(_09571_),
    .C(_09575_),
    .Y(_09576_));
 sg13g2_nor2_1 _18933_ (.A(net127),
    .B(_09576_),
    .Y(_09577_));
 sg13g2_o21ai_1 _18934_ (.B1(net181),
    .Y(_09578_),
    .A1(_07964_),
    .A2(_07997_));
 sg13g2_inv_1 _18935_ (.Y(_09579_),
    .A(_09578_));
 sg13g2_inv_1 _18936_ (.Y(_09580_),
    .A(_09564_));
 sg13g2_nor2_1 _18937_ (.A(_09580_),
    .B(_09541_),
    .Y(_09581_));
 sg13g2_nor2_1 _18938_ (.A(_09579_),
    .B(_09581_),
    .Y(_09582_));
 sg13g2_xor2_1 _18939_ (.B(_08911_),
    .A(_08030_),
    .X(_09583_));
 sg13g2_inv_1 _18940_ (.Y(_09584_),
    .A(_09583_));
 sg13g2_a21oi_1 _18941_ (.A1(_09582_),
    .A2(_09584_),
    .Y(_09585_),
    .B1(_09458_));
 sg13g2_o21ai_1 _18942_ (.B1(_09585_),
    .Y(_09586_),
    .A1(_09582_),
    .A2(_09584_));
 sg13g2_a22oi_1 _18943_ (.Y(_00486_),
    .B1(_09577_),
    .B2(_09586_),
    .A2(_09423_),
    .A1(_08059_));
 sg13g2_inv_1 _18944_ (.Y(_09587_),
    .A(_09567_));
 sg13g2_nand2_1 _18945_ (.Y(_09588_),
    .A(_09573_),
    .B(_09587_));
 sg13g2_nor2_1 _18946_ (.A(net219),
    .B(_06372_),
    .Y(_09589_));
 sg13g2_nor2_1 _18947_ (.A(net181),
    .B(_06364_),
    .Y(_09590_));
 sg13g2_nor2_1 _18948_ (.A(_09589_),
    .B(_09590_),
    .Y(_09591_));
 sg13g2_nor3_1 _18949_ (.A(_09547_),
    .B(_09574_),
    .C(_09572_),
    .Y(_09592_));
 sg13g2_nor3_1 _18950_ (.A(_09588_),
    .B(_09591_),
    .C(_09592_),
    .Y(_09593_));
 sg13g2_nor2_1 _18951_ (.A(_09588_),
    .B(_09592_),
    .Y(_09594_));
 sg13g2_nor2b_1 _18952_ (.A(_09594_),
    .B_N(_09591_),
    .Y(_09595_));
 sg13g2_nor3_1 _18953_ (.A(net159),
    .B(_09593_),
    .C(_09595_),
    .Y(_09596_));
 sg13g2_nor2_1 _18954_ (.A(_09556_),
    .B(_09596_),
    .Y(_09597_));
 sg13g2_xor2_1 _18955_ (.B(_08911_),
    .A(_08056_),
    .X(_09598_));
 sg13g2_nor2_1 _18956_ (.A(_09580_),
    .B(_09584_),
    .Y(_09599_));
 sg13g2_nand2_1 _18957_ (.Y(_09600_),
    .A(_09558_),
    .B(_09599_));
 sg13g2_a21oi_1 _18958_ (.A1(_09545_),
    .A2(_08059_),
    .Y(_09601_),
    .B1(_06372_));
 sg13g2_a21oi_1 _18959_ (.A1(_09599_),
    .A2(_09561_),
    .Y(_09602_),
    .B1(_09601_));
 sg13g2_o21ai_1 _18960_ (.B1(_09602_),
    .Y(_09603_),
    .A1(_09600_),
    .A2(_09523_));
 sg13g2_a21oi_1 _18961_ (.A1(_09603_),
    .A2(_09598_),
    .Y(_09604_),
    .B1(_09458_));
 sg13g2_o21ai_1 _18962_ (.B1(_09604_),
    .Y(_09605_),
    .A1(_09598_),
    .A2(_09603_));
 sg13g2_a22oi_1 _18963_ (.Y(_00487_),
    .B1(_09597_),
    .B2(_09605_),
    .A2(_09423_),
    .A1(_08090_));
 sg13g2_xor2_1 _18964_ (.B(_09386_),
    .A(_09357_),
    .X(_09606_));
 sg13g2_nand2_1 _18965_ (.Y(_09607_),
    .A(_06975_),
    .B(net157));
 sg13g2_nand2_1 _18966_ (.Y(_09608_),
    .A(net128),
    .B(_08083_));
 sg13g2_o21ai_1 _18967_ (.B1(_09608_),
    .Y(_00488_),
    .A1(_09606_),
    .A2(_09607_));
 sg13g2_xnor2_1 _18968_ (.Y(_09609_),
    .A(net218),
    .B(net181));
 sg13g2_nor2_1 _18969_ (.A(_09589_),
    .B(_09575_),
    .Y(_09610_));
 sg13g2_o21ai_1 _18970_ (.B1(_09587_),
    .Y(_09611_),
    .A1(_09590_),
    .A2(_09610_));
 sg13g2_or2_1 _18971_ (.X(_09612_),
    .B(_09611_),
    .A(_09609_));
 sg13g2_a21oi_1 _18972_ (.A1(_09611_),
    .A2(_09609_),
    .Y(_09613_),
    .B1(_09546_));
 sg13g2_xor2_1 _18973_ (.B(net181),
    .A(_08087_),
    .X(_09614_));
 sg13g2_nor2b_1 _18974_ (.A(_09584_),
    .B_N(_09598_),
    .Y(_09615_));
 sg13g2_a22oi_1 _18975_ (.Y(_09616_),
    .B1(_09579_),
    .B2(_09615_),
    .A2(net181),
    .A1(_08030_));
 sg13g2_o21ai_1 _18976_ (.B1(_09616_),
    .Y(_09617_),
    .A1(_08090_),
    .A2(_06372_));
 sg13g2_a21oi_1 _18977_ (.A1(_09581_),
    .A2(_09615_),
    .Y(_09618_),
    .B1(_09617_));
 sg13g2_xnor2_1 _18978_ (.Y(_09619_),
    .A(_09614_),
    .B(_09618_));
 sg13g2_a221oi_1 _18979_ (.B2(_09365_),
    .C1(net129),
    .B1(_09619_),
    .A1(_09612_),
    .Y(_09620_),
    .A2(_09613_));
 sg13g2_a21oi_1 _18980_ (.A1(_08111_),
    .A2(net114),
    .Y(_00489_),
    .B1(_09620_));
 sg13g2_inv_1 _18981_ (.Y(_09621_),
    .A(\vgadonut.donut.ycA[21] ));
 sg13g2_nand2_1 _18982_ (.Y(_09622_),
    .A(_09595_),
    .B(_09609_));
 sg13g2_a21oi_1 _18983_ (.A1(net219),
    .A2(net218),
    .Y(_09623_),
    .B1(_06372_));
 sg13g2_nor2_1 _18984_ (.A(_09623_),
    .B(net159),
    .Y(_09624_));
 sg13g2_a21oi_1 _18985_ (.A1(_09622_),
    .A2(_09624_),
    .Y(_09625_),
    .B1(_09556_));
 sg13g2_and3_1 _18986_ (.X(_09626_),
    .A(_09599_),
    .B(_09598_),
    .C(_09614_));
 sg13g2_nand3_1 _18987_ (.B(_09598_),
    .C(_09614_),
    .A(_09601_),
    .Y(_09627_));
 sg13g2_o21ai_1 _18988_ (.B1(net181),
    .Y(_09628_),
    .A1(_08056_),
    .A2(_08087_));
 sg13g2_nand2_1 _18989_ (.Y(_09629_),
    .A(_09627_),
    .B(_09628_));
 sg13g2_a21oi_1 _18990_ (.A1(_09563_),
    .A2(_09626_),
    .Y(_09630_),
    .B1(_09629_));
 sg13g2_xnor2_1 _18991_ (.Y(_09631_),
    .A(\vgadonut.donut.ycA[21] ),
    .B(_08912_));
 sg13g2_buf_1 _18992_ (.A(net168),
    .X(_09632_));
 sg13g2_a21oi_1 _18993_ (.A1(_09630_),
    .A2(_09631_),
    .Y(_09633_),
    .B1(_09632_));
 sg13g2_o21ai_1 _18994_ (.B1(_09633_),
    .Y(_09634_),
    .A1(_09630_),
    .A2(_09631_));
 sg13g2_a22oi_1 _18995_ (.Y(_00490_),
    .B1(_09625_),
    .B2(_09634_),
    .A2(net114),
    .A1(_09621_));
 sg13g2_xnor2_1 _18996_ (.Y(_09635_),
    .A(_09393_),
    .B(_09389_));
 sg13g2_nand2_1 _18997_ (.Y(_09636_),
    .A(net128),
    .B(_07680_));
 sg13g2_o21ai_1 _18998_ (.B1(_09636_),
    .Y(_00491_),
    .A1(_09635_),
    .A2(_09607_));
 sg13g2_inv_1 _18999_ (.Y(_09638_),
    .A(_07681_));
 sg13g2_nand2b_1 _19000_ (.Y(_09639_),
    .B(_09441_),
    .A_N(_09442_));
 sg13g2_nand3_1 _19001_ (.B(_06977_),
    .C(_09639_),
    .A(_09443_),
    .Y(_09640_));
 sg13g2_o21ai_1 _19002_ (.B1(_09640_),
    .Y(_00492_),
    .A1(_09638_),
    .A2(_06975_));
 sg13g2_xnor2_1 _19003_ (.Y(_09641_),
    .A(_09398_),
    .B(_09397_));
 sg13g2_a22oi_1 _19004_ (.Y(_09642_),
    .B1(net157),
    .B2(_09641_),
    .A2(_09361_),
    .A1(_06978_));
 sg13g2_a21o_1 _19005_ (.A2(net128),
    .A1(_07663_),
    .B1(_09642_),
    .X(_00493_));
 sg13g2_a21oi_1 _19006_ (.A1(_06252_),
    .A2(net158),
    .Y(_09643_),
    .B1(net127));
 sg13g2_a21oi_1 _19007_ (.A1(_09444_),
    .A2(_09445_),
    .Y(_09644_),
    .B1(_09632_));
 sg13g2_o21ai_1 _19008_ (.B1(_09644_),
    .Y(_09646_),
    .A1(_09445_),
    .A2(_09444_));
 sg13g2_a22oi_1 _19009_ (.Y(_00494_),
    .B1(_09643_),
    .B2(_09646_),
    .A2(net114),
    .A1(_07670_));
 sg13g2_a21oi_1 _19010_ (.A1(_06276_),
    .A2(net158),
    .Y(_09647_),
    .B1(net127));
 sg13g2_nand2b_1 _19011_ (.Y(_09648_),
    .B(_09383_),
    .A_N(_09403_));
 sg13g2_nand3_1 _19012_ (.B(_09356_),
    .C(_09404_),
    .A(_09648_),
    .Y(_09649_));
 sg13g2_a22oi_1 _19013_ (.Y(_00495_),
    .B1(_09647_),
    .B2(_09649_),
    .A2(net114),
    .A1(_07643_));
 sg13g2_o21ai_1 _19014_ (.B1(_06975_),
    .Y(_09650_),
    .A1(_06284_),
    .A2(_09356_));
 sg13g2_or2_1 _19015_ (.X(_09651_),
    .B(_09448_),
    .A(_09449_));
 sg13g2_a21oi_1 _19016_ (.A1(_09651_),
    .A2(_09450_),
    .Y(_09652_),
    .B1(net158));
 sg13g2_nand2_1 _19017_ (.Y(_09653_),
    .A(_09424_),
    .B(_07581_));
 sg13g2_o21ai_1 _19018_ (.B1(_09653_),
    .Y(_00496_),
    .A1(_09650_),
    .A2(_09652_));
 sg13g2_xor2_1 _19019_ (.B(_06260_),
    .A(_06292_),
    .X(_09655_));
 sg13g2_a21oi_1 _19020_ (.A1(_09491_),
    .A2(_09655_),
    .Y(_09656_),
    .B1(_09422_));
 sg13g2_nand2b_1 _19021_ (.Y(_09657_),
    .B(_09380_),
    .A_N(_09409_));
 sg13g2_nand3_1 _19022_ (.B(net159),
    .C(_09410_),
    .A(_09657_),
    .Y(_09658_));
 sg13g2_a22oi_1 _19023_ (.Y(_00497_),
    .B1(_09656_),
    .B2(_09658_),
    .A2(net114),
    .A1(_07597_));
 sg13g2_buf_1 _19024_ (.A(net129),
    .X(_09659_));
 sg13g2_xnor2_1 _19025_ (.Y(_09660_),
    .A(_09370_),
    .B(_09371_));
 sg13g2_a21oi_1 _19026_ (.A1(net158),
    .A2(_09660_),
    .Y(_09661_),
    .B1(_09422_));
 sg13g2_a21oi_1 _19027_ (.A1(_09453_),
    .A2(_09454_),
    .Y(_09662_),
    .B1(net156));
 sg13g2_o21ai_1 _19028_ (.B1(_09662_),
    .Y(_09664_),
    .A1(_09454_),
    .A2(_09453_));
 sg13g2_a22oi_1 _19029_ (.Y(_00498_),
    .B1(_09661_),
    .B2(_09664_),
    .A2(_09659_),
    .A1(_07624_));
 sg13g2_nand2_1 _19030_ (.Y(_09665_),
    .A(\vgadonut.donut.ysA[0] ),
    .B(_08851_));
 sg13g2_nand2_1 _19031_ (.Y(_09666_),
    .A(net159),
    .B(_09665_));
 sg13g2_nor2_1 _19032_ (.A(_08852_),
    .B(_06976_),
    .Y(_09667_));
 sg13g2_inv_1 _19033_ (.Y(_09668_),
    .A(_09667_));
 sg13g2_a22oi_1 _19034_ (.Y(_00499_),
    .B1(_08186_),
    .B2(_09668_),
    .A2(_06975_),
    .A1(_09666_));
 sg13g2_nor2_1 _19035_ (.A(net223),
    .B(_08823_),
    .Y(_09669_));
 sg13g2_nor2_1 _19036_ (.A(net215),
    .B(_06255_),
    .Y(_09670_));
 sg13g2_inv_1 _19037_ (.Y(_09671_),
    .A(_09670_));
 sg13g2_nand2b_1 _19038_ (.Y(_09673_),
    .B(_09671_),
    .A_N(_09669_));
 sg13g2_inv_1 _19039_ (.Y(_09674_),
    .A(_08856_));
 sg13g2_nor2_1 _19040_ (.A(_06262_),
    .B(_08852_),
    .Y(_09675_));
 sg13g2_xnor2_1 _19041_ (.Y(_09676_),
    .A(_08856_),
    .B(net195));
 sg13g2_nor2b_1 _19042_ (.A(_09675_),
    .B_N(_09676_),
    .Y(_09677_));
 sg13g2_a21oi_1 _19043_ (.A1(_09674_),
    .A2(_06258_),
    .Y(_09678_),
    .B1(_09677_));
 sg13g2_xnor2_1 _19044_ (.Y(_09679_),
    .A(_09673_),
    .B(_09678_));
 sg13g2_nor2_1 _19045_ (.A(_08281_),
    .B(net224),
    .Y(_09680_));
 sg13g2_nand2_1 _19046_ (.Y(_09681_),
    .A(_08281_),
    .B(net224));
 sg13g2_nor2b_1 _19047_ (.A(_09680_),
    .B_N(_09681_),
    .Y(_09682_));
 sg13g2_nor2_1 _19048_ (.A(_08263_),
    .B(net221),
    .Y(_09684_));
 sg13g2_nor2_1 _19049_ (.A(_08245_),
    .B(net193),
    .Y(_09685_));
 sg13g2_nor2_1 _19050_ (.A(_08305_),
    .B(net195),
    .Y(_09686_));
 sg13g2_nor2_1 _19051_ (.A(_08330_),
    .B(net198),
    .Y(_09687_));
 sg13g2_xor2_1 _19052_ (.B(_08856_),
    .A(_08701_),
    .X(_09688_));
 sg13g2_inv_1 _19053_ (.Y(_09689_),
    .A(_09688_));
 sg13g2_nand2_1 _19054_ (.Y(_09690_),
    .A(_08701_),
    .B(_08856_));
 sg13g2_o21ai_1 _19055_ (.B1(_09690_),
    .Y(_09691_),
    .A1(_09665_),
    .A2(_09689_));
 sg13g2_nor2_1 _19056_ (.A(_08341_),
    .B(net215),
    .Y(_09692_));
 sg13g2_nand2_1 _19057_ (.Y(_09693_),
    .A(_08341_),
    .B(net215));
 sg13g2_nor2b_1 _19058_ (.A(_09692_),
    .B_N(_09693_),
    .Y(_09695_));
 sg13g2_nand2_1 _19059_ (.Y(_09696_),
    .A(_08330_),
    .B(net198));
 sg13g2_nand2_1 _19060_ (.Y(_09697_),
    .A(_09696_),
    .B(_09693_));
 sg13g2_a21oi_1 _19061_ (.A1(_09691_),
    .A2(_09695_),
    .Y(_09698_),
    .B1(_09697_));
 sg13g2_nor2_1 _19062_ (.A(_09687_),
    .B(_09698_),
    .Y(_09699_));
 sg13g2_xor2_1 _19063_ (.B(net194),
    .A(_08317_),
    .X(_09700_));
 sg13g2_nand2_1 _19064_ (.Y(_09701_),
    .A(_09699_),
    .B(_09700_));
 sg13g2_nand2_1 _19065_ (.Y(_09702_),
    .A(_08305_),
    .B(net195));
 sg13g2_nand2_1 _19066_ (.Y(_09703_),
    .A(_08317_),
    .B(net194));
 sg13g2_nand3_1 _19067_ (.B(_09702_),
    .C(_09703_),
    .A(_09701_),
    .Y(_09704_));
 sg13g2_nor2b_1 _19068_ (.A(_09686_),
    .B_N(_09704_),
    .Y(_09706_));
 sg13g2_nor2_1 _19069_ (.A(_08298_),
    .B(net223),
    .Y(_09707_));
 sg13g2_nand2_1 _19070_ (.Y(_09708_),
    .A(_08298_),
    .B(_06251_));
 sg13g2_nor2b_1 _19071_ (.A(_09707_),
    .B_N(_09708_),
    .Y(_09709_));
 sg13g2_nand2_1 _19072_ (.Y(_09710_),
    .A(_08245_),
    .B(net193));
 sg13g2_nand2_1 _19073_ (.Y(_09711_),
    .A(_09708_),
    .B(_09710_));
 sg13g2_a21oi_1 _19074_ (.A1(_09706_),
    .A2(_09709_),
    .Y(_09712_),
    .B1(_09711_));
 sg13g2_nor2_1 _19075_ (.A(_09685_),
    .B(_09712_),
    .Y(_09713_));
 sg13g2_nor2_1 _19076_ (.A(_08249_),
    .B(net222),
    .Y(_09714_));
 sg13g2_nand2_1 _19077_ (.Y(_09715_),
    .A(_08249_),
    .B(net222));
 sg13g2_nor2b_1 _19078_ (.A(_09714_),
    .B_N(_09715_),
    .Y(_09717_));
 sg13g2_nand2_1 _19079_ (.Y(_09718_),
    .A(_08263_),
    .B(net221));
 sg13g2_nand2_1 _19080_ (.Y(_09719_),
    .A(_09715_),
    .B(_09718_));
 sg13g2_a21oi_1 _19081_ (.A1(_09713_),
    .A2(_09717_),
    .Y(_09720_),
    .B1(_09719_));
 sg13g2_nor2_1 _19082_ (.A(_09684_),
    .B(_09720_),
    .Y(_09721_));
 sg13g2_a21oi_1 _19083_ (.A1(_09721_),
    .A2(_09682_),
    .Y(_09722_),
    .B1(net168));
 sg13g2_o21ai_1 _19084_ (.B1(_09722_),
    .Y(_09723_),
    .A1(_09682_),
    .A2(_09721_));
 sg13g2_o21ai_1 _19085_ (.B1(_09723_),
    .Y(_09724_),
    .A1(_06340_),
    .A2(_09679_));
 sg13g2_nand2_1 _19086_ (.Y(_09725_),
    .A(_09724_),
    .B(net143));
 sg13g2_o21ai_1 _19087_ (.B1(_09725_),
    .Y(_00500_),
    .A1(_08282_),
    .A2(net144));
 sg13g2_nor2_1 _19088_ (.A(net198),
    .B(_06279_),
    .Y(_09727_));
 sg13g2_inv_1 _19089_ (.Y(_09728_),
    .A(_09727_));
 sg13g2_nor2_1 _19090_ (.A(net193),
    .B(_06264_),
    .Y(_09729_));
 sg13g2_inv_1 _19091_ (.Y(_09730_),
    .A(_09729_));
 sg13g2_o21ai_1 _19092_ (.B1(_09671_),
    .Y(_09731_),
    .A1(_09669_),
    .A2(_09678_));
 sg13g2_a21oi_1 _19093_ (.A1(_09728_),
    .A2(_09730_),
    .Y(_09732_),
    .B1(_09731_));
 sg13g2_nand2_1 _19094_ (.Y(_09733_),
    .A(_09731_),
    .B(_09730_));
 sg13g2_nor2_1 _19095_ (.A(_09727_),
    .B(_09733_),
    .Y(_09734_));
 sg13g2_nor3_1 _19096_ (.A(_09355_),
    .B(_09732_),
    .C(_09734_),
    .Y(_09735_));
 sg13g2_nor2_1 _19097_ (.A(net127),
    .B(_09735_),
    .Y(_09736_));
 sg13g2_nor2_1 _19098_ (.A(_08405_),
    .B(_06244_),
    .Y(_09738_));
 sg13g2_nand2_1 _19099_ (.Y(_09739_),
    .A(_08405_),
    .B(net226));
 sg13g2_nor2b_1 _19100_ (.A(_09738_),
    .B_N(_09739_),
    .Y(_09740_));
 sg13g2_inv_1 _19101_ (.Y(_09741_),
    .A(_09691_));
 sg13g2_o21ai_1 _19102_ (.B1(_09693_),
    .Y(_09742_),
    .A1(_09692_),
    .A2(_09741_));
 sg13g2_nor2b_1 _19103_ (.A(_09687_),
    .B_N(_09696_),
    .Y(_09743_));
 sg13g2_nand2_1 _19104_ (.Y(_09744_),
    .A(_09703_),
    .B(_09696_));
 sg13g2_a21oi_1 _19105_ (.A1(_09742_),
    .A2(_09743_),
    .Y(_09745_),
    .B1(_09744_));
 sg13g2_a21oi_1 _19106_ (.A1(_08318_),
    .A2(_06263_),
    .Y(_09746_),
    .B1(_09745_));
 sg13g2_nor2b_1 _19107_ (.A(_09686_),
    .B_N(_09702_),
    .Y(_09747_));
 sg13g2_nand2_1 _19108_ (.Y(_09749_),
    .A(_09708_),
    .B(_09702_));
 sg13g2_a21oi_1 _19109_ (.A1(_09746_),
    .A2(_09747_),
    .Y(_09750_),
    .B1(_09749_));
 sg13g2_nor2_1 _19110_ (.A(_09707_),
    .B(_09750_),
    .Y(_09751_));
 sg13g2_nor2b_1 _19111_ (.A(_09685_),
    .B_N(_09710_),
    .Y(_09752_));
 sg13g2_nand2_1 _19112_ (.Y(_09753_),
    .A(_09715_),
    .B(_09710_));
 sg13g2_a21oi_1 _19113_ (.A1(_09751_),
    .A2(_09752_),
    .Y(_09754_),
    .B1(_09753_));
 sg13g2_nor2_1 _19114_ (.A(_09714_),
    .B(_09754_),
    .Y(_09755_));
 sg13g2_nor2b_1 _19115_ (.A(_09684_),
    .B_N(_09718_),
    .Y(_09756_));
 sg13g2_nand2_1 _19116_ (.Y(_09757_),
    .A(_09681_),
    .B(_09718_));
 sg13g2_a21oi_1 _19117_ (.A1(_09755_),
    .A2(_09756_),
    .Y(_09758_),
    .B1(_09757_));
 sg13g2_nor2_1 _19118_ (.A(_09680_),
    .B(_09758_),
    .Y(_09760_));
 sg13g2_a21oi_1 _19119_ (.A1(_09760_),
    .A2(_09740_),
    .Y(_09761_),
    .B1(net156));
 sg13g2_o21ai_1 _19120_ (.B1(_09761_),
    .Y(_09762_),
    .A1(_09740_),
    .A2(_09760_));
 sg13g2_a22oi_1 _19121_ (.Y(_00501_),
    .B1(_09736_),
    .B2(_09762_),
    .A2(net113),
    .A1(_08406_));
 sg13g2_nor2_1 _19122_ (.A(net222),
    .B(_06263_),
    .Y(_09763_));
 sg13g2_nor2_1 _19123_ (.A(_06262_),
    .B(_06288_),
    .Y(_09764_));
 sg13g2_inv_1 _19124_ (.Y(_09765_),
    .A(_09764_));
 sg13g2_nand2b_1 _19125_ (.Y(_09766_),
    .B(_09765_),
    .A_N(_09763_));
 sg13g2_nand2_1 _19126_ (.Y(_09767_),
    .A(_09733_),
    .B(_09728_));
 sg13g2_xor2_1 _19127_ (.B(_09767_),
    .A(_09766_),
    .X(_09768_));
 sg13g2_nor2_1 _19128_ (.A(_08428_),
    .B(_06237_),
    .Y(_09770_));
 sg13g2_nand2_1 _19129_ (.Y(_09771_),
    .A(_08428_),
    .B(_06237_));
 sg13g2_nor2b_1 _19130_ (.A(_09770_),
    .B_N(_09771_),
    .Y(_09772_));
 sg13g2_nand2_1 _19131_ (.Y(_09773_),
    .A(_09681_),
    .B(_09739_));
 sg13g2_a21oi_1 _19132_ (.A1(_09721_),
    .A2(_09682_),
    .Y(_09774_),
    .B1(_09773_));
 sg13g2_nor2_1 _19133_ (.A(_09738_),
    .B(_09774_),
    .Y(_09775_));
 sg13g2_a21oi_1 _19134_ (.A1(_09775_),
    .A2(_09772_),
    .Y(_09776_),
    .B1(net168));
 sg13g2_o21ai_1 _19135_ (.B1(_09776_),
    .Y(_09777_),
    .A1(_09772_),
    .A2(_09775_));
 sg13g2_o21ai_1 _19136_ (.B1(_09777_),
    .Y(_09778_),
    .A1(_06340_),
    .A2(_09768_));
 sg13g2_nand2_1 _19137_ (.Y(_09779_),
    .A(_09778_),
    .B(_09363_));
 sg13g2_o21ai_1 _19138_ (.B1(_09779_),
    .Y(_00502_),
    .A1(_08429_),
    .A2(net144));
 sg13g2_nor2_1 _19139_ (.A(net221),
    .B(_06259_),
    .Y(_09781_));
 sg13g2_nor2_1 _19140_ (.A(_06258_),
    .B(_06295_),
    .Y(_09782_));
 sg13g2_inv_1 _19141_ (.Y(_09783_),
    .A(_09782_));
 sg13g2_nand2b_1 _19142_ (.Y(_09784_),
    .B(_09783_),
    .A_N(_09781_));
 sg13g2_inv_1 _19143_ (.Y(_09785_),
    .A(_09767_));
 sg13g2_a21oi_1 _19144_ (.A1(_09785_),
    .A2(_09765_),
    .Y(_09786_),
    .B1(_09763_));
 sg13g2_xor2_1 _19145_ (.B(_09786_),
    .A(_09784_),
    .X(_09787_));
 sg13g2_nor2_1 _19146_ (.A(_08474_),
    .B(net192),
    .Y(_09788_));
 sg13g2_nand2_1 _19147_ (.Y(_09789_),
    .A(_08474_),
    .B(net192));
 sg13g2_nor2b_1 _19148_ (.A(_09788_),
    .B_N(_09789_),
    .Y(_09791_));
 sg13g2_nand2_1 _19149_ (.Y(_09792_),
    .A(_09739_),
    .B(_09771_));
 sg13g2_a21oi_1 _19150_ (.A1(_09760_),
    .A2(_09740_),
    .Y(_09793_),
    .B1(_09792_));
 sg13g2_nor2_1 _19151_ (.A(_09770_),
    .B(_09793_),
    .Y(_09794_));
 sg13g2_a21oi_1 _19152_ (.A1(_09794_),
    .A2(_09791_),
    .Y(_09795_),
    .B1(net168));
 sg13g2_o21ai_1 _19153_ (.B1(_09795_),
    .Y(_09796_),
    .A1(_09791_),
    .A2(_09794_));
 sg13g2_o21ai_1 _19154_ (.B1(_09796_),
    .Y(_09797_),
    .A1(_06340_),
    .A2(_09787_));
 sg13g2_nand2_1 _19155_ (.Y(_09798_),
    .A(_09797_),
    .B(_09363_));
 sg13g2_o21ai_1 _19156_ (.B1(_09798_),
    .Y(_00503_),
    .A1(_08475_),
    .A2(net144));
 sg13g2_nor2_1 _19157_ (.A(_06251_),
    .B(_06249_),
    .Y(_09799_));
 sg13g2_nor2_1 _19158_ (.A(net224),
    .B(_06255_),
    .Y(_09801_));
 sg13g2_nor2_1 _19159_ (.A(_09799_),
    .B(_09801_),
    .Y(_09802_));
 sg13g2_inv_1 _19160_ (.Y(_09803_),
    .A(_09786_));
 sg13g2_a21oi_1 _19161_ (.A1(_09803_),
    .A2(_09783_),
    .Y(_09804_),
    .B1(_09781_));
 sg13g2_o21ai_1 _19162_ (.B1(net168),
    .Y(_09805_),
    .A1(_09802_),
    .A2(_09804_));
 sg13g2_a21oi_1 _19163_ (.A1(_09802_),
    .A2(_09804_),
    .Y(_09806_),
    .B1(_09805_));
 sg13g2_nor2_1 _19164_ (.A(net127),
    .B(_09806_),
    .Y(_09807_));
 sg13g2_nand2_1 _19165_ (.Y(_09808_),
    .A(_09771_),
    .B(_09789_));
 sg13g2_a21oi_1 _19166_ (.A1(_09775_),
    .A2(_09772_),
    .Y(_09809_),
    .B1(_09808_));
 sg13g2_xor2_1 _19167_ (.B(_06310_),
    .A(_08501_),
    .X(_09810_));
 sg13g2_inv_1 _19168_ (.Y(_09812_),
    .A(_09810_));
 sg13g2_o21ai_1 _19169_ (.B1(_09812_),
    .Y(_09813_),
    .A1(_09788_),
    .A2(_09809_));
 sg13g2_nor2_1 _19170_ (.A(_09788_),
    .B(_09809_),
    .Y(_09814_));
 sg13g2_nand2_1 _19171_ (.Y(_09815_),
    .A(_09814_),
    .B(_09810_));
 sg13g2_nand3_1 _19172_ (.B(net157),
    .C(_09815_),
    .A(_09813_),
    .Y(_09816_));
 sg13g2_a22oi_1 _19173_ (.Y(_00504_),
    .B1(_09807_),
    .B2(_09816_),
    .A2(net113),
    .A1(_08502_));
 sg13g2_nor2_1 _19174_ (.A(net226),
    .B(_06279_),
    .Y(_09817_));
 sg13g2_nor2_1 _19175_ (.A(_06275_),
    .B(_08896_),
    .Y(_09818_));
 sg13g2_inv_1 _19176_ (.Y(_09819_),
    .A(_09818_));
 sg13g2_nand2b_1 _19177_ (.Y(_09820_),
    .B(_09819_),
    .A_N(_09817_));
 sg13g2_nor2_1 _19178_ (.A(_09799_),
    .B(_09804_),
    .Y(_09822_));
 sg13g2_nor2_1 _19179_ (.A(_09801_),
    .B(_09822_),
    .Y(_09823_));
 sg13g2_xor2_1 _19180_ (.B(_09823_),
    .A(_09820_),
    .X(_09824_));
 sg13g2_nor2b_1 _19181_ (.A(_09812_),
    .B_N(_09791_),
    .Y(_09825_));
 sg13g2_o21ai_1 _19182_ (.B1(net180),
    .Y(_09826_),
    .A1(_08474_),
    .A2(_08501_));
 sg13g2_inv_1 _19183_ (.Y(_09827_),
    .A(_09826_));
 sg13g2_a21oi_1 _19184_ (.A1(_09794_),
    .A2(_09825_),
    .Y(_09828_),
    .B1(_09827_));
 sg13g2_xor2_1 _19185_ (.B(_06310_),
    .A(_08539_),
    .X(_09829_));
 sg13g2_inv_1 _19186_ (.Y(_09830_),
    .A(_09829_));
 sg13g2_a21oi_1 _19187_ (.A1(_09828_),
    .A2(_09830_),
    .Y(_09831_),
    .B1(net168));
 sg13g2_o21ai_1 _19188_ (.B1(_09831_),
    .Y(_09833_),
    .A1(_09828_),
    .A2(_09830_));
 sg13g2_o21ai_1 _19189_ (.B1(_09833_),
    .Y(_09834_),
    .A1(_06340_),
    .A2(_09824_));
 sg13g2_nand2_1 _19190_ (.Y(_09835_),
    .A(_09834_),
    .B(_09363_));
 sg13g2_o21ai_1 _19191_ (.B1(_09835_),
    .Y(_00505_),
    .A1(_08540_),
    .A2(net144));
 sg13g2_nor2_1 _19192_ (.A(_06283_),
    .B(_06238_),
    .Y(_09836_));
 sg13g2_nor2_1 _19193_ (.A(net196),
    .B(_06288_),
    .Y(_09837_));
 sg13g2_nor2_1 _19194_ (.A(_09836_),
    .B(_09837_),
    .Y(_09838_));
 sg13g2_inv_1 _19195_ (.Y(_09839_),
    .A(_09823_));
 sg13g2_a21oi_1 _19196_ (.A1(_09839_),
    .A2(_09819_),
    .Y(_09840_),
    .B1(_09817_));
 sg13g2_xnor2_1 _19197_ (.Y(_09841_),
    .A(_09838_),
    .B(_09840_));
 sg13g2_xor2_1 _19198_ (.B(net180),
    .A(_08568_),
    .X(_09843_));
 sg13g2_inv_1 _19199_ (.Y(_09844_),
    .A(_09843_));
 sg13g2_o21ai_1 _19200_ (.B1(net180),
    .Y(_09845_),
    .A1(_08501_),
    .A2(_08539_));
 sg13g2_o21ai_1 _19201_ (.B1(_09845_),
    .Y(_09846_),
    .A1(_09830_),
    .A2(_09815_));
 sg13g2_inv_1 _19202_ (.Y(_09847_),
    .A(_09846_));
 sg13g2_nor2_1 _19203_ (.A(_09844_),
    .B(_09847_),
    .Y(_09848_));
 sg13g2_inv_1 _19204_ (.Y(_09849_),
    .A(_09848_));
 sg13g2_nand2_1 _19205_ (.Y(_09850_),
    .A(_09847_),
    .B(_09844_));
 sg13g2_nand3_1 _19206_ (.B(_09850_),
    .C(_09355_),
    .A(_09849_),
    .Y(_09851_));
 sg13g2_o21ai_1 _19207_ (.B1(_09851_),
    .Y(_09852_),
    .A1(_06340_),
    .A2(_09841_));
 sg13g2_nand2_1 _19208_ (.Y(_09854_),
    .A(_09852_),
    .B(_09363_));
 sg13g2_o21ai_1 _19209_ (.B1(_09854_),
    .Y(_00506_),
    .A1(_08569_),
    .A2(net143));
 sg13g2_nor2_1 _19210_ (.A(_09836_),
    .B(_09840_),
    .Y(_09855_));
 sg13g2_nor2_1 _19211_ (.A(_09837_),
    .B(_09855_),
    .Y(_09856_));
 sg13g2_inv_1 _19212_ (.Y(_09857_),
    .A(_09856_));
 sg13g2_nor2_1 _19213_ (.A(net221),
    .B(_06312_),
    .Y(_09858_));
 sg13g2_nor2_1 _19214_ (.A(net180),
    .B(_06295_),
    .Y(_09859_));
 sg13g2_nor2_1 _19215_ (.A(_09858_),
    .B(_09859_),
    .Y(_09860_));
 sg13g2_inv_1 _19216_ (.Y(_09861_),
    .A(_09860_));
 sg13g2_nand2_1 _19217_ (.Y(_09862_),
    .A(_09857_),
    .B(_09861_));
 sg13g2_nor2_1 _19218_ (.A(_09861_),
    .B(_09857_),
    .Y(_09864_));
 sg13g2_nor2_1 _19219_ (.A(net157),
    .B(_09864_),
    .Y(_09865_));
 sg13g2_xor2_1 _19220_ (.B(net180),
    .A(_08611_),
    .X(_09866_));
 sg13g2_inv_1 _19221_ (.Y(_09867_),
    .A(_09866_));
 sg13g2_nor2_1 _19222_ (.A(_09830_),
    .B(_09844_),
    .Y(_09868_));
 sg13g2_nand3_1 _19223_ (.B(_09825_),
    .C(_09868_),
    .A(_09794_),
    .Y(_09869_));
 sg13g2_o21ai_1 _19224_ (.B1(_08916_),
    .Y(_09870_),
    .A1(_08539_),
    .A2(_08568_));
 sg13g2_inv_1 _19225_ (.Y(_09871_),
    .A(_09870_));
 sg13g2_a21oi_1 _19226_ (.A1(_09868_),
    .A2(_09827_),
    .Y(_09872_),
    .B1(_09871_));
 sg13g2_nand2_1 _19227_ (.Y(_09873_),
    .A(_09869_),
    .B(_09872_));
 sg13g2_xnor2_1 _19228_ (.Y(_09875_),
    .A(_09867_),
    .B(_09873_));
 sg13g2_a221oi_1 _19229_ (.B2(net169),
    .C1(net129),
    .B1(_09875_),
    .A1(_09862_),
    .Y(_09876_),
    .A2(_09865_));
 sg13g2_a21oi_1 _19230_ (.A1(_08612_),
    .A2(net114),
    .Y(_00507_),
    .B1(_09876_));
 sg13g2_nor2_1 _19231_ (.A(_06248_),
    .B(_06312_),
    .Y(_09877_));
 sg13g2_nor2_1 _19232_ (.A(net180),
    .B(_06249_),
    .Y(_09878_));
 sg13g2_nor2_1 _19233_ (.A(_09877_),
    .B(_09878_),
    .Y(_09879_));
 sg13g2_nor2_1 _19234_ (.A(_09859_),
    .B(_09857_),
    .Y(_09880_));
 sg13g2_nor3_1 _19235_ (.A(_09858_),
    .B(_09879_),
    .C(_09880_),
    .Y(_09881_));
 sg13g2_nor2_1 _19236_ (.A(_09858_),
    .B(_09880_),
    .Y(_09882_));
 sg13g2_nor2b_1 _19237_ (.A(_09882_),
    .B_N(_09879_),
    .Y(_09883_));
 sg13g2_nor3_1 _19238_ (.A(net157),
    .B(_09881_),
    .C(_09883_),
    .Y(_09885_));
 sg13g2_nor2_1 _19239_ (.A(net127),
    .B(_09885_),
    .Y(_09886_));
 sg13g2_xor2_1 _19240_ (.B(_08916_),
    .A(_08642_),
    .X(_09887_));
 sg13g2_o21ai_1 _19241_ (.B1(net177),
    .Y(_09888_),
    .A1(_08568_),
    .A2(_08611_));
 sg13g2_inv_1 _19242_ (.Y(_09889_),
    .A(_09888_));
 sg13g2_nor2_1 _19243_ (.A(_09867_),
    .B(_09849_),
    .Y(_09890_));
 sg13g2_nor2_1 _19244_ (.A(_09889_),
    .B(_09890_),
    .Y(_09891_));
 sg13g2_xnor2_1 _19245_ (.Y(_09892_),
    .A(_09887_),
    .B(_09891_));
 sg13g2_nand2_1 _19246_ (.Y(_09893_),
    .A(_09892_),
    .B(net169));
 sg13g2_a22oi_1 _19247_ (.Y(_00508_),
    .B1(_09886_),
    .B2(_09893_),
    .A2(net113),
    .A1(_08678_));
 sg13g2_inv_1 _19248_ (.Y(_09895_),
    .A(_08681_));
 sg13g2_nor2_1 _19249_ (.A(_06244_),
    .B(_06312_),
    .Y(_09896_));
 sg13g2_nor2_1 _19250_ (.A(net177),
    .B(_08896_),
    .Y(_09897_));
 sg13g2_nor2_1 _19251_ (.A(_09896_),
    .B(_09897_),
    .Y(_09898_));
 sg13g2_inv_1 _19252_ (.Y(_09899_),
    .A(_09877_));
 sg13g2_a21oi_1 _19253_ (.A1(_09882_),
    .A2(_09899_),
    .Y(_09900_),
    .B1(_09878_));
 sg13g2_o21ai_1 _19254_ (.B1(_09491_),
    .Y(_09901_),
    .A1(_09898_),
    .A2(_09900_));
 sg13g2_a21oi_1 _19255_ (.A1(_09898_),
    .A2(_09900_),
    .Y(_09902_),
    .B1(_09901_));
 sg13g2_nor2_1 _19256_ (.A(net127),
    .B(_09902_),
    .Y(_09903_));
 sg13g2_xor2_1 _19257_ (.B(net180),
    .A(_08681_),
    .X(_09904_));
 sg13g2_inv_1 _19258_ (.Y(_09906_),
    .A(_09887_));
 sg13g2_nor2_1 _19259_ (.A(_09867_),
    .B(_09906_),
    .Y(_09907_));
 sg13g2_nand2_1 _19260_ (.Y(_09908_),
    .A(_09868_),
    .B(_09907_));
 sg13g2_o21ai_1 _19261_ (.B1(net177),
    .Y(_09909_),
    .A1(_08611_),
    .A2(_08642_));
 sg13g2_inv_1 _19262_ (.Y(_09910_),
    .A(_09909_));
 sg13g2_a21oi_1 _19263_ (.A1(_09907_),
    .A2(_09871_),
    .Y(_09911_),
    .B1(_09910_));
 sg13g2_o21ai_1 _19264_ (.B1(_09911_),
    .Y(_09912_),
    .A1(_09908_),
    .A2(_09828_));
 sg13g2_a21oi_1 _19265_ (.A1(_09912_),
    .A2(_09904_),
    .Y(_09913_),
    .B1(net156));
 sg13g2_o21ai_1 _19266_ (.B1(_09913_),
    .Y(_09914_),
    .A1(_09904_),
    .A2(_09912_));
 sg13g2_a22oi_1 _19267_ (.Y(_00509_),
    .B1(_09903_),
    .B2(_09914_),
    .A2(net113),
    .A1(_09895_));
 sg13g2_xor2_1 _19268_ (.B(_09688_),
    .A(_09665_),
    .X(_09916_));
 sg13g2_nand2_1 _19269_ (.Y(_09917_),
    .A(net128),
    .B(_08701_));
 sg13g2_o21ai_1 _19270_ (.B1(_09917_),
    .Y(_00510_),
    .A1(_09916_),
    .A2(_09607_));
 sg13g2_xnor2_1 _19271_ (.Y(_09918_),
    .A(net196),
    .B(net177));
 sg13g2_nor2_1 _19272_ (.A(_09896_),
    .B(_09883_),
    .Y(_09919_));
 sg13g2_nor2_1 _19273_ (.A(_09897_),
    .B(_09919_),
    .Y(_09920_));
 sg13g2_nor2_1 _19274_ (.A(_09877_),
    .B(_09920_),
    .Y(_09921_));
 sg13g2_xor2_1 _19275_ (.B(_09921_),
    .A(_09918_),
    .X(_09922_));
 sg13g2_xor2_1 _19276_ (.B(net177),
    .A(_08718_),
    .X(_09923_));
 sg13g2_nand2_1 _19277_ (.Y(_09924_),
    .A(_09887_),
    .B(_09904_));
 sg13g2_inv_1 _19278_ (.Y(_09926_),
    .A(_09924_));
 sg13g2_o21ai_1 _19279_ (.B1(net177),
    .Y(_09927_),
    .A1(_08642_),
    .A2(_08681_));
 sg13g2_o21ai_1 _19280_ (.B1(_09927_),
    .Y(_09928_),
    .A1(_09888_),
    .A2(_09924_));
 sg13g2_a21oi_1 _19281_ (.A1(_09890_),
    .A2(_09926_),
    .Y(_09929_),
    .B1(_09928_));
 sg13g2_xnor2_1 _19282_ (.Y(_09930_),
    .A(_09923_),
    .B(_09929_));
 sg13g2_nand2_1 _19283_ (.Y(_09931_),
    .A(_09930_),
    .B(_06340_));
 sg13g2_o21ai_1 _19284_ (.B1(_09931_),
    .Y(_09932_),
    .A1(net169),
    .A2(_09922_));
 sg13g2_mux2_1 _19285_ (.A0(_08718_),
    .A1(_09932_),
    .S(net143),
    .X(_00511_));
 sg13g2_inv_1 _19286_ (.Y(_09933_),
    .A(\vgadonut.donut.ysA[21] ));
 sg13g2_nand2_1 _19287_ (.Y(_09934_),
    .A(_09904_),
    .B(_09923_));
 sg13g2_nor3_1 _19288_ (.A(_09867_),
    .B(_09906_),
    .C(_09934_),
    .Y(_09936_));
 sg13g2_o21ai_1 _19289_ (.B1(_08917_),
    .Y(_09937_),
    .A1(_08681_),
    .A2(_08718_));
 sg13g2_o21ai_1 _19290_ (.B1(_09937_),
    .Y(_09938_),
    .A1(_09909_),
    .A2(_09934_));
 sg13g2_a21oi_1 _19291_ (.A1(_09873_),
    .A2(_09936_),
    .Y(_09939_),
    .B1(_09938_));
 sg13g2_xnor2_1 _19292_ (.Y(_09940_),
    .A(\vgadonut.donut.ysA[21] ),
    .B(_08917_));
 sg13g2_a21oi_1 _19293_ (.A1(_09939_),
    .A2(_09940_),
    .Y(_09941_),
    .B1(net156));
 sg13g2_o21ai_1 _19294_ (.B1(_09941_),
    .Y(_09942_),
    .A1(_09939_),
    .A2(_09940_));
 sg13g2_a22oi_1 _19295_ (.Y(_09943_),
    .B1(_09898_),
    .B2(_09900_),
    .A2(net177),
    .A1(_06238_));
 sg13g2_a21oi_1 _19296_ (.A1(net196),
    .A2(_06312_),
    .Y(_09944_),
    .B1(_09943_));
 sg13g2_nor3_1 _19297_ (.A(net159),
    .B(_09896_),
    .C(_09944_),
    .Y(_09945_));
 sg13g2_nor2_1 _19298_ (.A(net128),
    .B(_09945_),
    .Y(_09947_));
 sg13g2_a22oi_1 _19299_ (.Y(_00512_),
    .B1(_09942_),
    .B2(_09947_),
    .A2(_09659_),
    .A1(_09933_));
 sg13g2_xnor2_1 _19300_ (.Y(_09948_),
    .A(_09695_),
    .B(_09691_));
 sg13g2_nand2_1 _19301_ (.Y(_09949_),
    .A(net128),
    .B(_08341_));
 sg13g2_o21ai_1 _19302_ (.B1(_09949_),
    .Y(_00513_),
    .A1(_09948_),
    .A2(_09607_));
 sg13g2_a21oi_1 _19303_ (.A1(_09742_),
    .A2(_09743_),
    .Y(_09950_),
    .B1(_06978_));
 sg13g2_o21ai_1 _19304_ (.B1(_09950_),
    .Y(_09951_),
    .A1(_09743_),
    .A2(_09742_));
 sg13g2_o21ai_1 _19305_ (.B1(_09951_),
    .Y(_00514_),
    .A1(_08331_),
    .A2(_09420_));
 sg13g2_xnor2_1 _19306_ (.Y(_09952_),
    .A(_09700_),
    .B(_09699_));
 sg13g2_a22oi_1 _19307_ (.Y(_09953_),
    .B1(net157),
    .B2(_09952_),
    .A2(_09668_),
    .A1(_06978_));
 sg13g2_a21o_1 _19308_ (.A2(net128),
    .A1(_08317_),
    .B1(_09953_),
    .X(_00515_));
 sg13g2_a21oi_1 _19309_ (.A1(_08856_),
    .A2(net158),
    .Y(_09955_),
    .B1(net129));
 sg13g2_a21oi_1 _19310_ (.A1(_09746_),
    .A2(_09747_),
    .Y(_09956_),
    .B1(net156));
 sg13g2_o21ai_1 _19311_ (.B1(_09956_),
    .Y(_09957_),
    .A1(_09747_),
    .A2(_09746_));
 sg13g2_a22oi_1 _19312_ (.Y(_00516_),
    .B1(_09955_),
    .B2(_09957_),
    .A2(net113),
    .A1(_08306_));
 sg13g2_inv_1 _19313_ (.Y(_09958_),
    .A(_08298_));
 sg13g2_a21oi_1 _19314_ (.A1(_08821_),
    .A2(net158),
    .Y(_09959_),
    .B1(net129));
 sg13g2_a21oi_1 _19315_ (.A1(_09706_),
    .A2(_09709_),
    .Y(_09960_),
    .B1(net156));
 sg13g2_o21ai_1 _19316_ (.B1(_09960_),
    .Y(_09961_),
    .A1(_09709_),
    .A2(_09706_));
 sg13g2_a22oi_1 _19317_ (.Y(_00517_),
    .B1(_09959_),
    .B2(_09961_),
    .A2(net113),
    .A1(_09958_));
 sg13g2_xnor2_1 _19318_ (.Y(_09963_),
    .A(_09752_),
    .B(_09751_));
 sg13g2_o21ai_1 _19319_ (.B1(_06975_),
    .Y(_09964_),
    .A1(_06027_),
    .A2(_09355_));
 sg13g2_a21oi_1 _19320_ (.A1(_09963_),
    .A2(net157),
    .Y(_09965_),
    .B1(_09964_));
 sg13g2_a21o_1 _19321_ (.A2(net128),
    .A1(_08245_),
    .B1(_09965_),
    .X(_00518_));
 sg13g2_xor2_1 _19322_ (.B(_08851_),
    .A(net194),
    .X(_09966_));
 sg13g2_a21oi_1 _19323_ (.A1(_09491_),
    .A2(_09966_),
    .Y(_09967_),
    .B1(net129));
 sg13g2_a21oi_1 _19324_ (.A1(_09713_),
    .A2(_09717_),
    .Y(_09968_),
    .B1(net156));
 sg13g2_o21ai_1 _19325_ (.B1(_09968_),
    .Y(_09969_),
    .A1(_09717_),
    .A2(_09713_));
 sg13g2_a22oi_1 _19326_ (.Y(_00519_),
    .B1(_09967_),
    .B2(_09969_),
    .A2(net113),
    .A1(_08250_));
 sg13g2_xnor2_1 _19327_ (.Y(_09970_),
    .A(_09675_),
    .B(_09676_));
 sg13g2_a21oi_1 _19328_ (.A1(net158),
    .A2(_09970_),
    .Y(_09972_),
    .B1(net129));
 sg13g2_a21oi_1 _19329_ (.A1(_09755_),
    .A2(_09756_),
    .Y(_09973_),
    .B1(net156));
 sg13g2_o21ai_1 _19330_ (.B1(_09973_),
    .Y(_09974_),
    .A1(_09756_),
    .A2(_09755_));
 sg13g2_a22oi_1 _19331_ (.Y(_00520_),
    .B1(_09972_),
    .B2(_09974_),
    .A2(net113),
    .A1(_08264_));
 sg13g2_nor2_1 _19332_ (.A(_05970_),
    .B(_09355_),
    .Y(_09975_));
 sg13g2_inv_1 _19333_ (.Y(_09976_),
    .A(_09975_));
 sg13g2_nor2_1 _19334_ (.A(_10004_),
    .B(_09976_),
    .Y(_09977_));
 sg13g2_mux2_1 _19335_ (.A0(_09811_),
    .A1(_00184_),
    .S(_09977_),
    .X(_00521_));
 sg13g2_nand2_1 _19336_ (.Y(_09978_),
    .A(_09977_),
    .B(_09811_));
 sg13g2_xnor2_1 _19337_ (.Y(_00522_),
    .A(\vgadonut.frame[1] ),
    .B(_09978_));
 sg13g2_inv_1 _19338_ (.Y(_09980_),
    .A(\vgadonut.frame[2] ));
 sg13g2_inv_1 _19339_ (.Y(_09981_),
    .A(\vgadonut.frame[1] ));
 sg13g2_nor2_1 _19340_ (.A(_09981_),
    .B(_09978_),
    .Y(_09982_));
 sg13g2_xnor2_1 _19341_ (.Y(_00523_),
    .A(_09980_),
    .B(_09982_));
 sg13g2_inv_1 _19342_ (.Y(_09983_),
    .A(\vgadonut.frame[3] ));
 sg13g2_inv_1 _19343_ (.Y(_09984_),
    .A(_09982_));
 sg13g2_nor2_1 _19344_ (.A(_09980_),
    .B(_09984_),
    .Y(_09985_));
 sg13g2_xnor2_1 _19345_ (.Y(_00524_),
    .A(_09983_),
    .B(_09985_));
 sg13g2_inv_1 _19346_ (.Y(_09986_),
    .A(\vgadonut.frame[4] ));
 sg13g2_nor3_1 _19347_ (.A(_09983_),
    .B(_09980_),
    .C(_09984_),
    .Y(_09987_));
 sg13g2_xnor2_1 _19348_ (.Y(_00525_),
    .A(_09986_),
    .B(_09987_));
 sg13g2_buf_1 _19349_ (.A(\vgadonut.frame[5] ),
    .X(_09989_));
 sg13g2_nand2_1 _19350_ (.Y(_09990_),
    .A(_09987_),
    .B(\vgadonut.frame[4] ));
 sg13g2_xnor2_1 _19351_ (.Y(_00526_),
    .A(_09989_),
    .B(_09990_));
 sg13g2_buf_1 _19352_ (.A(\vgadonut.frame[6] ),
    .X(_09991_));
 sg13g2_inv_1 _19353_ (.Y(_09992_),
    .A(_09991_));
 sg13g2_inv_1 _19354_ (.Y(_09993_),
    .A(_09989_));
 sg13g2_nor2_1 _19355_ (.A(_09993_),
    .B(_09990_),
    .Y(_09994_));
 sg13g2_xnor2_1 _19356_ (.Y(_00527_),
    .A(_09992_),
    .B(_09994_));
 sg13g2_nand2_1 _19357_ (.Y(_09995_),
    .A(_09994_),
    .B(_09991_));
 sg13g2_xnor2_1 _19358_ (.Y(_00528_),
    .A(\vgadonut.frame[7] ),
    .B(_09995_));
 sg13g2_nand3_1 _19359_ (.B(net159),
    .C(_00096_),
    .A(_05971_),
    .Y(_09997_));
 sg13g2_o21ai_1 _19360_ (.B1(_09997_),
    .Y(_00533_),
    .A1(_09863_),
    .A2(_05994_));
 sg13g2_nand2_1 _19361_ (.Y(_09998_),
    .A(_09894_),
    .B(_09832_));
 sg13g2_nand2_1 _19362_ (.Y(_09999_),
    .A(_06218_),
    .B(_09998_));
 sg13g2_nor2_1 _19363_ (.A(_09894_),
    .B(_05971_),
    .Y(_10000_));
 sg13g2_a21oi_1 _19364_ (.A1(_05971_),
    .A2(_09999_),
    .Y(_00534_),
    .B1(_10000_));
 sg13g2_nor2_1 _19365_ (.A(_09998_),
    .B(_05976_),
    .Y(_10001_));
 sg13g2_nor2_1 _19366_ (.A(_06000_),
    .B(_10001_),
    .Y(_10002_));
 sg13g2_inv_1 _19367_ (.Y(_10003_),
    .A(_06000_));
 sg13g2_inv_1 _19368_ (.Y(_10005_),
    .A(_10001_));
 sg13g2_nor2_1 _19369_ (.A(_10003_),
    .B(_10005_),
    .Y(_10006_));
 sg13g2_nor3_1 _19370_ (.A(_09975_),
    .B(_10002_),
    .C(_10006_),
    .Y(_00535_));
 sg13g2_nor2_1 _19371_ (.A(_06215_),
    .B(_10005_),
    .Y(_10007_));
 sg13g2_nor2_1 _19372_ (.A(_06002_),
    .B(_10006_),
    .Y(_10008_));
 sg13g2_nor3_1 _19373_ (.A(_09975_),
    .B(_10007_),
    .C(_10008_),
    .Y(_00536_));
 sg13g2_xnor2_1 _19374_ (.Y(_00537_),
    .A(_06214_),
    .B(_10007_));
 sg13g2_inv_1 _19375_ (.Y(_10009_),
    .A(_10007_));
 sg13g2_nor2_1 _19376_ (.A(_06214_),
    .B(_10009_),
    .Y(_10010_));
 sg13g2_xnor2_1 _19377_ (.Y(_00538_),
    .A(_06005_),
    .B(_10010_));
 sg13g2_nand2_1 _19378_ (.Y(_10012_),
    .A(_06004_),
    .B(_06009_));
 sg13g2_nor4_1 _19379_ (.A(_06337_),
    .B(_06215_),
    .C(_10012_),
    .D(_10005_),
    .Y(_10013_));
 sg13g2_nor2_1 _19380_ (.A(_10012_),
    .B(_10009_),
    .Y(_10014_));
 sg13g2_nor2_1 _19381_ (.A(_06008_),
    .B(_10014_),
    .Y(_10015_));
 sg13g2_nor2_1 _19382_ (.A(_10013_),
    .B(_10015_),
    .Y(_00539_));
 sg13g2_nand2_1 _19383_ (.Y(_10016_),
    .A(_10014_),
    .B(_06008_));
 sg13g2_o21ai_1 _19384_ (.B1(_09976_),
    .Y(_10017_),
    .A1(_06336_),
    .A2(_10016_));
 sg13g2_a21oi_1 _19385_ (.A1(_06336_),
    .A2(_10016_),
    .Y(_00540_),
    .B1(_10017_));
 sg13g2_nor3_1 _19386_ (.A(_06336_),
    .B(_06337_),
    .C(_06010_),
    .Y(_10018_));
 sg13g2_nand2_1 _19387_ (.Y(_10019_),
    .A(_10013_),
    .B(_06007_));
 sg13g2_a221oi_1 _19388_ (.B2(_06010_),
    .C1(_09975_),
    .B1(_10019_),
    .A1(_10014_),
    .Y(_00541_),
    .A2(_10018_));
 sg13g2_inv_1 _19389_ (.Y(_10021_),
    .A(\vgadonut.donut.v_count[9] ));
 sg13g2_nor4_1 _19390_ (.A(_06001_),
    .B(_00096_),
    .C(_06215_),
    .D(_10012_),
    .Y(_10022_));
 sg13g2_nand3_1 _19391_ (.B(_10018_),
    .C(_10022_),
    .A(_05977_),
    .Y(_10023_));
 sg13g2_xnor2_1 _19392_ (.Y(_10024_),
    .A(_10021_),
    .B(_10023_));
 sg13g2_a21oi_1 _19393_ (.A1(_05977_),
    .A2(_09491_),
    .Y(_00542_),
    .B1(_10024_));
 sg13g2_nand2_1 _19394_ (.Y(_10025_),
    .A(_03937_),
    .B(_03809_));
 sg13g2_inv_1 _19395_ (.Y(_10026_),
    .A(_10025_));
 sg13g2_inv_1 _19396_ (.Y(_10027_),
    .A(_03937_));
 sg13g2_a21oi_1 _19397_ (.A1(_10027_),
    .A2(_03954_),
    .Y(_10028_),
    .B1(_03818_));
 sg13g2_nor2_1 _19398_ (.A(_10026_),
    .B(_10028_),
    .Y(_10030_));
 sg13g2_o21ai_1 _19399_ (.B1(_10030_),
    .Y(_10031_),
    .A1(_03938_),
    .A2(_04009_));
 sg13g2_buf_1 _19400_ (.A(net52),
    .X(_10032_));
 sg13g2_buf_1 _19401_ (.A(_03792_),
    .X(_10033_));
 sg13g2_mux2_1 _19402_ (.A0(_03915_),
    .A1(_03911_),
    .S(net43),
    .X(_10034_));
 sg13g2_xnor2_1 _19403_ (.Y(_10035_),
    .A(_10032_),
    .B(_10034_));
 sg13g2_a21oi_1 _19404_ (.A1(_03768_),
    .A2(_03802_),
    .Y(_10036_),
    .B1(_03805_));
 sg13g2_a21oi_1 _19405_ (.A1(_03918_),
    .A2(_03907_),
    .Y(_10037_),
    .B1(_03928_));
 sg13g2_o21ai_1 _19406_ (.B1(_10037_),
    .Y(_10038_),
    .A1(_03810_),
    .A2(_10036_));
 sg13g2_nand2_1 _19407_ (.Y(_10039_),
    .A(_10038_),
    .B(_03920_));
 sg13g2_xnor2_1 _19408_ (.Y(_10041_),
    .A(_10035_),
    .B(_10039_));
 sg13g2_xnor2_1 _19409_ (.Y(_10042_),
    .A(_03808_),
    .B(_10041_));
 sg13g2_nand2_1 _19410_ (.Y(_10043_),
    .A(_10042_),
    .B(_03936_));
 sg13g2_inv_1 _19411_ (.Y(_10044_),
    .A(_10043_));
 sg13g2_or2_1 _19412_ (.X(_10045_),
    .B(_10042_),
    .A(_03936_));
 sg13g2_nor2b_1 _19413_ (.A(_10044_),
    .B_N(_10045_),
    .Y(_10046_));
 sg13g2_nand2_1 _19414_ (.Y(_10047_),
    .A(_10031_),
    .B(_10046_));
 sg13g2_a21oi_1 _19415_ (.A1(_03480_),
    .A2(_03494_),
    .Y(_10048_),
    .B1(_10033_));
 sg13g2_nand3_1 _19416_ (.B(_03418_),
    .C(_10033_),
    .A(_03417_),
    .Y(_10049_));
 sg13g2_nand2b_1 _19417_ (.Y(_10050_),
    .B(_10049_),
    .A_N(_10048_));
 sg13g2_o21ai_1 _19418_ (.B1(_03929_),
    .Y(_10052_),
    .A1(_03810_),
    .A2(_03731_));
 sg13g2_nand2_1 _19419_ (.Y(_10053_),
    .A(_10052_),
    .B(_03920_));
 sg13g2_nand2_1 _19420_ (.Y(_10054_),
    .A(_10053_),
    .B(_03921_));
 sg13g2_mux2_1 _19421_ (.A0(_10032_),
    .A1(_10034_),
    .S(_10054_),
    .X(_10055_));
 sg13g2_xnor2_1 _19422_ (.Y(_10056_),
    .A(_10050_),
    .B(_10055_));
 sg13g2_xor2_1 _19423_ (.B(_10056_),
    .A(_03933_),
    .X(_10057_));
 sg13g2_nand2_1 _19424_ (.Y(_10058_),
    .A(_10041_),
    .B(_03808_));
 sg13g2_nand2b_1 _19425_ (.Y(_10059_),
    .B(_10058_),
    .A_N(_10057_));
 sg13g2_nand3_1 _19426_ (.B(_10059_),
    .C(_10043_),
    .A(_10047_),
    .Y(_10060_));
 sg13g2_nand2b_1 _19427_ (.Y(_10061_),
    .B(_10057_),
    .A_N(_10058_));
 sg13g2_nand2_1 _19428_ (.Y(_10063_),
    .A(_10060_),
    .B(_10061_));
 sg13g2_inv_1 _19429_ (.Y(_10064_),
    .A(_10041_));
 sg13g2_nor2_1 _19430_ (.A(_03933_),
    .B(_10064_),
    .Y(_10065_));
 sg13g2_a21o_1 _19431_ (.A2(_10065_),
    .A1(_10063_),
    .B1(_10056_),
    .X(_10066_));
 sg13g2_nor2_1 _19432_ (.A(\vgadonut.donut.donuthit.t[15] ),
    .B(_10066_),
    .Y(_10067_));
 sg13g2_and2_1 _19433_ (.A(_10066_),
    .B(\vgadonut.donut.donuthit.t[15] ),
    .X(_10068_));
 sg13g2_nor2_1 _19434_ (.A(_10067_),
    .B(_10068_),
    .Y(_10069_));
 sg13g2_nor2b_1 _19435_ (.A(_10056_),
    .B_N(_03933_),
    .Y(_10070_));
 sg13g2_xnor2_1 _19436_ (.Y(_10071_),
    .A(_10064_),
    .B(_10070_));
 sg13g2_inv_1 _19437_ (.Y(_10072_),
    .A(_10071_));
 sg13g2_nand2b_1 _19438_ (.Y(_10074_),
    .B(_10046_),
    .A_N(_03957_));
 sg13g2_a21oi_1 _19439_ (.A1(_10045_),
    .A2(_10026_),
    .Y(_10075_),
    .B1(_10044_));
 sg13g2_nand2_1 _19440_ (.Y(_10076_),
    .A(_10074_),
    .B(_10075_));
 sg13g2_nand2b_1 _19441_ (.Y(_10077_),
    .B(_10059_),
    .A_N(_10076_));
 sg13g2_nand2_1 _19442_ (.Y(_10078_),
    .A(_10077_),
    .B(_10061_));
 sg13g2_nand2_1 _19443_ (.Y(_10079_),
    .A(_10056_),
    .B(_10064_));
 sg13g2_o21ai_1 _19444_ (.B1(_10079_),
    .Y(_10080_),
    .A1(_10072_),
    .A2(_10078_));
 sg13g2_nand2b_1 _19445_ (.Y(_10081_),
    .B(_10041_),
    .A_N(_10056_));
 sg13g2_nand2_1 _19446_ (.Y(_10082_),
    .A(_10080_),
    .B(_10081_));
 sg13g2_nor2_1 _19447_ (.A(_03933_),
    .B(_10081_),
    .Y(_10083_));
 sg13g2_nand2_1 _19448_ (.Y(_10085_),
    .A(_10078_),
    .B(_10083_));
 sg13g2_nand2_1 _19449_ (.Y(_10086_),
    .A(_10082_),
    .B(_10085_));
 sg13g2_xnor2_1 _19450_ (.Y(_10087_),
    .A(\vgadonut.donut.donuthit.t[14] ),
    .B(_10086_));
 sg13g2_xnor2_1 _19451_ (.Y(_10088_),
    .A(_10072_),
    .B(_10063_));
 sg13g2_inv_1 _19452_ (.Y(_10089_),
    .A(\vgadonut.donut.donuthit.t[13] ));
 sg13g2_nand2_1 _19453_ (.Y(_10090_),
    .A(_10088_),
    .B(_10089_));
 sg13g2_nand2b_1 _19454_ (.Y(_10091_),
    .B(_10090_),
    .A_N(_10087_));
 sg13g2_inv_1 _19455_ (.Y(_10092_),
    .A(\vgadonut.donut.donuthit.t[11] ));
 sg13g2_xnor2_1 _19456_ (.Y(_10093_),
    .A(_10046_),
    .B(_10031_));
 sg13g2_nor2_1 _19457_ (.A(_10092_),
    .B(_10093_),
    .Y(_10094_));
 sg13g2_nand2_1 _19458_ (.Y(_10096_),
    .A(_04007_),
    .B(\vgadonut.donut.donuthit.t[9] ));
 sg13g2_inv_1 _19459_ (.Y(_10097_),
    .A(\vgadonut.donut.donuthit.t[10] ));
 sg13g2_nor2_1 _19460_ (.A(_10097_),
    .B(_04139_),
    .Y(_10098_));
 sg13g2_inv_1 _19461_ (.Y(_10099_),
    .A(_10098_));
 sg13g2_nand2_1 _19462_ (.Y(_10100_),
    .A(_10096_),
    .B(_10099_));
 sg13g2_xnor2_1 _19463_ (.Y(_10101_),
    .A(\vgadonut.donut.donuthit.t[3] ),
    .B(_04018_));
 sg13g2_inv_1 _19464_ (.Y(_10102_),
    .A(\vgadonut.donut.donuthit.t[2] ));
 sg13g2_nor2_1 _19465_ (.A(_10102_),
    .B(_04052_),
    .Y(_10103_));
 sg13g2_inv_1 _19466_ (.Y(_10104_),
    .A(\vgadonut.donut.donuthit.t[1] ));
 sg13g2_nor2_1 _19467_ (.A(_10104_),
    .B(_04073_),
    .Y(_10105_));
 sg13g2_xnor2_1 _19468_ (.Y(_10107_),
    .A(_10104_),
    .B(_04073_));
 sg13g2_inv_1 _19469_ (.Y(_10108_),
    .A(\vgadonut.donut.donuthit.t[0] ));
 sg13g2_nor2_1 _19470_ (.A(_10108_),
    .B(_04082_),
    .Y(_10109_));
 sg13g2_nand2b_1 _19471_ (.Y(_10110_),
    .B(_10109_),
    .A_N(_10107_));
 sg13g2_nor2b_1 _19472_ (.A(_10105_),
    .B_N(_10110_),
    .Y(_10111_));
 sg13g2_xnor2_1 _19473_ (.Y(_10112_),
    .A(_10102_),
    .B(_04052_));
 sg13g2_or2_1 _19474_ (.X(_10113_),
    .B(_10112_),
    .A(_10111_));
 sg13g2_nor2b_1 _19475_ (.A(_10103_),
    .B_N(_10113_),
    .Y(_10114_));
 sg13g2_inv_1 _19476_ (.Y(_10115_),
    .A(_10114_));
 sg13g2_nand2b_1 _19477_ (.Y(_10116_),
    .B(_10115_),
    .A_N(_10101_));
 sg13g2_nand2_1 _19478_ (.Y(_10118_),
    .A(_04018_),
    .B(\vgadonut.donut.donuthit.t[3] ));
 sg13g2_nand2_1 _19479_ (.Y(_10119_),
    .A(_10116_),
    .B(_10118_));
 sg13g2_xor2_1 _19480_ (.B(_03979_),
    .A(\vgadonut.donut.donuthit.t[4] ),
    .X(_10120_));
 sg13g2_nand2_1 _19481_ (.Y(_10121_),
    .A(_10119_),
    .B(_10120_));
 sg13g2_nand2_1 _19482_ (.Y(_10122_),
    .A(_03979_),
    .B(\vgadonut.donut.donuthit.t[4] ));
 sg13g2_nand2_1 _19483_ (.Y(_10123_),
    .A(_10121_),
    .B(_10122_));
 sg13g2_xor2_1 _19484_ (.B(_03974_),
    .A(\vgadonut.donut.donuthit.t[5] ),
    .X(_10124_));
 sg13g2_nand2_1 _19485_ (.Y(_10125_),
    .A(_10123_),
    .B(_10124_));
 sg13g2_nand2_1 _19486_ (.Y(_10126_),
    .A(_03974_),
    .B(\vgadonut.donut.donuthit.t[5] ));
 sg13g2_nand2_1 _19487_ (.Y(_10127_),
    .A(_10125_),
    .B(_10126_));
 sg13g2_xnor2_1 _19488_ (.Y(_10129_),
    .A(\vgadonut.donut.donuthit.t[6] ),
    .B(_03985_));
 sg13g2_nand2_1 _19489_ (.Y(_10130_),
    .A(_10127_),
    .B(_10129_));
 sg13g2_nand2_1 _19490_ (.Y(_10131_),
    .A(_04068_),
    .B(\vgadonut.donut.donuthit.t[6] ));
 sg13g2_nand2_1 _19491_ (.Y(_10132_),
    .A(_10130_),
    .B(_10131_));
 sg13g2_nand2b_1 _19492_ (.Y(_10133_),
    .B(_03993_),
    .A_N(\vgadonut.donut.donuthit.t[7] ));
 sg13g2_nand2_1 _19493_ (.Y(_10134_),
    .A(_10132_),
    .B(_10133_));
 sg13g2_nand2_1 _19494_ (.Y(_10135_),
    .A(_03992_),
    .B(\vgadonut.donut.donuthit.t[7] ));
 sg13g2_nand2_1 _19495_ (.Y(_10136_),
    .A(_10134_),
    .B(_10135_));
 sg13g2_or2_1 _19496_ (.X(_10137_),
    .B(_04000_),
    .A(\vgadonut.donut.donuthit.t[8] ));
 sg13g2_nand2_1 _19497_ (.Y(_10138_),
    .A(_10136_),
    .B(_10137_));
 sg13g2_nand2_1 _19498_ (.Y(_10140_),
    .A(_04000_),
    .B(\vgadonut.donut.donuthit.t[8] ));
 sg13g2_nand2b_1 _19499_ (.Y(_10141_),
    .B(_04011_),
    .A_N(\vgadonut.donut.donuthit.t[9] ));
 sg13g2_nand2_1 _19500_ (.Y(_10142_),
    .A(_10096_),
    .B(_10141_));
 sg13g2_a21oi_1 _19501_ (.A1(_10138_),
    .A2(_10140_),
    .Y(_10143_),
    .B1(_10142_));
 sg13g2_nand2_1 _19502_ (.Y(_10144_),
    .A(_04139_),
    .B(_10097_));
 sg13g2_o21ai_1 _19503_ (.B1(_10144_),
    .Y(_10145_),
    .A1(_10100_),
    .A2(_10143_));
 sg13g2_nand2_1 _19504_ (.Y(_10146_),
    .A(_10093_),
    .B(_10092_));
 sg13g2_nor2b_1 _19505_ (.A(_10094_),
    .B_N(_10146_),
    .Y(_10147_));
 sg13g2_nand2b_1 _19506_ (.Y(_10148_),
    .B(_10147_),
    .A_N(_10145_));
 sg13g2_nand2_1 _19507_ (.Y(_10149_),
    .A(_10059_),
    .B(_10061_));
 sg13g2_xnor2_1 _19508_ (.Y(_10151_),
    .A(_10076_),
    .B(_10149_));
 sg13g2_nand2_1 _19509_ (.Y(_10152_),
    .A(_10151_),
    .B(\vgadonut.donut.donuthit.t[12] ));
 sg13g2_nand3b_1 _19510_ (.B(_10148_),
    .C(_10152_),
    .Y(_10153_),
    .A_N(_10094_));
 sg13g2_or2_1 _19511_ (.X(_10154_),
    .B(_10151_),
    .A(\vgadonut.donut.donuthit.t[12] ));
 sg13g2_buf_1 _19512_ (.A(_10154_),
    .X(_10155_));
 sg13g2_nor2_1 _19513_ (.A(_10089_),
    .B(_10088_),
    .Y(_10156_));
 sg13g2_a21oi_1 _19514_ (.A1(_10153_),
    .A2(_10155_),
    .Y(_10157_),
    .B1(_10156_));
 sg13g2_nand2_1 _19515_ (.Y(_10158_),
    .A(_10086_),
    .B(\vgadonut.donut.donuthit.t[14] ));
 sg13g2_o21ai_1 _19516_ (.B1(_10158_),
    .Y(_10159_),
    .A1(_10091_),
    .A2(_10157_));
 sg13g2_xnor2_1 _19517_ (.Y(_10160_),
    .A(_10069_),
    .B(_10159_));
 sg13g2_nand2_1 _19518_ (.Y(_10162_),
    .A(_10155_),
    .B(_10152_));
 sg13g2_nand3_1 _19519_ (.B(_10140_),
    .C(_10096_),
    .A(_10138_),
    .Y(_10163_));
 sg13g2_nand4_1 _19520_ (.B(_10144_),
    .C(_10141_),
    .A(_10163_),
    .Y(_10164_),
    .D(_10099_));
 sg13g2_nand2b_1 _19521_ (.Y(_10165_),
    .B(_10147_),
    .A_N(_10164_));
 sg13g2_a21oi_1 _19522_ (.A1(_10146_),
    .A2(_10098_),
    .Y(_10166_),
    .B1(_10094_));
 sg13g2_nand2_1 _19523_ (.Y(_10167_),
    .A(_10165_),
    .B(_10166_));
 sg13g2_nand2b_1 _19524_ (.Y(_10168_),
    .B(_10167_),
    .A_N(_10162_));
 sg13g2_inv_1 _19525_ (.Y(_10169_),
    .A(_10156_));
 sg13g2_nand3_1 _19526_ (.B(_10169_),
    .C(_10152_),
    .A(_10168_),
    .Y(_10170_));
 sg13g2_nand3b_1 _19527_ (.B(_10170_),
    .C(_10090_),
    .Y(_10171_),
    .A_N(_10087_));
 sg13g2_buf_1 _19528_ (.A(_10171_),
    .X(_10173_));
 sg13g2_nand2_1 _19529_ (.Y(_10174_),
    .A(_10170_),
    .B(_10090_));
 sg13g2_nand2_1 _19530_ (.Y(_10175_),
    .A(_10174_),
    .B(_10087_));
 sg13g2_nand2_1 _19531_ (.Y(_10176_),
    .A(_10169_),
    .B(_10090_));
 sg13g2_nand2_1 _19532_ (.Y(_10177_),
    .A(_10153_),
    .B(_10155_));
 sg13g2_xnor2_1 _19533_ (.Y(_10178_),
    .A(_10176_),
    .B(_10177_));
 sg13g2_xnor2_1 _19534_ (.Y(_10179_),
    .A(_10147_),
    .B(_10145_));
 sg13g2_xnor2_1 _19535_ (.Y(_10180_),
    .A(_10162_),
    .B(_10167_));
 sg13g2_nor2_1 _19536_ (.A(_10179_),
    .B(_10180_),
    .Y(_10181_));
 sg13g2_nand2_1 _19537_ (.Y(_10182_),
    .A(_10178_),
    .B(_10181_));
 sg13g2_a21oi_1 _19538_ (.A1(_10173_),
    .A2(_10175_),
    .Y(_10184_),
    .B1(_10182_));
 sg13g2_nand2_1 _19539_ (.Y(_10185_),
    .A(_10160_),
    .B(_10184_));
 sg13g2_a21oi_1 _19540_ (.A1(_10086_),
    .A2(\vgadonut.donut.donuthit.t[14] ),
    .Y(_10186_),
    .B1(_10067_));
 sg13g2_a21oi_1 _19541_ (.A1(_10173_),
    .A2(_10186_),
    .Y(_10187_),
    .B1(_10068_));
 sg13g2_nand2_1 _19542_ (.Y(_10188_),
    .A(_10185_),
    .B(_10187_));
 sg13g2_nand2_1 _19543_ (.Y(_10189_),
    .A(_10188_),
    .B(\vgadonut.donut.donuthit.hit ));
 sg13g2_nand2_1 _19544_ (.Y(_00297_),
    .A(_10189_),
    .B(_06918_));
 sg13g2_nor2_1 _19545_ (.A(\vgadonut.donut.donuthit.t[0] ),
    .B(_04080_),
    .Y(_10190_));
 sg13g2_nor3_1 _19546_ (.A(net110),
    .B(_10190_),
    .C(_10109_),
    .Y(_00331_));
 sg13g2_a22oi_1 _19547_ (.Y(_10191_),
    .B1(_10141_),
    .B2(_10163_),
    .A2(_10099_),
    .A1(_10144_));
 sg13g2_nand2_1 _19548_ (.Y(_10193_),
    .A(_10164_),
    .B(net120));
 sg13g2_nor2_1 _19549_ (.A(_10191_),
    .B(_10193_),
    .Y(_00332_));
 sg13g2_nor2b_1 _19550_ (.A(net110),
    .B_N(_10179_),
    .Y(_00333_));
 sg13g2_nor2b_1 _19551_ (.A(net110),
    .B_N(_10180_),
    .Y(_00334_));
 sg13g2_nor2_1 _19552_ (.A(net110),
    .B(_10178_),
    .Y(_00335_));
 sg13g2_and3_1 _19553_ (.X(_00336_),
    .A(_10173_),
    .B(_10175_),
    .C(_04741_));
 sg13g2_nor2_1 _19554_ (.A(_04667_),
    .B(_10160_),
    .Y(_00337_));
 sg13g2_inv_1 _19555_ (.Y(_10194_),
    .A(_10109_));
 sg13g2_nand2_1 _19556_ (.Y(_10195_),
    .A(_10110_),
    .B(net116));
 sg13g2_a21oi_1 _19557_ (.A1(_10194_),
    .A2(_10107_),
    .Y(_00338_),
    .B1(_10195_));
 sg13g2_nand2_1 _19558_ (.Y(_10197_),
    .A(_10113_),
    .B(_06959_));
 sg13g2_a21oi_1 _19559_ (.A1(_10111_),
    .A2(_10112_),
    .Y(_00339_),
    .B1(_10197_));
 sg13g2_nand2_1 _19560_ (.Y(_10198_),
    .A(_10116_),
    .B(_06959_));
 sg13g2_a21oi_1 _19561_ (.A1(_10101_),
    .A2(_10114_),
    .Y(_00340_),
    .B1(_10198_));
 sg13g2_nor2_1 _19562_ (.A(_10120_),
    .B(_10119_),
    .Y(_10199_));
 sg13g2_nand2_1 _19563_ (.Y(_10200_),
    .A(_10121_),
    .B(net120));
 sg13g2_nor2_1 _19564_ (.A(_10199_),
    .B(_10200_),
    .Y(_00341_));
 sg13g2_nor2_1 _19565_ (.A(_10124_),
    .B(_10123_),
    .Y(_10201_));
 sg13g2_nand2_1 _19566_ (.Y(_10202_),
    .A(_10125_),
    .B(_06919_));
 sg13g2_nor2_1 _19567_ (.A(_10201_),
    .B(_10202_),
    .Y(_00342_));
 sg13g2_nor2_1 _19568_ (.A(_10129_),
    .B(_10127_),
    .Y(_10204_));
 sg13g2_nand2_1 _19569_ (.Y(_10205_),
    .A(_10130_),
    .B(_06919_));
 sg13g2_nor2_1 _19570_ (.A(_10204_),
    .B(_10205_),
    .Y(_00343_));
 sg13g2_inv_1 _19571_ (.Y(_10206_),
    .A(_10132_));
 sg13g2_nand2_1 _19572_ (.Y(_10207_),
    .A(_10133_),
    .B(_10135_));
 sg13g2_o21ai_1 _19573_ (.B1(_04191_),
    .Y(_10208_),
    .A1(_10207_),
    .A2(_10206_));
 sg13g2_a21oi_1 _19574_ (.A1(_10206_),
    .A2(_10207_),
    .Y(_00344_),
    .B1(_10208_));
 sg13g2_a21oi_1 _19575_ (.A1(_10140_),
    .A2(_10137_),
    .Y(_10209_),
    .B1(_10136_));
 sg13g2_nor2b_1 _19576_ (.A(_10138_),
    .B_N(_10140_),
    .Y(_10210_));
 sg13g2_nor3_1 _19577_ (.A(net110),
    .B(_10209_),
    .C(_10210_),
    .Y(_00345_));
 sg13g2_and3_1 _19578_ (.X(_10211_),
    .A(_10138_),
    .B(_10140_),
    .C(_10142_));
 sg13g2_o21ai_1 _19579_ (.B1(_06918_),
    .Y(_00346_),
    .A1(_10143_),
    .A2(_10211_));
 sg13g2_a21oi_1 _19580_ (.A1(_01870_),
    .A2(net84),
    .Y(_00226_),
    .B1(net86));
 sg13g2_inv_1 _19581_ (.Y(_00227_),
    .A(_01863_));
 sg13g2_a21oi_1 _19582_ (.A1(_01263_),
    .A2(_00781_),
    .Y(_00229_),
    .B1(net86));
 sg13g2_nor2_2 _19583_ (.A(_00033_),
    .B(net182),
    .Y(_10212_));
 sg13g2_xor2_1 _19584_ (.B(\vgadonut.frame[7] ),
    .A(_06004_),
    .X(_10213_));
 sg13g2_nor2_1 _19585_ (.A(_06000_),
    .B(\vgadonut.frame[4] ),
    .Y(_10214_));
 sg13g2_a22oi_1 _19586_ (.Y(_10215_),
    .B1(_06214_),
    .B2(_09992_),
    .A2(_09993_),
    .A1(_06003_));
 sg13g2_nand2_1 _19587_ (.Y(_10216_),
    .A(_09894_),
    .B(\vgadonut.frame[3] ));
 sg13g2_o21ai_1 _19588_ (.B1(_10216_),
    .Y(_10218_),
    .A1(_09863_),
    .A2(_09980_));
 sg13g2_nand2_1 _19589_ (.Y(_10219_),
    .A(_06001_),
    .B(_09983_));
 sg13g2_nand3_1 _19590_ (.B(_10218_),
    .C(_10219_),
    .A(_10215_),
    .Y(_10220_));
 sg13g2_nand2_1 _19591_ (.Y(_10221_),
    .A(_06002_),
    .B(_09989_));
 sg13g2_o21ai_1 _19592_ (.B1(_10221_),
    .Y(_10222_),
    .A1(_10003_),
    .A2(_09986_));
 sg13g2_a22oi_1 _19593_ (.Y(_10223_),
    .B1(_10222_),
    .B2(_10215_),
    .A2(_09991_),
    .A1(_06009_));
 sg13g2_o21ai_1 _19594_ (.B1(_10223_),
    .Y(_10224_),
    .A1(_10214_),
    .A2(_10220_));
 sg13g2_xnor2_1 _19595_ (.Y(_10225_),
    .A(_10213_),
    .B(_10224_));
 sg13g2_xor2_1 _19596_ (.B(_09991_),
    .A(net255),
    .X(_10226_));
 sg13g2_nand2_1 _19597_ (.Y(_10227_),
    .A(_09694_),
    .B(_09989_));
 sg13g2_o21ai_1 _19598_ (.B1(_10227_),
    .Y(_10229_),
    .A1(_05974_),
    .A2(_09986_));
 sg13g2_inv_1 _19599_ (.Y(_10230_),
    .A(_10229_));
 sg13g2_a22oi_1 _19600_ (.Y(_10231_),
    .B1(_09853_),
    .B2(_09980_),
    .A2(_09981_),
    .A1(_10073_));
 sg13g2_nand2_1 _19601_ (.Y(_10232_),
    .A(_09884_),
    .B(_09811_));
 sg13g2_o21ai_1 _19602_ (.B1(_10232_),
    .Y(_10233_),
    .A1(_10073_),
    .A2(_09981_));
 sg13g2_nand2_1 _19603_ (.Y(_10234_),
    .A(_10231_),
    .B(_10233_));
 sg13g2_nand2_1 _19604_ (.Y(_10235_),
    .A(_09716_),
    .B(\vgadonut.frame[3] ));
 sg13g2_nand2_1 _19605_ (.Y(_10236_),
    .A(net254),
    .B(\vgadonut.frame[2] ));
 sg13g2_nand3_1 _19606_ (.B(_10235_),
    .C(_10236_),
    .A(_10234_),
    .Y(_10237_));
 sg13g2_nand2_1 _19607_ (.Y(_10238_),
    .A(_05974_),
    .B(_09986_));
 sg13g2_nand2b_1 _19608_ (.Y(_10240_),
    .B(_09983_),
    .A_N(_09716_));
 sg13g2_nand3_1 _19609_ (.B(_10238_),
    .C(_10240_),
    .A(_10237_),
    .Y(_10241_));
 sg13g2_a22oi_1 _19610_ (.Y(_10242_),
    .B1(_10230_),
    .B2(_10241_),
    .A2(_09993_),
    .A1(_09705_));
 sg13g2_xnor2_1 _19611_ (.Y(_10243_),
    .A(_10226_),
    .B(_10242_));
 sg13g2_xnor2_1 _19612_ (.Y(_10244_),
    .A(_10225_),
    .B(_10243_));
 sg13g2_nand2_1 _19613_ (.Y(_10245_),
    .A(_10244_),
    .B(_06915_));
 sg13g2_buf_1 _19614_ (.A(_10245_),
    .X(_10246_));
 sg13g2_o21ai_1 _19615_ (.B1(_10246_),
    .Y(_10247_),
    .A1(_06915_),
    .A2(_00032_));
 sg13g2_buf_1 _19616_ (.A(_10247_),
    .X(_10248_));
 sg13g2_inv_1 _19617_ (.Y(_10249_),
    .A(_10248_));
 sg13g2_xor2_1 _19618_ (.B(_09811_),
    .A(_09884_),
    .X(_10251_));
 sg13g2_buf_2 _19619_ (.A(_10251_),
    .X(_10252_));
 sg13g2_xnor2_1 _19620_ (.Y(_10253_),
    .A(_00096_),
    .B(_10252_));
 sg13g2_buf_2 _19621_ (.A(_10253_),
    .X(_10254_));
 sg13g2_nand2_1 _19622_ (.Y(_10255_),
    .A(_10249_),
    .B(_10254_));
 sg13g2_inv_1 _19623_ (.Y(_10256_),
    .A(_10254_));
 sg13g2_nand2_1 _19624_ (.Y(_10257_),
    .A(_10248_),
    .B(_10256_));
 sg13g2_inv_1 _19625_ (.Y(_10258_),
    .A(_10212_));
 sg13g2_nand2_1 _19626_ (.Y(_10259_),
    .A(_10257_),
    .B(_10258_));
 sg13g2_inv_1 _19627_ (.Y(_10260_),
    .A(_10259_));
 sg13g2_a21oi_1 _19628_ (.A1(_10212_),
    .A2(_10255_),
    .Y(_10262_),
    .B1(_10260_));
 sg13g2_o21ai_1 _19629_ (.B1(_10246_),
    .Y(_10263_),
    .A1(net182),
    .A2(_00030_));
 sg13g2_buf_1 _19630_ (.A(_10263_),
    .X(_10264_));
 sg13g2_xnor2_1 _19631_ (.Y(_10265_),
    .A(net254),
    .B(_09811_));
 sg13g2_inv_1 _19632_ (.Y(_10266_),
    .A(_10265_));
 sg13g2_nor2_1 _19633_ (.A(_00029_),
    .B(net182),
    .Y(_10267_));
 sg13g2_inv_1 _19634_ (.Y(_10268_),
    .A(_10267_));
 sg13g2_a21oi_1 _19635_ (.A1(_10266_),
    .A2(_10258_),
    .Y(_10269_),
    .B1(_10268_));
 sg13g2_a21oi_1 _19636_ (.A1(_10212_),
    .A2(_10265_),
    .Y(_10270_),
    .B1(_10269_));
 sg13g2_inv_1 _19637_ (.Y(_10271_),
    .A(_10270_));
 sg13g2_o21ai_1 _19638_ (.B1(_10246_),
    .Y(_10272_),
    .A1(net182),
    .A2(_00028_));
 sg13g2_xnor2_1 _19639_ (.Y(_10273_),
    .A(_09925_),
    .B(_10272_));
 sg13g2_nor2_1 _19640_ (.A(_10267_),
    .B(_10273_),
    .Y(_10274_));
 sg13g2_a21oi_1 _19641_ (.A1(_10264_),
    .A2(_10271_),
    .Y(_10275_),
    .B1(_10274_));
 sg13g2_nand2_1 _19642_ (.Y(_10276_),
    .A(_10273_),
    .B(_10267_));
 sg13g2_nand2_1 _19643_ (.Y(_10277_),
    .A(_10275_),
    .B(_10276_));
 sg13g2_o21ai_1 _19644_ (.B1(_10277_),
    .Y(_10278_),
    .A1(_10264_),
    .A2(_10271_));
 sg13g2_nor2_1 _19645_ (.A(_09925_),
    .B(_10272_),
    .Y(_10279_));
 sg13g2_nor2_1 _19646_ (.A(_10279_),
    .B(_10274_),
    .Y(_10280_));
 sg13g2_nand2b_1 _19647_ (.Y(_10281_),
    .B(net216),
    .A_N(_00031_));
 sg13g2_buf_1 _19648_ (.A(_10281_),
    .X(_10283_));
 sg13g2_nor2_1 _19649_ (.A(_09946_),
    .B(_10264_),
    .Y(_10284_));
 sg13g2_nand2_1 _19650_ (.Y(_10285_),
    .A(_10264_),
    .B(_09946_));
 sg13g2_nor2b_1 _19651_ (.A(_10284_),
    .B_N(_10285_),
    .Y(_10286_));
 sg13g2_xnor2_1 _19652_ (.Y(_10287_),
    .A(_10283_),
    .B(_10286_));
 sg13g2_nor2_1 _19653_ (.A(_10280_),
    .B(_10287_),
    .Y(_10288_));
 sg13g2_nand2_1 _19654_ (.Y(_10289_),
    .A(_10255_),
    .B(_10257_));
 sg13g2_xnor2_1 _19655_ (.Y(_10290_),
    .A(_10212_),
    .B(_10289_));
 sg13g2_xor2_1 _19656_ (.B(_10252_),
    .A(_10283_),
    .X(_10291_));
 sg13g2_inv_1 _19657_ (.Y(_10292_),
    .A(_10252_));
 sg13g2_nor2b_1 _19658_ (.A(_10292_),
    .B_N(_10283_),
    .Y(_10294_));
 sg13g2_a21o_1 _19659_ (.A2(_10291_),
    .A1(_10249_),
    .B1(_10294_),
    .X(_10295_));
 sg13g2_nand2b_1 _19660_ (.Y(_10296_),
    .B(_10295_),
    .A_N(_10290_));
 sg13g2_nand2b_1 _19661_ (.Y(_10297_),
    .B(_10290_),
    .A_N(_10295_));
 sg13g2_xnor2_1 _19662_ (.Y(_10298_),
    .A(_10291_),
    .B(_10248_));
 sg13g2_a21oi_1 _19663_ (.A1(_10285_),
    .A2(_10283_),
    .Y(_10299_),
    .B1(_10284_));
 sg13g2_xnor2_1 _19664_ (.Y(_10300_),
    .A(_10298_),
    .B(_10299_));
 sg13g2_nand3_1 _19665_ (.B(_10297_),
    .C(_10300_),
    .A(_10296_),
    .Y(_10301_));
 sg13g2_a21oi_1 _19666_ (.A1(_10280_),
    .A2(_10287_),
    .Y(_10302_),
    .B1(_10301_));
 sg13g2_o21ai_1 _19667_ (.B1(_10302_),
    .Y(_10303_),
    .A1(_10278_),
    .A2(_10288_));
 sg13g2_inv_1 _19668_ (.Y(_10305_),
    .A(_10299_));
 sg13g2_nand4_1 _19669_ (.B(_10297_),
    .C(_10305_),
    .A(_10296_),
    .Y(_10306_),
    .D(_10298_));
 sg13g2_nand3_1 _19670_ (.B(_10296_),
    .C(_10306_),
    .A(_10303_),
    .Y(_10307_));
 sg13g2_nor2b_1 _19671_ (.A(_09748_),
    .B_N(_09637_),
    .Y(_10308_));
 sg13g2_nand3_1 _19672_ (.B(_09853_),
    .C(_09705_),
    .A(_06013_),
    .Y(_10309_));
 sg13g2_nand2_1 _19673_ (.Y(_10310_),
    .A(_10018_),
    .B(_06004_));
 sg13g2_nand3_1 _19674_ (.B(_10021_),
    .C(_06019_),
    .A(_10310_),
    .Y(_10311_));
 sg13g2_a21oi_2 _19675_ (.B1(_10311_),
    .Y(_10312_),
    .A2(_10309_),
    .A1(_10308_));
 sg13g2_o21ai_1 _19676_ (.B1(_10312_),
    .Y(_10313_),
    .A1(_10262_),
    .A2(_10307_));
 sg13g2_nand2_1 _19677_ (.Y(_10314_),
    .A(_10307_),
    .B(_10262_));
 sg13g2_nor2b_1 _19678_ (.A(_10313_),
    .B_N(_10314_),
    .Y(_00230_));
 sg13g2_inv_1 _19679_ (.Y(_10316_),
    .A(_10312_));
 sg13g2_a21oi_1 _19680_ (.A1(_10314_),
    .A2(_10259_),
    .Y(_00231_),
    .B1(_10316_));
 sg13g2_nand2_1 _19681_ (.Y(_10317_),
    .A(net216),
    .B(_00101_));
 sg13g2_nand2_1 _19682_ (.Y(_10318_),
    .A(_10246_),
    .B(_10317_));
 sg13g2_nand2_1 _19683_ (.Y(_10319_),
    .A(net216),
    .B(_00039_));
 sg13g2_nand2_1 _19684_ (.Y(_10320_),
    .A(_10246_),
    .B(_10319_));
 sg13g2_inv_1 _19685_ (.Y(_10321_),
    .A(_10320_));
 sg13g2_a21oi_1 _19686_ (.A1(_10318_),
    .A2(_10256_),
    .Y(_10322_),
    .B1(_10321_));
 sg13g2_inv_1 _19687_ (.Y(_10323_),
    .A(_10322_));
 sg13g2_o21ai_1 _19688_ (.B1(_10321_),
    .Y(_10325_),
    .A1(_10256_),
    .A2(_10318_));
 sg13g2_nand2_1 _19689_ (.Y(_10326_),
    .A(_10323_),
    .B(_10325_));
 sg13g2_buf_1 _19690_ (.A(_00102_),
    .X(_10327_));
 sg13g2_nor2_1 _19691_ (.A(_00103_),
    .B(_06915_),
    .Y(_10328_));
 sg13g2_nand2b_1 _19692_ (.Y(_10329_),
    .B(_10328_),
    .A_N(_10327_));
 sg13g2_nand3_1 _19693_ (.B(_10327_),
    .C(_00103_),
    .A(net216),
    .Y(_10330_));
 sg13g2_nand2_1 _19694_ (.Y(_10331_),
    .A(_10329_),
    .B(_10330_));
 sg13g2_xor2_1 _19695_ (.B(_09935_),
    .A(_10331_),
    .X(_10332_));
 sg13g2_nor2_1 _19696_ (.A(_00104_),
    .B(net182),
    .Y(_10333_));
 sg13g2_nor2_1 _19697_ (.A(_00034_),
    .B(net182),
    .Y(_10334_));
 sg13g2_a22oi_1 _19698_ (.Y(_10335_),
    .B1(_00104_),
    .B2(_10334_),
    .A2(_00034_),
    .A1(_10333_));
 sg13g2_inv_1 _19699_ (.Y(_10336_),
    .A(_10335_));
 sg13g2_nand2b_1 _19700_ (.Y(_10337_),
    .B(_06915_),
    .A_N(_10244_));
 sg13g2_nor2b_1 _19701_ (.A(_10328_),
    .B_N(_10337_),
    .Y(_10338_));
 sg13g2_nand2_1 _19702_ (.Y(_10339_),
    .A(_10333_),
    .B(_00034_));
 sg13g2_o21ai_1 _19703_ (.B1(_10339_),
    .Y(_10340_),
    .A1(_10336_),
    .A2(_10338_));
 sg13g2_nor2b_1 _19704_ (.A(_10332_),
    .B_N(_10340_),
    .Y(_10341_));
 sg13g2_nor2_1 _19705_ (.A(_10266_),
    .B(_10320_),
    .Y(_10342_));
 sg13g2_a21oi_1 _19706_ (.A1(_10244_),
    .A2(net182),
    .Y(_10343_),
    .B1(_10333_));
 sg13g2_o21ai_1 _19707_ (.B1(_10343_),
    .Y(_10344_),
    .A1(_10265_),
    .A2(_10321_));
 sg13g2_nand2b_1 _19708_ (.Y(_10346_),
    .B(_10344_),
    .A_N(_10342_));
 sg13g2_inv_1 _19709_ (.Y(_10347_),
    .A(_09925_));
 sg13g2_inv_1 _19710_ (.Y(_10348_),
    .A(_10346_));
 sg13g2_xnor2_1 _19711_ (.Y(_10349_),
    .A(_10335_),
    .B(_10338_));
 sg13g2_o21ai_1 _19712_ (.B1(_10349_),
    .Y(_10350_),
    .A1(_10347_),
    .A2(_10348_));
 sg13g2_o21ai_1 _19713_ (.B1(_10350_),
    .Y(_10351_),
    .A1(_09925_),
    .A2(_10346_));
 sg13g2_nor2b_1 _19714_ (.A(_10340_),
    .B_N(_10332_),
    .Y(_10352_));
 sg13g2_nor3_1 _19715_ (.A(_00101_),
    .B(_10327_),
    .C(net182),
    .Y(_10353_));
 sg13g2_nand3_1 _19716_ (.B(_00101_),
    .C(_10327_),
    .A(net216),
    .Y(_10354_));
 sg13g2_nand2b_1 _19717_ (.Y(_10355_),
    .B(_10354_),
    .A_N(_10353_));
 sg13g2_xnor2_1 _19718_ (.Y(_10357_),
    .A(_10252_),
    .B(_10355_));
 sg13g2_o21ai_1 _19719_ (.B1(_10329_),
    .Y(_10358_),
    .A1(_10331_),
    .A2(_09946_));
 sg13g2_nor2_1 _19720_ (.A(_10357_),
    .B(_10358_),
    .Y(_10359_));
 sg13g2_xnor2_1 _19721_ (.Y(_10360_),
    .A(_10318_),
    .B(_10320_));
 sg13g2_xnor2_1 _19722_ (.Y(_10361_),
    .A(_10254_),
    .B(_10360_));
 sg13g2_a21oi_1 _19723_ (.A1(_10252_),
    .A2(_10354_),
    .Y(_10362_),
    .B1(_10353_));
 sg13g2_nand2_1 _19724_ (.Y(_10363_),
    .A(_10361_),
    .B(_10362_));
 sg13g2_inv_1 _19725_ (.Y(_10364_),
    .A(_10363_));
 sg13g2_nor2_1 _19726_ (.A(_10359_),
    .B(_10364_),
    .Y(_10365_));
 sg13g2_or2_1 _19727_ (.X(_10366_),
    .B(_10361_),
    .A(_10362_));
 sg13g2_nand2_1 _19728_ (.Y(_10368_),
    .A(_10358_),
    .B(_10357_));
 sg13g2_nand3_1 _19729_ (.B(_10366_),
    .C(_10368_),
    .A(_10365_),
    .Y(_10369_));
 sg13g2_nor2_1 _19730_ (.A(_10352_),
    .B(_10369_),
    .Y(_10370_));
 sg13g2_o21ai_1 _19731_ (.B1(_10370_),
    .Y(_10371_),
    .A1(_10341_),
    .A2(_10351_));
 sg13g2_a21o_1 _19732_ (.A2(_10368_),
    .A1(_10366_),
    .B1(_10364_),
    .X(_10372_));
 sg13g2_nand2_1 _19733_ (.Y(_10373_),
    .A(_10371_),
    .B(_10372_));
 sg13g2_xor2_1 _19734_ (.B(_10373_),
    .A(_10326_),
    .X(_10374_));
 sg13g2_nor2_1 _19735_ (.A(_10316_),
    .B(_10374_),
    .Y(_00529_));
 sg13g2_nand3b_1 _19736_ (.B(_10370_),
    .C(_10351_),
    .Y(_10375_),
    .A_N(_10341_));
 sg13g2_nand2_1 _19737_ (.Y(_10376_),
    .A(_10372_),
    .B(_10323_));
 sg13g2_a21oi_1 _19738_ (.A1(_10341_),
    .A2(_10365_),
    .Y(_10378_),
    .B1(_10376_));
 sg13g2_nand2_1 _19739_ (.Y(_10379_),
    .A(_10325_),
    .B(_10312_));
 sg13g2_a21oi_1 _19740_ (.A1(_10375_),
    .A2(_10378_),
    .Y(_00530_),
    .B1(_10379_));
 sg13g2_nand2_2 _19741_ (.Y(_10380_),
    .A(net216),
    .B(_00044_));
 sg13g2_inv_1 _19742_ (.Y(_10381_),
    .A(_10380_));
 sg13g2_o21ai_1 _19743_ (.B1(_10246_),
    .Y(_10382_),
    .A1(_06915_),
    .A2(_00098_));
 sg13g2_buf_1 _19744_ (.A(_10382_),
    .X(_10383_));
 sg13g2_a21oi_1 _19745_ (.A1(_10254_),
    .A2(_10381_),
    .Y(_10384_),
    .B1(_10383_));
 sg13g2_o21ai_1 _19746_ (.B1(_10383_),
    .Y(_10385_),
    .A1(_10254_),
    .A2(_10381_));
 sg13g2_inv_1 _19747_ (.Y(_10386_),
    .A(_10385_));
 sg13g2_nor2_1 _19748_ (.A(_10384_),
    .B(_10386_),
    .Y(_10387_));
 sg13g2_inv_1 _19749_ (.Y(_10388_),
    .A(_00099_));
 sg13g2_o21ai_1 _19750_ (.B1(_10337_),
    .Y(_10389_),
    .A1(_06915_),
    .A2(_10388_));
 sg13g2_nand2_1 _19751_ (.Y(_10390_),
    .A(_10389_),
    .B(_10380_));
 sg13g2_a22oi_1 _19752_ (.Y(_10391_),
    .B1(_10252_),
    .B2(_10390_),
    .A2(_10381_),
    .A1(_10388_));
 sg13g2_xnor2_1 _19753_ (.Y(_10392_),
    .A(_10380_),
    .B(_10383_));
 sg13g2_xnor2_1 _19754_ (.Y(_10393_),
    .A(_10254_),
    .B(_10392_));
 sg13g2_nor2_1 _19755_ (.A(_10391_),
    .B(_10393_),
    .Y(_10394_));
 sg13g2_nand2_2 _19756_ (.Y(_10395_),
    .A(net216),
    .B(_00042_));
 sg13g2_nand2_1 _19757_ (.Y(_10396_),
    .A(_10389_),
    .B(_10395_));
 sg13g2_nor2_1 _19758_ (.A(_10395_),
    .B(_10389_),
    .Y(_10398_));
 sg13g2_a21oi_1 _19759_ (.A1(_10396_),
    .A2(_09935_),
    .Y(_10399_),
    .B1(_10398_));
 sg13g2_o21ai_1 _19760_ (.B1(_10390_),
    .Y(_10400_),
    .A1(_00099_),
    .A2(_10380_));
 sg13g2_xnor2_1 _19761_ (.Y(_10401_),
    .A(_10292_),
    .B(_10400_));
 sg13g2_nor2_1 _19762_ (.A(_10399_),
    .B(_10401_),
    .Y(_10402_));
 sg13g2_nor2b_1 _19763_ (.A(_10398_),
    .B_N(_10396_),
    .Y(_10403_));
 sg13g2_xnor2_1 _19764_ (.Y(_10404_),
    .A(_09935_),
    .B(_10403_));
 sg13g2_inv_1 _19765_ (.Y(_10405_),
    .A(_00100_));
 sg13g2_nand2_1 _19766_ (.Y(_10406_),
    .A(net216),
    .B(_00040_));
 sg13g2_inv_1 _19767_ (.Y(_10407_),
    .A(_10406_));
 sg13g2_inv_1 _19768_ (.Y(_10409_),
    .A(_10395_));
 sg13g2_o21ai_1 _19769_ (.B1(_10337_),
    .Y(_10410_),
    .A1(_06916_),
    .A2(_10405_));
 sg13g2_nand2_1 _19770_ (.Y(_10411_),
    .A(_10410_),
    .B(_10406_));
 sg13g2_a22oi_1 _19771_ (.Y(_10412_),
    .B1(_10409_),
    .B2(_10411_),
    .A2(_10407_),
    .A1(_10405_));
 sg13g2_nand2_1 _19772_ (.Y(_10413_),
    .A(_10404_),
    .B(_10412_));
 sg13g2_nand2_1 _19773_ (.Y(_10414_),
    .A(_10401_),
    .B(_10399_));
 sg13g2_nand2_1 _19774_ (.Y(_10415_),
    .A(_10393_),
    .B(_10391_));
 sg13g2_nand3_1 _19775_ (.B(_10414_),
    .C(_10415_),
    .A(_10413_),
    .Y(_10416_));
 sg13g2_nor3_1 _19776_ (.A(_10394_),
    .B(_10402_),
    .C(_10416_),
    .Y(_10417_));
 sg13g2_nor2_1 _19777_ (.A(_10412_),
    .B(_10404_),
    .Y(_10418_));
 sg13g2_nand2_1 _19778_ (.Y(_10420_),
    .A(_10417_),
    .B(_10418_));
 sg13g2_o21ai_1 _19779_ (.B1(_10411_),
    .Y(_10421_),
    .A1(_00100_),
    .A2(_10406_));
 sg13g2_xnor2_1 _19780_ (.Y(_10422_),
    .A(_10395_),
    .B(_10421_));
 sg13g2_inv_1 _19781_ (.Y(_10423_),
    .A(_10410_));
 sg13g2_nor2_1 _19782_ (.A(_10383_),
    .B(_10423_),
    .Y(_10424_));
 sg13g2_nand2_1 _19783_ (.Y(_10425_),
    .A(_10423_),
    .B(_10383_));
 sg13g2_o21ai_1 _19784_ (.B1(_10425_),
    .Y(_10426_),
    .A1(_10265_),
    .A2(_10424_));
 sg13g2_nand2_1 _19785_ (.Y(_10427_),
    .A(_10426_),
    .B(_10347_));
 sg13g2_nor2_1 _19786_ (.A(_10347_),
    .B(_10426_),
    .Y(_10428_));
 sg13g2_a21oi_1 _19787_ (.A1(_10422_),
    .A2(_10427_),
    .Y(_10429_),
    .B1(_10428_));
 sg13g2_nand2_1 _19788_ (.Y(_00544_),
    .A(_10417_),
    .B(_10429_));
 sg13g2_o21ai_1 _19789_ (.B1(_10415_),
    .Y(_00545_),
    .A1(_10394_),
    .A2(_10402_));
 sg13g2_nand3_1 _19790_ (.B(_00544_),
    .C(_00545_),
    .A(_10420_),
    .Y(_00546_));
 sg13g2_o21ai_1 _19791_ (.B1(_10312_),
    .Y(_00547_),
    .A1(_10387_),
    .A2(_00546_));
 sg13g2_a21oi_1 _19792_ (.A1(_10387_),
    .A2(_00546_),
    .Y(_00531_),
    .B1(_00547_));
 sg13g2_nand2_1 _19793_ (.Y(_00548_),
    .A(_10414_),
    .B(_10415_));
 sg13g2_nor2_1 _19794_ (.A(_10402_),
    .B(_10418_),
    .Y(_00549_));
 sg13g2_nor2_1 _19795_ (.A(_00548_),
    .B(_00549_),
    .Y(_00550_));
 sg13g2_nor2_1 _19796_ (.A(_10418_),
    .B(_00544_),
    .Y(_00551_));
 sg13g2_nor4_1 _19797_ (.A(_10386_),
    .B(_10394_),
    .C(_00550_),
    .D(_00551_),
    .Y(_00552_));
 sg13g2_nor3_1 _19798_ (.A(_10316_),
    .B(_10384_),
    .C(_00552_),
    .Y(_00532_));
 sg13g2_xnor2_1 _19799_ (.Y(_00553_),
    .A(net232),
    .B(_06274_));
 sg13g2_nor3_1 _19800_ (.A(net233),
    .B(net223),
    .C(_00553_),
    .Y(_00554_));
 sg13g2_inv_1 _19801_ (.Y(_00555_),
    .A(_00554_));
 sg13g2_o21ai_1 _19802_ (.B1(_00553_),
    .Y(_00556_),
    .A1(net233),
    .A2(net223));
 sg13g2_nand2_1 _19803_ (.Y(_00557_),
    .A(_00555_),
    .B(_00556_));
 sg13g2_inv_1 _19804_ (.Y(_00558_),
    .A(_00557_));
 sg13g2_xor2_1 _19805_ (.B(_08856_),
    .A(_05380_),
    .X(_00559_));
 sg13g2_a21oi_1 _19806_ (.A1(_05405_),
    .A2(_08852_),
    .Y(_00560_),
    .B1(_00559_));
 sg13g2_xor2_1 _19807_ (.B(_08851_),
    .A(_05390_),
    .X(_00561_));
 sg13g2_inv_1 _19808_ (.Y(_00563_),
    .A(_00561_));
 sg13g2_nand3_1 _19809_ (.B(_05396_),
    .C(_08843_),
    .A(_00563_),
    .Y(_00564_));
 sg13g2_xor2_1 _19810_ (.B(_08843_),
    .A(_05396_),
    .X(_00565_));
 sg13g2_nor3_1 _19811_ (.A(_05403_),
    .B(\vgadonut.donut.sA[0] ),
    .C(_00565_),
    .Y(_00566_));
 sg13g2_a21oi_1 _19812_ (.A1(_05396_),
    .A2(_08843_),
    .Y(_00567_),
    .B1(_00563_));
 sg13g2_a21oi_1 _19813_ (.A1(_00564_),
    .A2(_00566_),
    .Y(_00568_),
    .B1(_00567_));
 sg13g2_nand3_1 _19814_ (.B(_05405_),
    .C(_08852_),
    .A(_00559_),
    .Y(_00569_));
 sg13g2_o21ai_1 _19815_ (.B1(_00569_),
    .Y(_00570_),
    .A1(_00560_),
    .A2(_00568_));
 sg13g2_buf_1 _19816_ (.A(_00570_),
    .X(_00571_));
 sg13g2_xor2_1 _19817_ (.B(net215),
    .A(net236),
    .X(_00572_));
 sg13g2_a21oi_1 _19818_ (.A1(_05401_),
    .A2(_09674_),
    .Y(_00574_),
    .B1(_00572_));
 sg13g2_inv_1 _19819_ (.Y(_00575_),
    .A(_00574_));
 sg13g2_and3_1 _19820_ (.X(_00576_),
    .A(_00572_),
    .B(_05401_),
    .C(_09674_));
 sg13g2_buf_1 _19821_ (.A(_00576_),
    .X(_00577_));
 sg13g2_a21o_1 _19822_ (.A2(_00575_),
    .A1(_00571_),
    .B1(_00577_),
    .X(_00578_));
 sg13g2_nor2_1 _19823_ (.A(net237),
    .B(_06027_),
    .Y(_00579_));
 sg13g2_inv_1 _19824_ (.Y(_00580_),
    .A(_00579_));
 sg13g2_xor2_1 _19825_ (.B(_06261_),
    .A(net235),
    .X(_00581_));
 sg13g2_xnor2_1 _19826_ (.Y(_00582_),
    .A(_00580_),
    .B(_00581_));
 sg13g2_xor2_1 _19827_ (.B(_06026_),
    .A(_05381_),
    .X(_00583_));
 sg13g2_inv_1 _19828_ (.Y(_00585_),
    .A(_00583_));
 sg13g2_nor3_1 _19829_ (.A(_05384_),
    .B(net215),
    .C(_00585_),
    .Y(_00586_));
 sg13g2_o21ai_1 _19830_ (.B1(_00585_),
    .Y(_00587_),
    .A1(_05384_),
    .A2(net215));
 sg13g2_nor2b_1 _19831_ (.A(_00586_),
    .B_N(_00587_),
    .Y(_00588_));
 sg13g2_nand3_1 _19832_ (.B(_00582_),
    .C(_00588_),
    .A(_00578_),
    .Y(_00589_));
 sg13g2_nor2b_1 _19833_ (.A(_00580_),
    .B_N(_00581_),
    .Y(_00590_));
 sg13g2_a21oi_1 _19834_ (.A1(_00586_),
    .A2(_00581_),
    .Y(_00591_),
    .B1(_00590_));
 sg13g2_nand2_1 _19835_ (.Y(_00592_),
    .A(_00589_),
    .B(_00591_));
 sg13g2_xor2_1 _19836_ (.B(_06257_),
    .A(net234),
    .X(_00593_));
 sg13g2_a21oi_1 _19837_ (.A1(_06482_),
    .A2(_06263_),
    .Y(_00594_),
    .B1(_00593_));
 sg13g2_inv_1 _19838_ (.Y(_00596_),
    .A(_00593_));
 sg13g2_nor3_2 _19839_ (.A(net235),
    .B(net194),
    .C(_00596_),
    .Y(_00597_));
 sg13g2_nor2_2 _19840_ (.A(_00594_),
    .B(_00597_),
    .Y(_00598_));
 sg13g2_nand2_1 _19841_ (.Y(_00599_),
    .A(_00592_),
    .B(_00598_));
 sg13g2_inv_1 _19842_ (.Y(_00600_),
    .A(_00599_));
 sg13g2_xor2_1 _19843_ (.B(net223),
    .A(net233),
    .X(_00601_));
 sg13g2_a21oi_1 _19844_ (.A1(_06460_),
    .A2(_06259_),
    .Y(_00602_),
    .B1(_00601_));
 sg13g2_nand3_1 _19845_ (.B(_06460_),
    .C(_06259_),
    .A(_00601_),
    .Y(_00603_));
 sg13g2_inv_1 _19846_ (.Y(_00604_),
    .A(_00603_));
 sg13g2_nor2_1 _19847_ (.A(_00602_),
    .B(_00604_),
    .Y(_00605_));
 sg13g2_inv_1 _19848_ (.Y(_00607_),
    .A(_00597_));
 sg13g2_a21oi_1 _19849_ (.A1(_00607_),
    .A2(_00603_),
    .Y(_00608_),
    .B1(_00602_));
 sg13g2_a21oi_1 _19850_ (.A1(_00600_),
    .A2(_00605_),
    .Y(_00609_),
    .B1(_00608_));
 sg13g2_xnor2_1 _19851_ (.Y(_00610_),
    .A(_00558_),
    .B(_00609_));
 sg13g2_nor2_1 _19852_ (.A(net220),
    .B(_06485_),
    .Y(_00611_));
 sg13g2_nor2_1 _19853_ (.A(net239),
    .B(_09478_),
    .Y(_00612_));
 sg13g2_nor2_2 _19854_ (.A(_00611_),
    .B(_00612_),
    .Y(_00613_));
 sg13g2_nor2b_1 _19855_ (.A(_04826_),
    .B_N(\vgadonut.donut.cA[0] ),
    .Y(_00614_));
 sg13g2_inv_1 _19856_ (.Y(_00615_),
    .A(\vgadonut.donut.cA[1] ));
 sg13g2_nand2_1 _19857_ (.Y(_00616_),
    .A(_00615_),
    .B(_04824_));
 sg13g2_nor2_1 _19858_ (.A(_04824_),
    .B(_00615_),
    .Y(_00618_));
 sg13g2_a21oi_1 _19859_ (.A1(_00614_),
    .A2(_00616_),
    .Y(_00619_),
    .B1(_00618_));
 sg13g2_xnor2_1 _19860_ (.Y(_00620_),
    .A(_04823_),
    .B(_06260_));
 sg13g2_nand2_1 _19861_ (.Y(_00621_),
    .A(_00619_),
    .B(_00620_));
 sg13g2_o21ai_1 _19862_ (.B1(_00621_),
    .Y(_00622_),
    .A1(_09054_),
    .A2(_06260_));
 sg13g2_xnor2_1 _19863_ (.Y(_00623_),
    .A(_04820_),
    .B(_06252_));
 sg13g2_nand2_1 _19864_ (.Y(_00624_),
    .A(_00622_),
    .B(_00623_));
 sg13g2_o21ai_1 _19865_ (.B1(_00624_),
    .Y(_00625_),
    .A1(_09061_),
    .A2(_06252_));
 sg13g2_nand2_1 _19866_ (.Y(_00626_),
    .A(_09046_),
    .B(_06276_));
 sg13g2_nand2_1 _19867_ (.Y(_00627_),
    .A(_00625_),
    .B(_00626_));
 sg13g2_nor2_1 _19868_ (.A(_06276_),
    .B(_09046_),
    .Y(_00628_));
 sg13g2_inv_1 _19869_ (.Y(_00629_),
    .A(_00628_));
 sg13g2_nand2_1 _19870_ (.Y(_00630_),
    .A(_00627_),
    .B(_00629_));
 sg13g2_nor2_1 _19871_ (.A(net243),
    .B(_06285_),
    .Y(_00631_));
 sg13g2_inv_1 _19872_ (.Y(_00632_),
    .A(_00631_));
 sg13g2_nor2_1 _19873_ (.A(_06284_),
    .B(_09050_),
    .Y(_00633_));
 sg13g2_a21o_1 _19874_ (.A2(_00632_),
    .A1(_00630_),
    .B1(_00633_),
    .X(_00634_));
 sg13g2_nor2_1 _19875_ (.A(net244),
    .B(_06293_),
    .Y(_00635_));
 sg13g2_inv_1 _19876_ (.Y(_00636_),
    .A(_00635_));
 sg13g2_nor2_1 _19877_ (.A(_06292_),
    .B(_09034_),
    .Y(_00637_));
 sg13g2_a21oi_1 _19878_ (.A1(_00634_),
    .A2(_00636_),
    .Y(_00639_),
    .B1(_00637_));
 sg13g2_nor2_1 _19879_ (.A(net225),
    .B(_09028_),
    .Y(_00640_));
 sg13g2_nor2_1 _19880_ (.A(net242),
    .B(_06314_),
    .Y(_00641_));
 sg13g2_nor2_1 _19881_ (.A(_00640_),
    .B(_00641_),
    .Y(_00642_));
 sg13g2_nand2b_1 _19882_ (.Y(_00643_),
    .B(_00642_),
    .A_N(_00639_));
 sg13g2_nor2_1 _19883_ (.A(_06245_),
    .B(_09020_),
    .Y(_00644_));
 sg13g2_nor2_1 _19884_ (.A(_00640_),
    .B(_00644_),
    .Y(_00645_));
 sg13g2_nor2_1 _19885_ (.A(net241),
    .B(_06301_),
    .Y(_00646_));
 sg13g2_a21oi_1 _19886_ (.A1(_00643_),
    .A2(_00645_),
    .Y(_00647_),
    .B1(_00646_));
 sg13g2_nor2_1 _19887_ (.A(net240),
    .B(_06311_),
    .Y(_00648_));
 sg13g2_nor2_1 _19888_ (.A(net227),
    .B(_06478_),
    .Y(_00650_));
 sg13g2_nor2_1 _19889_ (.A(_00648_),
    .B(_00650_),
    .Y(_00651_));
 sg13g2_inv_1 _19890_ (.Y(_00652_),
    .A(_00651_));
 sg13g2_nor2_1 _19891_ (.A(_06235_),
    .B(_09004_),
    .Y(_00653_));
 sg13g2_nor2_1 _19892_ (.A(net207),
    .B(_06240_),
    .Y(_00654_));
 sg13g2_nor2_1 _19893_ (.A(_00653_),
    .B(_00654_),
    .Y(_00655_));
 sg13g2_inv_1 _19894_ (.Y(_00656_),
    .A(_00655_));
 sg13g2_nor2_1 _19895_ (.A(_00652_),
    .B(_00656_),
    .Y(_00657_));
 sg13g2_nor2_1 _19896_ (.A(_00650_),
    .B(_00653_),
    .Y(_00658_));
 sg13g2_nor2_1 _19897_ (.A(_00648_),
    .B(_00658_),
    .Y(_00659_));
 sg13g2_a21oi_1 _19898_ (.A1(_00647_),
    .A2(_00657_),
    .Y(_00661_),
    .B1(_00659_));
 sg13g2_xnor2_1 _19899_ (.Y(_00662_),
    .A(_00613_),
    .B(_00661_));
 sg13g2_xnor2_1 _19900_ (.Y(_00663_),
    .A(_06067_),
    .B(_00662_));
 sg13g2_inv_1 _19901_ (.Y(_00664_),
    .A(_00640_));
 sg13g2_o21ai_1 _19902_ (.B1(_00664_),
    .Y(_00665_),
    .A1(_00641_),
    .A2(_00639_));
 sg13g2_nor2_1 _19903_ (.A(_00646_),
    .B(_00644_),
    .Y(_00666_));
 sg13g2_nand2_1 _19904_ (.Y(_00667_),
    .A(_00665_),
    .B(_00666_));
 sg13g2_nor2_1 _19905_ (.A(_00653_),
    .B(_00644_),
    .Y(_00668_));
 sg13g2_a21oi_1 _19906_ (.A1(_00667_),
    .A2(_00668_),
    .Y(_00669_),
    .B1(_00654_));
 sg13g2_xnor2_1 _19907_ (.Y(_00670_),
    .A(_00652_),
    .B(_00669_));
 sg13g2_inv_1 _19908_ (.Y(_00672_),
    .A(_00670_));
 sg13g2_xnor2_1 _19909_ (.Y(_00673_),
    .A(_00656_),
    .B(_00647_));
 sg13g2_inv_1 _19910_ (.Y(_00674_),
    .A(_00673_));
 sg13g2_xnor2_1 _19911_ (.Y(_00675_),
    .A(_00666_),
    .B(_00665_));
 sg13g2_nor2_1 _19912_ (.A(_00637_),
    .B(_00635_),
    .Y(_00676_));
 sg13g2_xnor2_1 _19913_ (.Y(_00677_),
    .A(_00676_),
    .B(_00634_));
 sg13g2_nor2_1 _19914_ (.A(_00633_),
    .B(_00631_),
    .Y(_00678_));
 sg13g2_nand3b_1 _19915_ (.B(_00627_),
    .C(_00629_),
    .Y(_00679_),
    .A_N(_00678_));
 sg13g2_nand2_1 _19916_ (.Y(_00680_),
    .A(_00630_),
    .B(_00678_));
 sg13g2_nand2_1 _19917_ (.Y(_00681_),
    .A(_00679_),
    .B(_00680_));
 sg13g2_nand2_1 _19918_ (.Y(_00683_),
    .A(_00629_),
    .B(_00626_));
 sg13g2_xor2_1 _19919_ (.B(_00625_),
    .A(_00683_),
    .X(_00684_));
 sg13g2_xnor2_1 _19920_ (.Y(_00685_),
    .A(net252),
    .B(_00684_));
 sg13g2_xnor2_1 _19921_ (.Y(_00686_),
    .A(_00623_),
    .B(_00622_));
 sg13g2_xnor2_1 _19922_ (.Y(_00687_),
    .A(net250),
    .B(_00686_));
 sg13g2_xor2_1 _19923_ (.B(_00619_),
    .A(_00620_),
    .X(_00688_));
 sg13g2_inv_1 _19924_ (.Y(_00689_),
    .A(_00688_));
 sg13g2_nor2_1 _19925_ (.A(_06157_),
    .B(_00689_),
    .Y(_00690_));
 sg13g2_nand2_1 _19926_ (.Y(_00691_),
    .A(_00687_),
    .B(_00690_));
 sg13g2_o21ai_1 _19927_ (.B1(_00691_),
    .Y(_00692_),
    .A1(_06132_),
    .A2(_00686_));
 sg13g2_nand2_1 _19928_ (.Y(_00694_),
    .A(_00685_),
    .B(_00692_));
 sg13g2_o21ai_1 _19929_ (.B1(_00694_),
    .Y(_00695_),
    .A1(_06172_),
    .A2(_00684_));
 sg13g2_xnor2_1 _19930_ (.Y(_00696_),
    .A(net249),
    .B(_00681_));
 sg13g2_nand2_1 _19931_ (.Y(_00697_),
    .A(_00695_),
    .B(_00696_));
 sg13g2_o21ai_1 _19932_ (.B1(_00697_),
    .Y(_00698_),
    .A1(_06178_),
    .A2(_00681_));
 sg13g2_xnor2_1 _19933_ (.Y(_00699_),
    .A(net251),
    .B(_00677_));
 sg13g2_nand2_1 _19934_ (.Y(_00700_),
    .A(_00698_),
    .B(_00699_));
 sg13g2_o21ai_1 _19935_ (.B1(_00700_),
    .Y(_00701_),
    .A1(_00153_),
    .A2(_00677_));
 sg13g2_xnor2_1 _19936_ (.Y(_00702_),
    .A(_00642_),
    .B(_00639_));
 sg13g2_xnor2_1 _19937_ (.Y(_00703_),
    .A(_06039_),
    .B(_00702_));
 sg13g2_nand2_1 _19938_ (.Y(_00705_),
    .A(_00701_),
    .B(_00703_));
 sg13g2_nand2_1 _19939_ (.Y(_00706_),
    .A(_00702_),
    .B(_06129_));
 sg13g2_nand2_1 _19940_ (.Y(_00707_),
    .A(_00705_),
    .B(_00706_));
 sg13g2_xnor2_1 _19941_ (.Y(_00708_),
    .A(_04311_),
    .B(_00675_));
 sg13g2_nand2_1 _19942_ (.Y(_00709_),
    .A(_00707_),
    .B(_00708_));
 sg13g2_o21ai_1 _19943_ (.B1(_00709_),
    .Y(_00710_),
    .A1(_00151_),
    .A2(_00675_));
 sg13g2_xor2_1 _19944_ (.B(_00673_),
    .A(_04372_),
    .X(_00711_));
 sg13g2_nand2_1 _19945_ (.Y(_00712_),
    .A(_00710_),
    .B(_00711_));
 sg13g2_o21ai_1 _19946_ (.B1(_00712_),
    .Y(_00713_),
    .A1(_06192_),
    .A2(_00674_));
 sg13g2_xor2_1 _19947_ (.B(_00670_),
    .A(_04413_),
    .X(_00714_));
 sg13g2_nand2_1 _19948_ (.Y(_00716_),
    .A(_00713_),
    .B(_00714_));
 sg13g2_o21ai_1 _19949_ (.B1(_00716_),
    .Y(_00717_),
    .A1(_00149_),
    .A2(_00672_));
 sg13g2_xnor2_1 _19950_ (.Y(_00718_),
    .A(_00663_),
    .B(_00717_));
 sg13g2_buf_1 _19951_ (.A(net171),
    .X(_00719_));
 sg13g2_buf_1 _19952_ (.A(net155),
    .X(_00720_));
 sg13g2_nor2_1 _19953_ (.A(_06200_),
    .B(_00662_),
    .Y(_00721_));
 sg13g2_inv_1 _19954_ (.Y(_00722_),
    .A(_00662_));
 sg13g2_nor2b_1 _19955_ (.A(_00722_),
    .B_N(_06200_),
    .Y(_00723_));
 sg13g2_nor2_1 _19956_ (.A(_00721_),
    .B(_00723_),
    .Y(_00724_));
 sg13g2_inv_1 _19957_ (.Y(_00725_),
    .A(_00149_));
 sg13g2_nor2_1 _19958_ (.A(_00725_),
    .B(_00672_),
    .Y(_00727_));
 sg13g2_inv_1 _19959_ (.Y(_00728_),
    .A(_00153_));
 sg13g2_nor2_1 _19960_ (.A(_00728_),
    .B(_00677_),
    .Y(_00729_));
 sg13g2_xor2_1 _19961_ (.B(_00681_),
    .A(_06178_),
    .X(_00730_));
 sg13g2_inv_1 _19962_ (.Y(_00731_),
    .A(_06172_));
 sg13g2_xnor2_1 _19963_ (.Y(_00732_),
    .A(_06132_),
    .B(_00686_));
 sg13g2_nand2_1 _19964_ (.Y(_00733_),
    .A(_00689_),
    .B(_06136_));
 sg13g2_nor2b_1 _19965_ (.A(_00686_),
    .B_N(_06132_),
    .Y(_00734_));
 sg13g2_a21oi_1 _19966_ (.A1(_00732_),
    .A2(_00733_),
    .Y(_00735_),
    .B1(_00734_));
 sg13g2_xnor2_1 _19967_ (.Y(_00736_),
    .A(_06172_),
    .B(_00684_));
 sg13g2_nand2b_1 _19968_ (.Y(_00738_),
    .B(_00736_),
    .A_N(_00735_));
 sg13g2_o21ai_1 _19969_ (.B1(_00738_),
    .Y(_00739_),
    .A1(_00731_),
    .A2(_00684_));
 sg13g2_nand2b_1 _19970_ (.Y(_00740_),
    .B(_00739_),
    .A_N(_00730_));
 sg13g2_nand3_1 _19971_ (.B(_00680_),
    .C(_06178_),
    .A(_00679_),
    .Y(_00741_));
 sg13g2_nand2_1 _19972_ (.Y(_00742_),
    .A(_00740_),
    .B(_00741_));
 sg13g2_nand2_1 _19973_ (.Y(_00743_),
    .A(_00677_),
    .B(_00728_));
 sg13g2_o21ai_1 _19974_ (.B1(_00743_),
    .Y(_00744_),
    .A1(_00729_),
    .A2(_00742_));
 sg13g2_nand2_1 _19975_ (.Y(_00745_),
    .A(_00702_),
    .B(_00152_));
 sg13g2_nor2_1 _19976_ (.A(_00152_),
    .B(_00702_),
    .Y(_00746_));
 sg13g2_a21oi_2 _19977_ (.B1(_00746_),
    .Y(_00747_),
    .A2(_00745_),
    .A1(_00744_));
 sg13g2_inv_1 _19978_ (.Y(_00749_),
    .A(_00151_));
 sg13g2_nand2_1 _19979_ (.Y(_00750_),
    .A(_00675_),
    .B(_00749_));
 sg13g2_nor2_1 _19980_ (.A(_00749_),
    .B(_00675_),
    .Y(_00751_));
 sg13g2_a221oi_1 _19981_ (.B2(_00750_),
    .C1(_00751_),
    .B1(_00747_),
    .A1(_06192_),
    .Y(_00752_),
    .A2(_00673_));
 sg13g2_nand2b_1 _19982_ (.Y(_00753_),
    .B(_00674_),
    .A_N(_06192_));
 sg13g2_nor2b_1 _19983_ (.A(_00752_),
    .B_N(_00753_),
    .Y(_00754_));
 sg13g2_xnor2_1 _19984_ (.Y(_00755_),
    .A(_00725_),
    .B(_00670_));
 sg13g2_nand2_1 _19985_ (.Y(_00756_),
    .A(_00754_),
    .B(_00755_));
 sg13g2_nand2b_1 _19986_ (.Y(_00757_),
    .B(_00756_),
    .A_N(_00727_));
 sg13g2_xor2_1 _19987_ (.B(_00757_),
    .A(_00724_),
    .X(_00758_));
 sg13g2_nor2_1 _19988_ (.A(net142),
    .B(_00758_),
    .Y(_00760_));
 sg13g2_a21oi_1 _19989_ (.A1(_00718_),
    .A2(net142),
    .Y(_00761_),
    .B1(_00760_));
 sg13g2_xnor2_1 _19990_ (.Y(_00762_),
    .A(net83),
    .B(_00761_));
 sg13g2_xor2_1 _19991_ (.B(_00754_),
    .A(_00755_),
    .X(_00763_));
 sg13g2_xor2_1 _19992_ (.B(_00713_),
    .A(_00714_),
    .X(_00764_));
 sg13g2_buf_1 _19993_ (.A(net167),
    .X(_00765_));
 sg13g2_mux2_1 _19994_ (.A0(_00763_),
    .A1(_00764_),
    .S(net141),
    .X(_00766_));
 sg13g2_buf_1 _19995_ (.A(_00766_),
    .X(_00767_));
 sg13g2_nor2b_1 _19996_ (.A(_00762_),
    .B_N(_00767_),
    .Y(_00768_));
 sg13g2_nand2b_1 _19997_ (.Y(_00769_),
    .B(_00762_),
    .A_N(_00767_));
 sg13g2_nor2b_1 _19998_ (.A(_00768_),
    .B_N(_00769_),
    .Y(_00771_));
 sg13g2_xor2_1 _19999_ (.B(_00698_),
    .A(_00699_),
    .X(_00772_));
 sg13g2_nand2b_1 _20000_ (.Y(_00773_),
    .B(_00743_),
    .A_N(_00729_));
 sg13g2_xnor2_1 _20001_ (.Y(_00774_),
    .A(_00742_),
    .B(_00773_));
 sg13g2_inv_1 _20002_ (.Y(_00775_),
    .A(_00774_));
 sg13g2_nor2_1 _20003_ (.A(net171),
    .B(_00775_),
    .Y(_00776_));
 sg13g2_a21oi_1 _20004_ (.A1(net171),
    .A2(_00772_),
    .Y(_00777_),
    .B1(_00776_));
 sg13g2_xnor2_1 _20005_ (.Y(_00778_),
    .A(net83),
    .B(_00777_));
 sg13g2_inv_1 _20006_ (.Y(_00779_),
    .A(_00778_));
 sg13g2_xnor2_1 _20007_ (.Y(_00780_),
    .A(_00730_),
    .B(_00739_));
 sg13g2_xnor2_1 _20008_ (.Y(_00782_),
    .A(_00696_),
    .B(_00695_));
 sg13g2_nor2_1 _20009_ (.A(net171),
    .B(_00782_),
    .Y(_00783_));
 sg13g2_a21o_1 _20010_ (.A2(_00780_),
    .A1(_00719_),
    .B1(_00783_),
    .X(_00784_));
 sg13g2_inv_1 _20011_ (.Y(_00785_),
    .A(_00784_));
 sg13g2_nand2_1 _20012_ (.Y(_00786_),
    .A(_00779_),
    .B(_00785_));
 sg13g2_nor2_1 _20013_ (.A(net171),
    .B(_00780_),
    .Y(_00787_));
 sg13g2_a21oi_1 _20014_ (.A1(net171),
    .A2(_00782_),
    .Y(_00788_),
    .B1(_00787_));
 sg13g2_xnor2_1 _20015_ (.Y(_00789_),
    .A(_02391_),
    .B(_00788_));
 sg13g2_xor2_1 _20016_ (.B(_00685_),
    .A(_00692_),
    .X(_00790_));
 sg13g2_xor2_1 _20017_ (.B(_00736_),
    .A(_00735_),
    .X(_00791_));
 sg13g2_nor2_1 _20018_ (.A(net167),
    .B(_00791_),
    .Y(_00793_));
 sg13g2_a21o_1 _20019_ (.A2(_00790_),
    .A1(net167),
    .B1(_00793_),
    .X(_00794_));
 sg13g2_inv_1 _20020_ (.Y(_00795_),
    .A(_00794_));
 sg13g2_nand2_1 _20021_ (.Y(_00796_),
    .A(_00789_),
    .B(_00795_));
 sg13g2_nor2_1 _20022_ (.A(net167),
    .B(_00790_),
    .Y(_00797_));
 sg13g2_a21oi_1 _20023_ (.A1(net167),
    .A2(_00791_),
    .Y(_00798_),
    .B1(_00797_));
 sg13g2_xnor2_1 _20024_ (.Y(_00799_),
    .A(net102),
    .B(_00798_));
 sg13g2_xnor2_1 _20025_ (.Y(_00800_),
    .A(_00733_),
    .B(_00732_));
 sg13g2_inv_1 _20026_ (.Y(_00801_),
    .A(_00690_));
 sg13g2_xnor2_1 _20027_ (.Y(_00802_),
    .A(_00801_),
    .B(_00687_));
 sg13g2_nor2_1 _20028_ (.A(net171),
    .B(_00802_),
    .Y(_00804_));
 sg13g2_a21oi_1 _20029_ (.A1(net171),
    .A2(_00800_),
    .Y(_00805_),
    .B1(_00804_));
 sg13g2_nand2_1 _20030_ (.Y(_00806_),
    .A(_00799_),
    .B(_00805_));
 sg13g2_xnor2_1 _20031_ (.Y(_00807_),
    .A(_04205_),
    .B(_00688_));
 sg13g2_nor2_1 _20032_ (.A(net167),
    .B(_00802_),
    .Y(_00808_));
 sg13g2_a21oi_1 _20033_ (.A1(net167),
    .A2(_00800_),
    .Y(_00809_),
    .B1(_00808_));
 sg13g2_xnor2_1 _20034_ (.Y(_00810_),
    .A(net102),
    .B(_00809_));
 sg13g2_nand2b_1 _20035_ (.Y(_00811_),
    .B(_00810_),
    .A_N(_00807_));
 sg13g2_nor2_1 _20036_ (.A(_00805_),
    .B(_00799_),
    .Y(_00812_));
 sg13g2_a21oi_1 _20037_ (.A1(_00806_),
    .A2(_00811_),
    .Y(_00813_),
    .B1(_00812_));
 sg13g2_nor2_1 _20038_ (.A(_00795_),
    .B(_00789_),
    .Y(_00815_));
 sg13g2_a21oi_1 _20039_ (.A1(_00796_),
    .A2(_00813_),
    .Y(_00816_),
    .B1(_00815_));
 sg13g2_inv_1 _20040_ (.Y(_00817_),
    .A(_00816_));
 sg13g2_nor2_1 _20041_ (.A(_00785_),
    .B(_00779_),
    .Y(_00818_));
 sg13g2_a21oi_1 _20042_ (.A1(_00786_),
    .A2(_00817_),
    .Y(_00819_),
    .B1(_00818_));
 sg13g2_inv_1 _20043_ (.Y(_00820_),
    .A(_00819_));
 sg13g2_xnor2_1 _20044_ (.Y(_00821_),
    .A(_00703_),
    .B(_00701_));
 sg13g2_nor2b_1 _20045_ (.A(_00746_),
    .B_N(_00745_),
    .Y(_00822_));
 sg13g2_xnor2_1 _20046_ (.Y(_00823_),
    .A(_00744_),
    .B(_00822_));
 sg13g2_nor2_1 _20047_ (.A(net155),
    .B(_00823_),
    .Y(_00824_));
 sg13g2_a21oi_1 _20048_ (.A1(_00821_),
    .A2(net155),
    .Y(_00826_),
    .B1(_00824_));
 sg13g2_xnor2_1 _20049_ (.Y(_00827_),
    .A(_02391_),
    .B(_00826_));
 sg13g2_nand2_1 _20050_ (.Y(_00828_),
    .A(_00772_),
    .B(net167));
 sg13g2_o21ai_1 _20051_ (.B1(_00828_),
    .Y(_00829_),
    .A1(_00765_),
    .A2(_00775_));
 sg13g2_inv_1 _20052_ (.Y(_00830_),
    .A(_00829_));
 sg13g2_nand2_1 _20053_ (.Y(_00831_),
    .A(_00827_),
    .B(_00830_));
 sg13g2_nor2_1 _20054_ (.A(_00830_),
    .B(_00827_),
    .Y(_00832_));
 sg13g2_a21o_1 _20055_ (.A2(_00831_),
    .A1(_00820_),
    .B1(_00832_),
    .X(_00833_));
 sg13g2_nor2b_1 _20056_ (.A(_00751_),
    .B_N(_00750_),
    .Y(_00834_));
 sg13g2_xnor2_1 _20057_ (.Y(_00835_),
    .A(_00747_),
    .B(_00834_));
 sg13g2_xnor2_1 _20058_ (.Y(_00837_),
    .A(_00708_),
    .B(_00707_));
 sg13g2_mux2_1 _20059_ (.A0(_00835_),
    .A1(_00837_),
    .S(net155),
    .X(_00838_));
 sg13g2_xnor2_1 _20060_ (.Y(_00839_),
    .A(_02328_),
    .B(_00838_));
 sg13g2_nand2_1 _20061_ (.Y(_00840_),
    .A(_00823_),
    .B(net155));
 sg13g2_o21ai_1 _20062_ (.B1(_00840_),
    .Y(_00841_),
    .A1(net155),
    .A2(_00821_));
 sg13g2_inv_1 _20063_ (.Y(_00842_),
    .A(_00841_));
 sg13g2_nand2_1 _20064_ (.Y(_00843_),
    .A(_00839_),
    .B(_00842_));
 sg13g2_nor2_1 _20065_ (.A(_00842_),
    .B(_00839_),
    .Y(_00844_));
 sg13g2_a21o_1 _20066_ (.A2(_00843_),
    .A1(_00833_),
    .B1(_00844_),
    .X(_00845_));
 sg13g2_nand2_1 _20067_ (.Y(_00846_),
    .A(_00673_),
    .B(_06192_));
 sg13g2_nand2_1 _20068_ (.Y(_00848_),
    .A(_00753_),
    .B(_00846_));
 sg13g2_a21oi_1 _20069_ (.A1(_00747_),
    .A2(_00750_),
    .Y(_00849_),
    .B1(_00751_));
 sg13g2_xor2_1 _20070_ (.B(_00849_),
    .A(_00848_),
    .X(_00850_));
 sg13g2_xnor2_1 _20071_ (.Y(_00851_),
    .A(_00711_),
    .B(_00710_));
 sg13g2_nor2_1 _20072_ (.A(net141),
    .B(_00851_),
    .Y(_00852_));
 sg13g2_a21oi_1 _20073_ (.A1(net141),
    .A2(_00850_),
    .Y(_00853_),
    .B1(_00852_));
 sg13g2_xnor2_1 _20074_ (.Y(_00854_),
    .A(_02328_),
    .B(_00853_));
 sg13g2_nor2_1 _20075_ (.A(_00765_),
    .B(_00835_),
    .Y(_00855_));
 sg13g2_nand2b_1 _20076_ (.Y(_00856_),
    .B(net141),
    .A_N(_00837_));
 sg13g2_nand2b_1 _20077_ (.Y(_00857_),
    .B(_00856_),
    .A_N(_00855_));
 sg13g2_inv_1 _20078_ (.Y(_00859_),
    .A(_00857_));
 sg13g2_nand2_1 _20079_ (.Y(_00860_),
    .A(_00854_),
    .B(_00859_));
 sg13g2_nor2_1 _20080_ (.A(_00859_),
    .B(_00854_),
    .Y(_00861_));
 sg13g2_a21o_1 _20081_ (.A2(_00860_),
    .A1(_00845_),
    .B1(_00861_),
    .X(_00862_));
 sg13g2_buf_1 _20082_ (.A(_00862_),
    .X(_00863_));
 sg13g2_mux2_1 _20083_ (.A0(_00763_),
    .A1(_00764_),
    .S(_00719_),
    .X(_00864_));
 sg13g2_xnor2_1 _20084_ (.Y(_00865_),
    .A(net83),
    .B(_00864_));
 sg13g2_nand2_1 _20085_ (.Y(_00866_),
    .A(_00850_),
    .B(net155));
 sg13g2_o21ai_1 _20086_ (.B1(_00866_),
    .Y(_00867_),
    .A1(net155),
    .A2(_00851_));
 sg13g2_inv_1 _20087_ (.Y(_00868_),
    .A(_00867_));
 sg13g2_nand2_1 _20088_ (.Y(_00870_),
    .A(_00865_),
    .B(_00868_));
 sg13g2_nor2_1 _20089_ (.A(_00868_),
    .B(_00865_),
    .Y(_00871_));
 sg13g2_a21o_1 _20090_ (.A2(_00870_),
    .A1(_00863_),
    .B1(_00871_),
    .X(_00872_));
 sg13g2_xnor2_1 _20091_ (.Y(_00873_),
    .A(_00771_),
    .B(_00872_));
 sg13g2_xnor2_1 _20092_ (.Y(_00874_),
    .A(net70),
    .B(_00873_));
 sg13g2_xnor2_1 _20093_ (.Y(_00875_),
    .A(net185),
    .B(_00838_));
 sg13g2_nor2b_1 _20094_ (.A(_00874_),
    .B_N(_00875_),
    .Y(_00876_));
 sg13g2_xor2_1 _20095_ (.B(_00874_),
    .A(_00875_),
    .X(_00877_));
 sg13g2_buf_1 _20096_ (.A(net94),
    .X(_00878_));
 sg13g2_xnor2_1 _20097_ (.Y(_00879_),
    .A(_00878_),
    .B(_00867_));
 sg13g2_nor2b_1 _20098_ (.A(_00877_),
    .B_N(_00879_),
    .Y(_00881_));
 sg13g2_nor2_1 _20099_ (.A(_00876_),
    .B(_00881_),
    .Y(_00882_));
 sg13g2_xnor2_1 _20100_ (.Y(_00883_),
    .A(net82),
    .B(_00767_));
 sg13g2_xnor2_1 _20101_ (.Y(_00884_),
    .A(net178),
    .B(_00853_));
 sg13g2_nor2b_1 _20102_ (.A(_00871_),
    .B_N(_00870_),
    .Y(_00885_));
 sg13g2_nand3_1 _20103_ (.B(_00863_),
    .C(_00885_),
    .A(_00771_),
    .Y(_00886_));
 sg13g2_a21oi_1 _20104_ (.A1(_00769_),
    .A2(_00871_),
    .Y(_00887_),
    .B1(_00768_));
 sg13g2_nand2_1 _20105_ (.Y(_00888_),
    .A(_00886_),
    .B(_00887_));
 sg13g2_nand2_1 _20106_ (.Y(_00889_),
    .A(_00758_),
    .B(net142));
 sg13g2_o21ai_1 _20107_ (.B1(_00889_),
    .Y(_00890_),
    .A1(net142),
    .A2(_00718_));
 sg13g2_inv_1 _20108_ (.Y(_00892_),
    .A(_00890_));
 sg13g2_nor2_1 _20109_ (.A(net238),
    .B(_06331_),
    .Y(_00893_));
 sg13g2_nor2_1 _20110_ (.A(_06330_),
    .B(_06488_),
    .Y(_00894_));
 sg13g2_nor2_2 _20111_ (.A(_00893_),
    .B(_00894_),
    .Y(_00895_));
 sg13g2_inv_1 _20112_ (.Y(_00896_),
    .A(_00613_));
 sg13g2_nand2_1 _20113_ (.Y(_00897_),
    .A(_00669_),
    .B(_00651_));
 sg13g2_a21oi_1 _20114_ (.A1(_00613_),
    .A2(_00650_),
    .Y(_00898_),
    .B1(_00611_));
 sg13g2_o21ai_1 _20115_ (.B1(_00898_),
    .Y(_00899_),
    .A1(_00896_),
    .A2(_00897_));
 sg13g2_xnor2_1 _20116_ (.Y(_00900_),
    .A(_00895_),
    .B(_00899_));
 sg13g2_xnor2_1 _20117_ (.Y(_00901_),
    .A(_04495_),
    .B(_00900_));
 sg13g2_nand2_1 _20118_ (.Y(_00903_),
    .A(_00717_),
    .B(_00663_));
 sg13g2_o21ai_1 _20119_ (.B1(_00903_),
    .Y(_00904_),
    .A1(_06200_),
    .A2(_00722_));
 sg13g2_xor2_1 _20120_ (.B(_00904_),
    .A(_00901_),
    .X(_00905_));
 sg13g2_inv_1 _20121_ (.Y(_00906_),
    .A(_00905_));
 sg13g2_nor2b_1 _20122_ (.A(_00900_),
    .B_N(_06202_),
    .Y(_00907_));
 sg13g2_nor2b_1 _20123_ (.A(_06202_),
    .B_N(_00900_),
    .Y(_00908_));
 sg13g2_nor2_1 _20124_ (.A(_00907_),
    .B(_00908_),
    .Y(_00909_));
 sg13g2_nor2_1 _20125_ (.A(_00727_),
    .B(_00723_),
    .Y(_00910_));
 sg13g2_a21oi_1 _20126_ (.A1(_00756_),
    .A2(_00910_),
    .Y(_00911_),
    .B1(_00721_));
 sg13g2_xor2_1 _20127_ (.B(_00911_),
    .A(_00909_),
    .X(_00912_));
 sg13g2_nor2_1 _20128_ (.A(net142),
    .B(_00912_),
    .Y(_00914_));
 sg13g2_a21oi_1 _20129_ (.A1(_00906_),
    .A2(net142),
    .Y(_00915_),
    .B1(_00914_));
 sg13g2_xnor2_1 _20130_ (.Y(_00916_),
    .A(net83),
    .B(_00915_));
 sg13g2_nor2_1 _20131_ (.A(_00892_),
    .B(_00916_),
    .Y(_00917_));
 sg13g2_nand2_1 _20132_ (.Y(_00918_),
    .A(_00916_),
    .B(_00892_));
 sg13g2_inv_1 _20133_ (.Y(_00919_),
    .A(_00918_));
 sg13g2_nor2_1 _20134_ (.A(_00917_),
    .B(_00919_),
    .Y(_00920_));
 sg13g2_xnor2_1 _20135_ (.Y(_00921_),
    .A(_00888_),
    .B(_00920_));
 sg13g2_xnor2_1 _20136_ (.Y(_00922_),
    .A(net70),
    .B(_00921_));
 sg13g2_xnor2_1 _20137_ (.Y(_00923_),
    .A(_00884_),
    .B(_00922_));
 sg13g2_xor2_1 _20138_ (.B(_00923_),
    .A(_00883_),
    .X(_00924_));
 sg13g2_nor2_1 _20139_ (.A(_00882_),
    .B(_00924_),
    .Y(_00925_));
 sg13g2_nor2b_1 _20140_ (.A(_00832_),
    .B_N(_00831_),
    .Y(_00926_));
 sg13g2_xnor2_1 _20141_ (.Y(_00927_),
    .A(_00819_),
    .B(_00926_));
 sg13g2_xnor2_1 _20142_ (.Y(_00928_),
    .A(net71),
    .B(_00927_));
 sg13g2_xnor2_1 _20143_ (.Y(_00929_),
    .A(net178),
    .B(_00798_));
 sg13g2_nor2b_1 _20144_ (.A(_00928_),
    .B_N(_00929_),
    .Y(_00930_));
 sg13g2_xor2_1 _20145_ (.B(_00928_),
    .A(_00929_),
    .X(_00931_));
 sg13g2_xnor2_1 _20146_ (.Y(_00932_),
    .A(net94),
    .B(_00784_));
 sg13g2_nor2b_1 _20147_ (.A(_00931_),
    .B_N(_00932_),
    .Y(_00933_));
 sg13g2_nor2_1 _20148_ (.A(_00930_),
    .B(_00933_),
    .Y(_00935_));
 sg13g2_xnor2_1 _20149_ (.Y(_00936_),
    .A(net94),
    .B(_00829_));
 sg13g2_xnor2_1 _20150_ (.Y(_00937_),
    .A(net185),
    .B(_00788_));
 sg13g2_nor2b_1 _20151_ (.A(_00844_),
    .B_N(_00843_),
    .Y(_00938_));
 sg13g2_xnor2_1 _20152_ (.Y(_00939_),
    .A(_00833_),
    .B(_00938_));
 sg13g2_xnor2_1 _20153_ (.Y(_00940_),
    .A(_02645_),
    .B(_00939_));
 sg13g2_xnor2_1 _20154_ (.Y(_00941_),
    .A(_00937_),
    .B(_00940_));
 sg13g2_xor2_1 _20155_ (.B(_00941_),
    .A(_00936_),
    .X(_00942_));
 sg13g2_xor2_1 _20156_ (.B(_00931_),
    .A(_00932_),
    .X(_00943_));
 sg13g2_nor2b_1 _20157_ (.A(_00818_),
    .B_N(_00786_),
    .Y(_00944_));
 sg13g2_xnor2_1 _20158_ (.Y(_00946_),
    .A(_00817_),
    .B(_00944_));
 sg13g2_xnor2_1 _20159_ (.Y(_00947_),
    .A(net70),
    .B(_00946_));
 sg13g2_xnor2_1 _20160_ (.Y(_00948_),
    .A(_03228_),
    .B(_00809_));
 sg13g2_nor2b_1 _20161_ (.A(_00947_),
    .B_N(_00948_),
    .Y(_00949_));
 sg13g2_xor2_1 _20162_ (.B(_00947_),
    .A(_00948_),
    .X(_00950_));
 sg13g2_xnor2_1 _20163_ (.Y(_00951_),
    .A(_02785_),
    .B(_00794_));
 sg13g2_nor2b_1 _20164_ (.A(_00950_),
    .B_N(_00951_),
    .Y(_00952_));
 sg13g2_nor2_1 _20165_ (.A(_00949_),
    .B(_00952_),
    .Y(_00953_));
 sg13g2_nand2_1 _20166_ (.Y(_00954_),
    .A(_00943_),
    .B(_00953_));
 sg13g2_xor2_1 _20167_ (.B(_00950_),
    .A(_00951_),
    .X(_00955_));
 sg13g2_xnor2_1 _20168_ (.Y(_00957_),
    .A(net185),
    .B(_00807_));
 sg13g2_xnor2_1 _20169_ (.Y(_00958_),
    .A(_02785_),
    .B(_00805_));
 sg13g2_nor2_1 _20170_ (.A(_00957_),
    .B(_00958_),
    .Y(_00959_));
 sg13g2_nand2b_1 _20171_ (.Y(_00960_),
    .B(_00796_),
    .A_N(_00815_));
 sg13g2_xnor2_1 _20172_ (.Y(_00961_),
    .A(_00813_),
    .B(_00960_));
 sg13g2_xnor2_1 _20173_ (.Y(_00962_),
    .A(_02627_),
    .B(_00961_));
 sg13g2_nand2_1 _20174_ (.Y(_00963_),
    .A(_00958_),
    .B(_00957_));
 sg13g2_o21ai_1 _20175_ (.B1(_00963_),
    .Y(_00964_),
    .A1(_00959_),
    .A2(_00962_));
 sg13g2_nor2b_1 _20176_ (.A(_00955_),
    .B_N(_00964_),
    .Y(_00965_));
 sg13g2_nor2_1 _20177_ (.A(_00953_),
    .B(_00943_),
    .Y(_00966_));
 sg13g2_a21oi_1 _20178_ (.A1(_00954_),
    .A2(_00965_),
    .Y(_00968_),
    .B1(_00966_));
 sg13g2_inv_1 _20179_ (.Y(_00969_),
    .A(_00935_));
 sg13g2_xnor2_1 _20180_ (.Y(_00970_),
    .A(_00969_),
    .B(_00942_));
 sg13g2_nand2b_1 _20181_ (.Y(_00971_),
    .B(_00970_),
    .A_N(_00968_));
 sg13g2_o21ai_1 _20182_ (.B1(_00971_),
    .Y(_00972_),
    .A1(_00935_),
    .A2(_00942_));
 sg13g2_xnor2_1 _20183_ (.Y(_00973_),
    .A(net82),
    .B(_00841_));
 sg13g2_xnor2_1 _20184_ (.Y(_00974_),
    .A(net185),
    .B(_00777_));
 sg13g2_nand2b_1 _20185_ (.Y(_00975_),
    .B(_00860_),
    .A_N(_00861_));
 sg13g2_xnor2_1 _20186_ (.Y(_00976_),
    .A(_02627_),
    .B(_00845_));
 sg13g2_xnor2_1 _20187_ (.Y(_00977_),
    .A(_00975_),
    .B(_00976_));
 sg13g2_xor2_1 _20188_ (.B(_00977_),
    .A(_00974_),
    .X(_00979_));
 sg13g2_xor2_1 _20189_ (.B(_00979_),
    .A(_00973_),
    .X(_00980_));
 sg13g2_nand2_1 _20190_ (.Y(_00981_),
    .A(_00940_),
    .B(_00937_));
 sg13g2_nor2_1 _20191_ (.A(_00937_),
    .B(_00940_),
    .Y(_00982_));
 sg13g2_a21oi_1 _20192_ (.A1(_00981_),
    .A2(_00936_),
    .Y(_00983_),
    .B1(_00982_));
 sg13g2_nand2_1 _20193_ (.Y(_00984_),
    .A(_00980_),
    .B(_00983_));
 sg13g2_nand2_1 _20194_ (.Y(_00985_),
    .A(_00972_),
    .B(_00984_));
 sg13g2_or2_1 _20195_ (.X(_00986_),
    .B(_00980_),
    .A(_00983_));
 sg13g2_nand2_1 _20196_ (.Y(_00987_),
    .A(_00985_),
    .B(_00986_));
 sg13g2_xnor2_1 _20197_ (.Y(_00988_),
    .A(_00878_),
    .B(_00857_));
 sg13g2_xnor2_1 _20198_ (.Y(_00990_),
    .A(net185),
    .B(_00826_));
 sg13g2_xnor2_1 _20199_ (.Y(_00991_),
    .A(_00863_),
    .B(_00885_));
 sg13g2_xnor2_1 _20200_ (.Y(_00992_),
    .A(net70),
    .B(_00991_));
 sg13g2_xnor2_1 _20201_ (.Y(_00993_),
    .A(_00990_),
    .B(_00992_));
 sg13g2_xor2_1 _20202_ (.B(_00993_),
    .A(_00988_),
    .X(_00994_));
 sg13g2_nor2b_1 _20203_ (.A(_00977_),
    .B_N(_00974_),
    .Y(_00995_));
 sg13g2_nor2b_1 _20204_ (.A(_00979_),
    .B_N(_00973_),
    .Y(_00996_));
 sg13g2_nor2_1 _20205_ (.A(_00995_),
    .B(_00996_),
    .Y(_00997_));
 sg13g2_nand2_1 _20206_ (.Y(_00998_),
    .A(_00994_),
    .B(_00997_));
 sg13g2_nor2_1 _20207_ (.A(_00997_),
    .B(_00994_),
    .Y(_00999_));
 sg13g2_a21o_1 _20208_ (.A2(_00998_),
    .A1(_00987_),
    .B1(_00999_),
    .X(_01001_));
 sg13g2_xor2_1 _20209_ (.B(_00877_),
    .A(_00879_),
    .X(_01002_));
 sg13g2_nand2_1 _20210_ (.Y(_01003_),
    .A(_00992_),
    .B(_00990_));
 sg13g2_nor2_1 _20211_ (.A(_00990_),
    .B(_00992_),
    .Y(_01004_));
 sg13g2_a21oi_1 _20212_ (.A1(_01003_),
    .A2(_00988_),
    .Y(_01005_),
    .B1(_01004_));
 sg13g2_nand2_1 _20213_ (.Y(_01006_),
    .A(_01002_),
    .B(_01005_));
 sg13g2_nor2_1 _20214_ (.A(_01005_),
    .B(_01002_),
    .Y(_01007_));
 sg13g2_a21oi_1 _20215_ (.A1(_01001_),
    .A2(_01006_),
    .Y(_01008_),
    .B1(_01007_));
 sg13g2_nand2_1 _20216_ (.Y(_01009_),
    .A(_00924_),
    .B(_00882_));
 sg13g2_nand2b_1 _20217_ (.Y(_01010_),
    .B(_01009_),
    .A_N(_01008_));
 sg13g2_nand2b_1 _20218_ (.Y(_01012_),
    .B(_01010_),
    .A_N(_00925_));
 sg13g2_nand2_1 _20219_ (.Y(_01013_),
    .A(_00922_),
    .B(_00884_));
 sg13g2_nor2_1 _20220_ (.A(_00884_),
    .B(_00922_),
    .Y(_01014_));
 sg13g2_a21oi_1 _20221_ (.A1(_01013_),
    .A2(_00883_),
    .Y(_01015_),
    .B1(_01014_));
 sg13g2_xnor2_1 _20222_ (.Y(_01016_),
    .A(net82),
    .B(_00890_));
 sg13g2_xnor2_1 _20223_ (.Y(_01017_),
    .A(net185),
    .B(_00864_));
 sg13g2_nor2_1 _20224_ (.A(_00768_),
    .B(_00917_),
    .Y(_01018_));
 sg13g2_nand2_1 _20225_ (.Y(_01019_),
    .A(_00872_),
    .B(_00771_));
 sg13g2_a21oi_1 _20226_ (.A1(_01018_),
    .A2(_01019_),
    .Y(_01020_),
    .B1(_00919_));
 sg13g2_nand2_1 _20227_ (.Y(_01021_),
    .A(_00912_),
    .B(net142));
 sg13g2_o21ai_1 _20228_ (.B1(_01021_),
    .Y(_01023_),
    .A1(net142),
    .A2(_00906_));
 sg13g2_buf_1 _20229_ (.A(_01023_),
    .X(_01024_));
 sg13g2_inv_1 _20230_ (.Y(_01025_),
    .A(_06115_));
 sg13g2_xnor2_1 _20231_ (.Y(_01026_),
    .A(_05094_),
    .B(net219));
 sg13g2_nand2_1 _20232_ (.Y(_01027_),
    .A(_00613_),
    .B(_00895_));
 sg13g2_a21oi_1 _20233_ (.A1(_00895_),
    .A2(_00611_),
    .Y(_01028_),
    .B1(_00894_));
 sg13g2_o21ai_1 _20234_ (.B1(_01028_),
    .Y(_01029_),
    .A1(_01027_),
    .A2(_00661_));
 sg13g2_xnor2_1 _20235_ (.Y(_01030_),
    .A(_01026_),
    .B(_01029_));
 sg13g2_nor2_1 _20236_ (.A(_01025_),
    .B(_01030_),
    .Y(_01031_));
 sg13g2_nand2_1 _20237_ (.Y(_01032_),
    .A(_01030_),
    .B(_01025_));
 sg13g2_nor2b_1 _20238_ (.A(_01031_),
    .B_N(_01032_),
    .Y(_01034_));
 sg13g2_inv_1 _20239_ (.Y(_01035_),
    .A(_01034_));
 sg13g2_nand2_1 _20240_ (.Y(_01036_),
    .A(_00757_),
    .B(_00724_));
 sg13g2_nor2_1 _20241_ (.A(_00723_),
    .B(_00907_),
    .Y(_01037_));
 sg13g2_a21oi_1 _20242_ (.A1(_01036_),
    .A2(_01037_),
    .Y(_01038_),
    .B1(_00908_));
 sg13g2_xnor2_1 _20243_ (.Y(_01039_),
    .A(_01035_),
    .B(_01038_));
 sg13g2_nand2_1 _20244_ (.Y(_01040_),
    .A(_00904_),
    .B(_00901_));
 sg13g2_o21ai_1 _20245_ (.B1(_01040_),
    .Y(_01041_),
    .A1(_06202_),
    .A2(_00900_));
 sg13g2_xnor2_1 _20246_ (.Y(_01042_),
    .A(_01035_),
    .B(_01041_));
 sg13g2_nor2_1 _20247_ (.A(net141),
    .B(_01042_),
    .Y(_01043_));
 sg13g2_a21oi_1 _20248_ (.A1(_01039_),
    .A2(net141),
    .Y(_01045_),
    .B1(_01043_));
 sg13g2_xnor2_1 _20249_ (.Y(_01046_),
    .A(net102),
    .B(_01045_));
 sg13g2_xnor2_1 _20250_ (.Y(_01047_),
    .A(_01024_),
    .B(_01046_));
 sg13g2_xnor2_1 _20251_ (.Y(_01048_),
    .A(_01020_),
    .B(_01047_));
 sg13g2_xnor2_1 _20252_ (.Y(_01049_),
    .A(net70),
    .B(_01048_));
 sg13g2_xnor2_1 _20253_ (.Y(_01050_),
    .A(_01017_),
    .B(_01049_));
 sg13g2_xor2_1 _20254_ (.B(_01050_),
    .A(_01016_),
    .X(_01051_));
 sg13g2_nor2_1 _20255_ (.A(_01015_),
    .B(_01051_),
    .Y(_01052_));
 sg13g2_nand2_1 _20256_ (.Y(_01053_),
    .A(_01051_),
    .B(_01015_));
 sg13g2_nor2b_1 _20257_ (.A(_01052_),
    .B_N(_01053_),
    .Y(_01054_));
 sg13g2_xor2_1 _20258_ (.B(_01054_),
    .A(_01012_),
    .X(_01056_));
 sg13g2_inv_1 _20259_ (.Y(_01057_),
    .A(_01056_));
 sg13g2_nand2_1 _20260_ (.Y(_01058_),
    .A(_01049_),
    .B(_01017_));
 sg13g2_nor2_1 _20261_ (.A(_01017_),
    .B(_01049_),
    .Y(_01059_));
 sg13g2_a21oi_2 _20262_ (.B1(_01059_),
    .Y(_01060_),
    .A2(_01016_),
    .A1(_01058_));
 sg13g2_xnor2_1 _20263_ (.Y(_01061_),
    .A(net82),
    .B(_01024_));
 sg13g2_xnor2_1 _20264_ (.Y(_01062_),
    .A(net178),
    .B(_00761_));
 sg13g2_inv_1 _20265_ (.Y(_01063_),
    .A(_01024_));
 sg13g2_nand2_1 _20266_ (.Y(_01064_),
    .A(_00920_),
    .B(_00888_));
 sg13g2_nor2_1 _20267_ (.A(_01063_),
    .B(_01046_),
    .Y(_01065_));
 sg13g2_nor2_1 _20268_ (.A(_00917_),
    .B(_01065_),
    .Y(_01067_));
 sg13g2_a22oi_1 _20269_ (.Y(_01068_),
    .B1(_01064_),
    .B2(_01067_),
    .A2(_01063_),
    .A1(_01046_));
 sg13g2_buf_1 _20270_ (.A(_00720_),
    .X(_01069_));
 sg13g2_nand2_1 _20271_ (.Y(_01070_),
    .A(_01039_),
    .B(_00720_));
 sg13g2_o21ai_1 _20272_ (.B1(_01070_),
    .Y(_01071_),
    .A1(net139),
    .A2(_01042_));
 sg13g2_inv_1 _20273_ (.Y(_01072_),
    .A(_01071_));
 sg13g2_xnor2_1 _20274_ (.Y(_01073_),
    .A(_05134_),
    .B(net218));
 sg13g2_nand2_1 _20275_ (.Y(_01074_),
    .A(_00895_),
    .B(_01026_));
 sg13g2_inv_1 _20276_ (.Y(_01075_),
    .A(_00899_));
 sg13g2_nor2_1 _20277_ (.A(net219),
    .B(_06496_),
    .Y(_01076_));
 sg13g2_a21oi_1 _20278_ (.A1(_01026_),
    .A2(_00894_),
    .Y(_01078_),
    .B1(_01076_));
 sg13g2_o21ai_1 _20279_ (.B1(_01078_),
    .Y(_01079_),
    .A1(_01074_),
    .A2(_01075_));
 sg13g2_xnor2_1 _20280_ (.Y(_01080_),
    .A(_01073_),
    .B(_01079_));
 sg13g2_buf_1 _20281_ (.A(_01080_),
    .X(_01081_));
 sg13g2_xnor2_1 _20282_ (.Y(_01082_),
    .A(_00145_),
    .B(_01081_));
 sg13g2_nand3_1 _20283_ (.B(_01034_),
    .C(_00909_),
    .A(_00911_),
    .Y(_01083_));
 sg13g2_o21ai_1 _20284_ (.B1(_01032_),
    .Y(_01084_),
    .A1(_01031_),
    .A2(_00907_));
 sg13g2_nand2_1 _20285_ (.Y(_01085_),
    .A(_01083_),
    .B(_01084_));
 sg13g2_xor2_1 _20286_ (.B(_01085_),
    .A(_01082_),
    .X(_01086_));
 sg13g2_xnor2_1 _20287_ (.Y(_01087_),
    .A(_04573_),
    .B(_01081_));
 sg13g2_nand2_1 _20288_ (.Y(_01089_),
    .A(_01041_),
    .B(_01035_));
 sg13g2_o21ai_1 _20289_ (.B1(_01089_),
    .Y(_01090_),
    .A1(_06115_),
    .A2(_01030_));
 sg13g2_xnor2_1 _20290_ (.Y(_01091_),
    .A(_01087_),
    .B(_01090_));
 sg13g2_nor2_1 _20291_ (.A(net141),
    .B(_01091_),
    .Y(_01092_));
 sg13g2_a21oi_2 _20292_ (.B1(_01092_),
    .Y(_01093_),
    .A2(_01086_),
    .A1(net141));
 sg13g2_xnor2_1 _20293_ (.Y(_01094_),
    .A(net102),
    .B(_01093_));
 sg13g2_nor2_1 _20294_ (.A(_01072_),
    .B(_01094_),
    .Y(_01095_));
 sg13g2_nand2_1 _20295_ (.Y(_01096_),
    .A(_01094_),
    .B(_01072_));
 sg13g2_nand2b_1 _20296_ (.Y(_01097_),
    .B(_01096_),
    .A_N(_01095_));
 sg13g2_xnor2_1 _20297_ (.Y(_01098_),
    .A(_01068_),
    .B(_01097_));
 sg13g2_xnor2_1 _20298_ (.Y(_01100_),
    .A(net71),
    .B(_01098_));
 sg13g2_xor2_1 _20299_ (.B(_01100_),
    .A(_01062_),
    .X(_01101_));
 sg13g2_xor2_1 _20300_ (.B(_01101_),
    .A(_01061_),
    .X(_01102_));
 sg13g2_nand2_1 _20301_ (.Y(_01103_),
    .A(_01054_),
    .B(_01012_));
 sg13g2_nor2_1 _20302_ (.A(_01060_),
    .B(_01102_),
    .Y(_01104_));
 sg13g2_nor2_1 _20303_ (.A(_01052_),
    .B(_01104_),
    .Y(_01105_));
 sg13g2_a22oi_1 _20304_ (.Y(_01106_),
    .B1(_01103_),
    .B2(_01105_),
    .A2(_01102_),
    .A1(_01060_));
 sg13g2_nor2b_1 _20305_ (.A(_01100_),
    .B_N(_01062_),
    .Y(_01107_));
 sg13g2_nor2b_1 _20306_ (.A(_01101_),
    .B_N(_01061_),
    .Y(_01108_));
 sg13g2_nor2_1 _20307_ (.A(_01107_),
    .B(_01108_),
    .Y(_01109_));
 sg13g2_xnor2_1 _20308_ (.Y(_01111_),
    .A(net82),
    .B(_01071_));
 sg13g2_xnor2_1 _20309_ (.Y(_01112_),
    .A(net178),
    .B(_00915_));
 sg13g2_a21o_1 _20310_ (.A2(_01096_),
    .A1(_01068_),
    .B1(_01095_),
    .X(_01113_));
 sg13g2_nand2_1 _20311_ (.Y(_01114_),
    .A(_01086_),
    .B(_01069_));
 sg13g2_o21ai_1 _20312_ (.B1(_01114_),
    .Y(_01115_),
    .A1(_01069_),
    .A2(_01091_));
 sg13g2_inv_1 _20313_ (.Y(_01116_),
    .A(_01115_));
 sg13g2_xor2_1 _20314_ (.B(_06371_),
    .A(_05168_),
    .X(_01117_));
 sg13g2_a221oi_1 _20315_ (.B2(_01026_),
    .C1(_01076_),
    .B1(_01029_),
    .A1(_05134_),
    .Y(_01118_),
    .A2(_06361_));
 sg13g2_a21oi_1 _20316_ (.A1(_09173_),
    .A2(net218),
    .Y(_01119_),
    .B1(_01118_));
 sg13g2_xor2_1 _20317_ (.B(_01119_),
    .A(_01117_),
    .X(_01120_));
 sg13g2_or2_1 _20318_ (.X(_01122_),
    .B(_01120_),
    .A(_00106_));
 sg13g2_nand2_1 _20319_ (.Y(_01123_),
    .A(_01120_),
    .B(_00106_));
 sg13g2_nand2_1 _20320_ (.Y(_01124_),
    .A(_01122_),
    .B(_01123_));
 sg13g2_nor2_1 _20321_ (.A(_06206_),
    .B(_01081_),
    .Y(_01125_));
 sg13g2_nor2_1 _20322_ (.A(_01031_),
    .B(_01125_),
    .Y(_01126_));
 sg13g2_nand2_1 _20323_ (.Y(_01127_),
    .A(_01038_),
    .B(_01034_));
 sg13g2_a22oi_1 _20324_ (.Y(_01128_),
    .B1(_01126_),
    .B2(_01127_),
    .A2(_01081_),
    .A1(_06206_));
 sg13g2_xnor2_1 _20325_ (.Y(_01129_),
    .A(_01124_),
    .B(_01128_));
 sg13g2_inv_1 _20326_ (.Y(_01130_),
    .A(_01081_));
 sg13g2_a22oi_1 _20327_ (.Y(_01131_),
    .B1(_01087_),
    .B2(_01090_),
    .A2(_01130_),
    .A1(_06206_));
 sg13g2_xnor2_1 _20328_ (.Y(_01133_),
    .A(_01124_),
    .B(_01131_));
 sg13g2_mux2_1 _20329_ (.A0(_01129_),
    .A1(_01133_),
    .S(net139),
    .X(_01134_));
 sg13g2_xnor2_1 _20330_ (.Y(_01135_),
    .A(net102),
    .B(_01134_));
 sg13g2_nor2_1 _20331_ (.A(_01116_),
    .B(_01135_),
    .Y(_01136_));
 sg13g2_nand2_1 _20332_ (.Y(_01137_),
    .A(_01135_),
    .B(_01116_));
 sg13g2_nor2b_1 _20333_ (.A(_01136_),
    .B_N(_01137_),
    .Y(_01138_));
 sg13g2_xnor2_1 _20334_ (.Y(_01139_),
    .A(_01113_),
    .B(_01138_));
 sg13g2_xnor2_1 _20335_ (.Y(_01140_),
    .A(net70),
    .B(_01139_));
 sg13g2_xor2_1 _20336_ (.B(_01140_),
    .A(_01112_),
    .X(_01141_));
 sg13g2_xor2_1 _20337_ (.B(_01141_),
    .A(_01111_),
    .X(_01142_));
 sg13g2_xnor2_1 _20338_ (.Y(_01144_),
    .A(_01109_),
    .B(_01142_));
 sg13g2_xor2_1 _20339_ (.B(_01144_),
    .A(_01106_),
    .X(_01145_));
 sg13g2_buf_1 _20340_ (.A(_01145_),
    .X(_01146_));
 sg13g2_nor2_1 _20341_ (.A(_01057_),
    .B(_01146_),
    .Y(_01147_));
 sg13g2_nand2_1 _20342_ (.Y(_01148_),
    .A(_01146_),
    .B(_01057_));
 sg13g2_nand2b_1 _20343_ (.Y(_01149_),
    .B(_01148_),
    .A_N(_01147_));
 sg13g2_nor2b_1 _20344_ (.A(_00925_),
    .B_N(_01009_),
    .Y(_01150_));
 sg13g2_xnor2_1 _20345_ (.Y(_01151_),
    .A(_01008_),
    .B(_01150_));
 sg13g2_a21oi_1 _20346_ (.A1(_01012_),
    .A2(_01053_),
    .Y(_01152_),
    .B1(_01052_));
 sg13g2_xnor2_1 _20347_ (.Y(_01153_),
    .A(_01060_),
    .B(_01102_));
 sg13g2_xor2_1 _20348_ (.B(_01153_),
    .A(_01152_),
    .X(_01155_));
 sg13g2_xnor2_1 _20349_ (.Y(_01156_),
    .A(_01151_),
    .B(_01155_));
 sg13g2_nor2b_1 _20350_ (.A(_01007_),
    .B_N(_01006_),
    .Y(_01157_));
 sg13g2_xor2_1 _20351_ (.B(_01157_),
    .A(_01001_),
    .X(_01158_));
 sg13g2_inv_1 _20352_ (.Y(_01159_),
    .A(_01158_));
 sg13g2_nor2_1 _20353_ (.A(_01159_),
    .B(_01057_),
    .Y(_01160_));
 sg13g2_nand2b_1 _20354_ (.Y(_01161_),
    .B(_00998_),
    .A_N(_00999_));
 sg13g2_xnor2_1 _20355_ (.Y(_01162_),
    .A(_00987_),
    .B(_01161_));
 sg13g2_inv_1 _20356_ (.Y(_01163_),
    .A(_01162_));
 sg13g2_inv_1 _20357_ (.Y(_01164_),
    .A(_01151_));
 sg13g2_nor2_1 _20358_ (.A(_01163_),
    .B(_01164_),
    .Y(_01165_));
 sg13g2_nand2_1 _20359_ (.Y(_01166_),
    .A(_00986_),
    .B(_00984_));
 sg13g2_xor2_1 _20360_ (.B(_01166_),
    .A(_00972_),
    .X(_01167_));
 sg13g2_nor2_1 _20361_ (.A(_01167_),
    .B(_01159_),
    .Y(_01168_));
 sg13g2_xnor2_1 _20362_ (.Y(_01169_),
    .A(_00968_),
    .B(_00970_));
 sg13g2_inv_1 _20363_ (.Y(_01170_),
    .A(_01167_));
 sg13g2_xnor2_1 _20364_ (.Y(_01171_),
    .A(_00953_),
    .B(_00943_));
 sg13g2_xnor2_1 _20365_ (.Y(_01172_),
    .A(_00965_),
    .B(_01171_));
 sg13g2_xor2_1 _20366_ (.B(_01167_),
    .A(_01172_),
    .X(_01173_));
 sg13g2_xnor2_1 _20367_ (.Y(_01174_),
    .A(_00964_),
    .B(_00955_));
 sg13g2_inv_1 _20368_ (.Y(_01176_),
    .A(_01174_));
 sg13g2_inv_1 _20369_ (.Y(_01177_),
    .A(_01169_));
 sg13g2_nor2_1 _20370_ (.A(_01176_),
    .B(_01177_),
    .Y(_01178_));
 sg13g2_nor2b_1 _20371_ (.A(_01173_),
    .B_N(_01178_),
    .Y(_01179_));
 sg13g2_a21oi_1 _20372_ (.A1(_01170_),
    .A2(_01172_),
    .Y(_01180_),
    .B1(_01179_));
 sg13g2_xnor2_1 _20373_ (.Y(_01181_),
    .A(_01177_),
    .B(_01162_));
 sg13g2_nor2b_1 _20374_ (.A(_01180_),
    .B_N(_01181_),
    .Y(_01182_));
 sg13g2_a21oi_1 _20375_ (.A1(_01162_),
    .A2(_01169_),
    .Y(_01183_),
    .B1(_01182_));
 sg13g2_xnor2_1 _20376_ (.Y(_01184_),
    .A(_01167_),
    .B(_01158_));
 sg13g2_nand2b_1 _20377_ (.Y(_01185_),
    .B(_01184_),
    .A_N(_01183_));
 sg13g2_nor2b_1 _20378_ (.A(_01168_),
    .B_N(_01185_),
    .Y(_01187_));
 sg13g2_inv_1 _20379_ (.Y(_01188_),
    .A(_01187_));
 sg13g2_nand2_1 _20380_ (.Y(_01189_),
    .A(_01164_),
    .B(_01163_));
 sg13g2_o21ai_1 _20381_ (.B1(_01189_),
    .Y(_01190_),
    .A1(_01165_),
    .A2(_01188_));
 sg13g2_inv_1 _20382_ (.Y(_01191_),
    .A(_01190_));
 sg13g2_nand2_1 _20383_ (.Y(_01192_),
    .A(_01057_),
    .B(_01159_));
 sg13g2_o21ai_1 _20384_ (.B1(_01192_),
    .Y(_01193_),
    .A1(_01160_),
    .A2(_01191_));
 sg13g2_inv_1 _20385_ (.Y(_01194_),
    .A(_01155_));
 sg13g2_nor2_1 _20386_ (.A(_01164_),
    .B(_01194_),
    .Y(_01195_));
 sg13g2_inv_1 _20387_ (.Y(_01196_),
    .A(_01195_));
 sg13g2_o21ai_1 _20388_ (.B1(_01196_),
    .Y(_01198_),
    .A1(_01156_),
    .A2(_01193_));
 sg13g2_xor2_1 _20389_ (.B(_01198_),
    .A(_01149_),
    .X(_01199_));
 sg13g2_nor2_1 _20390_ (.A(_00610_),
    .B(_01199_),
    .Y(_01200_));
 sg13g2_inv_1 _20391_ (.Y(_01201_),
    .A(_00610_));
 sg13g2_nor2_1 _20392_ (.A(_01201_),
    .B(_01199_),
    .Y(_01202_));
 sg13g2_nand2_1 _20393_ (.Y(_01203_),
    .A(_01199_),
    .B(_01201_));
 sg13g2_nand2b_1 _20394_ (.Y(_01204_),
    .B(_01203_),
    .A_N(_01202_));
 sg13g2_nand3_1 _20395_ (.B(_00588_),
    .C(_00575_),
    .A(_00571_),
    .Y(_01205_));
 sg13g2_a21oi_1 _20396_ (.A1(_00577_),
    .A2(_00587_),
    .Y(_01206_),
    .B1(_00586_));
 sg13g2_nand2_1 _20397_ (.Y(_01207_),
    .A(_01205_),
    .B(_01206_));
 sg13g2_nand3_1 _20398_ (.B(_00582_),
    .C(_00598_),
    .A(_01207_),
    .Y(_01209_));
 sg13g2_a21oi_1 _20399_ (.A1(_00598_),
    .A2(_00590_),
    .Y(_01210_),
    .B1(_00597_));
 sg13g2_nand2_1 _20400_ (.Y(_01211_),
    .A(_01209_),
    .B(_01210_));
 sg13g2_xor2_1 _20401_ (.B(_01211_),
    .A(_00605_),
    .X(_01212_));
 sg13g2_xnor2_1 _20402_ (.Y(_01213_),
    .A(_01156_),
    .B(_01193_));
 sg13g2_nor2_1 _20403_ (.A(_01212_),
    .B(_01213_),
    .Y(_01214_));
 sg13g2_xor2_1 _20404_ (.B(_00592_),
    .A(_00598_),
    .X(_01215_));
 sg13g2_inv_1 _20405_ (.Y(_01216_),
    .A(_01160_));
 sg13g2_nand2_1 _20406_ (.Y(_01217_),
    .A(_01216_),
    .B(_01192_));
 sg13g2_xnor2_1 _20407_ (.Y(_01218_),
    .A(_01217_),
    .B(_01190_));
 sg13g2_xor2_1 _20408_ (.B(_01218_),
    .A(_01215_),
    .X(_01220_));
 sg13g2_xor2_1 _20409_ (.B(_01207_),
    .A(_00582_),
    .X(_01221_));
 sg13g2_nand2b_1 _20410_ (.Y(_01222_),
    .B(_01189_),
    .A_N(_01165_));
 sg13g2_xnor2_1 _20411_ (.Y(_01223_),
    .A(_01222_),
    .B(_01187_));
 sg13g2_inv_1 _20412_ (.Y(_01224_),
    .A(_01221_));
 sg13g2_xnor2_1 _20413_ (.Y(_01225_),
    .A(_01224_),
    .B(_01223_));
 sg13g2_xor2_1 _20414_ (.B(_00578_),
    .A(_00588_),
    .X(_01226_));
 sg13g2_xor2_1 _20415_ (.B(_01183_),
    .A(_01184_),
    .X(_01227_));
 sg13g2_xor2_1 _20416_ (.B(_01227_),
    .A(_01226_),
    .X(_01228_));
 sg13g2_xnor2_1 _20417_ (.Y(_01229_),
    .A(_01178_),
    .B(_01173_));
 sg13g2_nand2b_1 _20418_ (.Y(_01231_),
    .B(_00569_),
    .A_N(_00560_));
 sg13g2_xnor2_1 _20419_ (.Y(_01232_),
    .A(_01231_),
    .B(_00568_));
 sg13g2_inv_1 _20420_ (.Y(_01233_),
    .A(_01232_));
 sg13g2_xnor2_1 _20421_ (.Y(_01234_),
    .A(_01233_),
    .B(_01229_));
 sg13g2_nand2_1 _20422_ (.Y(_01235_),
    .A(_01177_),
    .B(_01176_));
 sg13g2_nor2b_1 _20423_ (.A(_01178_),
    .B_N(_01235_),
    .Y(_01236_));
 sg13g2_nand2b_1 _20424_ (.Y(_01237_),
    .B(_00564_),
    .A_N(_00567_));
 sg13g2_xnor2_1 _20425_ (.Y(_01238_),
    .A(_00566_),
    .B(_01237_));
 sg13g2_nand2b_1 _20426_ (.Y(_01239_),
    .B(_01238_),
    .A_N(_01236_));
 sg13g2_and2_1 _20427_ (.A(_01234_),
    .B(_01239_),
    .X(_01240_));
 sg13g2_a21oi_1 _20428_ (.A1(_01229_),
    .A2(_01232_),
    .Y(_01242_),
    .B1(_01240_));
 sg13g2_nor2_1 _20429_ (.A(_00574_),
    .B(_00577_),
    .Y(_01243_));
 sg13g2_xor2_1 _20430_ (.B(_00571_),
    .A(_01243_),
    .X(_01244_));
 sg13g2_inv_1 _20431_ (.Y(_01245_),
    .A(_01244_));
 sg13g2_xor2_1 _20432_ (.B(_01181_),
    .A(_01180_),
    .X(_01246_));
 sg13g2_xnor2_1 _20433_ (.Y(_01247_),
    .A(_01245_),
    .B(_01246_));
 sg13g2_inv_1 _20434_ (.Y(_01248_),
    .A(_01247_));
 sg13g2_nand2b_1 _20435_ (.Y(_01249_),
    .B(_01245_),
    .A_N(_01246_));
 sg13g2_o21ai_1 _20436_ (.B1(_01249_),
    .Y(_01250_),
    .A1(_01242_),
    .A2(_01248_));
 sg13g2_nand2_1 _20437_ (.Y(_01251_),
    .A(_01228_),
    .B(_01250_));
 sg13g2_o21ai_1 _20438_ (.B1(_01251_),
    .Y(_01253_),
    .A1(_01226_),
    .A2(_01227_));
 sg13g2_nand2_1 _20439_ (.Y(_01254_),
    .A(_01225_),
    .B(_01253_));
 sg13g2_o21ai_1 _20440_ (.B1(_01254_),
    .Y(_01255_),
    .A1(_01221_),
    .A2(_01223_));
 sg13g2_nand2_1 _20441_ (.Y(_01256_),
    .A(_01220_),
    .B(_01255_));
 sg13g2_o21ai_1 _20442_ (.B1(_01256_),
    .Y(_01257_),
    .A1(_01215_),
    .A2(_01218_));
 sg13g2_nor2_1 _20443_ (.A(_01214_),
    .B(_01257_),
    .Y(_01258_));
 sg13g2_a21oi_1 _20444_ (.A1(_01212_),
    .A2(_01213_),
    .Y(_01259_),
    .B1(_01258_));
 sg13g2_nand2_1 _20445_ (.Y(_01260_),
    .A(_01204_),
    .B(_01259_));
 sg13g2_nand2b_1 _20446_ (.Y(_01261_),
    .B(_01260_),
    .A_N(_01200_));
 sg13g2_nor2_1 _20447_ (.A(net232),
    .B(_06275_),
    .Y(_01262_));
 sg13g2_inv_1 _20448_ (.Y(_01264_),
    .A(_01262_));
 sg13g2_xor2_1 _20449_ (.B(net222),
    .A(net203),
    .X(_01265_));
 sg13g2_xnor2_1 _20450_ (.Y(_01266_),
    .A(_01264_),
    .B(_01265_));
 sg13g2_nand3_1 _20451_ (.B(_00558_),
    .C(_00605_),
    .A(_01211_),
    .Y(_01267_));
 sg13g2_a21oi_1 _20452_ (.A1(_00604_),
    .A2(_00556_),
    .Y(_01268_),
    .B1(_00554_));
 sg13g2_nand2_1 _20453_ (.Y(_01269_),
    .A(_01267_),
    .B(_01268_));
 sg13g2_xor2_1 _20454_ (.B(_01269_),
    .A(_01266_),
    .X(_01270_));
 sg13g2_nand2b_1 _20455_ (.Y(_01271_),
    .B(_01106_),
    .A_N(_01144_));
 sg13g2_nor2_1 _20456_ (.A(_01109_),
    .B(_01142_),
    .Y(_01272_));
 sg13g2_inv_1 _20457_ (.Y(_01273_),
    .A(_01272_));
 sg13g2_nand2_1 _20458_ (.Y(_01275_),
    .A(_01271_),
    .B(_01273_));
 sg13g2_nor2b_1 _20459_ (.A(_01140_),
    .B_N(_01112_),
    .Y(_01276_));
 sg13g2_nand2b_1 _20460_ (.Y(_01277_),
    .B(_01111_),
    .A_N(_01141_));
 sg13g2_nor2b_1 _20461_ (.A(_01276_),
    .B_N(_01277_),
    .Y(_01278_));
 sg13g2_xnor2_1 _20462_ (.Y(_01279_),
    .A(net82),
    .B(_01115_));
 sg13g2_xnor2_1 _20463_ (.Y(_01280_),
    .A(net185),
    .B(_01045_));
 sg13g2_nand2b_1 _20464_ (.Y(_01281_),
    .B(net139),
    .A_N(_01129_));
 sg13g2_o21ai_1 _20465_ (.B1(_01281_),
    .Y(_01282_),
    .A1(net139),
    .A2(_01133_));
 sg13g2_inv_1 _20466_ (.Y(_01283_),
    .A(_01282_));
 sg13g2_o21ai_1 _20467_ (.B1(_01123_),
    .Y(_01284_),
    .A1(_01124_),
    .A2(_01131_));
 sg13g2_inv_1 _20468_ (.Y(_01286_),
    .A(_01284_));
 sg13g2_nor2_1 _20469_ (.A(_04602_),
    .B(_01120_),
    .Y(_01287_));
 sg13g2_inv_1 _20470_ (.Y(_01288_),
    .A(_01125_));
 sg13g2_a221oi_1 _20471_ (.B2(_01123_),
    .C1(_01287_),
    .B1(_01122_),
    .A1(_01085_),
    .Y(_01289_),
    .A2(_01082_));
 sg13g2_a22oi_1 _20472_ (.Y(_01290_),
    .B1(_01288_),
    .B2(_01289_),
    .A2(_01287_),
    .A1(_00106_));
 sg13g2_nor2_1 _20473_ (.A(net139),
    .B(_01290_),
    .Y(_01291_));
 sg13g2_a21oi_1 _20474_ (.A1(_01286_),
    .A2(net139),
    .Y(_01292_),
    .B1(_01291_));
 sg13g2_xnor2_1 _20475_ (.Y(_01293_),
    .A(net83),
    .B(_01292_));
 sg13g2_inv_1 _20476_ (.Y(_01294_),
    .A(_01293_));
 sg13g2_nor2_1 _20477_ (.A(_01283_),
    .B(_01294_),
    .Y(_01295_));
 sg13g2_nand2_1 _20478_ (.Y(_01297_),
    .A(_01294_),
    .B(_01283_));
 sg13g2_nand2b_1 _20479_ (.Y(_01298_),
    .B(_01297_),
    .A_N(_01295_));
 sg13g2_a21o_1 _20480_ (.A2(_01137_),
    .A1(_01113_),
    .B1(_01136_),
    .X(_01299_));
 sg13g2_xnor2_1 _20481_ (.Y(_01300_),
    .A(_01298_),
    .B(_01299_));
 sg13g2_xnor2_1 _20482_ (.Y(_01301_),
    .A(net71),
    .B(_01300_));
 sg13g2_xor2_1 _20483_ (.B(_01301_),
    .A(_01280_),
    .X(_01302_));
 sg13g2_xor2_1 _20484_ (.B(_01302_),
    .A(_01279_),
    .X(_01303_));
 sg13g2_or2_1 _20485_ (.X(_01304_),
    .B(_01303_),
    .A(_01278_));
 sg13g2_buf_1 _20486_ (.A(_01304_),
    .X(_01305_));
 sg13g2_nand2_1 _20487_ (.Y(_01306_),
    .A(_01303_),
    .B(_01278_));
 sg13g2_nand2_1 _20488_ (.Y(_01308_),
    .A(_01305_),
    .B(_01306_));
 sg13g2_xnor2_1 _20489_ (.Y(_01309_),
    .A(_01275_),
    .B(_01308_));
 sg13g2_inv_1 _20490_ (.Y(_01310_),
    .A(_01309_));
 sg13g2_nor2_1 _20491_ (.A(_01194_),
    .B(_01310_),
    .Y(_01311_));
 sg13g2_nand2_1 _20492_ (.Y(_01312_),
    .A(_01310_),
    .B(_01194_));
 sg13g2_nor2b_1 _20493_ (.A(_01311_),
    .B_N(_01312_),
    .Y(_01313_));
 sg13g2_a21o_1 _20494_ (.A2(_01148_),
    .A1(_01198_),
    .B1(_01147_),
    .X(_01314_));
 sg13g2_buf_1 _20495_ (.A(_01314_),
    .X(_01315_));
 sg13g2_xnor2_1 _20496_ (.Y(_01316_),
    .A(_01313_),
    .B(_01315_));
 sg13g2_nor2_1 _20497_ (.A(_01270_),
    .B(_01316_),
    .Y(_01317_));
 sg13g2_nand2_1 _20498_ (.Y(_01319_),
    .A(_01316_),
    .B(_01270_));
 sg13g2_nor2b_1 _20499_ (.A(_01317_),
    .B_N(_01319_),
    .Y(_01320_));
 sg13g2_xnor2_1 _20500_ (.Y(_01321_),
    .A(_01261_),
    .B(_01320_));
 sg13g2_inv_1 _20501_ (.Y(_01322_),
    .A(_01212_));
 sg13g2_xnor2_1 _20502_ (.Y(_01323_),
    .A(_01212_),
    .B(_01213_));
 sg13g2_inv_1 _20503_ (.Y(_01324_),
    .A(_01225_));
 sg13g2_nand2_1 _20504_ (.Y(_01325_),
    .A(_01236_),
    .B(_01238_));
 sg13g2_nor2_1 _20505_ (.A(_01325_),
    .B(_01234_),
    .Y(_01326_));
 sg13g2_a21oi_1 _20506_ (.A1(_01229_),
    .A2(_01233_),
    .Y(_01327_),
    .B1(_01326_));
 sg13g2_inv_1 _20507_ (.Y(_01328_),
    .A(_01327_));
 sg13g2_nor2_1 _20508_ (.A(_01245_),
    .B(_01246_),
    .Y(_01330_));
 sg13g2_a21oi_1 _20509_ (.A1(_01248_),
    .A2(_01328_),
    .Y(_01331_),
    .B1(_01330_));
 sg13g2_nand2b_1 _20510_ (.Y(_01332_),
    .B(_01226_),
    .A_N(_01227_));
 sg13g2_o21ai_1 _20511_ (.B1(_01332_),
    .Y(_01333_),
    .A1(_01331_),
    .A2(_01228_));
 sg13g2_nor2_1 _20512_ (.A(_01224_),
    .B(_01223_),
    .Y(_01334_));
 sg13g2_a21oi_1 _20513_ (.A1(_01324_),
    .A2(_01333_),
    .Y(_01335_),
    .B1(_01334_));
 sg13g2_nand2b_1 _20514_ (.Y(_01336_),
    .B(_01215_),
    .A_N(_01218_));
 sg13g2_o21ai_1 _20515_ (.B1(_01336_),
    .Y(_01337_),
    .A1(_01335_),
    .A2(_01220_));
 sg13g2_nand2_1 _20516_ (.Y(_01338_),
    .A(_01323_),
    .B(_01337_));
 sg13g2_o21ai_1 _20517_ (.B1(_01338_),
    .Y(_01339_),
    .A1(_01322_),
    .A2(_01213_));
 sg13g2_a21o_1 _20518_ (.A2(_01203_),
    .A1(_01339_),
    .B1(_01202_),
    .X(_01341_));
 sg13g2_xor2_1 _20519_ (.B(_01320_),
    .A(_01341_),
    .X(_01342_));
 sg13g2_buf_1 _20520_ (.A(net46),
    .X(_01343_));
 sg13g2_mux2_1 _20521_ (.A0(_01321_),
    .A1(_01342_),
    .S(net44),
    .X(_01344_));
 sg13g2_xnor2_1 _20522_ (.Y(_01345_),
    .A(net51),
    .B(_01344_));
 sg13g2_xnor2_1 _20523_ (.Y(_01346_),
    .A(net202),
    .B(net221));
 sg13g2_nor3_1 _20524_ (.A(net203),
    .B(net222),
    .C(_01346_),
    .Y(_01347_));
 sg13g2_inv_1 _20525_ (.Y(_01348_),
    .A(_01347_));
 sg13g2_o21ai_1 _20526_ (.B1(_01346_),
    .Y(_01349_),
    .A1(net203),
    .A2(net222));
 sg13g2_nand2_1 _20527_ (.Y(_01350_),
    .A(_01348_),
    .B(_01349_));
 sg13g2_inv_1 _20528_ (.Y(_01352_),
    .A(_01350_));
 sg13g2_inv_1 _20529_ (.Y(_01353_),
    .A(_00609_));
 sg13g2_nand2_1 _20530_ (.Y(_01354_),
    .A(_00558_),
    .B(_01266_));
 sg13g2_inv_1 _20531_ (.Y(_01355_),
    .A(_01354_));
 sg13g2_inv_1 _20532_ (.Y(_01356_),
    .A(_01265_));
 sg13g2_a21oi_1 _20533_ (.A1(_00555_),
    .A2(_01264_),
    .Y(_01357_),
    .B1(_01356_));
 sg13g2_a21oi_1 _20534_ (.A1(_01353_),
    .A2(_01355_),
    .Y(_01358_),
    .B1(_01357_));
 sg13g2_xnor2_1 _20535_ (.Y(_01359_),
    .A(_01352_),
    .B(_01358_));
 sg13g2_nor2b_1 _20536_ (.A(_01301_),
    .B_N(_01280_),
    .Y(_01360_));
 sg13g2_nor2b_1 _20537_ (.A(_01302_),
    .B_N(_01279_),
    .Y(_01361_));
 sg13g2_nor2_1 _20538_ (.A(_01360_),
    .B(_01361_),
    .Y(_01362_));
 sg13g2_xnor2_1 _20539_ (.Y(_01363_),
    .A(net82),
    .B(_01282_));
 sg13g2_xnor2_1 _20540_ (.Y(_01364_),
    .A(net178),
    .B(_01093_));
 sg13g2_nor2_1 _20541_ (.A(net139),
    .B(_01286_),
    .Y(_01365_));
 sg13g2_a21oi_2 _20542_ (.B1(_01365_),
    .Y(_01366_),
    .A2(_01290_),
    .A1(net139));
 sg13g2_xnor2_1 _20543_ (.Y(_01367_),
    .A(_01366_),
    .B(_01293_));
 sg13g2_xnor2_1 _20544_ (.Y(_01368_),
    .A(net70),
    .B(_01367_));
 sg13g2_a21o_1 _20545_ (.A2(_01297_),
    .A1(_01299_),
    .B1(_01295_),
    .X(_01369_));
 sg13g2_xnor2_1 _20546_ (.Y(_01370_),
    .A(_01368_),
    .B(_01369_));
 sg13g2_xor2_1 _20547_ (.B(_01370_),
    .A(_01364_),
    .X(_01371_));
 sg13g2_xor2_1 _20548_ (.B(_01371_),
    .A(_01363_),
    .X(_01373_));
 sg13g2_nor2_1 _20549_ (.A(_01362_),
    .B(_01373_),
    .Y(_01374_));
 sg13g2_inv_1 _20550_ (.Y(_01375_),
    .A(_01374_));
 sg13g2_nand2_1 _20551_ (.Y(_01376_),
    .A(_01373_),
    .B(_01362_));
 sg13g2_nand2_1 _20552_ (.Y(_01377_),
    .A(_01375_),
    .B(_01376_));
 sg13g2_inv_1 _20553_ (.Y(_01378_),
    .A(_01306_));
 sg13g2_inv_1 _20554_ (.Y(_01379_),
    .A(_01275_));
 sg13g2_o21ai_1 _20555_ (.B1(_01305_),
    .Y(_01380_),
    .A1(_01378_),
    .A2(_01379_));
 sg13g2_xor2_1 _20556_ (.B(_01380_),
    .A(_01377_),
    .X(_01381_));
 sg13g2_buf_1 _20557_ (.A(_01381_),
    .X(_01382_));
 sg13g2_xor2_1 _20558_ (.B(_01382_),
    .A(_01146_),
    .X(_01384_));
 sg13g2_a21oi_1 _20559_ (.A1(_01315_),
    .A2(_01312_),
    .Y(_01385_),
    .B1(_01311_));
 sg13g2_xor2_1 _20560_ (.B(_01385_),
    .A(_01384_),
    .X(_01386_));
 sg13g2_nor2_1 _20561_ (.A(_01359_),
    .B(_01386_),
    .Y(_01387_));
 sg13g2_nand2_1 _20562_ (.Y(_01388_),
    .A(_01386_),
    .B(_01359_));
 sg13g2_nand2b_1 _20563_ (.Y(_01389_),
    .B(_01388_),
    .A_N(_01387_));
 sg13g2_inv_1 _20564_ (.Y(_01390_),
    .A(_01270_));
 sg13g2_inv_1 _20565_ (.Y(_01391_),
    .A(_01320_));
 sg13g2_nand2_1 _20566_ (.Y(_01392_),
    .A(_01391_),
    .B(_01341_));
 sg13g2_o21ai_1 _20567_ (.B1(_01392_),
    .Y(_01393_),
    .A1(_01390_),
    .A2(_01316_));
 sg13g2_xnor2_1 _20568_ (.Y(_01395_),
    .A(_01389_),
    .B(_01393_));
 sg13g2_a21o_1 _20569_ (.A2(_01319_),
    .A1(_01261_),
    .B1(_01317_),
    .X(_01396_));
 sg13g2_xor2_1 _20570_ (.B(_01389_),
    .A(_01396_),
    .X(_01397_));
 sg13g2_nor2b_1 _20571_ (.A(net43),
    .B_N(_01397_),
    .Y(_01398_));
 sg13g2_a21oi_1 _20572_ (.A1(net43),
    .A2(_01395_),
    .Y(_01399_),
    .B1(_01398_));
 sg13g2_xnor2_1 _20573_ (.Y(_01400_),
    .A(net38),
    .B(_01399_));
 sg13g2_nand2b_1 _20574_ (.Y(_01401_),
    .B(_01400_),
    .A_N(_01345_));
 sg13g2_xnor2_1 _20575_ (.Y(_01402_),
    .A(_01323_),
    .B(_01257_));
 sg13g2_xnor2_1 _20576_ (.Y(_01403_),
    .A(_01337_),
    .B(_01323_));
 sg13g2_nand2_1 _20577_ (.Y(_01404_),
    .A(_01403_),
    .B(_01343_));
 sg13g2_o21ai_1 _20578_ (.B1(_01404_),
    .Y(_01406_),
    .A1(net44),
    .A2(_01402_));
 sg13g2_xnor2_1 _20579_ (.Y(_01407_),
    .A(net51),
    .B(_01406_));
 sg13g2_buf_8 _20580_ (.A(net40),
    .X(_01408_));
 sg13g2_xnor2_1 _20581_ (.Y(_01409_),
    .A(_01259_),
    .B(_01204_));
 sg13g2_xor2_1 _20582_ (.B(_01204_),
    .A(_01339_),
    .X(_01410_));
 sg13g2_mux2_1 _20583_ (.A0(_01409_),
    .A1(_01410_),
    .S(net43),
    .X(_01411_));
 sg13g2_xnor2_1 _20584_ (.Y(_01412_),
    .A(net39),
    .B(_01411_));
 sg13g2_nor2b_1 _20585_ (.A(_01407_),
    .B_N(_01412_),
    .Y(_01413_));
 sg13g2_xnor2_1 _20586_ (.Y(_01414_),
    .A(_01335_),
    .B(_01220_));
 sg13g2_xnor2_1 _20587_ (.Y(_01415_),
    .A(_01255_),
    .B(_01220_));
 sg13g2_mux2_1 _20588_ (.A0(_01414_),
    .A1(_01415_),
    .S(net45),
    .X(_01417_));
 sg13g2_xnor2_1 _20589_ (.Y(_01418_),
    .A(net51),
    .B(_01417_));
 sg13g2_nand2_1 _20590_ (.Y(_01419_),
    .A(_01403_),
    .B(net45));
 sg13g2_o21ai_1 _20591_ (.B1(_01419_),
    .Y(_01420_),
    .A1(net43),
    .A2(_01402_));
 sg13g2_xnor2_1 _20592_ (.Y(_01421_),
    .A(net39),
    .B(_01420_));
 sg13g2_xor2_1 _20593_ (.B(_01421_),
    .A(_01418_),
    .X(_01422_));
 sg13g2_xnor2_1 _20594_ (.Y(_01423_),
    .A(_01250_),
    .B(_01228_));
 sg13g2_xnor2_1 _20595_ (.Y(_01424_),
    .A(_01331_),
    .B(_01228_));
 sg13g2_mux2_1 _20596_ (.A0(_01423_),
    .A1(_01424_),
    .S(net46),
    .X(_01425_));
 sg13g2_xnor2_1 _20597_ (.Y(_01426_),
    .A(net52),
    .B(_01425_));
 sg13g2_xnor2_1 _20598_ (.Y(_01428_),
    .A(_01253_),
    .B(_01225_));
 sg13g2_xor2_1 _20599_ (.B(_01225_),
    .A(_01333_),
    .X(_01429_));
 sg13g2_mux2_1 _20600_ (.A0(_01428_),
    .A1(_01429_),
    .S(net45),
    .X(_01430_));
 sg13g2_xnor2_1 _20601_ (.Y(_01431_),
    .A(net39),
    .B(_01430_));
 sg13g2_xnor2_1 _20602_ (.Y(_01432_),
    .A(_01426_),
    .B(_01431_));
 sg13g2_xor2_1 _20603_ (.B(_01242_),
    .A(_01247_),
    .X(_01433_));
 sg13g2_xor2_1 _20604_ (.B(_01247_),
    .A(_01327_),
    .X(_01434_));
 sg13g2_nor2_1 _20605_ (.A(net45),
    .B(_01434_),
    .Y(_01435_));
 sg13g2_a21oi_1 _20606_ (.A1(net45),
    .A2(_01433_),
    .Y(_01436_),
    .B1(_01435_));
 sg13g2_xnor2_1 _20607_ (.Y(_01437_),
    .A(net53),
    .B(_01436_));
 sg13g2_mux2_1 _20608_ (.A0(_01423_),
    .A1(_01424_),
    .S(net45),
    .X(_01439_));
 sg13g2_xnor2_1 _20609_ (.Y(_01440_),
    .A(net39),
    .B(_01439_));
 sg13g2_nor2b_1 _20610_ (.A(_01437_),
    .B_N(_01440_),
    .Y(_01441_));
 sg13g2_xor2_1 _20611_ (.B(_01234_),
    .A(_01325_),
    .X(_01442_));
 sg13g2_xnor2_1 _20612_ (.Y(_01443_),
    .A(_01239_),
    .B(_01234_));
 sg13g2_nand2_1 _20613_ (.Y(_01444_),
    .A(_01443_),
    .B(net45));
 sg13g2_o21ai_1 _20614_ (.B1(_01444_),
    .Y(_01445_),
    .A1(net45),
    .A2(_01442_));
 sg13g2_xnor2_1 _20615_ (.Y(_01446_),
    .A(net52),
    .B(_01445_));
 sg13g2_nor2_1 _20616_ (.A(net46),
    .B(_01434_),
    .Y(_01447_));
 sg13g2_a21oi_1 _20617_ (.A1(net46),
    .A2(_01433_),
    .Y(_01448_),
    .B1(_01447_));
 sg13g2_xor2_1 _20618_ (.B(_01448_),
    .A(_01408_),
    .X(_01450_));
 sg13g2_nor2b_1 _20619_ (.A(_01446_),
    .B_N(_01450_),
    .Y(_01451_));
 sg13g2_nor2_1 _20620_ (.A(net46),
    .B(_01442_),
    .Y(_01452_));
 sg13g2_a21oi_1 _20621_ (.A1(net46),
    .A2(_01443_),
    .Y(_01453_),
    .B1(_01452_));
 sg13g2_nand2b_1 _20622_ (.Y(_01454_),
    .B(net38),
    .A_N(_01453_));
 sg13g2_nand2_1 _20623_ (.Y(_01455_),
    .A(_01408_),
    .B(_01453_));
 sg13g2_xnor2_1 _20624_ (.Y(_01456_),
    .A(_01238_),
    .B(_01236_));
 sg13g2_xnor2_1 _20625_ (.Y(_01457_),
    .A(_01456_),
    .B(net53));
 sg13g2_nand3_1 _20626_ (.B(_01455_),
    .C(_01457_),
    .A(_01454_),
    .Y(_01458_));
 sg13g2_xor2_1 _20627_ (.B(_01450_),
    .A(_01446_),
    .X(_01459_));
 sg13g2_nor2_1 _20628_ (.A(_01458_),
    .B(_01459_),
    .Y(_01461_));
 sg13g2_nor2_1 _20629_ (.A(_01451_),
    .B(_01461_),
    .Y(_01462_));
 sg13g2_xnor2_1 _20630_ (.Y(_01463_),
    .A(_01437_),
    .B(_01440_));
 sg13g2_nor2b_1 _20631_ (.A(_01462_),
    .B_N(_01463_),
    .Y(_01464_));
 sg13g2_nor2_1 _20632_ (.A(_01441_),
    .B(_01464_),
    .Y(_01465_));
 sg13g2_inv_1 _20633_ (.Y(_01466_),
    .A(_01465_));
 sg13g2_nor2b_1 _20634_ (.A(_01426_),
    .B_N(_01431_),
    .Y(_01467_));
 sg13g2_a21oi_1 _20635_ (.A1(_01432_),
    .A2(_01466_),
    .Y(_01468_),
    .B1(_01467_));
 sg13g2_mux2_1 _20636_ (.A0(_01428_),
    .A1(_01429_),
    .S(net44),
    .X(_01469_));
 sg13g2_xnor2_1 _20637_ (.Y(_01470_),
    .A(net52),
    .B(_01469_));
 sg13g2_mux2_1 _20638_ (.A0(_01414_),
    .A1(_01415_),
    .S(_01343_),
    .X(_01472_));
 sg13g2_xnor2_1 _20639_ (.Y(_01473_),
    .A(net39),
    .B(_01472_));
 sg13g2_xnor2_1 _20640_ (.Y(_01474_),
    .A(_01470_),
    .B(_01473_));
 sg13g2_nand2b_1 _20641_ (.Y(_01475_),
    .B(_01474_),
    .A_N(_01468_));
 sg13g2_nand2b_1 _20642_ (.Y(_01476_),
    .B(_01473_),
    .A_N(_01470_));
 sg13g2_nand2_1 _20643_ (.Y(_01477_),
    .A(_01475_),
    .B(_01476_));
 sg13g2_nand2b_1 _20644_ (.Y(_01478_),
    .B(_01477_),
    .A_N(_01422_));
 sg13g2_nand2b_1 _20645_ (.Y(_01479_),
    .B(_01421_),
    .A_N(_01418_));
 sg13g2_nand2_1 _20646_ (.Y(_01480_),
    .A(_01478_),
    .B(_01479_));
 sg13g2_nand2b_1 _20647_ (.Y(_01481_),
    .B(_01407_),
    .A_N(_01412_));
 sg13g2_o21ai_1 _20648_ (.B1(_01481_),
    .Y(_01482_),
    .A1(_01413_),
    .A2(_01480_));
 sg13g2_mux2_1 _20649_ (.A0(_01409_),
    .A1(_01410_),
    .S(net44),
    .X(_01483_));
 sg13g2_xnor2_1 _20650_ (.Y(_01484_),
    .A(net51),
    .B(_01483_));
 sg13g2_mux2_1 _20651_ (.A0(_01321_),
    .A1(_01342_),
    .S(net43),
    .X(_01485_));
 sg13g2_xnor2_1 _20652_ (.Y(_01486_),
    .A(net39),
    .B(_01485_));
 sg13g2_xnor2_1 _20653_ (.Y(_01487_),
    .A(_01484_),
    .B(_01486_));
 sg13g2_nand2b_1 _20654_ (.Y(_01488_),
    .B(_01487_),
    .A_N(_01482_));
 sg13g2_nand2b_1 _20655_ (.Y(_01489_),
    .B(_01486_),
    .A_N(_01484_));
 sg13g2_nand3_1 _20656_ (.B(_01488_),
    .C(_01489_),
    .A(_01401_),
    .Y(_01490_));
 sg13g2_nand2b_1 _20657_ (.Y(_01491_),
    .B(_01345_),
    .A_N(_01400_));
 sg13g2_nand2_1 _20658_ (.Y(_01493_),
    .A(_01490_),
    .B(_01491_));
 sg13g2_buf_1 _20659_ (.A(net44),
    .X(_01494_));
 sg13g2_nor2b_1 _20660_ (.A(net44),
    .B_N(_01397_),
    .Y(_01495_));
 sg13g2_a21oi_1 _20661_ (.A1(net42),
    .A2(_01395_),
    .Y(_01496_),
    .B1(_01495_));
 sg13g2_xnor2_1 _20662_ (.Y(_01497_),
    .A(net53),
    .B(_01496_));
 sg13g2_nor2_1 _20663_ (.A(net202),
    .B(net221),
    .Y(_01498_));
 sg13g2_inv_1 _20664_ (.Y(_01499_),
    .A(_01498_));
 sg13g2_xor2_1 _20665_ (.B(net224),
    .A(net201),
    .X(_01500_));
 sg13g2_xnor2_1 _20666_ (.Y(_01501_),
    .A(_01499_),
    .B(_01500_));
 sg13g2_nand3_1 _20667_ (.B(_01352_),
    .C(_01266_),
    .A(_01269_),
    .Y(_01502_));
 sg13g2_nand3_1 _20668_ (.B(_01265_),
    .C(_01262_),
    .A(_01352_),
    .Y(_01504_));
 sg13g2_nand3_1 _20669_ (.B(_01348_),
    .C(_01504_),
    .A(_01502_),
    .Y(_01505_));
 sg13g2_xor2_1 _20670_ (.B(_01505_),
    .A(_01501_),
    .X(_01506_));
 sg13g2_inv_1 _20671_ (.Y(_01507_),
    .A(_01506_));
 sg13g2_nor2b_1 _20672_ (.A(_01364_),
    .B_N(_01370_),
    .Y(_01508_));
 sg13g2_nor2b_1 _20673_ (.A(_01371_),
    .B_N(_01363_),
    .Y(_01509_));
 sg13g2_nor2_1 _20674_ (.A(_01508_),
    .B(_01509_),
    .Y(_01510_));
 sg13g2_xnor2_1 _20675_ (.Y(_01511_),
    .A(net82),
    .B(_01366_));
 sg13g2_buf_1 _20676_ (.A(_01511_),
    .X(_01512_));
 sg13g2_xnor2_1 _20677_ (.Y(_01513_),
    .A(net178),
    .B(_01134_));
 sg13g2_nand2b_1 _20678_ (.Y(_01515_),
    .B(_01369_),
    .A_N(_01367_));
 sg13g2_o21ai_1 _20679_ (.B1(_01515_),
    .Y(_01516_),
    .A1(_01293_),
    .A2(_01366_));
 sg13g2_xnor2_1 _20680_ (.Y(_01517_),
    .A(net70),
    .B(_01516_));
 sg13g2_buf_1 _20681_ (.A(_01517_),
    .X(_01518_));
 sg13g2_xnor2_1 _20682_ (.Y(_01519_),
    .A(_01513_),
    .B(_01518_));
 sg13g2_xor2_1 _20683_ (.B(_01519_),
    .A(_01512_),
    .X(_01520_));
 sg13g2_or2_1 _20684_ (.X(_01521_),
    .B(_01520_),
    .A(_01510_));
 sg13g2_buf_1 _20685_ (.A(_01521_),
    .X(_01522_));
 sg13g2_nand2_1 _20686_ (.Y(_01523_),
    .A(_01520_),
    .B(_01510_));
 sg13g2_nand2_1 _20687_ (.Y(_01524_),
    .A(_01522_),
    .B(_01523_));
 sg13g2_nand2_1 _20688_ (.Y(_01525_),
    .A(_01375_),
    .B(_01305_));
 sg13g2_nor2_1 _20689_ (.A(_01308_),
    .B(_01379_),
    .Y(_01526_));
 sg13g2_o21ai_1 _20690_ (.B1(_01376_),
    .Y(_01527_),
    .A1(_01525_),
    .A2(_01526_));
 sg13g2_xor2_1 _20691_ (.B(_01527_),
    .A(_01524_),
    .X(_01528_));
 sg13g2_nor2_1 _20692_ (.A(_01309_),
    .B(_01528_),
    .Y(_01529_));
 sg13g2_nor2b_1 _20693_ (.A(_01310_),
    .B_N(_01528_),
    .Y(_01530_));
 sg13g2_nor2_1 _20694_ (.A(_01529_),
    .B(_01530_),
    .Y(_01531_));
 sg13g2_nor2_1 _20695_ (.A(_01146_),
    .B(_01382_),
    .Y(_01532_));
 sg13g2_nor2_1 _20696_ (.A(_01311_),
    .B(_01532_),
    .Y(_01533_));
 sg13g2_nand2_1 _20697_ (.Y(_01534_),
    .A(_01315_),
    .B(_01313_));
 sg13g2_a22oi_1 _20698_ (.Y(_01536_),
    .B1(_01533_),
    .B2(_01534_),
    .A2(_01146_),
    .A1(_01382_));
 sg13g2_xnor2_1 _20699_ (.Y(_01537_),
    .A(_01531_),
    .B(_01536_));
 sg13g2_nor2_1 _20700_ (.A(_01507_),
    .B(_01537_),
    .Y(_01538_));
 sg13g2_nand2_1 _20701_ (.Y(_01539_),
    .A(_01537_),
    .B(_01507_));
 sg13g2_nor2b_1 _20702_ (.A(_01538_),
    .B_N(_01539_),
    .Y(_01540_));
 sg13g2_inv_1 _20703_ (.Y(_01541_),
    .A(_01540_));
 sg13g2_a21o_1 _20704_ (.A2(_01388_),
    .A1(_01396_),
    .B1(_01387_),
    .X(_01542_));
 sg13g2_xnor2_1 _20705_ (.Y(_01543_),
    .A(_01541_),
    .B(_01542_));
 sg13g2_nor2b_1 _20706_ (.A(_01386_),
    .B_N(_01359_),
    .Y(_01544_));
 sg13g2_nand2_1 _20707_ (.Y(_01545_),
    .A(_01393_),
    .B(_01389_));
 sg13g2_nand2b_1 _20708_ (.Y(_01547_),
    .B(_01545_),
    .A_N(_01544_));
 sg13g2_xnor2_1 _20709_ (.Y(_01548_),
    .A(_01540_),
    .B(_01547_));
 sg13g2_mux2_1 _20710_ (.A0(_01543_),
    .A1(_01548_),
    .S(net43),
    .X(_01549_));
 sg13g2_xnor2_1 _20711_ (.Y(_01550_),
    .A(net39),
    .B(_01549_));
 sg13g2_nor2b_1 _20712_ (.A(_01497_),
    .B_N(_01550_),
    .Y(_01551_));
 sg13g2_nand2b_1 _20713_ (.Y(_01552_),
    .B(_01497_),
    .A_N(_01550_));
 sg13g2_nor2b_1 _20714_ (.A(_01551_),
    .B_N(_01552_),
    .Y(_01553_));
 sg13g2_xnor2_1 _20715_ (.Y(_01554_),
    .A(_01493_),
    .B(_01553_));
 sg13g2_inv_1 _20716_ (.Y(_01555_),
    .A(_01554_));
 sg13g2_nor2_1 _20717_ (.A(net201),
    .B(net224),
    .Y(_01556_));
 sg13g2_inv_1 _20718_ (.Y(_01558_),
    .A(_01556_));
 sg13g2_xor2_1 _20719_ (.B(net226),
    .A(net200),
    .X(_01559_));
 sg13g2_xnor2_1 _20720_ (.Y(_01560_),
    .A(_01558_),
    .B(_01559_));
 sg13g2_inv_1 _20721_ (.Y(_01561_),
    .A(_01500_));
 sg13g2_a21oi_1 _20722_ (.A1(_01348_),
    .A2(_01499_),
    .Y(_01562_),
    .B1(_01561_));
 sg13g2_nand2_1 _20723_ (.Y(_01563_),
    .A(_01352_),
    .B(_01501_));
 sg13g2_nor2_1 _20724_ (.A(_01563_),
    .B(_01358_),
    .Y(_01564_));
 sg13g2_nor2_1 _20725_ (.A(_01562_),
    .B(_01564_),
    .Y(_01565_));
 sg13g2_xnor2_1 _20726_ (.Y(_01566_),
    .A(_01560_),
    .B(_01565_));
 sg13g2_inv_1 _20727_ (.Y(_01567_),
    .A(_01566_));
 sg13g2_nand2_1 _20728_ (.Y(_01568_),
    .A(_01518_),
    .B(_01513_));
 sg13g2_nor2_1 _20729_ (.A(_01513_),
    .B(_01518_),
    .Y(_01569_));
 sg13g2_a21oi_1 _20730_ (.A1(_01568_),
    .A2(_01512_),
    .Y(_01570_),
    .B1(_01569_));
 sg13g2_xnor2_1 _20731_ (.Y(_01571_),
    .A(net185),
    .B(_01292_));
 sg13g2_inv_1 _20732_ (.Y(_01572_),
    .A(_01571_));
 sg13g2_nor2_1 _20733_ (.A(_01572_),
    .B(_01518_),
    .Y(_01573_));
 sg13g2_nand2_1 _20734_ (.Y(_01574_),
    .A(_01518_),
    .B(_01572_));
 sg13g2_nor2b_1 _20735_ (.A(_01573_),
    .B_N(_01574_),
    .Y(_01575_));
 sg13g2_xnor2_1 _20736_ (.Y(_01576_),
    .A(_01512_),
    .B(_01575_));
 sg13g2_or2_1 _20737_ (.X(_01577_),
    .B(_01576_),
    .A(_01570_));
 sg13g2_nand2_1 _20738_ (.Y(_01579_),
    .A(_01576_),
    .B(_01570_));
 sg13g2_nand2_1 _20739_ (.Y(_01580_),
    .A(_01577_),
    .B(_01579_));
 sg13g2_nand2_1 _20740_ (.Y(_01581_),
    .A(_01522_),
    .B(_01375_));
 sg13g2_nor2b_1 _20741_ (.A(_01377_),
    .B_N(_01380_),
    .Y(_01582_));
 sg13g2_o21ai_1 _20742_ (.B1(_01523_),
    .Y(_01583_),
    .A1(_01581_),
    .A2(_01582_));
 sg13g2_xnor2_1 _20743_ (.Y(_01584_),
    .A(_01580_),
    .B(_01583_));
 sg13g2_nor2_1 _20744_ (.A(_01382_),
    .B(_01584_),
    .Y(_01585_));
 sg13g2_nand2_1 _20745_ (.Y(_01586_),
    .A(_01584_),
    .B(_01382_));
 sg13g2_inv_1 _20746_ (.Y(_01587_),
    .A(_01586_));
 sg13g2_nor2_1 _20747_ (.A(_01585_),
    .B(_01587_),
    .Y(_01588_));
 sg13g2_nand2b_1 _20748_ (.Y(_01590_),
    .B(_01384_),
    .A_N(_01385_));
 sg13g2_nor2_1 _20749_ (.A(_01532_),
    .B(_01530_),
    .Y(_01591_));
 sg13g2_a21oi_1 _20750_ (.A1(_01590_),
    .A2(_01591_),
    .Y(_01592_),
    .B1(_01529_));
 sg13g2_xnor2_1 _20751_ (.Y(_01593_),
    .A(_01588_),
    .B(_01592_));
 sg13g2_nor2_1 _20752_ (.A(_01567_),
    .B(_01593_),
    .Y(_01594_));
 sg13g2_nand2_1 _20753_ (.Y(_01595_),
    .A(_01593_),
    .B(_01567_));
 sg13g2_nor2b_1 _20754_ (.A(_01594_),
    .B_N(_01595_),
    .Y(_01596_));
 sg13g2_buf_1 _20755_ (.A(_01596_),
    .X(_01597_));
 sg13g2_inv_1 _20756_ (.Y(_01598_),
    .A(_01597_));
 sg13g2_nand2_1 _20757_ (.Y(_01599_),
    .A(_01542_),
    .B(_01541_));
 sg13g2_o21ai_1 _20758_ (.B1(_01599_),
    .Y(_01601_),
    .A1(_01537_),
    .A2(_01506_));
 sg13g2_xnor2_1 _20759_ (.Y(_01602_),
    .A(_01598_),
    .B(_01601_));
 sg13g2_buf_1 _20760_ (.A(net43),
    .X(_01603_));
 sg13g2_o21ai_1 _20761_ (.B1(_01539_),
    .Y(_01604_),
    .A1(_01544_),
    .A2(_01538_));
 sg13g2_o21ai_1 _20762_ (.B1(_01604_),
    .Y(_01605_),
    .A1(_01541_),
    .A2(_01545_));
 sg13g2_xnor2_1 _20763_ (.Y(_01606_),
    .A(_01597_),
    .B(_01605_));
 sg13g2_nor2b_1 _20764_ (.A(net41),
    .B_N(_01606_),
    .Y(_01607_));
 sg13g2_a21oi_1 _20765_ (.A1(_01602_),
    .A2(net41),
    .Y(_01608_),
    .B1(_01607_));
 sg13g2_xnor2_1 _20766_ (.Y(_01609_),
    .A(net53),
    .B(_01608_));
 sg13g2_nor2_1 _20767_ (.A(net200),
    .B(net226),
    .Y(_01610_));
 sg13g2_xor2_1 _20768_ (.B(_06236_),
    .A(_05772_),
    .X(_01612_));
 sg13g2_xor2_1 _20769_ (.B(_01612_),
    .A(_01610_),
    .X(_01613_));
 sg13g2_nand3_1 _20770_ (.B(_01560_),
    .C(_01501_),
    .A(_01505_),
    .Y(_01614_));
 sg13g2_nor2_1 _20771_ (.A(_01499_),
    .B(_01561_),
    .Y(_01615_));
 sg13g2_nor2b_1 _20772_ (.A(_01558_),
    .B_N(_01559_),
    .Y(_01616_));
 sg13g2_a21oi_1 _20773_ (.A1(_01615_),
    .A2(_01559_),
    .Y(_01617_),
    .B1(_01616_));
 sg13g2_nand2_1 _20774_ (.Y(_01618_),
    .A(_01614_),
    .B(_01617_));
 sg13g2_xnor2_1 _20775_ (.Y(_01619_),
    .A(_01613_),
    .B(_01618_));
 sg13g2_inv_1 _20776_ (.Y(_01620_),
    .A(_01619_));
 sg13g2_nor2_1 _20777_ (.A(_01512_),
    .B(_01574_),
    .Y(_01621_));
 sg13g2_nand2_1 _20778_ (.Y(_01623_),
    .A(_01577_),
    .B(_01522_));
 sg13g2_nor2_1 _20779_ (.A(_01524_),
    .B(_01527_),
    .Y(_01624_));
 sg13g2_nor2_1 _20780_ (.A(_01623_),
    .B(_01624_),
    .Y(_01625_));
 sg13g2_nor2b_1 _20781_ (.A(_01625_),
    .B_N(_01579_),
    .Y(_01626_));
 sg13g2_nand2_1 _20782_ (.Y(_01627_),
    .A(_01573_),
    .B(_01512_));
 sg13g2_o21ai_1 _20783_ (.B1(_01627_),
    .Y(_01628_),
    .A1(_01621_),
    .A2(_01626_));
 sg13g2_buf_2 _20784_ (.A(_01628_),
    .X(_01629_));
 sg13g2_nor2_1 _20785_ (.A(_01528_),
    .B(_01629_),
    .Y(_01630_));
 sg13g2_nand2_1 _20786_ (.Y(_01631_),
    .A(_01629_),
    .B(_01528_));
 sg13g2_inv_1 _20787_ (.Y(_01632_),
    .A(_01631_));
 sg13g2_nor2_1 _20788_ (.A(_01630_),
    .B(_01632_),
    .Y(_01634_));
 sg13g2_nor2_1 _20789_ (.A(_01530_),
    .B(_01585_),
    .Y(_01635_));
 sg13g2_nand2_1 _20790_ (.Y(_01636_),
    .A(_01536_),
    .B(_01531_));
 sg13g2_a21oi_1 _20791_ (.A1(_01635_),
    .A2(_01636_),
    .Y(_01637_),
    .B1(_01587_));
 sg13g2_xor2_1 _20792_ (.B(_01637_),
    .A(_01634_),
    .X(_01638_));
 sg13g2_nor2_1 _20793_ (.A(_01620_),
    .B(_01638_),
    .Y(_01639_));
 sg13g2_nand2_1 _20794_ (.Y(_01640_),
    .A(_01638_),
    .B(_01620_));
 sg13g2_inv_1 _20795_ (.Y(_01641_),
    .A(_01640_));
 sg13g2_nor2_2 _20796_ (.A(_01639_),
    .B(_01641_),
    .Y(_01642_));
 sg13g2_inv_1 _20797_ (.Y(_01643_),
    .A(_01642_));
 sg13g2_nand2_1 _20798_ (.Y(_01645_),
    .A(_01601_),
    .B(_01598_));
 sg13g2_o21ai_1 _20799_ (.B1(_01645_),
    .Y(_01646_),
    .A1(_01593_),
    .A2(_01566_));
 sg13g2_xnor2_1 _20800_ (.Y(_01647_),
    .A(_01643_),
    .B(_01646_));
 sg13g2_nand3_1 _20801_ (.B(_01540_),
    .C(_01547_),
    .A(_01597_),
    .Y(_01648_));
 sg13g2_o21ai_1 _20802_ (.B1(_01595_),
    .Y(_01649_),
    .A1(_01538_),
    .A2(_01594_));
 sg13g2_nand2_1 _20803_ (.Y(_01650_),
    .A(_01648_),
    .B(_01649_));
 sg13g2_xnor2_1 _20804_ (.Y(_01651_),
    .A(_01642_),
    .B(_01650_));
 sg13g2_nor2b_1 _20805_ (.A(net44),
    .B_N(_01651_),
    .Y(_01652_));
 sg13g2_a21oi_1 _20806_ (.A1(_01647_),
    .A2(net42),
    .Y(_01653_),
    .B1(_01652_));
 sg13g2_xnor2_1 _20807_ (.Y(_01654_),
    .A(net38),
    .B(_01653_));
 sg13g2_nor2b_1 _20808_ (.A(_01609_),
    .B_N(_01654_),
    .Y(_01656_));
 sg13g2_inv_1 _20809_ (.Y(_01657_),
    .A(_01656_));
 sg13g2_nand2b_1 _20810_ (.Y(_01658_),
    .B(_01609_),
    .A_N(_01654_));
 sg13g2_nand2_1 _20811_ (.Y(_01659_),
    .A(_01657_),
    .B(_01658_));
 sg13g2_inv_1 _20812_ (.Y(_01660_),
    .A(_01659_));
 sg13g2_mux2_1 _20813_ (.A0(_01543_),
    .A1(_01548_),
    .S(net42),
    .X(_01661_));
 sg13g2_xnor2_1 _20814_ (.Y(_01662_),
    .A(net51),
    .B(_01661_));
 sg13g2_nor2b_1 _20815_ (.A(net44),
    .B_N(_01606_),
    .Y(_01663_));
 sg13g2_a21oi_1 _20816_ (.A1(_01602_),
    .A2(net42),
    .Y(_01664_),
    .B1(_01663_));
 sg13g2_xnor2_1 _20817_ (.Y(_01665_),
    .A(net38),
    .B(_01664_));
 sg13g2_nor2b_1 _20818_ (.A(_01662_),
    .B_N(_01665_),
    .Y(_01667_));
 sg13g2_nand2b_1 _20819_ (.Y(_01668_),
    .B(_01662_),
    .A_N(_01665_));
 sg13g2_nor2b_1 _20820_ (.A(_01667_),
    .B_N(_01668_),
    .Y(_01669_));
 sg13g2_nand2_1 _20821_ (.Y(_01670_),
    .A(_01669_),
    .B(_01553_));
 sg13g2_a21oi_1 _20822_ (.A1(_01668_),
    .A2(_01551_),
    .Y(_01671_),
    .B1(_01667_));
 sg13g2_o21ai_1 _20823_ (.B1(_01671_),
    .Y(_01672_),
    .A1(_01493_),
    .A2(_01670_));
 sg13g2_xnor2_1 _20824_ (.Y(_01673_),
    .A(_01660_),
    .B(_01672_));
 sg13g2_nor2_1 _20825_ (.A(_01555_),
    .B(_01673_),
    .Y(_01674_));
 sg13g2_inv_1 _20826_ (.Y(_01675_),
    .A(_01674_));
 sg13g2_nand2_1 _20827_ (.Y(_01676_),
    .A(_01673_),
    .B(_01555_));
 sg13g2_nand2_1 _20828_ (.Y(_01677_),
    .A(_01675_),
    .B(_01676_));
 sg13g2_nand2_1 _20829_ (.Y(_01678_),
    .A(_01488_),
    .B(_01489_));
 sg13g2_nand2_1 _20830_ (.Y(_01679_),
    .A(_01491_),
    .B(_01401_));
 sg13g2_xor2_1 _20831_ (.B(_01679_),
    .A(_01678_),
    .X(_01680_));
 sg13g2_inv_1 _20832_ (.Y(_01681_),
    .A(_01680_));
 sg13g2_nor2b_1 _20833_ (.A(_01413_),
    .B_N(_01481_),
    .Y(_01682_));
 sg13g2_xnor2_1 _20834_ (.Y(_01683_),
    .A(_01480_),
    .B(_01682_));
 sg13g2_inv_1 _20835_ (.Y(_01684_),
    .A(_01683_));
 sg13g2_xnor2_1 _20836_ (.Y(_01685_),
    .A(_01482_),
    .B(_01487_));
 sg13g2_inv_1 _20837_ (.Y(_01686_),
    .A(_01685_));
 sg13g2_nor2_1 _20838_ (.A(_01686_),
    .B(_01555_),
    .Y(_01688_));
 sg13g2_a21oi_1 _20839_ (.A1(_01681_),
    .A2(_01684_),
    .Y(_01689_),
    .B1(_01688_));
 sg13g2_xnor2_1 _20840_ (.Y(_01690_),
    .A(_01477_),
    .B(_01422_));
 sg13g2_inv_1 _20841_ (.Y(_01691_),
    .A(_01690_));
 sg13g2_xor2_1 _20842_ (.B(_01474_),
    .A(_01468_),
    .X(_01692_));
 sg13g2_xnor2_1 _20843_ (.Y(_01693_),
    .A(_01458_),
    .B(_01459_));
 sg13g2_xnor2_1 _20844_ (.Y(_01694_),
    .A(_01466_),
    .B(_01432_));
 sg13g2_a21oi_1 _20845_ (.A1(_01691_),
    .A2(_01693_),
    .Y(_01695_),
    .B1(_01694_));
 sg13g2_xor2_1 _20846_ (.B(_01463_),
    .A(_01462_),
    .X(_01696_));
 sg13g2_a21oi_1 _20847_ (.A1(_01691_),
    .A2(_01694_),
    .Y(_01697_),
    .B1(_01696_));
 sg13g2_nor3_1 _20848_ (.A(_01695_),
    .B(_01697_),
    .C(_01684_),
    .Y(_01699_));
 sg13g2_nand2_1 _20849_ (.Y(_01700_),
    .A(_01691_),
    .B(_01696_));
 sg13g2_nand3_1 _20850_ (.B(_01695_),
    .C(_01700_),
    .A(_01684_),
    .Y(_01701_));
 sg13g2_o21ai_1 _20851_ (.B1(_01701_),
    .Y(_01702_),
    .A1(_01692_),
    .A2(_01699_));
 sg13g2_o21ai_1 _20852_ (.B1(_01702_),
    .Y(_01703_),
    .A1(_01685_),
    .A2(_01690_));
 sg13g2_o21ai_1 _20853_ (.B1(_01703_),
    .Y(_01704_),
    .A1(_01686_),
    .A2(_01691_));
 sg13g2_o21ai_1 _20854_ (.B1(_01704_),
    .Y(_01705_),
    .A1(_01681_),
    .A2(_01684_));
 sg13g2_nand2_1 _20855_ (.Y(_01706_),
    .A(_01689_),
    .B(_01705_));
 sg13g2_nand2b_1 _20856_ (.Y(_01707_),
    .B(_01552_),
    .A_N(_01493_));
 sg13g2_nand2b_1 _20857_ (.Y(_01708_),
    .B(_01707_),
    .A_N(_01551_));
 sg13g2_xor2_1 _20858_ (.B(_01669_),
    .A(_01708_),
    .X(_01710_));
 sg13g2_nor2_1 _20859_ (.A(_01681_),
    .B(_01710_),
    .Y(_01711_));
 sg13g2_nand2_1 _20860_ (.Y(_01712_),
    .A(_01711_),
    .B(_01688_));
 sg13g2_nand2_1 _20861_ (.Y(_01713_),
    .A(_01706_),
    .B(_01712_));
 sg13g2_a21oi_1 _20862_ (.A1(_01555_),
    .A2(_01686_),
    .Y(_01714_),
    .B1(_01711_));
 sg13g2_nand2_1 _20863_ (.Y(_01715_),
    .A(_01710_),
    .B(_01681_));
 sg13g2_a21oi_1 _20864_ (.A1(_01714_),
    .A2(_01715_),
    .Y(_01716_),
    .B1(_01688_));
 sg13g2_o21ai_1 _20865_ (.B1(_01715_),
    .Y(_01717_),
    .A1(_01713_),
    .A2(_01716_));
 sg13g2_nand2b_1 _20866_ (.Y(_01718_),
    .B(_01717_),
    .A_N(_01677_));
 sg13g2_inv_1 _20867_ (.Y(_01719_),
    .A(_01710_));
 sg13g2_nand2_1 _20868_ (.Y(_01721_),
    .A(_06695_),
    .B(_06238_));
 sg13g2_xnor2_1 _20869_ (.Y(_01722_),
    .A(_05807_),
    .B(_06232_));
 sg13g2_xnor2_1 _20870_ (.Y(_01723_),
    .A(_01721_),
    .B(_01722_));
 sg13g2_nand2_1 _20871_ (.Y(_01724_),
    .A(_01613_),
    .B(_01560_));
 sg13g2_o21ai_1 _20872_ (.B1(_01612_),
    .Y(_01725_),
    .A1(_01610_),
    .A2(_01616_));
 sg13g2_o21ai_1 _20873_ (.B1(_01725_),
    .Y(_01726_),
    .A1(_01724_),
    .A2(_01565_));
 sg13g2_xnor2_1 _20874_ (.Y(_01727_),
    .A(_01723_),
    .B(_01726_));
 sg13g2_buf_1 _20875_ (.A(_01727_),
    .X(_01728_));
 sg13g2_inv_1 _20876_ (.Y(_01729_),
    .A(_01728_));
 sg13g2_xnor2_1 _20877_ (.Y(_01730_),
    .A(_01584_),
    .B(_01629_));
 sg13g2_nand2_1 _20878_ (.Y(_01732_),
    .A(_01592_),
    .B(_01588_));
 sg13g2_nor2_1 _20879_ (.A(_01585_),
    .B(_01632_),
    .Y(_01733_));
 sg13g2_a21oi_1 _20880_ (.A1(_01732_),
    .A2(_01733_),
    .Y(_01734_),
    .B1(_01630_));
 sg13g2_xnor2_1 _20881_ (.Y(_01735_),
    .A(_01730_),
    .B(_01734_));
 sg13g2_nor2_1 _20882_ (.A(_01729_),
    .B(_01735_),
    .Y(_01736_));
 sg13g2_nor2b_1 _20883_ (.A(_01728_),
    .B_N(_01735_),
    .Y(_01737_));
 sg13g2_or2_1 _20884_ (.X(_01738_),
    .B(_01737_),
    .A(_01736_));
 sg13g2_buf_1 _20885_ (.A(_01738_),
    .X(_01739_));
 sg13g2_inv_1 _20886_ (.Y(_01740_),
    .A(_01638_));
 sg13g2_nand2_1 _20887_ (.Y(_01741_),
    .A(_01646_),
    .B(_01643_));
 sg13g2_o21ai_1 _20888_ (.B1(_01741_),
    .Y(_01743_),
    .A1(_01740_),
    .A2(_01620_));
 sg13g2_xor2_1 _20889_ (.B(_01743_),
    .A(_01739_),
    .X(_01744_));
 sg13g2_a21oi_1 _20890_ (.A1(_01642_),
    .A2(_01594_),
    .Y(_01745_),
    .B1(_01641_));
 sg13g2_nand3_1 _20891_ (.B(_01605_),
    .C(_01597_),
    .A(_01642_),
    .Y(_01746_));
 sg13g2_nand2_1 _20892_ (.Y(_01747_),
    .A(_01745_),
    .B(_01746_));
 sg13g2_xnor2_1 _20893_ (.Y(_01748_),
    .A(_01747_),
    .B(_01739_));
 sg13g2_inv_1 _20894_ (.Y(_01749_),
    .A(_01748_));
 sg13g2_nand2_1 _20895_ (.Y(_01750_),
    .A(_01749_),
    .B(net41));
 sg13g2_o21ai_1 _20896_ (.B1(_01750_),
    .Y(_01751_),
    .A1(net41),
    .A2(_01744_));
 sg13g2_xnor2_1 _20897_ (.Y(_01752_),
    .A(net39),
    .B(_01751_));
 sg13g2_nor2b_1 _20898_ (.A(net41),
    .B_N(_01651_),
    .Y(_01754_));
 sg13g2_a21oi_1 _20899_ (.A1(_01647_),
    .A2(net41),
    .Y(_01755_),
    .B1(_01754_));
 sg13g2_xnor2_1 _20900_ (.Y(_01756_),
    .A(net53),
    .B(_01755_));
 sg13g2_nand2b_1 _20901_ (.Y(_01757_),
    .B(_01756_),
    .A_N(_01752_));
 sg13g2_nand2b_1 _20902_ (.Y(_01758_),
    .B(_01752_),
    .A_N(_01756_));
 sg13g2_nand2_1 _20903_ (.Y(_01759_),
    .A(_01757_),
    .B(_01758_));
 sg13g2_nand3_1 _20904_ (.B(_01669_),
    .C(_01708_),
    .A(_01660_),
    .Y(_01760_));
 sg13g2_a21oi_1 _20905_ (.A1(_01658_),
    .A2(_01667_),
    .Y(_01761_),
    .B1(_01656_));
 sg13g2_nand2_1 _20906_ (.Y(_01762_),
    .A(_01760_),
    .B(_01761_));
 sg13g2_xor2_1 _20907_ (.B(_01762_),
    .A(_01759_),
    .X(_01763_));
 sg13g2_nor2_1 _20908_ (.A(_01719_),
    .B(_01763_),
    .Y(_01764_));
 sg13g2_inv_1 _20909_ (.Y(_01765_),
    .A(_01764_));
 sg13g2_nand3_1 _20910_ (.B(_01675_),
    .C(_01765_),
    .A(_01718_),
    .Y(_01766_));
 sg13g2_nand2_1 _20911_ (.Y(_01767_),
    .A(_01763_),
    .B(_01719_));
 sg13g2_nand2_1 _20912_ (.Y(_01768_),
    .A(_01672_),
    .B(_01660_));
 sg13g2_nand3_1 _20913_ (.B(_01657_),
    .C(_01758_),
    .A(_01768_),
    .Y(_01769_));
 sg13g2_nand2_1 _20914_ (.Y(_01770_),
    .A(_01749_),
    .B(net42));
 sg13g2_o21ai_1 _20915_ (.B1(_01770_),
    .Y(_01771_),
    .A1(net42),
    .A2(_01744_));
 sg13g2_xnor2_1 _20916_ (.Y(_01772_),
    .A(net51),
    .B(_01771_));
 sg13g2_inv_1 _20917_ (.Y(_01773_),
    .A(_01584_));
 sg13g2_nand3_1 _20918_ (.B(_01730_),
    .C(_01634_),
    .A(_01637_),
    .Y(_01775_));
 sg13g2_nand2_1 _20919_ (.Y(_01776_),
    .A(_01775_),
    .B(_01631_));
 sg13g2_a21oi_1 _20920_ (.A1(_01773_),
    .A2(_01629_),
    .Y(_01777_),
    .B1(_01776_));
 sg13g2_xnor2_1 _20921_ (.Y(_01778_),
    .A(_01728_),
    .B(_01777_));
 sg13g2_nand2_1 _20922_ (.Y(_01779_),
    .A(_01743_),
    .B(_01739_));
 sg13g2_o21ai_1 _20923_ (.B1(_01779_),
    .Y(_01780_),
    .A1(_01728_),
    .A2(_01735_));
 sg13g2_xnor2_1 _20924_ (.Y(_01781_),
    .A(_01778_),
    .B(_01780_));
 sg13g2_nand2_1 _20925_ (.Y(_01782_),
    .A(_01650_),
    .B(_01642_));
 sg13g2_nor2_1 _20926_ (.A(_01641_),
    .B(_01736_),
    .Y(_01783_));
 sg13g2_a21oi_1 _20927_ (.A1(_01782_),
    .A2(_01783_),
    .Y(_01784_),
    .B1(_01737_));
 sg13g2_xnor2_1 _20928_ (.Y(_01786_),
    .A(_01778_),
    .B(_01784_));
 sg13g2_nand2_1 _20929_ (.Y(_01787_),
    .A(_01786_),
    .B(_01603_));
 sg13g2_o21ai_1 _20930_ (.B1(_01787_),
    .Y(_01788_),
    .A1(net41),
    .A2(_01781_));
 sg13g2_xnor2_1 _20931_ (.Y(_01789_),
    .A(net38),
    .B(_01788_));
 sg13g2_nor2_1 _20932_ (.A(_01772_),
    .B(_01789_),
    .Y(_01790_));
 sg13g2_nand2_1 _20933_ (.Y(_01791_),
    .A(_01789_),
    .B(_01772_));
 sg13g2_nor2b_1 _20934_ (.A(_01790_),
    .B_N(_01791_),
    .Y(_01792_));
 sg13g2_a21oi_1 _20935_ (.A1(_01757_),
    .A2(_01769_),
    .Y(_01793_),
    .B1(_01792_));
 sg13g2_nand3_1 _20936_ (.B(_01757_),
    .C(_01769_),
    .A(_01792_),
    .Y(_01794_));
 sg13g2_nand2b_1 _20937_ (.Y(_01795_),
    .B(_01794_),
    .A_N(_01793_));
 sg13g2_buf_1 _20938_ (.A(_01795_),
    .X(_01797_));
 sg13g2_nor2_1 _20939_ (.A(_01673_),
    .B(_01797_),
    .Y(_01798_));
 sg13g2_nand2_1 _20940_ (.Y(_01799_),
    .A(_01797_),
    .B(_01673_));
 sg13g2_nor2b_1 _20941_ (.A(_01798_),
    .B_N(_01799_),
    .Y(_01800_));
 sg13g2_a21oi_1 _20942_ (.A1(_01766_),
    .A2(_01767_),
    .Y(_01801_),
    .B1(_01800_));
 sg13g2_nand3_1 _20943_ (.B(_01767_),
    .C(_01766_),
    .A(_01800_),
    .Y(_01802_));
 sg13g2_nor2b_1 _20944_ (.A(_01801_),
    .B_N(_01802_),
    .Y(\vgadonut.donut.donuthit.cordicxz.x2out[10] ));
 sg13g2_nand2_1 _20945_ (.Y(_01803_),
    .A(_01786_),
    .B(net42));
 sg13g2_o21ai_1 _20946_ (.B1(_01803_),
    .Y(_01804_),
    .A1(net42),
    .A2(_01781_));
 sg13g2_xnor2_1 _20947_ (.Y(_01805_),
    .A(net51),
    .B(_01804_));
 sg13g2_nor2b_1 _20948_ (.A(_01739_),
    .B_N(_01778_),
    .Y(_01807_));
 sg13g2_a21oi_1 _20949_ (.A1(_01777_),
    .A2(_01735_),
    .Y(_01808_),
    .B1(_01729_));
 sg13g2_a21o_1 _20950_ (.A2(_01747_),
    .A1(_01807_),
    .B1(_01808_),
    .X(_01809_));
 sg13g2_xnor2_1 _20951_ (.Y(_01810_),
    .A(_01729_),
    .B(_01629_));
 sg13g2_nor2_1 _20952_ (.A(_01728_),
    .B(_01629_),
    .Y(_01811_));
 sg13g2_a21oi_1 _20953_ (.A1(_01809_),
    .A2(_01810_),
    .Y(_01812_),
    .B1(_01811_));
 sg13g2_a21o_1 _20954_ (.A2(_01735_),
    .A1(_01777_),
    .B1(_01728_),
    .X(_01813_));
 sg13g2_o21ai_1 _20955_ (.B1(_01813_),
    .Y(_01814_),
    .A1(_01778_),
    .A2(_01779_));
 sg13g2_xor2_1 _20956_ (.B(_01814_),
    .A(_01810_),
    .X(_01815_));
 sg13g2_nand2_1 _20957_ (.Y(_01816_),
    .A(_01815_),
    .B(_01494_));
 sg13g2_o21ai_1 _20958_ (.B1(_01816_),
    .Y(_01817_),
    .A1(_01494_),
    .A2(_01812_));
 sg13g2_xnor2_1 _20959_ (.Y(_01818_),
    .A(net38),
    .B(_01817_));
 sg13g2_or2_1 _20960_ (.X(_01819_),
    .B(_01818_),
    .A(_01805_));
 sg13g2_nand2_1 _20961_ (.Y(_01820_),
    .A(_01818_),
    .B(_01805_));
 sg13g2_nand2_1 _20962_ (.Y(_01821_),
    .A(_01819_),
    .B(_01820_));
 sg13g2_a21oi_1 _20963_ (.A1(_01760_),
    .A2(_01761_),
    .Y(_01822_),
    .B1(_01759_));
 sg13g2_inv_1 _20964_ (.Y(_01823_),
    .A(_01790_));
 sg13g2_nand2_1 _20965_ (.Y(_01824_),
    .A(_01823_),
    .B(_01758_));
 sg13g2_o21ai_1 _20966_ (.B1(_01791_),
    .Y(_01825_),
    .A1(_01822_),
    .A2(_01824_));
 sg13g2_xor2_1 _20967_ (.B(_01825_),
    .A(_01821_),
    .X(_01826_));
 sg13g2_nor2b_1 _20968_ (.A(_01763_),
    .B_N(_01826_),
    .Y(_01828_));
 sg13g2_nand2b_1 _20969_ (.Y(_01829_),
    .B(_01763_),
    .A_N(_01826_));
 sg13g2_nor2b_1 _20970_ (.A(_01828_),
    .B_N(_01829_),
    .Y(_01830_));
 sg13g2_nand2_1 _20971_ (.Y(_01831_),
    .A(_01714_),
    .B(_01706_));
 sg13g2_nand3_1 _20972_ (.B(_01715_),
    .C(_01831_),
    .A(_01675_),
    .Y(_01832_));
 sg13g2_nand2_1 _20973_ (.Y(_01833_),
    .A(_01832_),
    .B(_01676_));
 sg13g2_nor2b_1 _20974_ (.A(_01764_),
    .B_N(_01767_),
    .Y(_01834_));
 sg13g2_nor2b_1 _20975_ (.A(_01833_),
    .B_N(_01834_),
    .Y(_01835_));
 sg13g2_o21ai_1 _20976_ (.B1(_01765_),
    .Y(_01836_),
    .A1(_01673_),
    .A2(_01797_));
 sg13g2_o21ai_1 _20977_ (.B1(_01799_),
    .Y(_01837_),
    .A1(_01835_),
    .A2(_01836_));
 sg13g2_xnor2_1 _20978_ (.Y(\vgadonut.donut.donuthit.cordicxz.x2out[11] ),
    .A(_01830_),
    .B(_01837_));
 sg13g2_nor2_1 _20979_ (.A(_01603_),
    .B(_01812_),
    .Y(_01839_));
 sg13g2_a21oi_1 _20980_ (.A1(_01815_),
    .A2(net41),
    .Y(_01840_),
    .B1(_01839_));
 sg13g2_xnor2_1 _20981_ (.Y(_01841_),
    .A(net51),
    .B(_01840_));
 sg13g2_xnor2_1 _20982_ (.Y(_01842_),
    .A(_01841_),
    .B(_01818_));
 sg13g2_nand3_1 _20983_ (.B(_01823_),
    .C(_01819_),
    .A(_01794_),
    .Y(_01843_));
 sg13g2_nand2_1 _20984_ (.Y(_01844_),
    .A(_01843_),
    .B(_01820_));
 sg13g2_xnor2_1 _20985_ (.Y(_01845_),
    .A(_01842_),
    .B(_01844_));
 sg13g2_nand2b_1 _20986_ (.Y(_01846_),
    .B(_01797_),
    .A_N(_01845_));
 sg13g2_nand2b_1 _20987_ (.Y(_01847_),
    .B(_01845_),
    .A_N(_01797_));
 sg13g2_nand2_1 _20988_ (.Y(_01848_),
    .A(_01846_),
    .B(_01847_));
 sg13g2_inv_1 _20989_ (.Y(_01849_),
    .A(_01828_));
 sg13g2_nand3b_1 _20990_ (.B(_01802_),
    .C(_01849_),
    .Y(_01850_),
    .A_N(_01798_));
 sg13g2_nand2_1 _20991_ (.Y(_01851_),
    .A(_01850_),
    .B(_01829_));
 sg13g2_xor2_1 _20992_ (.B(_01851_),
    .A(_01848_),
    .X(\vgadonut.donut.donuthit.cordicxz.x2out[12] ));
 sg13g2_xor2_1 _20993_ (.B(_01845_),
    .A(_01826_),
    .X(_01852_));
 sg13g2_nand2_1 _20994_ (.Y(_01853_),
    .A(_01847_),
    .B(_01849_));
 sg13g2_nor2b_1 _20995_ (.A(_01837_),
    .B_N(_01830_),
    .Y(_01854_));
 sg13g2_o21ai_1 _20996_ (.B1(_01846_),
    .Y(_01855_),
    .A1(_01853_),
    .A2(_01854_));
 sg13g2_xnor2_1 _20997_ (.Y(\vgadonut.donut.donuthit.cordicxz.x2out[13] ),
    .A(_01852_),
    .B(_01855_));
 sg13g2_xnor2_1 _20998_ (.Y(\vgadonut.donut.donuthit.cordicxz.x2out[8] ),
    .A(_01677_),
    .B(_01717_));
 sg13g2_xnor2_1 _20999_ (.Y(\vgadonut.donut.donuthit.cordicxz.x2out[9] ),
    .A(_01833_),
    .B(_01834_));
 sg13g2_dfrbp_1 _21000_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net299),
    .D(_00000_),
    .Q_N(_10653_),
    .Q(_00028_));
 sg13g2_dfrbp_1 _21001_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net300),
    .D(_00001_),
    .Q_N(_10654_),
    .Q(_00029_));
 sg13g2_dfrbp_1 _21002_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net301),
    .D(_00002_),
    .Q_N(_10655_),
    .Q(_00030_));
 sg13g2_dfrbp_1 _21003_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net302),
    .D(_00003_),
    .Q_N(_10656_),
    .Q(_00031_));
 sg13g2_dfrbp_1 _21004_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net303),
    .D(_00004_),
    .Q_N(_10657_),
    .Q(_00034_));
 sg13g2_dfrbp_1 _21005_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net304),
    .D(_00005_),
    .Q_N(_00104_),
    .Q(_00035_));
 sg13g2_dfrbp_1 _21006_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net305),
    .D(_00006_),
    .Q_N(_00103_),
    .Q(_00036_));
 sg13g2_dfrbp_1 _21007_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net306),
    .D(_00007_),
    .Q_N(_00102_),
    .Q(_00037_));
 sg13g2_dfrbp_1 _21008_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net307),
    .D(_00008_),
    .Q_N(_00101_),
    .Q(_00038_));
 sg13g2_dfrbp_1 _21009_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net308),
    .D(_00009_),
    .Q_N(_10658_),
    .Q(_00040_));
 sg13g2_dfrbp_1 _21010_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net309),
    .D(_00010_),
    .Q_N(_00100_),
    .Q(_00041_));
 sg13g2_dfrbp_1 _21011_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net310),
    .D(_00011_),
    .Q_N(_10659_),
    .Q(_00042_));
 sg13g2_dfrbp_1 _21012_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net311),
    .D(_00012_),
    .Q_N(_00099_),
    .Q(_00043_));
 sg13g2_dfrbp_1 _21013_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net312),
    .D(_00013_),
    .Q_N(_10652_),
    .Q(_00044_));
 sg13g2_dfrbp_1 _21014_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net313),
    .D(_00226_),
    .Q_N(_10651_),
    .Q(_00039_));
 sg13g2_dfrbp_1 _21015_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net314),
    .D(_00227_),
    .Q_N(_10650_),
    .Q(_00033_));
 sg13g2_dfrbp_1 _21016_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net315),
    .D(_00228_),
    .Q_N(_00098_),
    .Q(_00045_));
 sg13g2_dfrbp_1 _21017_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net316),
    .D(_00229_),
    .Q_N(_10649_),
    .Q(_00032_));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_tiehi _21000__299 (.L_HI(net299));
 sg13g2_buf_1 _21020_ (.A(net283),
    .X(uio_oe[0]));
 sg13g2_buf_1 _21021_ (.A(net284),
    .X(uio_oe[1]));
 sg13g2_buf_1 _21022_ (.A(net285),
    .X(uio_oe[2]));
 sg13g2_buf_1 _21023_ (.A(net286),
    .X(uio_oe[3]));
 sg13g2_buf_1 _21024_ (.A(net287),
    .X(uio_oe[4]));
 sg13g2_buf_1 _21025_ (.A(net288),
    .X(uio_oe[5]));
 sg13g2_buf_1 _21026_ (.A(net289),
    .X(uio_oe[6]));
 sg13g2_buf_1 _21027_ (.A(net290),
    .X(uio_oe[7]));
 sg13g2_buf_1 _21028_ (.A(net291),
    .X(uio_out[0]));
 sg13g2_buf_1 _21029_ (.A(net292),
    .X(uio_out[1]));
 sg13g2_buf_1 _21030_ (.A(net293),
    .X(uio_out[2]));
 sg13g2_buf_1 _21031_ (.A(net294),
    .X(uio_out[3]));
 sg13g2_buf_1 _21032_ (.A(net295),
    .X(uio_out[4]));
 sg13g2_buf_1 _21033_ (.A(net296),
    .X(uio_out[5]));
 sg13g2_buf_1 _21034_ (.A(net297),
    .X(uio_out[6]));
 sg13g2_buf_1 _21035_ (.A(net298),
    .X(uio_out[7]));
 sg13g2_buf_1 _21036_ (.A(\vgadonut.vsync ),
    .X(net5));
 sg13g2_buf_1 _21037_ (.A(hsync),
    .X(net9));
 sg13g2_dfrbp_1 \vgadonut.b_out[0]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net317),
    .D(_00230_),
    .Q_N(_10648_),
    .Q(net8));
 sg13g2_dfrbp_1 \vgadonut.b_out[1]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net318),
    .D(_00231_),
    .Q_N(_10647_),
    .Q(net4));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net259),
    .D(_00232_),
    .Q_N(\vgadonut.donut.cA[0] ),
    .Q(_00185_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[10]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net270),
    .D(_00233_),
    .Q_N(\vgadonut.donut.cA[10] ),
    .Q(_00186_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[11]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net270),
    .D(_00234_),
    .Q_N(\vgadonut.donut.cA[11] ),
    .Q(_00187_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net259),
    .D(_00235_),
    .Q_N(_10646_),
    .Q(\vgadonut.donut.cA[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[13]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net270),
    .D(_00236_),
    .Q_N(\vgadonut.donut.cA[13] ),
    .Q(_00188_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net260),
    .D(_00237_),
    .Q_N(_10645_),
    .Q(\vgadonut.donut.cA[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net275),
    .D(_00238_),
    .Q_N(_10644_),
    .Q(\vgadonut.donut.cA[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net260),
    .D(_00239_),
    .Q_N(\vgadonut.donut.cA[1] ),
    .Q(_00189_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net260),
    .D(_00240_),
    .Q_N(\vgadonut.donut.cA[2] ),
    .Q(_00190_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net260),
    .D(_00241_),
    .Q_N(\vgadonut.donut.cA[3] ),
    .Q(_00191_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net260),
    .D(_00242_),
    .Q_N(\vgadonut.donut.cA[4] ),
    .Q(_00192_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net270),
    .D(_00243_),
    .Q_N(\vgadonut.donut.cA[5] ),
    .Q(_00193_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net260),
    .D(_00244_),
    .Q_N(_10643_),
    .Q(\vgadonut.donut.cA[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net261),
    .D(_00245_),
    .Q_N(_10642_),
    .Q(\vgadonut.donut.cA[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[8]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net270),
    .D(_00246_),
    .Q_N(\vgadonut.donut.cA[8] ),
    .Q(_00194_));
 sg13g2_dfrbp_1 \vgadonut.donut.cA[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net261),
    .D(_00247_),
    .Q_N(_10641_),
    .Q(\vgadonut.donut.cA[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net263),
    .D(_00248_),
    .Q_N(\vgadonut.donut.cAcB[0] ),
    .Q(_00195_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[10]$_DFFE_PN1P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net261),
    .D(_00249_),
    .Q_N(\vgadonut.donut.cAcB[10] ),
    .Q(_00196_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[11]$_DFFE_PN1P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net261),
    .D(_00250_),
    .Q_N(\vgadonut.donut.cAcB[11] ),
    .Q(_00197_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net261),
    .D(_00251_),
    .Q_N(_10640_),
    .Q(\vgadonut.donut.cAcB[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[13]$_DFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net266),
    .D(_00252_),
    .Q_N(\vgadonut.donut.cAcB[13] ),
    .Q(_00198_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net261),
    .D(_00253_),
    .Q_N(_10639_),
    .Q(\vgadonut.donut.cAcB[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net264),
    .D(_00254_),
    .Q_N(_10638_),
    .Q(\vgadonut.donut.cAcB[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net264),
    .D(_00255_),
    .Q_N(\vgadonut.donut.cAcB[1] ),
    .Q(_00199_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net266),
    .D(_00256_),
    .Q_N(\vgadonut.donut.cAcB[2] ),
    .Q(_00200_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net266),
    .D(_00257_),
    .Q_N(\vgadonut.donut.cAcB[3] ),
    .Q(_00201_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net266),
    .D(_00258_),
    .Q_N(\vgadonut.donut.cAcB[4] ),
    .Q(_00202_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net266),
    .D(_00259_),
    .Q_N(\vgadonut.donut.cAcB[5] ),
    .Q(_00203_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net266),
    .D(_00260_),
    .Q_N(_10637_),
    .Q(\vgadonut.donut.cAcB[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net266),
    .D(_00261_),
    .Q_N(_10636_),
    .Q(\vgadonut.donut.cAcB[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[8]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net266),
    .D(_00262_),
    .Q_N(\vgadonut.donut.cAcB[8] ),
    .Q(_00204_));
 sg13g2_dfrbp_1 \vgadonut.donut.cAcB[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net267),
    .D(_00263_),
    .Q_N(_10635_),
    .Q(\vgadonut.donut.cAcB[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net281),
    .D(_00264_),
    .Q_N(_00108_),
    .Q(\vgadonut.donut.cAsB[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net263),
    .D(_00265_),
    .Q_N(_00115_),
    .Q(\vgadonut.donut.cAsB[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net264),
    .D(_00266_),
    .Q_N(_00116_),
    .Q(\vgadonut.donut.cAsB[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net264),
    .D(_00267_),
    .Q_N(_00117_),
    .Q(\vgadonut.donut.cAsB[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net264),
    .D(_00268_),
    .Q_N(_00118_),
    .Q(\vgadonut.donut.cAsB[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net264),
    .D(_00269_),
    .Q_N(_00119_),
    .Q(\vgadonut.donut.cAsB[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net275),
    .D(_00270_),
    .Q_N(_00120_),
    .Q(\vgadonut.donut.cAsB[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net281),
    .D(_00271_),
    .Q_N(_00097_),
    .Q(\vgadonut.donut.cAsB[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net263),
    .D(_00272_),
    .Q_N(_00105_),
    .Q(\vgadonut.donut.cAsB[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net263),
    .D(_00273_),
    .Q_N(_00107_),
    .Q(\vgadonut.donut.cAsB[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net281),
    .D(_00274_),
    .Q_N(_00109_),
    .Q(\vgadonut.donut.cAsB[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net281),
    .D(_00275_),
    .Q_N(_00110_),
    .Q(\vgadonut.donut.cAsB[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net263),
    .D(_00276_),
    .Q_N(_00111_),
    .Q(\vgadonut.donut.cAsB[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net263),
    .D(_00277_),
    .Q_N(_00112_),
    .Q(\vgadonut.donut.cAsB[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net263),
    .D(_00278_),
    .Q_N(_00113_),
    .Q(\vgadonut.donut.cAsB[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cAsB[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net263),
    .D(_00279_),
    .Q_N(_00114_),
    .Q(\vgadonut.donut.cAsB[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net277),
    .D(_00280_),
    .Q_N(_00133_),
    .Q(\vgadonut.donut.cB[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net276),
    .D(_00281_),
    .Q_N(_00140_),
    .Q(\vgadonut.donut.cB[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net276),
    .D(_00282_),
    .Q_N(_00141_),
    .Q(\vgadonut.donut.cB[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net278),
    .D(_00283_),
    .Q_N(_00142_),
    .Q(\vgadonut.donut.cB[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net278),
    .D(_00284_),
    .Q_N(_00143_),
    .Q(\vgadonut.donut.cB[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[14]$_DFFE_PN1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net278),
    .D(_00285_),
    .Q_N(\vgadonut.donut.cB[14] ),
    .Q(_00205_));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net278),
    .D(_00286_),
    .Q_N(_00144_),
    .Q(\vgadonut.donut.cB[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net280),
    .D(_00287_),
    .Q_N(_10634_),
    .Q(\vgadonut.donut.cB[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net277),
    .D(_00288_),
    .Q_N(_10633_),
    .Q(\vgadonut.donut.cB[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net277),
    .D(_00289_),
    .Q_N(_10632_),
    .Q(\vgadonut.donut.cB[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net277),
    .D(_00290_),
    .Q_N(_00134_),
    .Q(\vgadonut.donut.cB[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net277),
    .D(_00291_),
    .Q_N(_00135_),
    .Q(\vgadonut.donut.cB[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net277),
    .D(_00292_),
    .Q_N(_00136_),
    .Q(\vgadonut.donut.cB[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net276),
    .D(_00293_),
    .Q_N(_00137_),
    .Q(\vgadonut.donut.cB[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net276),
    .D(_00294_),
    .Q_N(_00138_),
    .Q(\vgadonut.donut.cB[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.cB[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net276),
    .D(_00295_),
    .Q_N(_00139_),
    .Q(\vgadonut.donut.cB[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donut_luma[0]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net319),
    .D(_00178_),
    .Q_N(_10631_),
    .Q(\vgadonut.donut.donut_luma[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donut_luma[1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net320),
    .D(_00177_),
    .Q_N(_10630_),
    .Q(\vgadonut.donut.donut_luma[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donut_luma[2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net321),
    .D(net87),
    .Q_N(_10629_),
    .Q(\vgadonut.donut.donut_luma[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donut_luma[3]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net322),
    .D(_00180_),
    .Q_N(_10628_),
    .Q(\vgadonut.donut.donut_luma[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donut_luma[4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net323),
    .D(_00173_),
    .Q_N(_10627_),
    .Q(\vgadonut.donut.donut_luma[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donut_luma[5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net324),
    .D(_00014_),
    .Q_N(_10626_),
    .Q(\vgadonut.donut.donut_luma[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donut_visible$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net325),
    .D(_00296_),
    .Q_N(_10625_),
    .Q(\vgadonut.donut.donut_visible ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.hit$_SDFF_PP1_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net326),
    .D(_00297_),
    .Q_N(_10660_),
    .Q(\vgadonut.donut.donuthit.hit ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.light[10]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net327),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[10] ),
    .Q_N(_10661_),
    .Q(\vgadonut.donut.donuthit.light[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.light[11]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net328),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[11] ),
    .Q_N(_10662_),
    .Q(\vgadonut.donut.donuthit.light[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.light[12]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net329),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[12] ),
    .Q_N(_10663_),
    .Q(\vgadonut.donut.donuthit.light[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.light[13]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net330),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[13] ),
    .Q_N(_00046_),
    .Q(\vgadonut.donut.donuthit.light[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.light[8]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net331),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[8] ),
    .Q_N(_10664_),
    .Q(\vgadonut.donut.donuthit.light[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.light[9]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net332),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[9] ),
    .Q_N(_10665_),
    .Q(\vgadonut.donut.donuthit.light[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[0]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net333),
    .D(_00047_),
    .Q_N(_10666_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[10]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net334),
    .D(_00048_),
    .Q_N(_10667_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[11]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net335),
    .D(_00049_),
    .Q_N(_10668_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[12]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net336),
    .D(_00050_),
    .Q_N(_10669_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[13]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net337),
    .D(_00051_),
    .Q_N(_00175_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[14]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net338),
    .D(_00052_),
    .Q_N(_00176_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[15]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net339),
    .D(_00053_),
    .Q_N(_10670_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[1]$_DFF_P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net340),
    .D(_00054_),
    .Q_N(_10671_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[2]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net341),
    .D(_00055_),
    .Q_N(_10672_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[3]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net342),
    .D(_00056_),
    .Q_N(_10673_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[4]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net343),
    .D(_00057_),
    .Q_N(_10674_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[5]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net344),
    .D(_00058_),
    .Q_N(_10675_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[6]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net345),
    .D(_00059_),
    .Q_N(_10676_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[7]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net346),
    .D(_00060_),
    .Q_N(_10677_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[8]$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net347),
    .D(_00061_),
    .Q_N(_10678_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.px[9]$_DFF_P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net348),
    .D(_00062_),
    .Q_N(_10679_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[0]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net349),
    .D(_00063_),
    .Q_N(_10680_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[10]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net350),
    .D(_00064_),
    .Q_N(_10681_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[11]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net351),
    .D(_00065_),
    .Q_N(_10682_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[12]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net352),
    .D(_00066_),
    .Q_N(_10683_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[13]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net353),
    .D(_00067_),
    .Q_N(_00182_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[14]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net354),
    .D(_00068_),
    .Q_N(_00183_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[15]$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net355),
    .D(_00069_),
    .Q_N(_10684_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[1]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net356),
    .D(_00070_),
    .Q_N(_10685_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[2]$_DFF_P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net357),
    .D(_00071_),
    .Q_N(_10686_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[3]$_DFF_P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net358),
    .D(_00072_),
    .Q_N(_10687_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[4]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net359),
    .D(_00073_),
    .Q_N(_10688_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[5]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net360),
    .D(_00074_),
    .Q_N(_10689_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[6]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net361),
    .D(_00075_),
    .Q_N(_10690_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[7]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net362),
    .D(_00076_),
    .Q_N(_10691_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[8]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net363),
    .D(_00077_),
    .Q_N(_10692_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.py[9]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net364),
    .D(_00078_),
    .Q_N(_10693_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[0]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net365),
    .D(_00079_),
    .Q_N(_00163_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[10]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net366),
    .D(_00080_),
    .Q_N(_00164_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[11]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net367),
    .D(_00081_),
    .Q_N(_00158_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[12]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net368),
    .D(_00082_),
    .Q_N(_00167_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[13]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net369),
    .D(_00083_),
    .Q_N(_00166_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[14]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net370),
    .D(_00084_),
    .Q_N(_00168_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[15]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net371),
    .D(_00085_),
    .Q_N(_00165_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[1]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net372),
    .D(_00086_),
    .Q_N(_10694_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[2]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net373),
    .D(_00087_),
    .Q_N(_00162_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[3]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net374),
    .D(_00088_),
    .Q_N(_00161_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[4]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net375),
    .D(_00089_),
    .Q_N(_10695_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[5]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net376),
    .D(_00090_),
    .Q_N(_00160_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[6]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net377),
    .D(_00091_),
    .Q_N(_10696_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[7]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net378),
    .D(_00092_),
    .Q_N(_00159_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[8]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net379),
    .D(_00093_),
    .Q_N(_10697_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.pz[9]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net380),
    .D(_00094_),
    .Q_N(_10624_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[10]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net381),
    .D(_00298_),
    .Q_N(_10623_),
    .Q(\vgadonut.donut.donuthit.rx[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[11]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net382),
    .D(_00299_),
    .Q_N(_10622_),
    .Q(\vgadonut.donut.donuthit.rx[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[12]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net383),
    .D(_00300_),
    .Q_N(_10621_),
    .Q(\vgadonut.donut.donuthit.rx[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[13]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net384),
    .D(_00301_),
    .Q_N(_10620_),
    .Q(\vgadonut.donut.donuthit.rx[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[14]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net385),
    .D(_00302_),
    .Q_N(_10619_),
    .Q(\vgadonut.donut.donuthit.rx[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[15]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net386),
    .D(_00303_),
    .Q_N(_10618_),
    .Q(\vgadonut.donut.donuthit.rx[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[5]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net387),
    .D(_00304_),
    .Q_N(_10617_),
    .Q(\vgadonut.donut.donuthit.rx[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net388),
    .D(_00305_),
    .Q_N(_10616_),
    .Q(\vgadonut.donut.donuthit.rx[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[7]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net389),
    .D(_00306_),
    .Q_N(_10615_),
    .Q(\vgadonut.donut.donuthit.rx[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[8]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net390),
    .D(_00307_),
    .Q_N(_10614_),
    .Q(\vgadonut.donut.donuthit.rx[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rx[9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net391),
    .D(_00308_),
    .Q_N(_10613_),
    .Q(\vgadonut.donut.donuthit.rx[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[10]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net392),
    .D(_00309_),
    .Q_N(_10612_),
    .Q(\vgadonut.donut.donuthit.ry[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net393),
    .D(_00310_),
    .Q_N(_10611_),
    .Q(\vgadonut.donut.donuthit.ry[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[12]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net394),
    .D(_00311_),
    .Q_N(_10610_),
    .Q(\vgadonut.donut.donuthit.ry[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[13]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net395),
    .D(_00312_),
    .Q_N(_10609_),
    .Q(\vgadonut.donut.donuthit.ry[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[14]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net396),
    .D(_00313_),
    .Q_N(_10608_),
    .Q(\vgadonut.donut.donuthit.ry[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[15]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net397),
    .D(_00314_),
    .Q_N(_10607_),
    .Q(\vgadonut.donut.donuthit.ry[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net398),
    .D(_00315_),
    .Q_N(_10606_),
    .Q(\vgadonut.donut.donuthit.ry[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[6]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net399),
    .D(_00316_),
    .Q_N(_10605_),
    .Q(\vgadonut.donut.donuthit.ry[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[7]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net400),
    .D(_00317_),
    .Q_N(_10604_),
    .Q(\vgadonut.donut.donuthit.ry[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net401),
    .D(_00318_),
    .Q_N(_10603_),
    .Q(\vgadonut.donut.donuthit.ry[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.ry[9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net402),
    .D(_00319_),
    .Q_N(_10602_),
    .Q(\vgadonut.donut.donuthit.ry[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[10]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net403),
    .D(_00320_),
    .Q_N(_10601_),
    .Q(\vgadonut.donut.donuthit.rz[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[11]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net404),
    .D(_00321_),
    .Q_N(_10600_),
    .Q(\vgadonut.donut.donuthit.rz[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[12]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net405),
    .D(_00322_),
    .Q_N(_10599_),
    .Q(\vgadonut.donut.donuthit.rz[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[13]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net406),
    .D(_00323_),
    .Q_N(_10598_),
    .Q(\vgadonut.donut.donuthit.rz[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[14]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net407),
    .D(_00324_),
    .Q_N(_10597_),
    .Q(\vgadonut.donut.donuthit.rz[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[15]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net408),
    .D(_00325_),
    .Q_N(_10596_),
    .Q(\vgadonut.donut.donuthit.rz[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[5]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net409),
    .D(_00326_),
    .Q_N(_10595_),
    .Q(\vgadonut.donut.donuthit.rz[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net410),
    .D(_00327_),
    .Q_N(_10594_),
    .Q(\vgadonut.donut.donuthit.rz[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net411),
    .D(_00328_),
    .Q_N(_10593_),
    .Q(\vgadonut.donut.donuthit.rz[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[8]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net412),
    .D(_00329_),
    .Q_N(_10592_),
    .Q(\vgadonut.donut.donuthit.rz[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.rz[9]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net413),
    .D(_00330_),
    .Q_N(_10591_),
    .Q(\vgadonut.donut.donuthit.rz[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[0]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net414),
    .D(_00331_),
    .Q_N(_10590_),
    .Q(\vgadonut.donut.donuthit.t[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[10]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net415),
    .D(_00332_),
    .Q_N(_10589_),
    .Q(\vgadonut.donut.donuthit.t[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[11]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net416),
    .D(_00333_),
    .Q_N(_10588_),
    .Q(\vgadonut.donut.donuthit.t[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[12]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net417),
    .D(_00334_),
    .Q_N(_10587_),
    .Q(\vgadonut.donut.donuthit.t[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[13]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net418),
    .D(_00335_),
    .Q_N(_10586_),
    .Q(\vgadonut.donut.donuthit.t[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[14]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net419),
    .D(_00336_),
    .Q_N(_10585_),
    .Q(\vgadonut.donut.donuthit.t[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[15]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net420),
    .D(_00337_),
    .Q_N(_10584_),
    .Q(\vgadonut.donut.donuthit.t[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[1]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net421),
    .D(_00338_),
    .Q_N(_10583_),
    .Q(\vgadonut.donut.donuthit.t[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[2]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net422),
    .D(_00339_),
    .Q_N(_10582_),
    .Q(\vgadonut.donut.donuthit.t[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[3]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net423),
    .D(_00340_),
    .Q_N(_10581_),
    .Q(\vgadonut.donut.donuthit.t[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[4]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net424),
    .D(_00341_),
    .Q_N(_10580_),
    .Q(\vgadonut.donut.donuthit.t[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[5]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net425),
    .D(_00342_),
    .Q_N(_10579_),
    .Q(\vgadonut.donut.donuthit.t[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[6]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net426),
    .D(_00343_),
    .Q_N(_10578_),
    .Q(\vgadonut.donut.donuthit.t[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[7]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net427),
    .D(_00344_),
    .Q_N(_10577_),
    .Q(\vgadonut.donut.donuthit.t[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[8]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net428),
    .D(_00345_),
    .Q_N(_10576_),
    .Q(\vgadonut.donut.donuthit.t[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.donuthit.t[9]$_SDFF_PP1_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net429),
    .D(_00346_),
    .Q_N(_10575_),
    .Q(\vgadonut.donut.donuthit.t[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net430),
    .D(_00347_),
    .Q_N(_10574_),
    .Q(\vgadonut.donut.rx6[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[10]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net431),
    .D(_00348_),
    .Q_N(_10573_),
    .Q(\vgadonut.donut.donuthit.rxin[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[11]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net432),
    .D(_00349_),
    .Q_N(_10572_),
    .Q(\vgadonut.donut.donuthit.rxin[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[12]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net433),
    .D(_00350_),
    .Q_N(_10571_),
    .Q(\vgadonut.donut.donuthit.rxin[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[13]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net434),
    .D(_00351_),
    .Q_N(_10570_),
    .Q(\vgadonut.donut.donuthit.rxin[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[14]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net435),
    .D(_00352_),
    .Q_N(_10569_),
    .Q(\vgadonut.donut.donuthit.rxin[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[15]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net436),
    .D(_00353_),
    .Q_N(_10568_),
    .Q(\vgadonut.donut.donuthit.rxin[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[16]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net437),
    .D(_00354_),
    .Q_N(_10567_),
    .Q(\vgadonut.donut.donuthit.rxin[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net438),
    .D(_00355_),
    .Q_N(_10566_),
    .Q(\vgadonut.donut.donuthit.rxin[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[18]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net439),
    .D(_00356_),
    .Q_N(_10565_),
    .Q(\vgadonut.donut.donuthit.rxin[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[19]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net440),
    .D(_00357_),
    .Q_N(_10564_),
    .Q(\vgadonut.donut.donuthit.rxin[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net441),
    .D(_00358_),
    .Q_N(_10563_),
    .Q(\vgadonut.donut.rx6[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[20]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net442),
    .D(_00359_),
    .Q_N(_10562_),
    .Q(\vgadonut.donut.donuthit.rxin[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[21]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net443),
    .D(_00360_),
    .Q_N(_00174_),
    .Q(\vgadonut.donut.donuthit.rxin[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net444),
    .D(_00361_),
    .Q_N(_10561_),
    .Q(\vgadonut.donut.rx6[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[3]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net445),
    .D(_00362_),
    .Q_N(_10560_),
    .Q(\vgadonut.donut.rx6[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net446),
    .D(_00363_),
    .Q_N(_10559_),
    .Q(\vgadonut.donut.rx6[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[5]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net447),
    .D(_00364_),
    .Q_N(_10558_),
    .Q(\vgadonut.donut.rx6[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[6]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net448),
    .D(_00365_),
    .Q_N(_10557_),
    .Q(\vgadonut.donut.donuthit.rxin[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[7]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net449),
    .D(_00366_),
    .Q_N(_10556_),
    .Q(\vgadonut.donut.donuthit.rxin[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[8]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net450),
    .D(_00367_),
    .Q_N(_10555_),
    .Q(\vgadonut.donut.donuthit.rxin[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rx6[9]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net451),
    .D(_00368_),
    .Q_N(_10554_),
    .Q(\vgadonut.donut.donuthit.rxin[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[0]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net452),
    .D(_00369_),
    .Q_N(_10553_),
    .Q(\vgadonut.donut.ry6[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[10]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net453),
    .D(_00370_),
    .Q_N(_10552_),
    .Q(\vgadonut.donut.donuthit.ryin[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[11]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net454),
    .D(_00371_),
    .Q_N(_00123_),
    .Q(\vgadonut.donut.donuthit.ryin[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[12]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net455),
    .D(_00372_),
    .Q_N(_00124_),
    .Q(\vgadonut.donut.donuthit.ryin[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net456),
    .D(_00373_),
    .Q_N(_00125_),
    .Q(\vgadonut.donut.donuthit.ryin[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net457),
    .D(_00374_),
    .Q_N(_00126_),
    .Q(\vgadonut.donut.donuthit.ryin[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[15]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net458),
    .D(_00375_),
    .Q_N(_00127_),
    .Q(\vgadonut.donut.donuthit.ryin[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[16]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net459),
    .D(_00376_),
    .Q_N(_00128_),
    .Q(\vgadonut.donut.donuthit.ryin[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[17]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net460),
    .D(_00377_),
    .Q_N(_00129_),
    .Q(\vgadonut.donut.donuthit.ryin[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[18]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net461),
    .D(_00378_),
    .Q_N(_00130_),
    .Q(\vgadonut.donut.donuthit.ryin[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[19]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net462),
    .D(_00379_),
    .Q_N(_00131_),
    .Q(\vgadonut.donut.donuthit.ryin[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[1]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net463),
    .D(_00380_),
    .Q_N(_10551_),
    .Q(\vgadonut.donut.ry6[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[20]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net464),
    .D(_00381_),
    .Q_N(_00132_),
    .Q(\vgadonut.donut.donuthit.ryin[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[21]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net465),
    .D(_00382_),
    .Q_N(_00181_),
    .Q(\vgadonut.donut.donuthit.ryin[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[2]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net466),
    .D(_00383_),
    .Q_N(_10550_),
    .Q(\vgadonut.donut.ry6[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[3]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net467),
    .D(_00384_),
    .Q_N(_10549_),
    .Q(\vgadonut.donut.ry6[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[4]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net468),
    .D(_00385_),
    .Q_N(_10548_),
    .Q(\vgadonut.donut.ry6[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[5]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net469),
    .D(_00386_),
    .Q_N(_10547_),
    .Q(\vgadonut.donut.ry6[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[6]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net470),
    .D(_00387_),
    .Q_N(_10546_),
    .Q(\vgadonut.donut.donuthit.ryin[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[7]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net471),
    .D(_00388_),
    .Q_N(_10545_),
    .Q(\vgadonut.donut.donuthit.ryin[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[8]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net472),
    .D(_00389_),
    .Q_N(_10544_),
    .Q(\vgadonut.donut.donuthit.ryin[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ry6[9]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net473),
    .D(_00390_),
    .Q_N(_10543_),
    .Q(\vgadonut.donut.donuthit.ryin[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[0]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net474),
    .D(_00391_),
    .Q_N(_10542_),
    .Q(\vgadonut.donut.rz6[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[10]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net475),
    .D(_00392_),
    .Q_N(_10541_),
    .Q(\vgadonut.donut.donuthit.rzin[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[11]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net476),
    .D(_00393_),
    .Q_N(_10540_),
    .Q(\vgadonut.donut.donuthit.rzin[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[12]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net477),
    .D(_00394_),
    .Q_N(_10539_),
    .Q(\vgadonut.donut.donuthit.rzin[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[13]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net478),
    .D(_00395_),
    .Q_N(_10538_),
    .Q(\vgadonut.donut.donuthit.rzin[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[14]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net479),
    .D(_00396_),
    .Q_N(_10537_),
    .Q(\vgadonut.donut.donuthit.rzin[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[15]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net480),
    .D(_00397_),
    .Q_N(_10536_),
    .Q(\vgadonut.donut.donuthit.rzin[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[16]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net481),
    .D(_00398_),
    .Q_N(_10535_),
    .Q(\vgadonut.donut.donuthit.rzin[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[17]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net482),
    .D(_00399_),
    .Q_N(_10534_),
    .Q(\vgadonut.donut.donuthit.rzin[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[18]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net483),
    .D(_00400_),
    .Q_N(_10533_),
    .Q(\vgadonut.donut.donuthit.rzin[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[19]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net484),
    .D(_00401_),
    .Q_N(_10532_),
    .Q(\vgadonut.donut.donuthit.rzin[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[1]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net485),
    .D(_00402_),
    .Q_N(_10531_),
    .Q(\vgadonut.donut.rz6[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[20]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net486),
    .D(_00403_),
    .Q_N(_10530_),
    .Q(\vgadonut.donut.donuthit.rzin[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[21]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net487),
    .D(_00404_),
    .Q_N(_00095_),
    .Q(\vgadonut.donut.donuthit.rzin[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[2]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net488),
    .D(_00405_),
    .Q_N(_10529_),
    .Q(\vgadonut.donut.rz6[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net489),
    .D(_00406_),
    .Q_N(_10528_),
    .Q(\vgadonut.donut.rz6[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[4]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net490),
    .D(_00407_),
    .Q_N(_10527_),
    .Q(\vgadonut.donut.rz6[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[5]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net491),
    .D(_00408_),
    .Q_N(_10526_),
    .Q(\vgadonut.donut.rz6[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net492),
    .D(_00409_),
    .Q_N(_10525_),
    .Q(\vgadonut.donut.donuthit.rzin[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net493),
    .D(_00410_),
    .Q_N(_10524_),
    .Q(\vgadonut.donut.donuthit.rzin[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[8]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net494),
    .D(_00411_),
    .Q_N(_10523_),
    .Q(\vgadonut.donut.donuthit.rzin[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.rz6[9]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net495),
    .D(_00412_),
    .Q_N(_10522_),
    .Q(\vgadonut.donut.donuthit.rzin[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net271),
    .D(_00413_),
    .Q_N(\vgadonut.donut.sA[0] ),
    .Q(_00206_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[10]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net271),
    .D(_00414_),
    .Q_N(\vgadonut.donut.sA[10] ),
    .Q(_00207_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[11]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net269),
    .D(_00415_),
    .Q_N(\vgadonut.donut.sA[11] ),
    .Q(_00208_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net271),
    .D(_00416_),
    .Q_N(_10521_),
    .Q(\vgadonut.donut.sA[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[13]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net271),
    .D(_00417_),
    .Q_N(\vgadonut.donut.sA[13] ),
    .Q(_00209_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net271),
    .D(_00418_),
    .Q_N(_10520_),
    .Q(\vgadonut.donut.sA[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net271),
    .D(_00419_),
    .Q_N(_10519_),
    .Q(\vgadonut.donut.sA[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net269),
    .D(_00420_),
    .Q_N(\vgadonut.donut.sA[1] ),
    .Q(_00210_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net268),
    .D(_00421_),
    .Q_N(\vgadonut.donut.sA[2] ),
    .Q(_00211_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net268),
    .D(_00422_),
    .Q_N(\vgadonut.donut.sA[3] ),
    .Q(_00212_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net268),
    .D(_00423_),
    .Q_N(\vgadonut.donut.sA[4] ),
    .Q(_00213_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net268),
    .D(_00424_),
    .Q_N(\vgadonut.donut.sA[5] ),
    .Q(_00214_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net268),
    .D(_00425_),
    .Q_N(_10518_),
    .Q(\vgadonut.donut.sA[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net268),
    .D(_00426_),
    .Q_N(_10517_),
    .Q(\vgadonut.donut.sA[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[8]$_DFFE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net268),
    .D(_00427_),
    .Q_N(\vgadonut.donut.sA[8] ),
    .Q(_00215_));
 sg13g2_dfrbp_1 \vgadonut.donut.sA[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net269),
    .D(_00428_),
    .Q_N(_10516_),
    .Q(\vgadonut.donut.sA[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net256),
    .D(_00429_),
    .Q_N(\vgadonut.donut.sAcB[0] ),
    .Q(_00216_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[10]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net256),
    .D(_00430_),
    .Q_N(\vgadonut.donut.sAcB[10] ),
    .Q(_00217_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[11]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net259),
    .D(_00431_),
    .Q_N(\vgadonut.donut.sAcB[11] ),
    .Q(_00218_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net259),
    .D(_00432_),
    .Q_N(_10515_),
    .Q(\vgadonut.donut.sAcB[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[13]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net259),
    .D(_00433_),
    .Q_N(\vgadonut.donut.sAcB[13] ),
    .Q(_00219_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net259),
    .D(_00434_),
    .Q_N(_10514_),
    .Q(\vgadonut.donut.sAcB[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net259),
    .D(_00435_),
    .Q_N(_10513_),
    .Q(\vgadonut.donut.sAcB[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net257),
    .D(_00436_),
    .Q_N(\vgadonut.donut.sAcB[1] ),
    .Q(_00220_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net257),
    .D(_00437_),
    .Q_N(\vgadonut.donut.sAcB[2] ),
    .Q(_00221_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net257),
    .D(_00438_),
    .Q_N(\vgadonut.donut.sAcB[3] ),
    .Q(_00222_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net258),
    .D(_00439_),
    .Q_N(\vgadonut.donut.sAcB[4] ),
    .Q(_00223_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net257),
    .D(_00440_),
    .Q_N(\vgadonut.donut.sAcB[5] ),
    .Q(_00224_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net265),
    .D(_00441_),
    .Q_N(_10512_),
    .Q(\vgadonut.donut.sAcB[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net265),
    .D(_00442_),
    .Q_N(_10511_),
    .Q(\vgadonut.donut.sAcB[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[8]$_DFFE_PN1P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net262),
    .D(_00443_),
    .Q_N(\vgadonut.donut.sAcB[8] ),
    .Q(_00225_));
 sg13g2_dfrbp_1 \vgadonut.donut.sAcB[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net259),
    .D(_00444_),
    .Q_N(_10510_),
    .Q(\vgadonut.donut.sAcB[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net264),
    .D(_00445_),
    .Q_N(_00121_),
    .Q(\vgadonut.donut.sAsB[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net258),
    .D(_00446_),
    .Q_N(_10509_),
    .Q(\vgadonut.donut.sAsB[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net256),
    .D(_00447_),
    .Q_N(_10508_),
    .Q(\vgadonut.donut.sAsB[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net258),
    .D(_00448_),
    .Q_N(_10507_),
    .Q(\vgadonut.donut.sAsB[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net258),
    .D(_00449_),
    .Q_N(_10506_),
    .Q(\vgadonut.donut.sAsB[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net258),
    .D(_00450_),
    .Q_N(_10505_),
    .Q(\vgadonut.donut.sAsB[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net265),
    .D(_00451_),
    .Q_N(_10504_),
    .Q(\vgadonut.donut.sAsB[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net258),
    .D(_00452_),
    .Q_N(_10503_),
    .Q(\vgadonut.donut.sAsB[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net262),
    .D(_00453_),
    .Q_N(_10502_),
    .Q(\vgadonut.donut.sAsB[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net256),
    .D(_00454_),
    .Q_N(_10501_),
    .Q(\vgadonut.donut.sAsB[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net256),
    .D(_00455_),
    .Q_N(_10500_),
    .Q(\vgadonut.donut.sAsB[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net256),
    .D(_00456_),
    .Q_N(_10499_),
    .Q(\vgadonut.donut.sAsB[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net256),
    .D(_00457_),
    .Q_N(_10498_),
    .Q(\vgadonut.donut.sAsB[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net256),
    .D(_00458_),
    .Q_N(_10497_),
    .Q(\vgadonut.donut.sAsB[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net262),
    .D(_00459_),
    .Q_N(_10496_),
    .Q(\vgadonut.donut.sAsB[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sAsB[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net265),
    .D(_00460_),
    .Q_N(_10495_),
    .Q(\vgadonut.donut.sAsB[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net277),
    .D(_00461_),
    .Q_N(_10494_),
    .Q(\vgadonut.donut.sB[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net279),
    .D(_00462_),
    .Q_N(_00149_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net278),
    .D(_00463_),
    .Q_N(_00148_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net278),
    .D(_00464_),
    .Q_N(_00147_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net279),
    .D(_00465_),
    .Q_N(_00146_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net279),
    .D(_00466_),
    .Q_N(_00145_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net282),
    .D(_00467_),
    .Q_N(_00106_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net276),
    .D(_00468_),
    .Q_N(_10493_),
    .Q(\vgadonut.donut.sB[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net276),
    .D(_00469_),
    .Q_N(_00157_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net280),
    .D(_00470_),
    .Q_N(_00156_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net276),
    .D(_00471_),
    .Q_N(_00155_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net278),
    .D(_00472_),
    .Q_N(_00154_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net279),
    .D(_00473_),
    .Q_N(_00153_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net279),
    .D(_00474_),
    .Q_N(_00152_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net278),
    .D(_00475_),
    .Q_N(_00151_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.sB[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net279),
    .D(_00476_),
    .Q_N(_00150_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net496),
    .D(_00477_),
    .Q_N(_10492_),
    .Q(\vgadonut.donut.ycA[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[10]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net497),
    .D(_00478_),
    .Q_N(_10491_),
    .Q(\vgadonut.donut.ycA[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[11]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net498),
    .D(_00479_),
    .Q_N(_10490_),
    .Q(\vgadonut.donut.ycA[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[12]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net499),
    .D(_00480_),
    .Q_N(_10489_),
    .Q(\vgadonut.donut.ycA[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[13]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net500),
    .D(_00481_),
    .Q_N(_10488_),
    .Q(\vgadonut.donut.ycA[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[14]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net501),
    .D(_00482_),
    .Q_N(_10487_),
    .Q(\vgadonut.donut.ycA[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[15]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net502),
    .D(_00483_),
    .Q_N(_10486_),
    .Q(\vgadonut.donut.ycA[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[16]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net503),
    .D(_00484_),
    .Q_N(_10485_),
    .Q(\vgadonut.donut.ycA[16] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[17]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net504),
    .D(_00485_),
    .Q_N(_10484_),
    .Q(\vgadonut.donut.ycA[17] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[18]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net505),
    .D(_00486_),
    .Q_N(_10483_),
    .Q(\vgadonut.donut.ycA[18] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[19]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net506),
    .D(_00487_),
    .Q_N(_10482_),
    .Q(\vgadonut.donut.ycA[19] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net507),
    .D(_00488_),
    .Q_N(_10481_),
    .Q(\vgadonut.donut.ycA[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[20]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net508),
    .D(_00489_),
    .Q_N(_10480_),
    .Q(\vgadonut.donut.ycA[20] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[21]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net509),
    .D(_00490_),
    .Q_N(_10479_),
    .Q(\vgadonut.donut.ycA[21] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net510),
    .D(_00491_),
    .Q_N(_10478_),
    .Q(\vgadonut.donut.ycA[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net511),
    .D(_00492_),
    .Q_N(_00122_),
    .Q(\vgadonut.donut.ycA[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[4]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net512),
    .D(_00493_),
    .Q_N(_10477_),
    .Q(\vgadonut.donut.ycA[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net513),
    .D(_00494_),
    .Q_N(_10476_),
    .Q(\vgadonut.donut.ycA[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[6]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net514),
    .D(_00495_),
    .Q_N(_10475_),
    .Q(\vgadonut.donut.ycA[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[7]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net515),
    .D(_00496_),
    .Q_N(_10474_),
    .Q(\vgadonut.donut.ycA[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[8]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net516),
    .D(_00497_),
    .Q_N(_10473_),
    .Q(\vgadonut.donut.ycA[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ycA[9]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net517),
    .D(_00498_),
    .Q_N(_10472_),
    .Q(\vgadonut.donut.ycA[9] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net518),
    .D(_00499_),
    .Q_N(_10471_),
    .Q(\vgadonut.donut.ysA[0] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[10]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net519),
    .D(_00500_),
    .Q_N(_10470_),
    .Q(\vgadonut.donut.ysA[10] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[11]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net520),
    .D(_00501_),
    .Q_N(_10469_),
    .Q(\vgadonut.donut.ysA[11] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[12]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net521),
    .D(_00502_),
    .Q_N(_10468_),
    .Q(\vgadonut.donut.ysA[12] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[13]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net522),
    .D(_00503_),
    .Q_N(_10467_),
    .Q(\vgadonut.donut.ysA[13] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[14]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net523),
    .D(_00504_),
    .Q_N(_10466_),
    .Q(\vgadonut.donut.ysA[14] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[15]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net524),
    .D(_00505_),
    .Q_N(_10465_),
    .Q(\vgadonut.donut.ysA[15] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[16]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net525),
    .D(_00506_),
    .Q_N(_10464_),
    .Q(\vgadonut.donut.ysA[16] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[17]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net526),
    .D(_00507_),
    .Q_N(_10463_),
    .Q(\vgadonut.donut.ysA[17] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[18]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net527),
    .D(_00508_),
    .Q_N(_10462_),
    .Q(\vgadonut.donut.ysA[18] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[19]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net528),
    .D(_00509_),
    .Q_N(_10461_),
    .Q(\vgadonut.donut.ysA[19] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net529),
    .D(_00510_),
    .Q_N(_10460_),
    .Q(\vgadonut.donut.ysA[1] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[20]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net530),
    .D(_00511_),
    .Q_N(_10459_),
    .Q(\vgadonut.donut.ysA[20] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[21]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net531),
    .D(_00512_),
    .Q_N(_10458_),
    .Q(\vgadonut.donut.ysA[21] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net532),
    .D(_00513_),
    .Q_N(_10457_),
    .Q(\vgadonut.donut.ysA[2] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net533),
    .D(_00514_),
    .Q_N(_10456_),
    .Q(\vgadonut.donut.ysA[3] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[4]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net534),
    .D(_00515_),
    .Q_N(_10455_),
    .Q(\vgadonut.donut.ysA[4] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net535),
    .D(_00516_),
    .Q_N(_10454_),
    .Q(\vgadonut.donut.ysA[5] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[6]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net536),
    .D(_00517_),
    .Q_N(_10453_),
    .Q(\vgadonut.donut.ysA[6] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[7]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net537),
    .D(_00518_),
    .Q_N(_10452_),
    .Q(\vgadonut.donut.ysA[7] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[8]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net538),
    .D(_00519_),
    .Q_N(_10451_),
    .Q(\vgadonut.donut.ysA[8] ));
 sg13g2_dfrbp_1 \vgadonut.donut.ysA[9]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net539),
    .D(_00520_),
    .Q_N(_10450_),
    .Q(\vgadonut.donut.ysA[9] ));
 sg13g2_dfrbp_1 \vgadonut.frame[0]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net540),
    .D(_00521_),
    .Q_N(_00184_),
    .Q(\vgadonut.donut.frame ));
 sg13g2_dfrbp_1 \vgadonut.frame[1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net541),
    .D(_00522_),
    .Q_N(_10449_),
    .Q(\vgadonut.frame[1] ));
 sg13g2_dfrbp_1 \vgadonut.frame[2]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net542),
    .D(_00523_),
    .Q_N(_10448_),
    .Q(\vgadonut.frame[2] ));
 sg13g2_dfrbp_1 \vgadonut.frame[3]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net543),
    .D(_00524_),
    .Q_N(_10447_),
    .Q(\vgadonut.frame[3] ));
 sg13g2_dfrbp_1 \vgadonut.frame[4]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net544),
    .D(_00525_),
    .Q_N(_10446_),
    .Q(\vgadonut.frame[4] ));
 sg13g2_dfrbp_1 \vgadonut.frame[5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net545),
    .D(_00526_),
    .Q_N(_10445_),
    .Q(\vgadonut.frame[5] ));
 sg13g2_dfrbp_1 \vgadonut.frame[6]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net546),
    .D(_00527_),
    .Q_N(_10444_),
    .Q(\vgadonut.frame[6] ));
 sg13g2_dfrbp_1 \vgadonut.frame[7]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net547),
    .D(_00528_),
    .Q_N(_10443_),
    .Q(\vgadonut.frame[7] ));
 sg13g2_dfrbp_1 \vgadonut.g_out[0]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net548),
    .D(_00529_),
    .Q_N(_10442_),
    .Q(net7));
 sg13g2_dfrbp_1 \vgadonut.g_out[1]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net549),
    .D(_00530_),
    .Q_N(_10698_),
    .Q(net3));
 sg13g2_dfrbp_1 \vgadonut.h_count[0]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net272),
    .D(_00015_),
    .Q_N(_10699_),
    .Q(\vgadonut.donut.h_count[0] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[10]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net272),
    .D(_00016_),
    .Q_N(_00169_),
    .Q(\vgadonut.donut.h_count[10] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[1]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net272),
    .D(_00017_),
    .Q_N(_10700_),
    .Q(\vgadonut.donut.h_count[1] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[2]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net273),
    .D(_00018_),
    .Q_N(_00171_),
    .Q(\vgadonut.donut.h_count[2] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[3]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net273),
    .D(_00019_),
    .Q_N(_00170_),
    .Q(\vgadonut.donut.h_count[3] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[4]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net273),
    .D(_00020_),
    .Q_N(_10701_),
    .Q(\vgadonut.donut.h_count[4] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[5]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net273),
    .D(_00021_),
    .Q_N(_10702_),
    .Q(\vgadonut.donut.h_count[5] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[6]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net274),
    .D(_00022_),
    .Q_N(_10703_),
    .Q(\vgadonut.donut.h_count[6] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[7]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net274),
    .D(_00023_),
    .Q_N(_10704_),
    .Q(\vgadonut.donut.h_count[7] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[8]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net272),
    .D(_00024_),
    .Q_N(_00172_),
    .Q(\vgadonut.donut.h_count[8] ));
 sg13g2_dfrbp_1 \vgadonut.h_count[9]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net274),
    .D(_00025_),
    .Q_N(_10705_),
    .Q(\vgadonut.donut.h_count[9] ));
 sg13g2_dfrbp_1 \vgadonut.hsync$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net550),
    .D(_00026_),
    .Q_N(_10441_),
    .Q(hsync));
 sg13g2_dfrbp_1 \vgadonut.r_out[0]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net551),
    .D(_00531_),
    .Q_N(_10440_),
    .Q(net6));
 sg13g2_dfrbp_1 \vgadonut.r_out[1]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net552),
    .D(_00532_),
    .Q_N(_10439_),
    .Q(net2));
 sg13g2_dfrbp_1 \vgadonut.v_count[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net272),
    .D(_00533_),
    .Q_N(_00096_),
    .Q(\vgadonut.bayer_j[0] ));
 sg13g2_dfrbp_1 \vgadonut.v_count[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net272),
    .D(_00534_),
    .Q_N(_10438_),
    .Q(\vgadonut.bayer_j[1] ));
 sg13g2_dfrbp_1 \vgadonut.v_count[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net272),
    .D(_00535_),
    .Q_N(_10437_),
    .Q(\vgadonut.donut.v_count[2] ));
 sg13g2_dfrbp_1 \vgadonut.v_count[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net272),
    .D(_00536_),
    .Q_N(_10436_),
    .Q(\vgadonut.donut.v_count[3] ));
 sg13g2_dfrbp_1 \vgadonut.v_count[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net268),
    .D(_00537_),
    .Q_N(_10435_),
    .Q(\vgadonut.donut.v_count[4] ));
 sg13g2_dfrbp_1 \vgadonut.v_count[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net269),
    .D(_00538_),
    .Q_N(_10434_),
    .Q(\vgadonut.donut.v_count[5] ));
 sg13g2_dfrbp_1 \vgadonut.v_count[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net269),
    .D(_00539_),
    .Q_N(_10433_),
    .Q(\vgadonut.donut.v_count[6] ));
 sg13g2_dfrbp_1 \vgadonut.v_count[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net269),
    .D(_00540_),
    .Q_N(_10432_),
    .Q(\vgadonut.donut.v_count[7] ));
 sg13g2_dfrbp_1 \vgadonut.v_count[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net274),
    .D(_00541_),
    .Q_N(_10431_),
    .Q(\vgadonut.donut.v_count[8] ));
 sg13g2_dfrbp_1 \vgadonut.v_count[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net274),
    .D(_00542_),
    .Q_N(_10706_),
    .Q(\vgadonut.donut.v_count[9] ));
 sg13g2_dfrbp_1 \vgadonut.vsync$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net553),
    .D(_00027_),
    .Q_N(_10430_),
    .Q(\vgadonut.vsync ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout10 (.A(_04178_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_04354_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_04325_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_04177_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_04291_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_04176_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_04271_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_04332_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_04024_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_05355_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_04757_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_04520_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_04147_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_04138_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_04136_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_04094_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_04031_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_04519_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_04146_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_04097_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_04017_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_04391_),
    .X(net31));
 sg13g2_buf_4 fanout32 (.X(net32),
    .A(_04139_));
 sg13g2_buf_4 fanout33 (.X(net33),
    .A(_04098_));
 sg13g2_buf_2 fanout34 (.A(_04015_),
    .X(net34));
 sg13g2_buf_4 fanout35 (.X(net35),
    .A(_03962_));
 sg13g2_buf_2 fanout36 (.A(_03961_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_03960_),
    .X(net37));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(_03675_));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(_01408_));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(_03499_));
 sg13g2_buf_2 fanout41 (.A(_01603_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_01494_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_10033_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_01343_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_03792_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_03703_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_03510_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_03613_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_03509_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_03508_),
    .X(net50));
 sg13g2_buf_4 fanout51 (.X(net51),
    .A(_10032_));
 sg13g2_buf_4 fanout52 (.X(net52),
    .A(_03518_));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(_03573_));
 sg13g2_buf_2 fanout54 (.A(_09180_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_09185_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_08923_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_06908_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_06868_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_06761_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_06452_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_06228_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_06832_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_06753_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_06345_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_06227_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_06818_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_06344_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_06731_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_09115_),
    .X(net69));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(_02645_));
 sg13g2_buf_2 fanout71 (.A(_02627_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_02632_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_02594_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_06571_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_06567_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_06120_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_06722_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_00180_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_00617_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_00173_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_00014_),
    .X(net81));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_00878_));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_02391_));
 sg13g2_buf_2 fanout84 (.A(_00902_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_00858_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_00803_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_00179_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_00177_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_08168_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_07885_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_07532_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_07367_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_06991_),
    .X(net93));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(_02785_));
 sg13g2_buf_2 fanout95 (.A(_08126_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_07956_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_07401_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_07271_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_07043_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_06990_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_02471_),
    .X(net101));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(_02328_));
 sg13g2_buf_2 fanout103 (.A(_02436_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_07517_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_06981_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_10161_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_06980_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_06930_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_06918_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_04667_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_04407_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_04195_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_09659_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_09423_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_08049_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_06959_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_06945_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_06941_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_06927_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_06919_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_04741_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_04531_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_04362_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_04306_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_04303_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_04191_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_09556_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_09424_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_09422_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_09191_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_08940_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_08909_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_06900_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_06743_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_06394_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_06230_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_04305_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_04190_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_01069_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_09334_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_00765_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_00720_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_09420_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_09364_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_09130_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_07522_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_07335_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_07273_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_07236_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_07200_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_07140_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_06878_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_06763_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_06343_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_00719_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_09632_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_09546_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_09458_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_09356_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_07521_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_07499_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_07235_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_07185_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_07042_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_06983_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_06342_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_02237_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_09416_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_09365_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_06982_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_02374_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_02236_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_02172_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_02177_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_02157_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_02128_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_08917_),
    .X(net177));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(_03228_));
 sg13g2_buf_2 fanout179 (.A(_02127_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_08916_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_08912_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_06916_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_06892_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_06507_),
    .X(net184));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(_03037_));
 sg13g2_buf_2 fanout186 (.A(_02461_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_02022_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_08911_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_08586_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_06901_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_06510_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_06310_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_06275_),
    .X(net193));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(_06262_));
 sg13g2_buf_2 fanout195 (.A(_06258_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_06237_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_06030_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_06027_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_05773_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_05730_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_05694_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_05643_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_05598_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_05169_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_05135_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_05095_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_04959_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_04603_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_04534_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_04496_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_04414_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_04373_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_04312_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_02096_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_08821_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_06914_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_06419_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_06360_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_06352_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_06307_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_06291_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_06283_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_06251_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_06248_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_06247_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_06244_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_06233_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_06108_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_06054_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_06040_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_06038_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_05553_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_05505_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_05421_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_05385_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_05384_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_05381_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_05062_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_05025_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_04990_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_04944_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_04842_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_04821_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_04816_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_04602_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_04573_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_04452_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_04223_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_04203_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_04202_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_04198_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_04197_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_01956_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_09769_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_09637_),
    .X(net255));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(net258));
 sg13g2_buf_2 fanout257 (.A(net258),
    .X(net257));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(net262));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(net261));
 sg13g2_buf_2 fanout260 (.A(net261),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(net262));
 sg13g2_buf_2 fanout262 (.A(net267),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net265));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(net265));
 sg13g2_buf_2 fanout265 (.A(net267),
    .X(net265));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(net267));
 sg13g2_buf_1 fanout267 (.A(net282),
    .X(net267));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(net269));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(net270));
 sg13g2_buf_2 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(net275));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(net274));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(net275),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(net282),
    .X(net275));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(net277));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(net280));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(net279));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(net280));
 sg13g2_buf_2 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(net282),
    .X(net281));
 sg13g2_buf_1 fanout282 (.A(net1),
    .X(net282));
 sg13g2_tielo _21020__283 (.L_LO(net283));
 sg13g2_tielo _21021__284 (.L_LO(net284));
 sg13g2_tielo _21022__285 (.L_LO(net285));
 sg13g2_tielo _21023__286 (.L_LO(net286));
 sg13g2_tielo _21024__287 (.L_LO(net287));
 sg13g2_tielo _21025__288 (.L_LO(net288));
 sg13g2_tielo _21026__289 (.L_LO(net289));
 sg13g2_tielo _21027__290 (.L_LO(net290));
 sg13g2_tielo _21028__291 (.L_LO(net291));
 sg13g2_tielo _21029__292 (.L_LO(net292));
 sg13g2_tielo _21030__293 (.L_LO(net293));
 sg13g2_tielo _21031__294 (.L_LO(net294));
 sg13g2_tielo _21032__295 (.L_LO(net295));
 sg13g2_tielo _21033__296 (.L_LO(net296));
 sg13g2_tielo _21034__297 (.L_LO(net297));
 sg13g2_tielo _21035__298 (.L_LO(net298));
 sg13g2_tiehi _21001__300 (.L_HI(net300));
 sg13g2_tiehi _21002__301 (.L_HI(net301));
 sg13g2_tiehi _21003__302 (.L_HI(net302));
 sg13g2_tiehi _21004__303 (.L_HI(net303));
 sg13g2_tiehi _21005__304 (.L_HI(net304));
 sg13g2_tiehi _21006__305 (.L_HI(net305));
 sg13g2_tiehi _21007__306 (.L_HI(net306));
 sg13g2_tiehi _21008__307 (.L_HI(net307));
 sg13g2_tiehi _21009__308 (.L_HI(net308));
 sg13g2_tiehi _21010__309 (.L_HI(net309));
 sg13g2_tiehi _21011__310 (.L_HI(net310));
 sg13g2_tiehi _21012__311 (.L_HI(net311));
 sg13g2_tiehi _21013__312 (.L_HI(net312));
 sg13g2_tiehi _21014__313 (.L_HI(net313));
 sg13g2_tiehi _21015__314 (.L_HI(net314));
 sg13g2_tiehi _21016__315 (.L_HI(net315));
 sg13g2_tiehi _21017__316 (.L_HI(net316));
 sg13g2_tiehi \vgadonut.b_out[0]$_SDFF_PN0__317  (.L_HI(net317));
 sg13g2_tiehi \vgadonut.b_out[1]$_SDFF_PN0__318  (.L_HI(net318));
 sg13g2_tiehi \vgadonut.donut.donut_luma[0]$_DFFE_PP__319  (.L_HI(net319));
 sg13g2_tiehi \vgadonut.donut.donut_luma[1]$_DFFE_PP__320  (.L_HI(net320));
 sg13g2_tiehi \vgadonut.donut.donut_luma[2]$_DFFE_PP__321  (.L_HI(net321));
 sg13g2_tiehi \vgadonut.donut.donut_luma[3]$_DFFE_PP__322  (.L_HI(net322));
 sg13g2_tiehi \vgadonut.donut.donut_luma[4]$_DFFE_PP__323  (.L_HI(net323));
 sg13g2_tiehi \vgadonut.donut.donut_luma[5]$_DFFE_PP__324  (.L_HI(net324));
 sg13g2_tiehi \vgadonut.donut.donut_visible$_DFFE_PP__325  (.L_HI(net325));
 sg13g2_tiehi \vgadonut.donut.donuthit.hit$_SDFF_PP1__326  (.L_HI(net326));
 sg13g2_tiehi \vgadonut.donut.donuthit.light[10]$_DFF_P__327  (.L_HI(net327));
 sg13g2_tiehi \vgadonut.donut.donuthit.light[11]$_DFF_P__328  (.L_HI(net328));
 sg13g2_tiehi \vgadonut.donut.donuthit.light[12]$_DFF_P__329  (.L_HI(net329));
 sg13g2_tiehi \vgadonut.donut.donuthit.light[13]$_DFF_P__330  (.L_HI(net330));
 sg13g2_tiehi \vgadonut.donut.donuthit.light[8]$_DFF_P__331  (.L_HI(net331));
 sg13g2_tiehi \vgadonut.donut.donuthit.light[9]$_DFF_P__332  (.L_HI(net332));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[0]$_DFF_P__333  (.L_HI(net333));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[10]$_DFF_P__334  (.L_HI(net334));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[11]$_DFF_P__335  (.L_HI(net335));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[12]$_DFF_P__336  (.L_HI(net336));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[13]$_DFF_P__337  (.L_HI(net337));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[14]$_DFF_P__338  (.L_HI(net338));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[15]$_DFF_P__339  (.L_HI(net339));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[1]$_DFF_P__340  (.L_HI(net340));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[2]$_DFF_P__341  (.L_HI(net341));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[3]$_DFF_P__342  (.L_HI(net342));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[4]$_DFF_P__343  (.L_HI(net343));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[5]$_DFF_P__344  (.L_HI(net344));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[6]$_DFF_P__345  (.L_HI(net345));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[7]$_DFF_P__346  (.L_HI(net346));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[8]$_DFF_P__347  (.L_HI(net347));
 sg13g2_tiehi \vgadonut.donut.donuthit.px[9]$_DFF_P__348  (.L_HI(net348));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[0]$_DFF_P__349  (.L_HI(net349));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[10]$_DFF_P__350  (.L_HI(net350));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[11]$_DFF_P__351  (.L_HI(net351));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[12]$_DFF_P__352  (.L_HI(net352));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[13]$_DFF_P__353  (.L_HI(net353));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[14]$_DFF_P__354  (.L_HI(net354));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[15]$_DFF_P__355  (.L_HI(net355));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[1]$_DFF_P__356  (.L_HI(net356));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[2]$_DFF_P__357  (.L_HI(net357));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[3]$_DFF_P__358  (.L_HI(net358));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[4]$_DFF_P__359  (.L_HI(net359));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[5]$_DFF_P__360  (.L_HI(net360));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[6]$_DFF_P__361  (.L_HI(net361));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[7]$_DFF_P__362  (.L_HI(net362));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[8]$_DFF_P__363  (.L_HI(net363));
 sg13g2_tiehi \vgadonut.donut.donuthit.py[9]$_DFF_P__364  (.L_HI(net364));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[0]$_DFF_P__365  (.L_HI(net365));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[10]$_DFF_P__366  (.L_HI(net366));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[11]$_DFF_P__367  (.L_HI(net367));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[12]$_DFF_P__368  (.L_HI(net368));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[13]$_DFF_P__369  (.L_HI(net369));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[14]$_DFF_P__370  (.L_HI(net370));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[15]$_DFF_P__371  (.L_HI(net371));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[1]$_DFF_P__372  (.L_HI(net372));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[2]$_DFF_P__373  (.L_HI(net373));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[3]$_DFF_P__374  (.L_HI(net374));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[4]$_DFF_P__375  (.L_HI(net375));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[5]$_DFF_P__376  (.L_HI(net376));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[6]$_DFF_P__377  (.L_HI(net377));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[7]$_DFF_P__378  (.L_HI(net378));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[8]$_DFF_P__379  (.L_HI(net379));
 sg13g2_tiehi \vgadonut.donut.donuthit.pz[9]$_DFF_P__380  (.L_HI(net380));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[10]$_DFFE_PP__381  (.L_HI(net381));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[11]$_DFFE_PP__382  (.L_HI(net382));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[12]$_DFFE_PP__383  (.L_HI(net383));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[13]$_DFFE_PP__384  (.L_HI(net384));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[14]$_DFFE_PP__385  (.L_HI(net385));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[15]$_DFFE_PP__386  (.L_HI(net386));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[5]$_DFFE_PP__387  (.L_HI(net387));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[6]$_DFFE_PP__388  (.L_HI(net388));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[7]$_DFFE_PP__389  (.L_HI(net389));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[8]$_DFFE_PP__390  (.L_HI(net390));
 sg13g2_tiehi \vgadonut.donut.donuthit.rx[9]$_DFFE_PP__391  (.L_HI(net391));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[10]$_DFFE_PP__392  (.L_HI(net392));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[11]$_DFFE_PP__393  (.L_HI(net393));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[12]$_DFFE_PP__394  (.L_HI(net394));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[13]$_DFFE_PP__395  (.L_HI(net395));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[14]$_DFFE_PP__396  (.L_HI(net396));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[15]$_DFFE_PP__397  (.L_HI(net397));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[5]$_DFFE_PP__398  (.L_HI(net398));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[6]$_DFFE_PP__399  (.L_HI(net399));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[7]$_DFFE_PP__400  (.L_HI(net400));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[8]$_DFFE_PP__401  (.L_HI(net401));
 sg13g2_tiehi \vgadonut.donut.donuthit.ry[9]$_DFFE_PP__402  (.L_HI(net402));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[10]$_DFFE_PP__403  (.L_HI(net403));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[11]$_DFFE_PP__404  (.L_HI(net404));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[12]$_DFFE_PP__405  (.L_HI(net405));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[13]$_DFFE_PP__406  (.L_HI(net406));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[14]$_DFFE_PP__407  (.L_HI(net407));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[15]$_DFFE_PP__408  (.L_HI(net408));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[5]$_DFFE_PP__409  (.L_HI(net409));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[6]$_DFFE_PP__410  (.L_HI(net410));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[7]$_DFFE_PP__411  (.L_HI(net411));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[8]$_DFFE_PP__412  (.L_HI(net412));
 sg13g2_tiehi \vgadonut.donut.donuthit.rz[9]$_DFFE_PP__413  (.L_HI(net413));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[0]$_SDFF_PP0__414  (.L_HI(net414));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[10]$_SDFF_PP0__415  (.L_HI(net415));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[11]$_SDFF_PP0__416  (.L_HI(net416));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[12]$_SDFF_PP0__417  (.L_HI(net417));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[13]$_SDFF_PP0__418  (.L_HI(net418));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[14]$_SDFF_PP0__419  (.L_HI(net419));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[15]$_SDFF_PP0__420  (.L_HI(net420));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[1]$_SDFF_PP0__421  (.L_HI(net421));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[2]$_SDFF_PP0__422  (.L_HI(net422));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[3]$_SDFF_PP0__423  (.L_HI(net423));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[4]$_SDFF_PP0__424  (.L_HI(net424));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[5]$_SDFF_PP0__425  (.L_HI(net425));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[6]$_SDFF_PP0__426  (.L_HI(net426));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[7]$_SDFF_PP0__427  (.L_HI(net427));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[8]$_SDFF_PP0__428  (.L_HI(net428));
 sg13g2_tiehi \vgadonut.donut.donuthit.t[9]$_SDFF_PP1__429  (.L_HI(net429));
 sg13g2_tiehi \vgadonut.donut.rx6[0]$_SDFFCE_PP0P__430  (.L_HI(net430));
 sg13g2_tiehi \vgadonut.donut.rx6[10]$_DFFE_PP__431  (.L_HI(net431));
 sg13g2_tiehi \vgadonut.donut.rx6[11]$_DFFE_PP__432  (.L_HI(net432));
 sg13g2_tiehi \vgadonut.donut.rx6[12]$_DFFE_PP__433  (.L_HI(net433));
 sg13g2_tiehi \vgadonut.donut.rx6[13]$_DFFE_PP__434  (.L_HI(net434));
 sg13g2_tiehi \vgadonut.donut.rx6[14]$_DFFE_PP__435  (.L_HI(net435));
 sg13g2_tiehi \vgadonut.donut.rx6[15]$_DFFE_PP__436  (.L_HI(net436));
 sg13g2_tiehi \vgadonut.donut.rx6[16]$_DFFE_PP__437  (.L_HI(net437));
 sg13g2_tiehi \vgadonut.donut.rx6[17]$_DFFE_PP__438  (.L_HI(net438));
 sg13g2_tiehi \vgadonut.donut.rx6[18]$_DFFE_PP__439  (.L_HI(net439));
 sg13g2_tiehi \vgadonut.donut.rx6[19]$_DFFE_PP__440  (.L_HI(net440));
 sg13g2_tiehi \vgadonut.donut.rx6[1]$_SDFFCE_PP0P__441  (.L_HI(net441));
 sg13g2_tiehi \vgadonut.donut.rx6[20]$_DFFE_PP__442  (.L_HI(net442));
 sg13g2_tiehi \vgadonut.donut.rx6[21]$_DFFE_PP__443  (.L_HI(net443));
 sg13g2_tiehi \vgadonut.donut.rx6[2]$_DFFE_PP__444  (.L_HI(net444));
 sg13g2_tiehi \vgadonut.donut.rx6[3]$_DFFE_PP__445  (.L_HI(net445));
 sg13g2_tiehi \vgadonut.donut.rx6[4]$_DFFE_PP__446  (.L_HI(net446));
 sg13g2_tiehi \vgadonut.donut.rx6[5]$_DFFE_PP__447  (.L_HI(net447));
 sg13g2_tiehi \vgadonut.donut.rx6[6]$_DFFE_PP__448  (.L_HI(net448));
 sg13g2_tiehi \vgadonut.donut.rx6[7]$_DFFE_PP__449  (.L_HI(net449));
 sg13g2_tiehi \vgadonut.donut.rx6[8]$_DFFE_PP__450  (.L_HI(net450));
 sg13g2_tiehi \vgadonut.donut.rx6[9]$_DFFE_PP__451  (.L_HI(net451));
 sg13g2_tiehi \vgadonut.donut.ry6[0]$_DFFE_PP__452  (.L_HI(net452));
 sg13g2_tiehi \vgadonut.donut.ry6[10]$_DFFE_PP__453  (.L_HI(net453));
 sg13g2_tiehi \vgadonut.donut.ry6[11]$_DFFE_PP__454  (.L_HI(net454));
 sg13g2_tiehi \vgadonut.donut.ry6[12]$_DFFE_PP__455  (.L_HI(net455));
 sg13g2_tiehi \vgadonut.donut.ry6[13]$_DFFE_PP__456  (.L_HI(net456));
 sg13g2_tiehi \vgadonut.donut.ry6[14]$_DFFE_PP__457  (.L_HI(net457));
 sg13g2_tiehi \vgadonut.donut.ry6[15]$_DFFE_PP__458  (.L_HI(net458));
 sg13g2_tiehi \vgadonut.donut.ry6[16]$_DFFE_PP__459  (.L_HI(net459));
 sg13g2_tiehi \vgadonut.donut.ry6[17]$_DFFE_PP__460  (.L_HI(net460));
 sg13g2_tiehi \vgadonut.donut.ry6[18]$_DFFE_PP__461  (.L_HI(net461));
 sg13g2_tiehi \vgadonut.donut.ry6[19]$_DFFE_PP__462  (.L_HI(net462));
 sg13g2_tiehi \vgadonut.donut.ry6[1]$_DFFE_PP__463  (.L_HI(net463));
 sg13g2_tiehi \vgadonut.donut.ry6[20]$_DFFE_PP__464  (.L_HI(net464));
 sg13g2_tiehi \vgadonut.donut.ry6[21]$_DFFE_PP__465  (.L_HI(net465));
 sg13g2_tiehi \vgadonut.donut.ry6[2]$_DFFE_PP__466  (.L_HI(net466));
 sg13g2_tiehi \vgadonut.donut.ry6[3]$_DFFE_PP__467  (.L_HI(net467));
 sg13g2_tiehi \vgadonut.donut.ry6[4]$_DFFE_PP__468  (.L_HI(net468));
 sg13g2_tiehi \vgadonut.donut.ry6[5]$_DFFE_PP__469  (.L_HI(net469));
 sg13g2_tiehi \vgadonut.donut.ry6[6]$_DFFE_PP__470  (.L_HI(net470));
 sg13g2_tiehi \vgadonut.donut.ry6[7]$_DFFE_PP__471  (.L_HI(net471));
 sg13g2_tiehi \vgadonut.donut.ry6[8]$_DFFE_PP__472  (.L_HI(net472));
 sg13g2_tiehi \vgadonut.donut.ry6[9]$_DFFE_PP__473  (.L_HI(net473));
 sg13g2_tiehi \vgadonut.donut.rz6[0]$_DFFE_PP__474  (.L_HI(net474));
 sg13g2_tiehi \vgadonut.donut.rz6[10]$_DFFE_PP__475  (.L_HI(net475));
 sg13g2_tiehi \vgadonut.donut.rz6[11]$_DFFE_PP__476  (.L_HI(net476));
 sg13g2_tiehi \vgadonut.donut.rz6[12]$_DFFE_PP__477  (.L_HI(net477));
 sg13g2_tiehi \vgadonut.donut.rz6[13]$_DFFE_PP__478  (.L_HI(net478));
 sg13g2_tiehi \vgadonut.donut.rz6[14]$_DFFE_PP__479  (.L_HI(net479));
 sg13g2_tiehi \vgadonut.donut.rz6[15]$_DFFE_PP__480  (.L_HI(net480));
 sg13g2_tiehi \vgadonut.donut.rz6[16]$_DFFE_PP__481  (.L_HI(net481));
 sg13g2_tiehi \vgadonut.donut.rz6[17]$_DFFE_PP__482  (.L_HI(net482));
 sg13g2_tiehi \vgadonut.donut.rz6[18]$_DFFE_PP__483  (.L_HI(net483));
 sg13g2_tiehi \vgadonut.donut.rz6[19]$_DFFE_PP__484  (.L_HI(net484));
 sg13g2_tiehi \vgadonut.donut.rz6[1]$_DFFE_PP__485  (.L_HI(net485));
 sg13g2_tiehi \vgadonut.donut.rz6[20]$_DFFE_PP__486  (.L_HI(net486));
 sg13g2_tiehi \vgadonut.donut.rz6[21]$_DFFE_PP__487  (.L_HI(net487));
 sg13g2_tiehi \vgadonut.donut.rz6[2]$_DFFE_PP__488  (.L_HI(net488));
 sg13g2_tiehi \vgadonut.donut.rz6[3]$_DFFE_PP__489  (.L_HI(net489));
 sg13g2_tiehi \vgadonut.donut.rz6[4]$_DFFE_PP__490  (.L_HI(net490));
 sg13g2_tiehi \vgadonut.donut.rz6[5]$_DFFE_PP__491  (.L_HI(net491));
 sg13g2_tiehi \vgadonut.donut.rz6[6]$_DFFE_PP__492  (.L_HI(net492));
 sg13g2_tiehi \vgadonut.donut.rz6[7]$_DFFE_PP__493  (.L_HI(net493));
 sg13g2_tiehi \vgadonut.donut.rz6[8]$_DFFE_PP__494  (.L_HI(net494));
 sg13g2_tiehi \vgadonut.donut.rz6[9]$_DFFE_PP__495  (.L_HI(net495));
 sg13g2_tiehi \vgadonut.donut.ycA[0]$_SDFFCE_PP0P__496  (.L_HI(net496));
 sg13g2_tiehi \vgadonut.donut.ycA[10]$_DFFE_PP__497  (.L_HI(net497));
 sg13g2_tiehi \vgadonut.donut.ycA[11]$_DFFE_PP__498  (.L_HI(net498));
 sg13g2_tiehi \vgadonut.donut.ycA[12]$_DFFE_PP__499  (.L_HI(net499));
 sg13g2_tiehi \vgadonut.donut.ycA[13]$_DFFE_PP__500  (.L_HI(net500));
 sg13g2_tiehi \vgadonut.donut.ycA[14]$_DFFE_PP__501  (.L_HI(net501));
 sg13g2_tiehi \vgadonut.donut.ycA[15]$_DFFE_PP__502  (.L_HI(net502));
 sg13g2_tiehi \vgadonut.donut.ycA[16]$_DFFE_PP__503  (.L_HI(net503));
 sg13g2_tiehi \vgadonut.donut.ycA[17]$_DFFE_PP__504  (.L_HI(net504));
 sg13g2_tiehi \vgadonut.donut.ycA[18]$_DFFE_PP__505  (.L_HI(net505));
 sg13g2_tiehi \vgadonut.donut.ycA[19]$_DFFE_PP__506  (.L_HI(net506));
 sg13g2_tiehi \vgadonut.donut.ycA[1]$_SDFFCE_PP0P__507  (.L_HI(net507));
 sg13g2_tiehi \vgadonut.donut.ycA[20]$_DFFE_PP__508  (.L_HI(net508));
 sg13g2_tiehi \vgadonut.donut.ycA[21]$_DFFE_PP__509  (.L_HI(net509));
 sg13g2_tiehi \vgadonut.donut.ycA[2]$_SDFFCE_PP0P__510  (.L_HI(net510));
 sg13g2_tiehi \vgadonut.donut.ycA[3]$_SDFFCE_PP0P__511  (.L_HI(net511));
 sg13g2_tiehi \vgadonut.donut.ycA[4]$_DFFE_PP__512  (.L_HI(net512));
 sg13g2_tiehi \vgadonut.donut.ycA[5]$_DFFE_PP__513  (.L_HI(net513));
 sg13g2_tiehi \vgadonut.donut.ycA[6]$_DFFE_PP__514  (.L_HI(net514));
 sg13g2_tiehi \vgadonut.donut.ycA[7]$_DFFE_PP__515  (.L_HI(net515));
 sg13g2_tiehi \vgadonut.donut.ycA[8]$_DFFE_PP__516  (.L_HI(net516));
 sg13g2_tiehi \vgadonut.donut.ycA[9]$_DFFE_PP__517  (.L_HI(net517));
 sg13g2_tiehi \vgadonut.donut.ysA[0]$_SDFFCE_PP0P__518  (.L_HI(net518));
 sg13g2_tiehi \vgadonut.donut.ysA[10]$_DFFE_PP__519  (.L_HI(net519));
 sg13g2_tiehi \vgadonut.donut.ysA[11]$_DFFE_PP__520  (.L_HI(net520));
 sg13g2_tiehi \vgadonut.donut.ysA[12]$_DFFE_PP__521  (.L_HI(net521));
 sg13g2_tiehi \vgadonut.donut.ysA[13]$_DFFE_PP__522  (.L_HI(net522));
 sg13g2_tiehi \vgadonut.donut.ysA[14]$_DFFE_PP__523  (.L_HI(net523));
 sg13g2_tiehi \vgadonut.donut.ysA[15]$_DFFE_PP__524  (.L_HI(net524));
 sg13g2_tiehi \vgadonut.donut.ysA[16]$_DFFE_PP__525  (.L_HI(net525));
 sg13g2_tiehi \vgadonut.donut.ysA[17]$_DFFE_PP__526  (.L_HI(net526));
 sg13g2_tiehi \vgadonut.donut.ysA[18]$_DFFE_PP__527  (.L_HI(net527));
 sg13g2_tiehi \vgadonut.donut.ysA[19]$_DFFE_PP__528  (.L_HI(net528));
 sg13g2_tiehi \vgadonut.donut.ysA[1]$_SDFFCE_PP0P__529  (.L_HI(net529));
 sg13g2_tiehi \vgadonut.donut.ysA[20]$_DFFE_PP__530  (.L_HI(net530));
 sg13g2_tiehi \vgadonut.donut.ysA[21]$_DFFE_PP__531  (.L_HI(net531));
 sg13g2_tiehi \vgadonut.donut.ysA[2]$_SDFFCE_PP0P__532  (.L_HI(net532));
 sg13g2_tiehi \vgadonut.donut.ysA[3]$_SDFFCE_PP0P__533  (.L_HI(net533));
 sg13g2_tiehi \vgadonut.donut.ysA[4]$_DFFE_PP__534  (.L_HI(net534));
 sg13g2_tiehi \vgadonut.donut.ysA[5]$_DFFE_PP__535  (.L_HI(net535));
 sg13g2_tiehi \vgadonut.donut.ysA[6]$_DFFE_PP__536  (.L_HI(net536));
 sg13g2_tiehi \vgadonut.donut.ysA[7]$_DFFE_PP__537  (.L_HI(net537));
 sg13g2_tiehi \vgadonut.donut.ysA[8]$_DFFE_PP__538  (.L_HI(net538));
 sg13g2_tiehi \vgadonut.donut.ysA[9]$_DFFE_PP__539  (.L_HI(net539));
 sg13g2_tiehi \vgadonut.frame[0]$_DFFE_PP__540  (.L_HI(net540));
 sg13g2_tiehi \vgadonut.frame[1]$_DFFE_PP__541  (.L_HI(net541));
 sg13g2_tiehi \vgadonut.frame[2]$_DFFE_PP__542  (.L_HI(net542));
 sg13g2_tiehi \vgadonut.frame[3]$_DFFE_PP__543  (.L_HI(net543));
 sg13g2_tiehi \vgadonut.frame[4]$_DFFE_PP__544  (.L_HI(net544));
 sg13g2_tiehi \vgadonut.frame[5]$_DFFE_PP__545  (.L_HI(net545));
 sg13g2_tiehi \vgadonut.frame[6]$_DFFE_PP__546  (.L_HI(net546));
 sg13g2_tiehi \vgadonut.frame[7]$_DFFE_PP__547  (.L_HI(net547));
 sg13g2_tiehi \vgadonut.g_out[0]$_SDFF_PN0__548  (.L_HI(net548));
 sg13g2_tiehi \vgadonut.g_out[1]$_SDFF_PN0__549  (.L_HI(net549));
 sg13g2_tiehi \vgadonut.hsync$_DFF_P__550  (.L_HI(net550));
 sg13g2_tiehi \vgadonut.r_out[0]$_SDFF_PN0__551  (.L_HI(net551));
 sg13g2_tiehi \vgadonut.r_out[1]$_SDFF_PN0__552  (.L_HI(net552));
 sg13g2_tiehi \vgadonut.vsync$_DFF_P__553  (.L_HI(net553));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_62_clk (.X(clknet_leaf_62_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_63_clk (.X(clknet_leaf_63_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_64_clk (.X(clknet_leaf_64_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_65_clk (.X(clknet_leaf_65_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_66_clk (.X(clknet_leaf_66_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_67_clk (.X(clknet_leaf_67_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_68_clk (.X(clknet_leaf_68_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_69_clk (.X(clknet_leaf_69_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkload6 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkload8 (.A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkload9 (.A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_67_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_leaf_68_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_69_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_4_clk));
 sg13g2_buf_16 clkload15 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_63_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_65_clk));
 sg13g2_buf_8 clkload18 (.A(clknet_leaf_66_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_leaf_59_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_leaf_60_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_61_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_5_clk));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_15_clk));
 sg13g2_buf_16 clkload25 (.A(clknet_leaf_17_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_21_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_34_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_9_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_10_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_20_clk));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_53_clk));
 sg13g2_inv_2 clkload33 (.A(clknet_leaf_54_clk));
 sg13g2_buf_8 clkload34 (.A(clknet_leaf_55_clk));
 sg13g2_inv_4 clkload35 (.A(clknet_leaf_56_clk));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_57_clk));
 sg13g2_buf_16 clkload37 (.A(clknet_leaf_58_clk));
 sg13g2_buf_16 clkload38 (.A(clknet_leaf_46_clk));
 sg13g2_buf_16 clkload39 (.A(clknet_leaf_48_clk));
 sg13g2_inv_1 clkload40 (.A(clknet_leaf_50_clk));
 sg13g2_buf_8 clkload41 (.A(clknet_leaf_38_clk));
 sg13g2_buf_16 clkload42 (.A(clknet_leaf_44_clk));
 sg13g2_inv_2 clkload43 (.A(clknet_leaf_45_clk));
 sg13g2_buf_16 clkload44 (.A(clknet_leaf_30_clk));
 sg13g2_inv_4 clkload45 (.A(clknet_leaf_33_clk));
 sg13g2_buf_8 clkload46 (.A(clknet_leaf_23_clk));
 sg13g2_inv_4 clkload47 (.A(clknet_leaf_25_clk));
 sg13g2_inv_4 clkload48 (.A(clknet_leaf_32_clk));
 sg13g2_buf_16 clkload49 (.A(clknet_leaf_40_clk));
 sg13g2_inv_4 clkload50 (.A(clknet_leaf_41_clk));
 sg13g2_inv_2 clkload51 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload52 (.A(clknet_leaf_29_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00530_));
 sg13g2_antennanp ANTENNA_2 (.A(_03792_));
 sg13g2_antennanp ANTENNA_3 (.A(_03792_));
 sg13g2_antennanp ANTENNA_4 (.A(_03792_));
 sg13g2_antennanp ANTENNA_5 (.A(_03792_));
 sg13g2_antennanp ANTENNA_6 (.A(_06224_));
 sg13g2_antennanp ANTENNA_7 (.A(_06224_));
 sg13g2_antennanp ANTENNA_8 (.A(_03792_));
 sg13g2_antennanp ANTENNA_9 (.A(_03792_));
 sg13g2_antennanp ANTENNA_10 (.A(_03792_));
 sg13g2_antennanp ANTENNA_11 (.A(_03792_));
 sg13g2_antennanp ANTENNA_12 (.A(_06224_));
 sg13g2_antennanp ANTENNA_13 (.A(_06224_));
 sg13g2_antennanp ANTENNA_14 (.A(_03792_));
 sg13g2_antennanp ANTENNA_15 (.A(_03792_));
 sg13g2_antennanp ANTENNA_16 (.A(_03792_));
 sg13g2_antennanp ANTENNA_17 (.A(_03792_));
 sg13g2_antennanp ANTENNA_18 (.A(_06224_));
 sg13g2_antennanp ANTENNA_19 (.A(_06224_));
 sg13g2_antennanp ANTENNA_20 (.A(_03792_));
 sg13g2_antennanp ANTENNA_21 (.A(_03792_));
 sg13g2_antennanp ANTENNA_22 (.A(_03792_));
 sg13g2_antennanp ANTENNA_23 (.A(_03792_));
 sg13g2_antennanp ANTENNA_24 (.A(_06224_));
 sg13g2_antennanp ANTENNA_25 (.A(_06224_));
 sg13g2_antennanp ANTENNA_26 (.A(_03792_));
 sg13g2_antennanp ANTENNA_27 (.A(_03792_));
 sg13g2_antennanp ANTENNA_28 (.A(_03792_));
 sg13g2_antennanp ANTENNA_29 (.A(_03792_));
 sg13g2_antennanp ANTENNA_30 (.A(_06224_));
 sg13g2_antennanp ANTENNA_31 (.A(_06224_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_4 FILLER_0_14 ();
 sg13g2_fill_2 FILLER_0_78 ();
 sg13g2_decap_4 FILLER_0_144 ();
 sg13g2_fill_2 FILLER_0_251 ();
 sg13g2_fill_1 FILLER_0_253 ();
 sg13g2_decap_4 FILLER_0_305 ();
 sg13g2_fill_2 FILLER_0_309 ();
 sg13g2_fill_1 FILLER_0_320 ();
 sg13g2_fill_1 FILLER_0_345 ();
 sg13g2_fill_2 FILLER_0_351 ();
 sg13g2_decap_4 FILLER_0_362 ();
 sg13g2_fill_1 FILLER_0_366 ();
 sg13g2_decap_4 FILLER_0_452 ();
 sg13g2_fill_1 FILLER_0_456 ();
 sg13g2_fill_2 FILLER_0_486 ();
 sg13g2_fill_1 FILLER_0_488 ();
 sg13g2_fill_2 FILLER_0_581 ();
 sg13g2_fill_1 FILLER_0_672 ();
 sg13g2_fill_2 FILLER_0_712 ();
 sg13g2_fill_2 FILLER_0_743 ();
 sg13g2_fill_2 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_772 ();
 sg13g2_decap_8 FILLER_0_779 ();
 sg13g2_decap_8 FILLER_0_786 ();
 sg13g2_decap_8 FILLER_0_793 ();
 sg13g2_decap_8 FILLER_0_800 ();
 sg13g2_decap_8 FILLER_0_807 ();
 sg13g2_decap_8 FILLER_0_814 ();
 sg13g2_decap_8 FILLER_0_821 ();
 sg13g2_decap_8 FILLER_0_828 ();
 sg13g2_decap_8 FILLER_0_835 ();
 sg13g2_decap_8 FILLER_0_842 ();
 sg13g2_decap_8 FILLER_0_849 ();
 sg13g2_decap_8 FILLER_0_856 ();
 sg13g2_decap_8 FILLER_0_863 ();
 sg13g2_decap_8 FILLER_0_870 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_7 ();
 sg13g2_fill_1 FILLER_1_62 ();
 sg13g2_fill_2 FILLER_1_66 ();
 sg13g2_fill_1 FILLER_1_92 ();
 sg13g2_fill_1 FILLER_1_122 ();
 sg13g2_fill_1 FILLER_1_127 ();
 sg13g2_fill_2 FILLER_1_211 ();
 sg13g2_fill_2 FILLER_1_217 ();
 sg13g2_fill_1 FILLER_1_270 ();
 sg13g2_fill_1 FILLER_1_292 ();
 sg13g2_fill_1 FILLER_1_300 ();
 sg13g2_fill_1 FILLER_1_309 ();
 sg13g2_fill_1 FILLER_1_340 ();
 sg13g2_fill_2 FILLER_1_345 ();
 sg13g2_fill_2 FILLER_1_480 ();
 sg13g2_fill_1 FILLER_1_513 ();
 sg13g2_fill_1 FILLER_1_577 ();
 sg13g2_fill_2 FILLER_1_586 ();
 sg13g2_fill_1 FILLER_1_656 ();
 sg13g2_decap_4 FILLER_1_771 ();
 sg13g2_fill_1 FILLER_1_775 ();
 sg13g2_fill_1 FILLER_1_795 ();
 sg13g2_fill_1 FILLER_1_800 ();
 sg13g2_decap_8 FILLER_1_810 ();
 sg13g2_decap_8 FILLER_1_817 ();
 sg13g2_decap_8 FILLER_1_824 ();
 sg13g2_decap_8 FILLER_1_831 ();
 sg13g2_decap_8 FILLER_1_838 ();
 sg13g2_decap_8 FILLER_1_845 ();
 sg13g2_decap_8 FILLER_1_852 ();
 sg13g2_decap_8 FILLER_1_859 ();
 sg13g2_decap_8 FILLER_1_866 ();
 sg13g2_decap_4 FILLER_1_873 ();
 sg13g2_fill_1 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_1 FILLER_2_45 ();
 sg13g2_fill_2 FILLER_2_66 ();
 sg13g2_fill_2 FILLER_2_97 ();
 sg13g2_fill_1 FILLER_2_103 ();
 sg13g2_fill_1 FILLER_2_131 ();
 sg13g2_fill_2 FILLER_2_174 ();
 sg13g2_fill_2 FILLER_2_184 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_fill_1 FILLER_2_219 ();
 sg13g2_fill_2 FILLER_2_240 ();
 sg13g2_fill_2 FILLER_2_281 ();
 sg13g2_fill_1 FILLER_2_283 ();
 sg13g2_decap_4 FILLER_2_287 ();
 sg13g2_fill_1 FILLER_2_291 ();
 sg13g2_fill_1 FILLER_2_329 ();
 sg13g2_fill_1 FILLER_2_356 ();
 sg13g2_fill_1 FILLER_2_365 ();
 sg13g2_fill_1 FILLER_2_371 ();
 sg13g2_fill_1 FILLER_2_381 ();
 sg13g2_fill_1 FILLER_2_399 ();
 sg13g2_fill_1 FILLER_2_405 ();
 sg13g2_fill_1 FILLER_2_411 ();
 sg13g2_fill_2 FILLER_2_430 ();
 sg13g2_fill_2 FILLER_2_448 ();
 sg13g2_decap_4 FILLER_2_455 ();
 sg13g2_fill_1 FILLER_2_521 ();
 sg13g2_fill_1 FILLER_2_540 ();
 sg13g2_fill_1 FILLER_2_549 ();
 sg13g2_fill_1 FILLER_2_648 ();
 sg13g2_fill_1 FILLER_2_667 ();
 sg13g2_fill_1 FILLER_2_718 ();
 sg13g2_fill_1 FILLER_2_723 ();
 sg13g2_fill_2 FILLER_2_754 ();
 sg13g2_fill_2 FILLER_2_773 ();
 sg13g2_fill_2 FILLER_2_779 ();
 sg13g2_fill_2 FILLER_2_784 ();
 sg13g2_fill_1 FILLER_2_786 ();
 sg13g2_fill_2 FILLER_2_790 ();
 sg13g2_decap_4 FILLER_2_821 ();
 sg13g2_fill_2 FILLER_2_825 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_4 FILLER_2_872 ();
 sg13g2_fill_2 FILLER_2_876 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_11 ();
 sg13g2_fill_1 FILLER_3_13 ();
 sg13g2_fill_1 FILLER_3_44 ();
 sg13g2_fill_1 FILLER_3_102 ();
 sg13g2_fill_1 FILLER_3_112 ();
 sg13g2_fill_2 FILLER_3_138 ();
 sg13g2_fill_1 FILLER_3_145 ();
 sg13g2_fill_1 FILLER_3_172 ();
 sg13g2_fill_2 FILLER_3_199 ();
 sg13g2_fill_2 FILLER_3_228 ();
 sg13g2_fill_1 FILLER_3_407 ();
 sg13g2_fill_2 FILLER_3_438 ();
 sg13g2_fill_1 FILLER_3_448 ();
 sg13g2_fill_2 FILLER_3_454 ();
 sg13g2_fill_2 FILLER_3_487 ();
 sg13g2_fill_1 FILLER_3_505 ();
 sg13g2_fill_1 FILLER_3_525 ();
 sg13g2_fill_1 FILLER_3_557 ();
 sg13g2_fill_2 FILLER_3_562 ();
 sg13g2_fill_1 FILLER_3_568 ();
 sg13g2_fill_1 FILLER_3_577 ();
 sg13g2_fill_1 FILLER_3_583 ();
 sg13g2_fill_1 FILLER_3_590 ();
 sg13g2_fill_1 FILLER_3_595 ();
 sg13g2_fill_1 FILLER_3_633 ();
 sg13g2_fill_1 FILLER_3_647 ();
 sg13g2_fill_2 FILLER_3_723 ();
 sg13g2_fill_2 FILLER_3_743 ();
 sg13g2_fill_1 FILLER_3_768 ();
 sg13g2_fill_1 FILLER_3_789 ();
 sg13g2_fill_1 FILLER_3_828 ();
 sg13g2_fill_2 FILLER_3_833 ();
 sg13g2_fill_2 FILLER_3_842 ();
 sg13g2_fill_1 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_851 ();
 sg13g2_decap_8 FILLER_3_858 ();
 sg13g2_decap_8 FILLER_3_865 ();
 sg13g2_decap_4 FILLER_3_872 ();
 sg13g2_fill_2 FILLER_3_876 ();
 sg13g2_fill_1 FILLER_4_50 ();
 sg13g2_fill_1 FILLER_4_77 ();
 sg13g2_fill_1 FILLER_4_107 ();
 sg13g2_fill_2 FILLER_4_129 ();
 sg13g2_fill_2 FILLER_4_135 ();
 sg13g2_fill_1 FILLER_4_145 ();
 sg13g2_fill_1 FILLER_4_151 ();
 sg13g2_fill_1 FILLER_4_156 ();
 sg13g2_fill_2 FILLER_4_162 ();
 sg13g2_fill_1 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_177 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_fill_2 FILLER_4_228 ();
 sg13g2_fill_1 FILLER_4_230 ();
 sg13g2_fill_1 FILLER_4_256 ();
 sg13g2_fill_1 FILLER_4_267 ();
 sg13g2_fill_2 FILLER_4_291 ();
 sg13g2_fill_1 FILLER_4_293 ();
 sg13g2_decap_4 FILLER_4_302 ();
 sg13g2_decap_4 FILLER_4_311 ();
 sg13g2_fill_1 FILLER_4_315 ();
 sg13g2_fill_2 FILLER_4_324 ();
 sg13g2_fill_1 FILLER_4_344 ();
 sg13g2_fill_1 FILLER_4_357 ();
 sg13g2_fill_2 FILLER_4_374 ();
 sg13g2_fill_1 FILLER_4_426 ();
 sg13g2_fill_2 FILLER_4_441 ();
 sg13g2_fill_1 FILLER_4_443 ();
 sg13g2_fill_1 FILLER_4_490 ();
 sg13g2_fill_1 FILLER_4_558 ();
 sg13g2_fill_1 FILLER_4_589 ();
 sg13g2_fill_1 FILLER_4_595 ();
 sg13g2_fill_1 FILLER_4_600 ();
 sg13g2_fill_1 FILLER_4_656 ();
 sg13g2_fill_2 FILLER_4_710 ();
 sg13g2_fill_1 FILLER_4_716 ();
 sg13g2_fill_1 FILLER_4_721 ();
 sg13g2_fill_1 FILLER_4_761 ();
 sg13g2_fill_2 FILLER_4_794 ();
 sg13g2_fill_1 FILLER_4_801 ();
 sg13g2_fill_1 FILLER_4_852 ();
 sg13g2_decap_8 FILLER_4_866 ();
 sg13g2_fill_2 FILLER_4_876 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_49 ();
 sg13g2_fill_2 FILLER_5_58 ();
 sg13g2_fill_1 FILLER_5_68 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_fill_2 FILLER_5_133 ();
 sg13g2_fill_1 FILLER_5_189 ();
 sg13g2_fill_1 FILLER_5_198 ();
 sg13g2_fill_1 FILLER_5_207 ();
 sg13g2_fill_1 FILLER_5_213 ();
 sg13g2_fill_1 FILLER_5_219 ();
 sg13g2_fill_2 FILLER_5_224 ();
 sg13g2_fill_1 FILLER_5_231 ();
 sg13g2_fill_2 FILLER_5_340 ();
 sg13g2_fill_1 FILLER_5_342 ();
 sg13g2_fill_1 FILLER_5_367 ();
 sg13g2_fill_1 FILLER_5_372 ();
 sg13g2_fill_1 FILLER_5_381 ();
 sg13g2_fill_1 FILLER_5_387 ();
 sg13g2_fill_2 FILLER_5_439 ();
 sg13g2_fill_1 FILLER_5_450 ();
 sg13g2_fill_1 FILLER_5_493 ();
 sg13g2_fill_1 FILLER_5_498 ();
 sg13g2_fill_1 FILLER_5_503 ();
 sg13g2_fill_1 FILLER_5_508 ();
 sg13g2_fill_1 FILLER_5_530 ();
 sg13g2_fill_1 FILLER_5_738 ();
 sg13g2_fill_1 FILLER_5_747 ();
 sg13g2_fill_2 FILLER_5_760 ();
 sg13g2_fill_1 FILLER_5_762 ();
 sg13g2_fill_1 FILLER_5_787 ();
 sg13g2_fill_1 FILLER_5_796 ();
 sg13g2_fill_1 FILLER_6_79 ();
 sg13g2_fill_2 FILLER_6_88 ();
 sg13g2_fill_2 FILLER_6_121 ();
 sg13g2_fill_1 FILLER_6_160 ();
 sg13g2_fill_2 FILLER_6_165 ();
 sg13g2_fill_2 FILLER_6_184 ();
 sg13g2_fill_2 FILLER_6_264 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_fill_2 FILLER_6_291 ();
 sg13g2_fill_2 FILLER_6_346 ();
 sg13g2_fill_1 FILLER_6_394 ();
 sg13g2_fill_1 FILLER_6_412 ();
 sg13g2_fill_1 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_431 ();
 sg13g2_fill_2 FILLER_6_471 ();
 sg13g2_fill_1 FILLER_6_482 ();
 sg13g2_fill_1 FILLER_6_492 ();
 sg13g2_fill_1 FILLER_6_500 ();
 sg13g2_fill_1 FILLER_6_535 ();
 sg13g2_fill_1 FILLER_6_540 ();
 sg13g2_fill_2 FILLER_6_549 ();
 sg13g2_fill_2 FILLER_6_584 ();
 sg13g2_fill_1 FILLER_6_602 ();
 sg13g2_fill_1 FILLER_6_634 ();
 sg13g2_fill_1 FILLER_6_669 ();
 sg13g2_fill_1 FILLER_6_695 ();
 sg13g2_fill_2 FILLER_6_727 ();
 sg13g2_fill_2 FILLER_6_768 ();
 sg13g2_fill_1 FILLER_6_778 ();
 sg13g2_fill_2 FILLER_6_804 ();
 sg13g2_fill_1 FILLER_6_825 ();
 sg13g2_fill_2 FILLER_6_876 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_8 ();
 sg13g2_fill_2 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_25 ();
 sg13g2_fill_2 FILLER_7_59 ();
 sg13g2_fill_1 FILLER_7_79 ();
 sg13g2_fill_1 FILLER_7_84 ();
 sg13g2_fill_2 FILLER_7_104 ();
 sg13g2_fill_1 FILLER_7_128 ();
 sg13g2_fill_1 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_183 ();
 sg13g2_fill_1 FILLER_7_185 ();
 sg13g2_fill_2 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_285 ();
 sg13g2_fill_1 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_377 ();
 sg13g2_fill_2 FILLER_7_386 ();
 sg13g2_fill_1 FILLER_7_400 ();
 sg13g2_fill_1 FILLER_7_411 ();
 sg13g2_fill_1 FILLER_7_421 ();
 sg13g2_fill_1 FILLER_7_425 ();
 sg13g2_fill_2 FILLER_7_430 ();
 sg13g2_fill_1 FILLER_7_457 ();
 sg13g2_fill_1 FILLER_7_513 ();
 sg13g2_fill_2 FILLER_7_578 ();
 sg13g2_fill_2 FILLER_7_610 ();
 sg13g2_fill_1 FILLER_7_612 ();
 sg13g2_fill_1 FILLER_7_617 ();
 sg13g2_fill_1 FILLER_7_623 ();
 sg13g2_fill_1 FILLER_7_679 ();
 sg13g2_fill_1 FILLER_7_725 ();
 sg13g2_fill_2 FILLER_7_733 ();
 sg13g2_fill_1 FILLER_7_735 ();
 sg13g2_fill_2 FILLER_7_740 ();
 sg13g2_fill_1 FILLER_7_746 ();
 sg13g2_fill_1 FILLER_7_752 ();
 sg13g2_fill_1 FILLER_7_761 ();
 sg13g2_fill_1 FILLER_7_767 ();
 sg13g2_fill_1 FILLER_7_780 ();
 sg13g2_fill_1 FILLER_7_794 ();
 sg13g2_fill_1 FILLER_7_799 ();
 sg13g2_fill_1 FILLER_7_820 ();
 sg13g2_fill_2 FILLER_7_837 ();
 sg13g2_fill_2 FILLER_7_872 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_57 ();
 sg13g2_fill_1 FILLER_8_67 ();
 sg13g2_fill_1 FILLER_8_82 ();
 sg13g2_fill_1 FILLER_8_88 ();
 sg13g2_fill_1 FILLER_8_149 ();
 sg13g2_fill_2 FILLER_8_154 ();
 sg13g2_fill_1 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_178 ();
 sg13g2_fill_1 FILLER_8_219 ();
 sg13g2_fill_1 FILLER_8_230 ();
 sg13g2_fill_1 FILLER_8_236 ();
 sg13g2_fill_1 FILLER_8_241 ();
 sg13g2_fill_2 FILLER_8_250 ();
 sg13g2_fill_1 FILLER_8_257 ();
 sg13g2_fill_1 FILLER_8_263 ();
 sg13g2_fill_1 FILLER_8_306 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_fill_1 FILLER_8_328 ();
 sg13g2_fill_1 FILLER_8_362 ();
 sg13g2_fill_1 FILLER_8_403 ();
 sg13g2_fill_1 FILLER_8_479 ();
 sg13g2_fill_1 FILLER_8_517 ();
 sg13g2_fill_2 FILLER_8_531 ();
 sg13g2_fill_1 FILLER_8_614 ();
 sg13g2_fill_2 FILLER_8_639 ();
 sg13g2_fill_1 FILLER_8_687 ();
 sg13g2_fill_2 FILLER_8_696 ();
 sg13g2_fill_2 FILLER_8_763 ();
 sg13g2_fill_1 FILLER_8_765 ();
 sg13g2_fill_1 FILLER_8_779 ();
 sg13g2_fill_2 FILLER_8_815 ();
 sg13g2_fill_2 FILLER_8_839 ();
 sg13g2_fill_1 FILLER_9_21 ();
 sg13g2_fill_1 FILLER_9_44 ();
 sg13g2_fill_1 FILLER_9_50 ();
 sg13g2_fill_1 FILLER_9_60 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_fill_1 FILLER_9_114 ();
 sg13g2_fill_1 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_135 ();
 sg13g2_fill_2 FILLER_9_157 ();
 sg13g2_fill_1 FILLER_9_184 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_237 ();
 sg13g2_fill_1 FILLER_9_243 ();
 sg13g2_fill_1 FILLER_9_252 ();
 sg13g2_fill_2 FILLER_9_337 ();
 sg13g2_fill_1 FILLER_9_339 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_388 ();
 sg13g2_fill_2 FILLER_9_422 ();
 sg13g2_fill_2 FILLER_9_429 ();
 sg13g2_fill_1 FILLER_9_431 ();
 sg13g2_fill_1 FILLER_9_457 ();
 sg13g2_fill_2 FILLER_9_466 ();
 sg13g2_fill_2 FILLER_9_476 ();
 sg13g2_fill_2 FILLER_9_497 ();
 sg13g2_fill_1 FILLER_9_513 ();
 sg13g2_fill_2 FILLER_9_547 ();
 sg13g2_fill_2 FILLER_9_685 ();
 sg13g2_fill_2 FILLER_9_710 ();
 sg13g2_fill_1 FILLER_9_733 ();
 sg13g2_fill_2 FILLER_9_756 ();
 sg13g2_fill_1 FILLER_9_766 ();
 sg13g2_fill_2 FILLER_9_805 ();
 sg13g2_fill_1 FILLER_9_840 ();
 sg13g2_fill_1 FILLER_9_877 ();
 sg13g2_fill_1 FILLER_10_29 ();
 sg13g2_fill_1 FILLER_10_38 ();
 sg13g2_fill_1 FILLER_10_56 ();
 sg13g2_fill_1 FILLER_10_78 ();
 sg13g2_fill_1 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_156 ();
 sg13g2_fill_2 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_fill_1 FILLER_10_282 ();
 sg13g2_fill_2 FILLER_10_331 ();
 sg13g2_fill_1 FILLER_10_374 ();
 sg13g2_fill_1 FILLER_10_395 ();
 sg13g2_decap_4 FILLER_10_425 ();
 sg13g2_fill_1 FILLER_10_434 ();
 sg13g2_fill_1 FILLER_10_442 ();
 sg13g2_fill_2 FILLER_10_446 ();
 sg13g2_fill_1 FILLER_10_448 ();
 sg13g2_fill_1 FILLER_10_456 ();
 sg13g2_fill_1 FILLER_10_527 ();
 sg13g2_fill_1 FILLER_10_532 ();
 sg13g2_fill_2 FILLER_10_567 ();
 sg13g2_fill_1 FILLER_10_613 ();
 sg13g2_fill_2 FILLER_10_671 ();
 sg13g2_fill_1 FILLER_10_677 ();
 sg13g2_fill_1 FILLER_10_682 ();
 sg13g2_fill_1 FILLER_10_688 ();
 sg13g2_fill_2 FILLER_10_763 ();
 sg13g2_fill_1 FILLER_10_783 ();
 sg13g2_fill_2 FILLER_10_876 ();
 sg13g2_fill_1 FILLER_11_29 ();
 sg13g2_fill_1 FILLER_11_91 ();
 sg13g2_fill_1 FILLER_11_109 ();
 sg13g2_fill_1 FILLER_11_190 ();
 sg13g2_fill_1 FILLER_11_252 ();
 sg13g2_fill_2 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_283 ();
 sg13g2_fill_2 FILLER_11_347 ();
 sg13g2_fill_1 FILLER_11_390 ();
 sg13g2_fill_1 FILLER_11_395 ();
 sg13g2_fill_2 FILLER_11_400 ();
 sg13g2_fill_1 FILLER_11_402 ();
 sg13g2_fill_1 FILLER_11_433 ();
 sg13g2_fill_2 FILLER_11_442 ();
 sg13g2_fill_1 FILLER_11_449 ();
 sg13g2_fill_1 FILLER_11_458 ();
 sg13g2_fill_2 FILLER_11_469 ();
 sg13g2_fill_2 FILLER_11_478 ();
 sg13g2_fill_1 FILLER_11_537 ();
 sg13g2_fill_2 FILLER_11_561 ();
 sg13g2_fill_1 FILLER_11_573 ();
 sg13g2_fill_1 FILLER_11_597 ();
 sg13g2_fill_1 FILLER_11_606 ();
 sg13g2_fill_1 FILLER_11_611 ();
 sg13g2_fill_1 FILLER_11_617 ();
 sg13g2_fill_2 FILLER_11_626 ();
 sg13g2_fill_1 FILLER_11_697 ();
 sg13g2_fill_1 FILLER_11_726 ();
 sg13g2_fill_2 FILLER_11_766 ();
 sg13g2_fill_1 FILLER_11_768 ();
 sg13g2_fill_1 FILLER_11_801 ();
 sg13g2_fill_2 FILLER_11_825 ();
 sg13g2_fill_1 FILLER_11_834 ();
 sg13g2_fill_1 FILLER_11_840 ();
 sg13g2_fill_2 FILLER_11_847 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_27 ();
 sg13g2_fill_1 FILLER_12_33 ();
 sg13g2_fill_1 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_75 ();
 sg13g2_fill_2 FILLER_12_113 ();
 sg13g2_fill_1 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_136 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_176 ();
 sg13g2_fill_2 FILLER_12_215 ();
 sg13g2_fill_1 FILLER_12_337 ();
 sg13g2_decap_4 FILLER_12_376 ();
 sg13g2_fill_1 FILLER_12_388 ();
 sg13g2_fill_1 FILLER_12_413 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_2 FILLER_12_444 ();
 sg13g2_fill_1 FILLER_12_446 ();
 sg13g2_fill_1 FILLER_12_461 ();
 sg13g2_fill_2 FILLER_12_467 ();
 sg13g2_fill_1 FILLER_12_484 ();
 sg13g2_fill_1 FILLER_12_507 ();
 sg13g2_fill_1 FILLER_12_548 ();
 sg13g2_fill_1 FILLER_12_558 ();
 sg13g2_fill_1 FILLER_12_577 ();
 sg13g2_fill_2 FILLER_12_581 ();
 sg13g2_decap_4 FILLER_12_685 ();
 sg13g2_fill_1 FILLER_12_689 ();
 sg13g2_fill_2 FILLER_12_762 ();
 sg13g2_fill_1 FILLER_12_769 ();
 sg13g2_fill_1 FILLER_12_778 ();
 sg13g2_fill_2 FILLER_12_833 ();
 sg13g2_fill_1 FILLER_13_13 ();
 sg13g2_fill_1 FILLER_13_24 ();
 sg13g2_fill_1 FILLER_13_117 ();
 sg13g2_fill_1 FILLER_13_172 ();
 sg13g2_fill_2 FILLER_13_193 ();
 sg13g2_fill_1 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_247 ();
 sg13g2_fill_2 FILLER_13_256 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_294 ();
 sg13g2_fill_1 FILLER_13_304 ();
 sg13g2_fill_2 FILLER_13_326 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_fill_2 FILLER_13_371 ();
 sg13g2_fill_2 FILLER_13_381 ();
 sg13g2_fill_1 FILLER_13_391 ();
 sg13g2_fill_2 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_415 ();
 sg13g2_fill_1 FILLER_13_417 ();
 sg13g2_fill_2 FILLER_13_434 ();
 sg13g2_fill_1 FILLER_13_460 ();
 sg13g2_fill_1 FILLER_13_471 ();
 sg13g2_fill_1 FILLER_13_484 ();
 sg13g2_fill_1 FILLER_13_506 ();
 sg13g2_fill_1 FILLER_13_520 ();
 sg13g2_fill_1 FILLER_13_529 ();
 sg13g2_fill_1 FILLER_13_542 ();
 sg13g2_fill_1 FILLER_13_576 ();
 sg13g2_fill_2 FILLER_13_638 ();
 sg13g2_fill_1 FILLER_13_644 ();
 sg13g2_fill_1 FILLER_13_692 ();
 sg13g2_fill_2 FILLER_13_701 ();
 sg13g2_fill_2 FILLER_13_711 ();
 sg13g2_fill_2 FILLER_13_717 ();
 sg13g2_fill_2 FILLER_13_755 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_55 ();
 sg13g2_fill_2 FILLER_14_60 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_86 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_fill_2 FILLER_14_109 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_fill_1 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_168 ();
 sg13g2_fill_2 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_220 ();
 sg13g2_fill_2 FILLER_14_225 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_fill_1 FILLER_14_324 ();
 sg13g2_fill_1 FILLER_14_351 ();
 sg13g2_fill_1 FILLER_14_357 ();
 sg13g2_fill_1 FILLER_14_363 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_382 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_14_416 ();
 sg13g2_fill_1 FILLER_14_421 ();
 sg13g2_fill_1 FILLER_14_431 ();
 sg13g2_fill_2 FILLER_14_436 ();
 sg13g2_fill_2 FILLER_14_442 ();
 sg13g2_fill_1 FILLER_14_456 ();
 sg13g2_fill_2 FILLER_14_469 ();
 sg13g2_fill_1 FILLER_14_479 ();
 sg13g2_fill_2 FILLER_14_510 ();
 sg13g2_fill_1 FILLER_14_527 ();
 sg13g2_decap_4 FILLER_14_540 ();
 sg13g2_fill_1 FILLER_14_571 ();
 sg13g2_fill_2 FILLER_14_585 ();
 sg13g2_fill_1 FILLER_14_595 ();
 sg13g2_fill_1 FILLER_14_654 ();
 sg13g2_fill_2 FILLER_14_711 ();
 sg13g2_fill_1 FILLER_14_747 ();
 sg13g2_fill_1 FILLER_14_752 ();
 sg13g2_fill_1 FILLER_14_757 ();
 sg13g2_fill_1 FILLER_14_828 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_fill_1 FILLER_15_74 ();
 sg13g2_fill_1 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_fill_2 FILLER_15_190 ();
 sg13g2_fill_2 FILLER_15_197 ();
 sg13g2_fill_2 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_343 ();
 sg13g2_fill_1 FILLER_15_370 ();
 sg13g2_fill_2 FILLER_15_397 ();
 sg13g2_fill_1 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_412 ();
 sg13g2_fill_2 FILLER_15_421 ();
 sg13g2_fill_1 FILLER_15_423 ();
 sg13g2_fill_2 FILLER_15_526 ();
 sg13g2_fill_1 FILLER_15_528 ();
 sg13g2_fill_2 FILLER_15_565 ();
 sg13g2_fill_1 FILLER_15_579 ();
 sg13g2_fill_1 FILLER_15_584 ();
 sg13g2_fill_2 FILLER_15_638 ();
 sg13g2_fill_1 FILLER_15_653 ();
 sg13g2_fill_2 FILLER_15_691 ();
 sg13g2_fill_2 FILLER_15_725 ();
 sg13g2_fill_2 FILLER_15_761 ();
 sg13g2_fill_1 FILLER_15_768 ();
 sg13g2_fill_1 FILLER_15_777 ();
 sg13g2_fill_2 FILLER_15_786 ();
 sg13g2_fill_1 FILLER_15_796 ();
 sg13g2_fill_1 FILLER_15_820 ();
 sg13g2_fill_2 FILLER_16_40 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_97 ();
 sg13g2_fill_1 FILLER_16_108 ();
 sg13g2_fill_1 FILLER_16_113 ();
 sg13g2_fill_1 FILLER_16_122 ();
 sg13g2_fill_2 FILLER_16_142 ();
 sg13g2_fill_1 FILLER_16_159 ();
 sg13g2_fill_1 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_173 ();
 sg13g2_fill_1 FILLER_16_178 ();
 sg13g2_fill_1 FILLER_16_213 ();
 sg13g2_fill_1 FILLER_16_227 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_1 FILLER_16_242 ();
 sg13g2_fill_1 FILLER_16_247 ();
 sg13g2_fill_1 FILLER_16_252 ();
 sg13g2_fill_1 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_263 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_363 ();
 sg13g2_fill_2 FILLER_16_390 ();
 sg13g2_fill_1 FILLER_16_395 ();
 sg13g2_fill_1 FILLER_16_400 ();
 sg13g2_fill_1 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_444 ();
 sg13g2_fill_2 FILLER_16_455 ();
 sg13g2_fill_1 FILLER_16_457 ();
 sg13g2_fill_1 FILLER_16_470 ();
 sg13g2_decap_8 FILLER_16_510 ();
 sg13g2_fill_1 FILLER_16_529 ();
 sg13g2_fill_1 FILLER_16_553 ();
 sg13g2_fill_1 FILLER_16_558 ();
 sg13g2_fill_2 FILLER_16_563 ();
 sg13g2_fill_1 FILLER_16_577 ();
 sg13g2_fill_1 FILLER_16_621 ();
 sg13g2_fill_2 FILLER_16_635 ();
 sg13g2_fill_1 FILLER_16_767 ();
 sg13g2_fill_1 FILLER_16_776 ();
 sg13g2_fill_1 FILLER_16_782 ();
 sg13g2_fill_1 FILLER_16_807 ();
 sg13g2_fill_2 FILLER_16_826 ();
 sg13g2_fill_1 FILLER_16_832 ();
 sg13g2_fill_1 FILLER_16_845 ();
 sg13g2_fill_1 FILLER_17_30 ();
 sg13g2_fill_2 FILLER_17_60 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_331 ();
 sg13g2_fill_2 FILLER_17_352 ();
 sg13g2_fill_1 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_363 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_fill_1 FILLER_17_381 ();
 sg13g2_fill_2 FILLER_17_398 ();
 sg13g2_fill_2 FILLER_17_424 ();
 sg13g2_decap_8 FILLER_17_436 ();
 sg13g2_decap_4 FILLER_17_443 ();
 sg13g2_fill_2 FILLER_17_447 ();
 sg13g2_fill_1 FILLER_17_479 ();
 sg13g2_fill_2 FILLER_17_523 ();
 sg13g2_fill_2 FILLER_17_536 ();
 sg13g2_decap_4 FILLER_17_568 ();
 sg13g2_fill_1 FILLER_17_572 ();
 sg13g2_fill_1 FILLER_17_580 ();
 sg13g2_fill_1 FILLER_17_624 ();
 sg13g2_fill_2 FILLER_17_673 ();
 sg13g2_fill_1 FILLER_17_696 ();
 sg13g2_fill_2 FILLER_17_745 ();
 sg13g2_fill_2 FILLER_17_796 ();
 sg13g2_fill_2 FILLER_17_813 ();
 sg13g2_fill_2 FILLER_17_831 ();
 sg13g2_fill_2 FILLER_18_36 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_209 ();
 sg13g2_fill_1 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_fill_2 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_281 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_fill_1 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_fill_2 FILLER_18_375 ();
 sg13g2_fill_2 FILLER_18_398 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_4 FILLER_18_414 ();
 sg13g2_fill_2 FILLER_18_422 ();
 sg13g2_fill_1 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_433 ();
 sg13g2_fill_2 FILLER_18_439 ();
 sg13g2_fill_1 FILLER_18_483 ();
 sg13g2_fill_1 FILLER_18_534 ();
 sg13g2_fill_1 FILLER_18_548 ();
 sg13g2_fill_2 FILLER_18_573 ();
 sg13g2_fill_2 FILLER_18_619 ();
 sg13g2_fill_1 FILLER_18_645 ();
 sg13g2_fill_1 FILLER_18_676 ();
 sg13g2_fill_2 FILLER_18_681 ();
 sg13g2_fill_2 FILLER_18_735 ();
 sg13g2_fill_2 FILLER_18_835 ();
 sg13g2_fill_1 FILLER_18_877 ();
 sg13g2_fill_2 FILLER_19_15 ();
 sg13g2_fill_1 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_fill_1 FILLER_19_260 ();
 sg13g2_fill_2 FILLER_19_284 ();
 sg13g2_fill_2 FILLER_19_354 ();
 sg13g2_fill_2 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_371 ();
 sg13g2_fill_1 FILLER_19_416 ();
 sg13g2_fill_1 FILLER_19_428 ();
 sg13g2_fill_1 FILLER_19_459 ();
 sg13g2_fill_1 FILLER_19_509 ();
 sg13g2_fill_1 FILLER_19_526 ();
 sg13g2_fill_1 FILLER_19_535 ();
 sg13g2_fill_2 FILLER_19_548 ();
 sg13g2_fill_1 FILLER_19_558 ();
 sg13g2_fill_1 FILLER_19_579 ();
 sg13g2_fill_2 FILLER_19_584 ();
 sg13g2_fill_2 FILLER_19_612 ();
 sg13g2_fill_1 FILLER_19_619 ();
 sg13g2_fill_2 FILLER_19_685 ();
 sg13g2_fill_1 FILLER_19_703 ();
 sg13g2_fill_1 FILLER_19_736 ();
 sg13g2_fill_1 FILLER_19_746 ();
 sg13g2_fill_2 FILLER_19_769 ();
 sg13g2_fill_1 FILLER_19_805 ();
 sg13g2_fill_1 FILLER_19_851 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_13 ();
 sg13g2_fill_2 FILLER_20_49 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_fill_2 FILLER_20_345 ();
 sg13g2_decap_4 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_484 ();
 sg13g2_fill_1 FILLER_20_511 ();
 sg13g2_fill_1 FILLER_20_520 ();
 sg13g2_fill_1 FILLER_20_543 ();
 sg13g2_fill_2 FILLER_20_552 ();
 sg13g2_fill_1 FILLER_20_578 ();
 sg13g2_fill_1 FILLER_20_599 ();
 sg13g2_fill_1 FILLER_20_617 ();
 sg13g2_fill_1 FILLER_20_733 ();
 sg13g2_fill_1 FILLER_20_743 ();
 sg13g2_fill_1 FILLER_20_771 ();
 sg13g2_fill_1 FILLER_20_775 ();
 sg13g2_fill_1 FILLER_20_782 ();
 sg13g2_fill_2 FILLER_20_789 ();
 sg13g2_fill_2 FILLER_20_810 ();
 sg13g2_fill_1 FILLER_20_838 ();
 sg13g2_fill_1 FILLER_20_843 ();
 sg13g2_fill_2 FILLER_20_849 ();
 sg13g2_fill_1 FILLER_20_877 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_fill_2 FILLER_21_156 ();
 sg13g2_fill_2 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_315 ();
 sg13g2_fill_1 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_348 ();
 sg13g2_fill_1 FILLER_21_407 ();
 sg13g2_fill_2 FILLER_21_420 ();
 sg13g2_fill_2 FILLER_21_443 ();
 sg13g2_fill_2 FILLER_21_506 ();
 sg13g2_fill_2 FILLER_21_518 ();
 sg13g2_fill_2 FILLER_21_533 ();
 sg13g2_fill_2 FILLER_21_555 ();
 sg13g2_fill_1 FILLER_21_557 ();
 sg13g2_fill_2 FILLER_21_574 ();
 sg13g2_fill_1 FILLER_21_698 ();
 sg13g2_fill_1 FILLER_21_720 ();
 sg13g2_fill_2 FILLER_21_734 ();
 sg13g2_fill_1 FILLER_21_744 ();
 sg13g2_fill_2 FILLER_21_789 ();
 sg13g2_fill_2 FILLER_21_798 ();
 sg13g2_fill_1 FILLER_21_826 ();
 sg13g2_fill_2 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_864 ();
 sg13g2_fill_2 FILLER_21_869 ();
 sg13g2_fill_1 FILLER_22_30 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_fill_2 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_406 ();
 sg13g2_decap_4 FILLER_22_432 ();
 sg13g2_fill_1 FILLER_22_436 ();
 sg13g2_fill_1 FILLER_22_442 ();
 sg13g2_fill_1 FILLER_22_447 ();
 sg13g2_fill_1 FILLER_22_452 ();
 sg13g2_fill_1 FILLER_22_457 ();
 sg13g2_fill_1 FILLER_22_463 ();
 sg13g2_fill_1 FILLER_22_475 ();
 sg13g2_fill_1 FILLER_22_495 ();
 sg13g2_fill_2 FILLER_22_525 ();
 sg13g2_fill_1 FILLER_22_527 ();
 sg13g2_fill_2 FILLER_22_536 ();
 sg13g2_fill_1 FILLER_22_538 ();
 sg13g2_fill_2 FILLER_22_551 ();
 sg13g2_fill_1 FILLER_22_606 ();
 sg13g2_fill_1 FILLER_22_760 ();
 sg13g2_fill_2 FILLER_22_771 ();
 sg13g2_fill_1 FILLER_22_793 ();
 sg13g2_fill_1 FILLER_22_813 ();
 sg13g2_fill_1 FILLER_22_830 ();
 sg13g2_fill_1 FILLER_22_849 ();
 sg13g2_fill_2 FILLER_22_876 ();
 sg13g2_fill_1 FILLER_23_38 ();
 sg13g2_fill_1 FILLER_23_52 ();
 sg13g2_fill_1 FILLER_23_58 ();
 sg13g2_fill_2 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_141 ();
 sg13g2_fill_1 FILLER_23_155 ();
 sg13g2_decap_4 FILLER_23_176 ();
 sg13g2_decap_4 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_fill_1 FILLER_23_287 ();
 sg13g2_fill_1 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_372 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_383 ();
 sg13g2_fill_2 FILLER_23_387 ();
 sg13g2_fill_2 FILLER_23_414 ();
 sg13g2_fill_1 FILLER_23_424 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_fill_1 FILLER_23_461 ();
 sg13g2_fill_2 FILLER_23_466 ();
 sg13g2_fill_1 FILLER_23_499 ();
 sg13g2_fill_2 FILLER_23_545 ();
 sg13g2_fill_1 FILLER_23_550 ();
 sg13g2_fill_1 FILLER_23_593 ();
 sg13g2_fill_1 FILLER_23_604 ();
 sg13g2_fill_1 FILLER_23_668 ();
 sg13g2_fill_1 FILLER_23_674 ();
 sg13g2_fill_1 FILLER_23_742 ();
 sg13g2_fill_2 FILLER_23_759 ();
 sg13g2_fill_1 FILLER_23_766 ();
 sg13g2_fill_1 FILLER_23_816 ();
 sg13g2_fill_1 FILLER_23_822 ();
 sg13g2_fill_2 FILLER_23_876 ();
 sg13g2_fill_1 FILLER_24_41 ();
 sg13g2_fill_1 FILLER_24_46 ();
 sg13g2_fill_2 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_145 ();
 sg13g2_fill_2 FILLER_24_155 ();
 sg13g2_fill_2 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_222 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_393 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_fill_1 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_fill_1 FILLER_24_438 ();
 sg13g2_fill_1 FILLER_24_447 ();
 sg13g2_fill_1 FILLER_24_453 ();
 sg13g2_fill_2 FILLER_24_500 ();
 sg13g2_fill_1 FILLER_24_510 ();
 sg13g2_fill_1 FILLER_24_519 ();
 sg13g2_fill_1 FILLER_24_532 ();
 sg13g2_fill_2 FILLER_24_559 ();
 sg13g2_fill_2 FILLER_24_566 ();
 sg13g2_fill_1 FILLER_24_572 ();
 sg13g2_fill_2 FILLER_24_627 ();
 sg13g2_fill_2 FILLER_24_648 ();
 sg13g2_fill_1 FILLER_24_738 ();
 sg13g2_fill_1 FILLER_24_743 ();
 sg13g2_fill_1 FILLER_24_769 ();
 sg13g2_fill_1 FILLER_24_845 ();
 sg13g2_fill_2 FILLER_24_876 ();
 sg13g2_fill_1 FILLER_25_72 ();
 sg13g2_fill_2 FILLER_25_92 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_2 FILLER_25_130 ();
 sg13g2_fill_2 FILLER_25_182 ();
 sg13g2_fill_2 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_204 ();
 sg13g2_fill_1 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_1 FILLER_25_300 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_1 FILLER_25_318 ();
 sg13g2_fill_1 FILLER_25_356 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_1 FILLER_25_387 ();
 sg13g2_fill_2 FILLER_25_397 ();
 sg13g2_fill_1 FILLER_25_437 ();
 sg13g2_fill_2 FILLER_25_466 ();
 sg13g2_fill_2 FILLER_25_498 ();
 sg13g2_fill_2 FILLER_25_516 ();
 sg13g2_fill_1 FILLER_25_518 ();
 sg13g2_fill_1 FILLER_25_529 ();
 sg13g2_fill_1 FILLER_25_543 ();
 sg13g2_fill_2 FILLER_25_587 ();
 sg13g2_fill_2 FILLER_25_610 ();
 sg13g2_fill_2 FILLER_25_620 ();
 sg13g2_fill_1 FILLER_25_630 ();
 sg13g2_fill_1 FILLER_25_657 ();
 sg13g2_fill_1 FILLER_25_676 ();
 sg13g2_fill_1 FILLER_25_687 ();
 sg13g2_fill_2 FILLER_25_709 ();
 sg13g2_fill_1 FILLER_25_737 ();
 sg13g2_fill_2 FILLER_25_742 ();
 sg13g2_fill_1 FILLER_25_748 ();
 sg13g2_fill_1 FILLER_25_779 ();
 sg13g2_fill_1 FILLER_25_795 ();
 sg13g2_fill_1 FILLER_25_848 ();
 sg13g2_fill_1 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_80 ();
 sg13g2_fill_1 FILLER_26_89 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_fill_1 FILLER_26_158 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_2 FILLER_26_243 ();
 sg13g2_fill_1 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_fill_2 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_1 FILLER_26_411 ();
 sg13g2_fill_2 FILLER_26_524 ();
 sg13g2_fill_2 FILLER_26_544 ();
 sg13g2_fill_1 FILLER_26_560 ();
 sg13g2_fill_1 FILLER_26_579 ();
 sg13g2_fill_2 FILLER_26_596 ();
 sg13g2_fill_2 FILLER_26_604 ();
 sg13g2_fill_1 FILLER_26_660 ();
 sg13g2_fill_1 FILLER_26_728 ();
 sg13g2_fill_2 FILLER_26_750 ();
 sg13g2_fill_2 FILLER_26_795 ();
 sg13g2_fill_2 FILLER_26_805 ();
 sg13g2_fill_1 FILLER_26_872 ();
 sg13g2_fill_1 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_117 ();
 sg13g2_fill_2 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_205 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_fill_1 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_344 ();
 sg13g2_fill_2 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_414 ();
 sg13g2_fill_1 FILLER_27_416 ();
 sg13g2_fill_1 FILLER_27_446 ();
 sg13g2_fill_2 FILLER_27_481 ();
 sg13g2_fill_2 FILLER_27_494 ();
 sg13g2_decap_4 FILLER_27_545 ();
 sg13g2_fill_2 FILLER_27_549 ();
 sg13g2_fill_1 FILLER_27_555 ();
 sg13g2_fill_2 FILLER_27_584 ();
 sg13g2_fill_2 FILLER_27_620 ();
 sg13g2_fill_2 FILLER_27_663 ();
 sg13g2_fill_2 FILLER_27_730 ();
 sg13g2_fill_1 FILLER_27_746 ();
 sg13g2_fill_1 FILLER_27_789 ();
 sg13g2_fill_1 FILLER_27_811 ();
 sg13g2_fill_1 FILLER_27_818 ();
 sg13g2_fill_1 FILLER_27_851 ();
 sg13g2_fill_1 FILLER_28_36 ();
 sg13g2_fill_1 FILLER_28_45 ();
 sg13g2_fill_1 FILLER_28_55 ();
 sg13g2_fill_2 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_95 ();
 sg13g2_fill_1 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_decap_4 FILLER_28_376 ();
 sg13g2_fill_2 FILLER_28_409 ();
 sg13g2_fill_1 FILLER_28_425 ();
 sg13g2_decap_4 FILLER_28_470 ();
 sg13g2_fill_1 FILLER_28_474 ();
 sg13g2_decap_8 FILLER_28_492 ();
 sg13g2_fill_1 FILLER_28_499 ();
 sg13g2_fill_2 FILLER_28_518 ();
 sg13g2_fill_1 FILLER_28_520 ();
 sg13g2_fill_2 FILLER_28_543 ();
 sg13g2_fill_1 FILLER_28_554 ();
 sg13g2_fill_2 FILLER_28_563 ();
 sg13g2_fill_2 FILLER_28_569 ();
 sg13g2_fill_2 FILLER_28_577 ();
 sg13g2_decap_4 FILLER_28_584 ();
 sg13g2_fill_1 FILLER_28_627 ();
 sg13g2_fill_2 FILLER_28_638 ();
 sg13g2_fill_2 FILLER_28_645 ();
 sg13g2_fill_2 FILLER_28_650 ();
 sg13g2_fill_1 FILLER_28_689 ();
 sg13g2_fill_2 FILLER_28_764 ();
 sg13g2_fill_2 FILLER_28_782 ();
 sg13g2_fill_2 FILLER_29_61 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_168 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_183 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_254 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_344 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_4 FILLER_29_500 ();
 sg13g2_fill_1 FILLER_29_504 ();
 sg13g2_fill_1 FILLER_29_536 ();
 sg13g2_fill_2 FILLER_29_599 ();
 sg13g2_fill_1 FILLER_29_611 ();
 sg13g2_fill_1 FILLER_29_686 ();
 sg13g2_fill_1 FILLER_29_691 ();
 sg13g2_fill_1 FILLER_29_709 ();
 sg13g2_fill_2 FILLER_29_739 ();
 sg13g2_fill_2 FILLER_29_758 ();
 sg13g2_fill_1 FILLER_29_764 ();
 sg13g2_fill_1 FILLER_29_808 ();
 sg13g2_fill_1 FILLER_29_817 ();
 sg13g2_fill_1 FILLER_29_851 ();
 sg13g2_fill_2 FILLER_30_44 ();
 sg13g2_fill_2 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_fill_1 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_185 ();
 sg13g2_fill_1 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_fill_2 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_413 ();
 sg13g2_fill_2 FILLER_30_425 ();
 sg13g2_fill_1 FILLER_30_436 ();
 sg13g2_fill_2 FILLER_30_456 ();
 sg13g2_fill_1 FILLER_30_465 ();
 sg13g2_fill_2 FILLER_30_474 ();
 sg13g2_fill_1 FILLER_30_489 ();
 sg13g2_fill_1 FILLER_30_613 ();
 sg13g2_fill_1 FILLER_30_628 ();
 sg13g2_fill_2 FILLER_30_637 ();
 sg13g2_fill_1 FILLER_30_712 ();
 sg13g2_fill_1 FILLER_30_826 ();
 sg13g2_fill_2 FILLER_31_34 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_fill_1 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_97 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_fill_2 FILLER_31_242 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_249 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_387 ();
 sg13g2_fill_1 FILLER_31_392 ();
 sg13g2_fill_1 FILLER_31_418 ();
 sg13g2_fill_1 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_444 ();
 sg13g2_fill_2 FILLER_31_479 ();
 sg13g2_fill_1 FILLER_31_484 ();
 sg13g2_fill_1 FILLER_31_526 ();
 sg13g2_fill_2 FILLER_31_530 ();
 sg13g2_fill_2 FILLER_31_545 ();
 sg13g2_fill_2 FILLER_31_552 ();
 sg13g2_fill_1 FILLER_31_562 ();
 sg13g2_fill_1 FILLER_31_586 ();
 sg13g2_fill_1 FILLER_31_628 ();
 sg13g2_fill_1 FILLER_31_651 ();
 sg13g2_fill_1 FILLER_31_657 ();
 sg13g2_fill_1 FILLER_31_662 ();
 sg13g2_fill_2 FILLER_31_667 ();
 sg13g2_fill_1 FILLER_31_677 ();
 sg13g2_fill_1 FILLER_31_687 ();
 sg13g2_fill_1 FILLER_31_692 ();
 sg13g2_fill_2 FILLER_31_712 ();
 sg13g2_fill_1 FILLER_31_719 ();
 sg13g2_fill_1 FILLER_31_779 ();
 sg13g2_fill_1 FILLER_31_789 ();
 sg13g2_fill_1 FILLER_31_795 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_115 ();
 sg13g2_fill_2 FILLER_32_169 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_198 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_239 ();
 sg13g2_fill_2 FILLER_32_266 ();
 sg13g2_fill_2 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_378 ();
 sg13g2_fill_1 FILLER_32_388 ();
 sg13g2_fill_1 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_402 ();
 sg13g2_fill_1 FILLER_32_411 ();
 sg13g2_fill_2 FILLER_32_416 ();
 sg13g2_fill_2 FILLER_32_423 ();
 sg13g2_fill_2 FILLER_32_433 ();
 sg13g2_fill_1 FILLER_32_435 ();
 sg13g2_fill_2 FILLER_32_470 ();
 sg13g2_fill_2 FILLER_32_513 ();
 sg13g2_fill_1 FILLER_32_515 ();
 sg13g2_fill_1 FILLER_32_519 ();
 sg13g2_fill_1 FILLER_32_599 ();
 sg13g2_fill_2 FILLER_32_619 ();
 sg13g2_fill_2 FILLER_32_652 ();
 sg13g2_fill_1 FILLER_32_745 ();
 sg13g2_fill_2 FILLER_32_829 ();
 sg13g2_fill_1 FILLER_32_831 ();
 sg13g2_fill_2 FILLER_32_849 ();
 sg13g2_fill_1 FILLER_32_851 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_fill_1 FILLER_33_39 ();
 sg13g2_fill_1 FILLER_33_48 ();
 sg13g2_fill_1 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_121 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_189 ();
 sg13g2_fill_1 FILLER_33_235 ();
 sg13g2_fill_1 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_1 FILLER_33_370 ();
 sg13g2_fill_1 FILLER_33_375 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_fill_1 FILLER_33_388 ();
 sg13g2_fill_2 FILLER_33_394 ();
 sg13g2_fill_1 FILLER_33_509 ();
 sg13g2_fill_2 FILLER_33_525 ();
 sg13g2_fill_1 FILLER_33_531 ();
 sg13g2_fill_2 FILLER_33_543 ();
 sg13g2_fill_2 FILLER_33_551 ();
 sg13g2_fill_2 FILLER_33_582 ();
 sg13g2_fill_1 FILLER_33_590 ();
 sg13g2_fill_2 FILLER_33_598 ();
 sg13g2_fill_2 FILLER_33_604 ();
 sg13g2_fill_1 FILLER_33_636 ();
 sg13g2_fill_1 FILLER_33_663 ();
 sg13g2_fill_1 FILLER_33_752 ();
 sg13g2_fill_2 FILLER_33_767 ();
 sg13g2_fill_1 FILLER_33_769 ();
 sg13g2_fill_1 FILLER_33_796 ();
 sg13g2_fill_2 FILLER_33_866 ();
 sg13g2_fill_2 FILLER_33_876 ();
 sg13g2_fill_2 FILLER_34_13 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_fill_2 FILLER_34_169 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_fill_2 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_385 ();
 sg13g2_fill_1 FILLER_34_391 ();
 sg13g2_fill_1 FILLER_34_395 ();
 sg13g2_fill_1 FILLER_34_401 ();
 sg13g2_fill_2 FILLER_34_414 ();
 sg13g2_decap_4 FILLER_34_438 ();
 sg13g2_fill_1 FILLER_34_472 ();
 sg13g2_fill_2 FILLER_34_504 ();
 sg13g2_fill_1 FILLER_34_514 ();
 sg13g2_fill_1 FILLER_34_528 ();
 sg13g2_fill_2 FILLER_34_534 ();
 sg13g2_fill_1 FILLER_34_541 ();
 sg13g2_fill_2 FILLER_34_553 ();
 sg13g2_fill_1 FILLER_34_617 ();
 sg13g2_fill_2 FILLER_34_696 ();
 sg13g2_fill_2 FILLER_34_730 ();
 sg13g2_fill_1 FILLER_34_835 ();
 sg13g2_fill_1 FILLER_35_23 ();
 sg13g2_fill_2 FILLER_35_68 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_90 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_fill_1 FILLER_35_144 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_317 ();
 sg13g2_fill_2 FILLER_35_405 ();
 sg13g2_fill_1 FILLER_35_426 ();
 sg13g2_fill_1 FILLER_35_431 ();
 sg13g2_fill_2 FILLER_35_440 ();
 sg13g2_fill_1 FILLER_35_446 ();
 sg13g2_fill_1 FILLER_35_453 ();
 sg13g2_fill_1 FILLER_35_457 ();
 sg13g2_fill_1 FILLER_35_462 ();
 sg13g2_fill_1 FILLER_35_466 ();
 sg13g2_fill_1 FILLER_35_511 ();
 sg13g2_fill_1 FILLER_35_523 ();
 sg13g2_fill_1 FILLER_35_536 ();
 sg13g2_fill_1 FILLER_35_545 ();
 sg13g2_fill_2 FILLER_35_563 ();
 sg13g2_fill_1 FILLER_35_702 ();
 sg13g2_fill_1 FILLER_35_716 ();
 sg13g2_fill_2 FILLER_35_755 ();
 sg13g2_fill_1 FILLER_35_801 ();
 sg13g2_fill_2 FILLER_35_811 ();
 sg13g2_fill_1 FILLER_35_831 ();
 sg13g2_fill_2 FILLER_35_853 ();
 sg13g2_fill_1 FILLER_35_871 ();
 sg13g2_fill_1 FILLER_35_877 ();
 sg13g2_fill_2 FILLER_36_24 ();
 sg13g2_fill_2 FILLER_36_41 ();
 sg13g2_fill_1 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_73 ();
 sg13g2_fill_1 FILLER_36_82 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_decap_4 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_116 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_185 ();
 sg13g2_fill_2 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_254 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_fill_1 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_426 ();
 sg13g2_fill_2 FILLER_36_432 ();
 sg13g2_fill_1 FILLER_36_434 ();
 sg13g2_fill_1 FILLER_36_512 ();
 sg13g2_fill_1 FILLER_36_536 ();
 sg13g2_fill_2 FILLER_36_542 ();
 sg13g2_fill_2 FILLER_36_653 ();
 sg13g2_fill_1 FILLER_36_655 ();
 sg13g2_fill_2 FILLER_36_692 ();
 sg13g2_fill_1 FILLER_36_694 ();
 sg13g2_fill_2 FILLER_36_737 ();
 sg13g2_fill_2 FILLER_36_747 ();
 sg13g2_fill_1 FILLER_36_775 ();
 sg13g2_fill_1 FILLER_36_801 ();
 sg13g2_fill_1 FILLER_36_807 ();
 sg13g2_fill_2 FILLER_36_858 ();
 sg13g2_fill_2 FILLER_36_876 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_97 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_275 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_fill_1 FILLER_37_312 ();
 sg13g2_fill_1 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_fill_1 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_389 ();
 sg13g2_fill_1 FILLER_37_419 ();
 sg13g2_fill_1 FILLER_37_424 ();
 sg13g2_decap_4 FILLER_37_430 ();
 sg13g2_fill_2 FILLER_37_439 ();
 sg13g2_fill_2 FILLER_37_444 ();
 sg13g2_fill_1 FILLER_37_457 ();
 sg13g2_fill_1 FILLER_37_477 ();
 sg13g2_fill_2 FILLER_37_483 ();
 sg13g2_fill_1 FILLER_37_575 ();
 sg13g2_fill_1 FILLER_37_812 ();
 sg13g2_fill_1 FILLER_37_856 ();
 sg13g2_fill_2 FILLER_38_50 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_78 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_88 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_fill_1 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_130 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_fill_2 FILLER_38_145 ();
 sg13g2_fill_2 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_158 ();
 sg13g2_fill_1 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_231 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_fill_2 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_347 ();
 sg13g2_fill_1 FILLER_38_353 ();
 sg13g2_fill_1 FILLER_38_358 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_4 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_384 ();
 sg13g2_fill_2 FILLER_38_393 ();
 sg13g2_fill_2 FILLER_38_447 ();
 sg13g2_fill_1 FILLER_38_465 ();
 sg13g2_fill_2 FILLER_38_470 ();
 sg13g2_fill_1 FILLER_38_480 ();
 sg13g2_fill_1 FILLER_38_486 ();
 sg13g2_fill_2 FILLER_38_519 ();
 sg13g2_fill_1 FILLER_38_529 ();
 sg13g2_fill_1 FILLER_38_549 ();
 sg13g2_fill_1 FILLER_38_595 ();
 sg13g2_fill_1 FILLER_38_609 ();
 sg13g2_fill_1 FILLER_38_614 ();
 sg13g2_fill_1 FILLER_38_620 ();
 sg13g2_fill_1 FILLER_38_647 ();
 sg13g2_fill_2 FILLER_38_678 ();
 sg13g2_fill_1 FILLER_38_717 ();
 sg13g2_fill_1 FILLER_38_736 ();
 sg13g2_fill_2 FILLER_38_793 ();
 sg13g2_fill_1 FILLER_38_851 ();
 sg13g2_fill_1 FILLER_38_857 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_6 ();
 sg13g2_decap_8 FILLER_39_30 ();
 sg13g2_fill_1 FILLER_39_37 ();
 sg13g2_fill_2 FILLER_39_91 ();
 sg13g2_fill_2 FILLER_39_139 ();
 sg13g2_fill_1 FILLER_39_141 ();
 sg13g2_fill_1 FILLER_39_147 ();
 sg13g2_fill_2 FILLER_39_156 ();
 sg13g2_fill_1 FILLER_39_199 ();
 sg13g2_fill_2 FILLER_39_325 ();
 sg13g2_fill_1 FILLER_39_335 ();
 sg13g2_fill_1 FILLER_39_360 ();
 sg13g2_fill_1 FILLER_39_365 ();
 sg13g2_fill_1 FILLER_39_370 ();
 sg13g2_fill_1 FILLER_39_392 ();
 sg13g2_fill_2 FILLER_39_415 ();
 sg13g2_fill_2 FILLER_39_440 ();
 sg13g2_fill_1 FILLER_39_442 ();
 sg13g2_fill_1 FILLER_39_453 ();
 sg13g2_fill_1 FILLER_39_457 ();
 sg13g2_fill_1 FILLER_39_473 ();
 sg13g2_fill_2 FILLER_39_529 ();
 sg13g2_fill_1 FILLER_39_536 ();
 sg13g2_fill_1 FILLER_39_542 ();
 sg13g2_fill_2 FILLER_39_547 ();
 sg13g2_fill_1 FILLER_39_579 ();
 sg13g2_fill_1 FILLER_39_619 ();
 sg13g2_fill_2 FILLER_39_625 ();
 sg13g2_fill_2 FILLER_39_631 ();
 sg13g2_fill_1 FILLER_39_640 ();
 sg13g2_fill_1 FILLER_39_654 ();
 sg13g2_fill_1 FILLER_39_668 ();
 sg13g2_fill_1 FILLER_39_673 ();
 sg13g2_fill_2 FILLER_39_678 ();
 sg13g2_fill_2 FILLER_39_721 ();
 sg13g2_fill_1 FILLER_39_737 ();
 sg13g2_fill_2 FILLER_39_769 ();
 sg13g2_fill_2 FILLER_39_789 ();
 sg13g2_fill_2 FILLER_39_864 ();
 sg13g2_fill_1 FILLER_40_30 ();
 sg13g2_fill_1 FILLER_40_39 ();
 sg13g2_fill_2 FILLER_40_66 ();
 sg13g2_fill_2 FILLER_40_114 ();
 sg13g2_fill_1 FILLER_40_120 ();
 sg13g2_fill_2 FILLER_40_126 ();
 sg13g2_fill_1 FILLER_40_132 ();
 sg13g2_fill_1 FILLER_40_146 ();
 sg13g2_fill_1 FILLER_40_151 ();
 sg13g2_fill_1 FILLER_40_177 ();
 sg13g2_fill_2 FILLER_40_189 ();
 sg13g2_fill_1 FILLER_40_232 ();
 sg13g2_fill_1 FILLER_40_236 ();
 sg13g2_fill_1 FILLER_40_247 ();
 sg13g2_fill_1 FILLER_40_261 ();
 sg13g2_fill_1 FILLER_40_266 ();
 sg13g2_fill_2 FILLER_40_272 ();
 sg13g2_fill_2 FILLER_40_287 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_fill_1 FILLER_40_317 ();
 sg13g2_fill_2 FILLER_40_323 ();
 sg13g2_fill_1 FILLER_40_333 ();
 sg13g2_fill_2 FILLER_40_342 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_decap_8 FILLER_40_377 ();
 sg13g2_fill_2 FILLER_40_392 ();
 sg13g2_fill_2 FILLER_40_419 ();
 sg13g2_fill_1 FILLER_40_426 ();
 sg13g2_fill_1 FILLER_40_440 ();
 sg13g2_fill_2 FILLER_40_487 ();
 sg13g2_fill_2 FILLER_40_519 ();
 sg13g2_decap_8 FILLER_40_577 ();
 sg13g2_fill_2 FILLER_40_584 ();
 sg13g2_fill_1 FILLER_40_599 ();
 sg13g2_fill_1 FILLER_40_604 ();
 sg13g2_fill_1 FILLER_40_612 ();
 sg13g2_fill_1 FILLER_40_618 ();
 sg13g2_fill_1 FILLER_40_658 ();
 sg13g2_fill_2 FILLER_40_685 ();
 sg13g2_fill_1 FILLER_40_703 ();
 sg13g2_fill_1 FILLER_40_708 ();
 sg13g2_fill_2 FILLER_40_746 ();
 sg13g2_fill_2 FILLER_40_773 ();
 sg13g2_fill_1 FILLER_40_782 ();
 sg13g2_decap_4 FILLER_40_787 ();
 sg13g2_fill_2 FILLER_40_795 ();
 sg13g2_fill_1 FILLER_40_797 ();
 sg13g2_fill_1 FILLER_40_803 ();
 sg13g2_fill_2 FILLER_40_847 ();
 sg13g2_fill_1 FILLER_40_872 ();
 sg13g2_fill_1 FILLER_40_877 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_decap_4 FILLER_41_5 ();
 sg13g2_fill_2 FILLER_41_9 ();
 sg13g2_fill_1 FILLER_41_26 ();
 sg13g2_fill_2 FILLER_41_32 ();
 sg13g2_fill_1 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_48 ();
 sg13g2_decap_4 FILLER_41_59 ();
 sg13g2_fill_2 FILLER_41_71 ();
 sg13g2_fill_1 FILLER_41_73 ();
 sg13g2_fill_1 FILLER_41_100 ();
 sg13g2_fill_1 FILLER_41_104 ();
 sg13g2_fill_1 FILLER_41_109 ();
 sg13g2_fill_1 FILLER_41_115 ();
 sg13g2_fill_1 FILLER_41_142 ();
 sg13g2_fill_2 FILLER_41_173 ();
 sg13g2_fill_2 FILLER_41_197 ();
 sg13g2_fill_2 FILLER_41_234 ();
 sg13g2_decap_8 FILLER_41_247 ();
 sg13g2_fill_2 FILLER_41_280 ();
 sg13g2_fill_1 FILLER_41_282 ();
 sg13g2_decap_8 FILLER_41_355 ();
 sg13g2_decap_8 FILLER_41_362 ();
 sg13g2_fill_1 FILLER_41_393 ();
 sg13g2_decap_4 FILLER_41_440 ();
 sg13g2_fill_2 FILLER_41_444 ();
 sg13g2_decap_4 FILLER_41_456 ();
 sg13g2_fill_1 FILLER_41_460 ();
 sg13g2_fill_1 FILLER_41_494 ();
 sg13g2_fill_2 FILLER_41_499 ();
 sg13g2_fill_1 FILLER_41_501 ();
 sg13g2_decap_4 FILLER_41_506 ();
 sg13g2_fill_2 FILLER_41_510 ();
 sg13g2_fill_2 FILLER_41_517 ();
 sg13g2_fill_1 FILLER_41_524 ();
 sg13g2_fill_2 FILLER_41_546 ();
 sg13g2_decap_8 FILLER_41_555 ();
 sg13g2_decap_4 FILLER_41_562 ();
 sg13g2_fill_1 FILLER_41_566 ();
 sg13g2_fill_1 FILLER_41_585 ();
 sg13g2_decap_4 FILLER_41_591 ();
 sg13g2_fill_1 FILLER_41_595 ();
 sg13g2_fill_2 FILLER_41_600 ();
 sg13g2_fill_1 FILLER_41_622 ();
 sg13g2_fill_1 FILLER_41_627 ();
 sg13g2_decap_8 FILLER_41_675 ();
 sg13g2_decap_8 FILLER_41_682 ();
 sg13g2_fill_2 FILLER_41_689 ();
 sg13g2_fill_1 FILLER_41_700 ();
 sg13g2_fill_1 FILLER_41_739 ();
 sg13g2_fill_1 FILLER_41_744 ();
 sg13g2_fill_1 FILLER_41_749 ();
 sg13g2_fill_1 FILLER_41_768 ();
 sg13g2_fill_1 FILLER_41_773 ();
 sg13g2_fill_1 FILLER_41_778 ();
 sg13g2_fill_1 FILLER_41_783 ();
 sg13g2_fill_2 FILLER_41_789 ();
 sg13g2_fill_1 FILLER_41_791 ();
 sg13g2_fill_2 FILLER_41_798 ();
 sg13g2_fill_2 FILLER_41_813 ();
 sg13g2_fill_1 FILLER_41_819 ();
 sg13g2_fill_1 FILLER_41_828 ();
 sg13g2_fill_2 FILLER_42_30 ();
 sg13g2_fill_1 FILLER_42_32 ();
 sg13g2_decap_4 FILLER_42_63 ();
 sg13g2_fill_1 FILLER_42_67 ();
 sg13g2_fill_1 FILLER_42_77 ();
 sg13g2_fill_1 FILLER_42_86 ();
 sg13g2_fill_2 FILLER_42_90 ();
 sg13g2_decap_8 FILLER_42_127 ();
 sg13g2_fill_2 FILLER_42_137 ();
 sg13g2_fill_1 FILLER_42_143 ();
 sg13g2_fill_1 FILLER_42_182 ();
 sg13g2_fill_1 FILLER_42_191 ();
 sg13g2_fill_1 FILLER_42_225 ();
 sg13g2_fill_1 FILLER_42_245 ();
 sg13g2_fill_1 FILLER_42_251 ();
 sg13g2_fill_1 FILLER_42_260 ();
 sg13g2_fill_2 FILLER_42_265 ();
 sg13g2_fill_2 FILLER_42_271 ();
 sg13g2_fill_1 FILLER_42_290 ();
 sg13g2_fill_1 FILLER_42_296 ();
 sg13g2_fill_2 FILLER_42_310 ();
 sg13g2_decap_4 FILLER_42_315 ();
 sg13g2_fill_1 FILLER_42_324 ();
 sg13g2_fill_2 FILLER_42_329 ();
 sg13g2_fill_1 FILLER_42_336 ();
 sg13g2_fill_2 FILLER_42_341 ();
 sg13g2_decap_8 FILLER_42_347 ();
 sg13g2_decap_4 FILLER_42_354 ();
 sg13g2_fill_1 FILLER_42_358 ();
 sg13g2_fill_1 FILLER_42_371 ();
 sg13g2_fill_1 FILLER_42_379 ();
 sg13g2_fill_1 FILLER_42_402 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_fill_2 FILLER_42_417 ();
 sg13g2_fill_1 FILLER_42_419 ();
 sg13g2_fill_2 FILLER_42_423 ();
 sg13g2_fill_1 FILLER_42_425 ();
 sg13g2_fill_1 FILLER_42_464 ();
 sg13g2_decap_8 FILLER_42_473 ();
 sg13g2_decap_8 FILLER_42_480 ();
 sg13g2_fill_2 FILLER_42_487 ();
 sg13g2_fill_1 FILLER_42_489 ();
 sg13g2_fill_2 FILLER_42_499 ();
 sg13g2_fill_2 FILLER_42_514 ();
 sg13g2_fill_1 FILLER_42_531 ();
 sg13g2_fill_2 FILLER_42_576 ();
 sg13g2_fill_1 FILLER_42_578 ();
 sg13g2_fill_1 FILLER_42_596 ();
 sg13g2_fill_2 FILLER_42_601 ();
 sg13g2_fill_1 FILLER_42_650 ();
 sg13g2_fill_2 FILLER_42_655 ();
 sg13g2_fill_2 FILLER_42_662 ();
 sg13g2_decap_8 FILLER_42_669 ();
 sg13g2_fill_1 FILLER_42_680 ();
 sg13g2_fill_2 FILLER_42_693 ();
 sg13g2_decap_4 FILLER_42_722 ();
 sg13g2_fill_1 FILLER_42_726 ();
 sg13g2_fill_1 FILLER_42_739 ();
 sg13g2_fill_1 FILLER_42_744 ();
 sg13g2_fill_1 FILLER_42_753 ();
 sg13g2_fill_1 FILLER_42_758 ();
 sg13g2_fill_2 FILLER_42_784 ();
 sg13g2_fill_2 FILLER_42_804 ();
 sg13g2_fill_1 FILLER_42_806 ();
 sg13g2_fill_1 FILLER_42_819 ();
 sg13g2_fill_1 FILLER_42_825 ();
 sg13g2_fill_1 FILLER_42_843 ();
 sg13g2_fill_2 FILLER_42_871 ();
 sg13g2_fill_2 FILLER_42_876 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_27 ();
 sg13g2_fill_1 FILLER_43_54 ();
 sg13g2_fill_1 FILLER_43_81 ();
 sg13g2_fill_1 FILLER_43_112 ();
 sg13g2_fill_1 FILLER_43_155 ();
 sg13g2_fill_1 FILLER_43_186 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_fill_2 FILLER_43_211 ();
 sg13g2_decap_4 FILLER_43_348 ();
 sg13g2_fill_1 FILLER_43_365 ();
 sg13g2_fill_2 FILLER_43_371 ();
 sg13g2_fill_1 FILLER_43_373 ();
 sg13g2_fill_1 FILLER_43_401 ();
 sg13g2_fill_2 FILLER_43_415 ();
 sg13g2_fill_1 FILLER_43_417 ();
 sg13g2_fill_1 FILLER_43_448 ();
 sg13g2_fill_2 FILLER_43_483 ();
 sg13g2_fill_1 FILLER_43_493 ();
 sg13g2_decap_4 FILLER_43_525 ();
 sg13g2_fill_1 FILLER_43_529 ();
 sg13g2_fill_1 FILLER_43_567 ();
 sg13g2_fill_1 FILLER_43_585 ();
 sg13g2_fill_1 FILLER_43_594 ();
 sg13g2_fill_2 FILLER_43_598 ();
 sg13g2_fill_2 FILLER_43_609 ();
 sg13g2_fill_1 FILLER_43_619 ();
 sg13g2_fill_1 FILLER_43_673 ();
 sg13g2_fill_1 FILLER_43_708 ();
 sg13g2_fill_2 FILLER_43_713 ();
 sg13g2_fill_1 FILLER_43_719 ();
 sg13g2_fill_2 FILLER_43_724 ();
 sg13g2_fill_1 FILLER_43_735 ();
 sg13g2_fill_1 FILLER_43_740 ();
 sg13g2_fill_1 FILLER_43_749 ();
 sg13g2_fill_2 FILLER_43_765 ();
 sg13g2_fill_1 FILLER_43_776 ();
 sg13g2_fill_1 FILLER_43_781 ();
 sg13g2_fill_1 FILLER_43_787 ();
 sg13g2_fill_1 FILLER_43_792 ();
 sg13g2_fill_1 FILLER_43_803 ();
 sg13g2_fill_1 FILLER_43_808 ();
 sg13g2_fill_1 FILLER_43_837 ();
 sg13g2_fill_2 FILLER_43_841 ();
 sg13g2_fill_2 FILLER_43_875 ();
 sg13g2_fill_1 FILLER_43_877 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_40 ();
 sg13g2_fill_1 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_62 ();
 sg13g2_fill_2 FILLER_44_69 ();
 sg13g2_fill_1 FILLER_44_75 ();
 sg13g2_fill_1 FILLER_44_80 ();
 sg13g2_fill_1 FILLER_44_101 ();
 sg13g2_fill_2 FILLER_44_106 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_fill_2 FILLER_44_126 ();
 sg13g2_fill_1 FILLER_44_136 ();
 sg13g2_fill_2 FILLER_44_141 ();
 sg13g2_fill_1 FILLER_44_161 ();
 sg13g2_fill_2 FILLER_44_229 ();
 sg13g2_fill_1 FILLER_44_235 ();
 sg13g2_fill_1 FILLER_44_241 ();
 sg13g2_fill_2 FILLER_44_314 ();
 sg13g2_fill_2 FILLER_44_343 ();
 sg13g2_fill_1 FILLER_44_345 ();
 sg13g2_fill_2 FILLER_44_350 ();
 sg13g2_fill_2 FILLER_44_383 ();
 sg13g2_fill_1 FILLER_44_393 ();
 sg13g2_fill_1 FILLER_44_399 ();
 sg13g2_fill_1 FILLER_44_404 ();
 sg13g2_fill_2 FILLER_44_418 ();
 sg13g2_decap_4 FILLER_44_428 ();
 sg13g2_fill_1 FILLER_44_432 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_fill_2 FILLER_44_448 ();
 sg13g2_fill_1 FILLER_44_450 ();
 sg13g2_fill_1 FILLER_44_470 ();
 sg13g2_fill_1 FILLER_44_507 ();
 sg13g2_fill_1 FILLER_44_534 ();
 sg13g2_fill_1 FILLER_44_539 ();
 sg13g2_fill_1 FILLER_44_544 ();
 sg13g2_fill_2 FILLER_44_583 ();
 sg13g2_fill_1 FILLER_44_597 ();
 sg13g2_fill_2 FILLER_44_614 ();
 sg13g2_fill_1 FILLER_44_632 ();
 sg13g2_fill_1 FILLER_44_655 ();
 sg13g2_fill_2 FILLER_44_680 ();
 sg13g2_fill_1 FILLER_44_682 ();
 sg13g2_fill_1 FILLER_44_725 ();
 sg13g2_fill_1 FILLER_44_734 ();
 sg13g2_decap_4 FILLER_44_739 ();
 sg13g2_fill_1 FILLER_44_776 ();
 sg13g2_fill_1 FILLER_44_784 ();
 sg13g2_fill_1 FILLER_44_804 ();
 sg13g2_fill_2 FILLER_44_821 ();
 sg13g2_decap_4 FILLER_44_837 ();
 sg13g2_fill_1 FILLER_44_841 ();
 sg13g2_fill_2 FILLER_44_861 ();
 sg13g2_fill_2 FILLER_44_876 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_5 ();
 sg13g2_fill_1 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_108 ();
 sg13g2_fill_1 FILLER_45_113 ();
 sg13g2_fill_1 FILLER_45_125 ();
 sg13g2_fill_1 FILLER_45_130 ();
 sg13g2_fill_1 FILLER_45_152 ();
 sg13g2_fill_2 FILLER_45_194 ();
 sg13g2_fill_1 FILLER_45_205 ();
 sg13g2_fill_1 FILLER_45_211 ();
 sg13g2_fill_1 FILLER_45_217 ();
 sg13g2_fill_1 FILLER_45_222 ();
 sg13g2_fill_1 FILLER_45_228 ();
 sg13g2_fill_1 FILLER_45_236 ();
 sg13g2_decap_4 FILLER_45_241 ();
 sg13g2_fill_1 FILLER_45_249 ();
 sg13g2_fill_2 FILLER_45_294 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_fill_1 FILLER_45_310 ();
 sg13g2_fill_2 FILLER_45_314 ();
 sg13g2_fill_1 FILLER_45_339 ();
 sg13g2_fill_2 FILLER_45_365 ();
 sg13g2_fill_1 FILLER_45_391 ();
 sg13g2_fill_2 FILLER_45_405 ();
 sg13g2_fill_1 FILLER_45_407 ();
 sg13g2_fill_1 FILLER_45_416 ();
 sg13g2_fill_1 FILLER_45_425 ();
 sg13g2_fill_1 FILLER_45_434 ();
 sg13g2_fill_1 FILLER_45_442 ();
 sg13g2_decap_4 FILLER_45_564 ();
 sg13g2_fill_1 FILLER_45_598 ();
 sg13g2_fill_1 FILLER_45_634 ();
 sg13g2_fill_1 FILLER_45_651 ();
 sg13g2_fill_2 FILLER_45_695 ();
 sg13g2_decap_4 FILLER_45_723 ();
 sg13g2_fill_2 FILLER_45_760 ();
 sg13g2_fill_1 FILLER_45_766 ();
 sg13g2_fill_2 FILLER_45_783 ();
 sg13g2_fill_1 FILLER_45_799 ();
 sg13g2_fill_1 FILLER_45_818 ();
 sg13g2_fill_1 FILLER_45_824 ();
 sg13g2_fill_2 FILLER_45_875 ();
 sg13g2_fill_1 FILLER_45_877 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_48 ();
 sg13g2_fill_2 FILLER_46_59 ();
 sg13g2_fill_2 FILLER_46_78 ();
 sg13g2_fill_1 FILLER_46_116 ();
 sg13g2_fill_1 FILLER_46_149 ();
 sg13g2_fill_1 FILLER_46_154 ();
 sg13g2_fill_1 FILLER_46_191 ();
 sg13g2_fill_1 FILLER_46_200 ();
 sg13g2_fill_1 FILLER_46_235 ();
 sg13g2_fill_2 FILLER_46_254 ();
 sg13g2_fill_2 FILLER_46_291 ();
 sg13g2_fill_1 FILLER_46_322 ();
 sg13g2_fill_1 FILLER_46_384 ();
 sg13g2_decap_4 FILLER_46_399 ();
 sg13g2_fill_2 FILLER_46_403 ();
 sg13g2_fill_2 FILLER_46_456 ();
 sg13g2_fill_1 FILLER_46_462 ();
 sg13g2_fill_2 FILLER_46_493 ();
 sg13g2_fill_1 FILLER_46_521 ();
 sg13g2_fill_1 FILLER_46_527 ();
 sg13g2_fill_1 FILLER_46_532 ();
 sg13g2_fill_1 FILLER_46_536 ();
 sg13g2_fill_1 FILLER_46_542 ();
 sg13g2_fill_1 FILLER_46_584 ();
 sg13g2_fill_2 FILLER_46_596 ();
 sg13g2_fill_1 FILLER_46_610 ();
 sg13g2_fill_1 FILLER_46_615 ();
 sg13g2_fill_1 FILLER_46_621 ();
 sg13g2_fill_1 FILLER_46_627 ();
 sg13g2_fill_1 FILLER_46_632 ();
 sg13g2_fill_1 FILLER_46_639 ();
 sg13g2_fill_2 FILLER_46_652 ();
 sg13g2_fill_2 FILLER_46_665 ();
 sg13g2_fill_2 FILLER_46_688 ();
 sg13g2_fill_1 FILLER_46_690 ();
 sg13g2_fill_2 FILLER_46_703 ();
 sg13g2_fill_1 FILLER_46_714 ();
 sg13g2_decap_4 FILLER_46_719 ();
 sg13g2_fill_1 FILLER_46_742 ();
 sg13g2_fill_2 FILLER_46_778 ();
 sg13g2_fill_2 FILLER_46_808 ();
 sg13g2_fill_1 FILLER_46_810 ();
 sg13g2_decap_4 FILLER_46_824 ();
 sg13g2_fill_2 FILLER_46_848 ();
 sg13g2_fill_2 FILLER_46_871 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_52 ();
 sg13g2_fill_1 FILLER_47_141 ();
 sg13g2_fill_1 FILLER_47_162 ();
 sg13g2_fill_2 FILLER_47_181 ();
 sg13g2_fill_2 FILLER_47_209 ();
 sg13g2_fill_1 FILLER_47_211 ();
 sg13g2_fill_1 FILLER_47_232 ();
 sg13g2_fill_2 FILLER_47_259 ();
 sg13g2_fill_1 FILLER_47_273 ();
 sg13g2_fill_1 FILLER_47_281 ();
 sg13g2_fill_2 FILLER_47_307 ();
 sg13g2_fill_1 FILLER_47_321 ();
 sg13g2_fill_1 FILLER_47_326 ();
 sg13g2_fill_1 FILLER_47_330 ();
 sg13g2_fill_1 FILLER_47_361 ();
 sg13g2_fill_1 FILLER_47_388 ();
 sg13g2_decap_4 FILLER_47_417 ();
 sg13g2_fill_2 FILLER_47_425 ();
 sg13g2_fill_1 FILLER_47_427 ();
 sg13g2_fill_2 FILLER_47_439 ();
 sg13g2_fill_1 FILLER_47_459 ();
 sg13g2_fill_1 FILLER_47_523 ();
 sg13g2_fill_1 FILLER_47_533 ();
 sg13g2_fill_1 FILLER_47_538 ();
 sg13g2_fill_2 FILLER_47_543 ();
 sg13g2_fill_2 FILLER_47_573 ();
 sg13g2_fill_1 FILLER_47_575 ();
 sg13g2_fill_1 FILLER_47_583 ();
 sg13g2_fill_1 FILLER_47_698 ();
 sg13g2_fill_2 FILLER_47_717 ();
 sg13g2_fill_2 FILLER_47_731 ();
 sg13g2_fill_1 FILLER_47_733 ();
 sg13g2_fill_1 FILLER_47_746 ();
 sg13g2_fill_1 FILLER_47_751 ();
 sg13g2_fill_1 FILLER_47_756 ();
 sg13g2_fill_1 FILLER_47_762 ();
 sg13g2_fill_2 FILLER_47_772 ();
 sg13g2_fill_2 FILLER_47_799 ();
 sg13g2_fill_1 FILLER_47_805 ();
 sg13g2_fill_1 FILLER_47_822 ();
 sg13g2_fill_2 FILLER_47_828 ();
 sg13g2_decap_4 FILLER_47_847 ();
 sg13g2_fill_1 FILLER_47_851 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_fill_2 FILLER_47_866 ();
 sg13g2_fill_1 FILLER_47_868 ();
 sg13g2_decap_4 FILLER_47_873 ();
 sg13g2_fill_1 FILLER_47_877 ();
 sg13g2_fill_2 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_57 ();
 sg13g2_fill_1 FILLER_48_69 ();
 sg13g2_fill_2 FILLER_48_106 ();
 sg13g2_fill_1 FILLER_48_114 ();
 sg13g2_fill_1 FILLER_48_135 ();
 sg13g2_fill_1 FILLER_48_163 ();
 sg13g2_fill_1 FILLER_48_169 ();
 sg13g2_fill_1 FILLER_48_177 ();
 sg13g2_fill_2 FILLER_48_187 ();
 sg13g2_fill_2 FILLER_48_220 ();
 sg13g2_fill_1 FILLER_48_222 ();
 sg13g2_fill_1 FILLER_48_227 ();
 sg13g2_fill_2 FILLER_48_241 ();
 sg13g2_fill_1 FILLER_48_243 ();
 sg13g2_fill_1 FILLER_48_274 ();
 sg13g2_fill_1 FILLER_48_279 ();
 sg13g2_fill_2 FILLER_48_333 ();
 sg13g2_fill_1 FILLER_48_390 ();
 sg13g2_fill_1 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_414 ();
 sg13g2_fill_2 FILLER_48_421 ();
 sg13g2_fill_1 FILLER_48_439 ();
 sg13g2_decap_4 FILLER_48_444 ();
 sg13g2_fill_1 FILLER_48_448 ();
 sg13g2_fill_1 FILLER_48_470 ();
 sg13g2_fill_1 FILLER_48_524 ();
 sg13g2_fill_2 FILLER_48_559 ();
 sg13g2_fill_1 FILLER_48_617 ();
 sg13g2_fill_1 FILLER_48_623 ();
 sg13g2_fill_1 FILLER_48_628 ();
 sg13g2_fill_1 FILLER_48_634 ();
 sg13g2_fill_2 FILLER_48_647 ();
 sg13g2_fill_1 FILLER_48_653 ();
 sg13g2_fill_1 FILLER_48_659 ();
 sg13g2_fill_2 FILLER_48_733 ();
 sg13g2_fill_1 FILLER_48_735 ();
 sg13g2_fill_1 FILLER_48_764 ();
 sg13g2_fill_2 FILLER_48_769 ();
 sg13g2_fill_1 FILLER_48_771 ();
 sg13g2_fill_1 FILLER_48_788 ();
 sg13g2_fill_1 FILLER_48_797 ();
 sg13g2_fill_1 FILLER_48_806 ();
 sg13g2_decap_4 FILLER_48_841 ();
 sg13g2_fill_2 FILLER_49_20 ();
 sg13g2_fill_1 FILLER_49_39 ();
 sg13g2_fill_1 FILLER_49_148 ();
 sg13g2_fill_1 FILLER_49_154 ();
 sg13g2_fill_1 FILLER_49_185 ();
 sg13g2_fill_1 FILLER_49_189 ();
 sg13g2_fill_1 FILLER_49_211 ();
 sg13g2_fill_2 FILLER_49_232 ();
 sg13g2_fill_1 FILLER_49_242 ();
 sg13g2_fill_1 FILLER_49_264 ();
 sg13g2_fill_2 FILLER_49_274 ();
 sg13g2_fill_2 FILLER_49_284 ();
 sg13g2_fill_2 FILLER_49_332 ();
 sg13g2_decap_4 FILLER_49_365 ();
 sg13g2_fill_2 FILLER_49_401 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_fill_1 FILLER_49_409 ();
 sg13g2_fill_1 FILLER_49_415 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_4 FILLER_49_427 ();
 sg13g2_fill_2 FILLER_49_443 ();
 sg13g2_decap_4 FILLER_49_458 ();
 sg13g2_fill_1 FILLER_49_462 ();
 sg13g2_fill_1 FILLER_49_479 ();
 sg13g2_fill_1 FILLER_49_509 ();
 sg13g2_fill_1 FILLER_49_518 ();
 sg13g2_fill_2 FILLER_49_545 ();
 sg13g2_fill_1 FILLER_49_547 ();
 sg13g2_decap_4 FILLER_49_551 ();
 sg13g2_fill_1 FILLER_49_555 ();
 sg13g2_fill_2 FILLER_49_596 ();
 sg13g2_fill_2 FILLER_49_608 ();
 sg13g2_fill_2 FILLER_49_639 ();
 sg13g2_fill_1 FILLER_49_645 ();
 sg13g2_fill_1 FILLER_49_650 ();
 sg13g2_fill_2 FILLER_49_655 ();
 sg13g2_fill_2 FILLER_49_666 ();
 sg13g2_fill_2 FILLER_49_714 ();
 sg13g2_fill_1 FILLER_49_716 ();
 sg13g2_decap_4 FILLER_49_722 ();
 sg13g2_fill_2 FILLER_49_760 ();
 sg13g2_fill_1 FILLER_49_785 ();
 sg13g2_fill_1 FILLER_49_791 ();
 sg13g2_fill_2 FILLER_49_815 ();
 sg13g2_fill_1 FILLER_49_843 ();
 sg13g2_fill_2 FILLER_49_852 ();
 sg13g2_decap_8 FILLER_49_870 ();
 sg13g2_fill_1 FILLER_49_877 ();
 sg13g2_fill_2 FILLER_50_30 ();
 sg13g2_fill_1 FILLER_50_54 ();
 sg13g2_fill_2 FILLER_50_86 ();
 sg13g2_decap_8 FILLER_50_114 ();
 sg13g2_decap_4 FILLER_50_121 ();
 sg13g2_fill_1 FILLER_50_169 ();
 sg13g2_fill_1 FILLER_50_202 ();
 sg13g2_decap_8 FILLER_50_235 ();
 sg13g2_fill_1 FILLER_50_258 ();
 sg13g2_fill_1 FILLER_50_299 ();
 sg13g2_fill_1 FILLER_50_311 ();
 sg13g2_fill_2 FILLER_50_323 ();
 sg13g2_fill_1 FILLER_50_333 ();
 sg13g2_fill_1 FILLER_50_342 ();
 sg13g2_fill_2 FILLER_50_351 ();
 sg13g2_fill_1 FILLER_50_353 ();
 sg13g2_fill_2 FILLER_50_382 ();
 sg13g2_fill_1 FILLER_50_389 ();
 sg13g2_fill_1 FILLER_50_394 ();
 sg13g2_fill_1 FILLER_50_399 ();
 sg13g2_fill_1 FILLER_50_405 ();
 sg13g2_fill_1 FILLER_50_425 ();
 sg13g2_fill_2 FILLER_50_436 ();
 sg13g2_fill_2 FILLER_50_492 ();
 sg13g2_fill_1 FILLER_50_497 ();
 sg13g2_fill_1 FILLER_50_506 ();
 sg13g2_decap_8 FILLER_50_511 ();
 sg13g2_fill_2 FILLER_50_518 ();
 sg13g2_fill_2 FILLER_50_523 ();
 sg13g2_fill_2 FILLER_50_550 ();
 sg13g2_fill_1 FILLER_50_552 ();
 sg13g2_fill_2 FILLER_50_559 ();
 sg13g2_fill_1 FILLER_50_561 ();
 sg13g2_fill_1 FILLER_50_612 ();
 sg13g2_fill_1 FILLER_50_646 ();
 sg13g2_fill_2 FILLER_50_650 ();
 sg13g2_fill_2 FILLER_50_678 ();
 sg13g2_fill_1 FILLER_50_680 ();
 sg13g2_decap_4 FILLER_50_689 ();
 sg13g2_fill_2 FILLER_50_693 ();
 sg13g2_fill_1 FILLER_50_704 ();
 sg13g2_fill_1 FILLER_50_735 ();
 sg13g2_fill_1 FILLER_50_749 ();
 sg13g2_fill_1 FILLER_50_754 ();
 sg13g2_fill_2 FILLER_50_760 ();
 sg13g2_fill_2 FILLER_50_775 ();
 sg13g2_fill_1 FILLER_50_777 ();
 sg13g2_fill_2 FILLER_50_782 ();
 sg13g2_fill_1 FILLER_50_784 ();
 sg13g2_fill_2 FILLER_50_790 ();
 sg13g2_fill_2 FILLER_50_796 ();
 sg13g2_decap_8 FILLER_50_813 ();
 sg13g2_decap_4 FILLER_50_833 ();
 sg13g2_fill_2 FILLER_50_841 ();
 sg13g2_decap_4 FILLER_50_865 ();
 sg13g2_fill_1 FILLER_50_877 ();
 sg13g2_fill_1 FILLER_51_58 ();
 sg13g2_fill_1 FILLER_51_80 ();
 sg13g2_fill_2 FILLER_51_137 ();
 sg13g2_fill_1 FILLER_51_143 ();
 sg13g2_fill_2 FILLER_51_152 ();
 sg13g2_fill_1 FILLER_51_209 ();
 sg13g2_fill_1 FILLER_51_222 ();
 sg13g2_decap_4 FILLER_51_231 ();
 sg13g2_fill_1 FILLER_51_264 ();
 sg13g2_fill_1 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_291 ();
 sg13g2_fill_1 FILLER_51_300 ();
 sg13g2_fill_2 FILLER_51_337 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_decap_4 FILLER_51_366 ();
 sg13g2_fill_2 FILLER_51_370 ();
 sg13g2_fill_1 FILLER_51_409 ();
 sg13g2_fill_1 FILLER_51_414 ();
 sg13g2_fill_1 FILLER_51_439 ();
 sg13g2_fill_1 FILLER_51_444 ();
 sg13g2_fill_1 FILLER_51_453 ();
 sg13g2_fill_1 FILLER_51_458 ();
 sg13g2_fill_1 FILLER_51_463 ();
 sg13g2_fill_1 FILLER_51_467 ();
 sg13g2_fill_1 FILLER_51_473 ();
 sg13g2_decap_8 FILLER_51_509 ();
 sg13g2_decap_4 FILLER_51_520 ();
 sg13g2_decap_4 FILLER_51_536 ();
 sg13g2_fill_1 FILLER_51_548 ();
 sg13g2_fill_2 FILLER_51_575 ();
 sg13g2_fill_1 FILLER_51_589 ();
 sg13g2_fill_2 FILLER_51_622 ();
 sg13g2_fill_2 FILLER_51_632 ();
 sg13g2_fill_1 FILLER_51_634 ();
 sg13g2_fill_2 FILLER_51_663 ();
 sg13g2_fill_2 FILLER_51_673 ();
 sg13g2_fill_2 FILLER_51_679 ();
 sg13g2_fill_1 FILLER_51_681 ();
 sg13g2_decap_4 FILLER_51_711 ();
 sg13g2_decap_4 FILLER_51_724 ();
 sg13g2_fill_1 FILLER_51_728 ();
 sg13g2_decap_8 FILLER_51_734 ();
 sg13g2_fill_1 FILLER_51_741 ();
 sg13g2_decap_8 FILLER_51_746 ();
 sg13g2_decap_4 FILLER_51_753 ();
 sg13g2_fill_2 FILLER_51_757 ();
 sg13g2_fill_1 FILLER_51_785 ();
 sg13g2_decap_4 FILLER_51_794 ();
 sg13g2_fill_2 FILLER_51_798 ();
 sg13g2_decap_4 FILLER_51_805 ();
 sg13g2_fill_2 FILLER_51_813 ();
 sg13g2_fill_1 FILLER_51_837 ();
 sg13g2_fill_1 FILLER_51_846 ();
 sg13g2_fill_1 FILLER_51_855 ();
 sg13g2_fill_2 FILLER_51_869 ();
 sg13g2_fill_2 FILLER_51_875 ();
 sg13g2_fill_1 FILLER_51_877 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_45 ();
 sg13g2_fill_1 FILLER_52_72 ();
 sg13g2_fill_2 FILLER_52_117 ();
 sg13g2_fill_1 FILLER_52_127 ();
 sg13g2_fill_2 FILLER_52_162 ();
 sg13g2_fill_1 FILLER_52_164 ();
 sg13g2_fill_2 FILLER_52_283 ();
 sg13g2_fill_1 FILLER_52_367 ();
 sg13g2_fill_1 FILLER_52_376 ();
 sg13g2_fill_1 FILLER_52_383 ();
 sg13g2_fill_1 FILLER_52_388 ();
 sg13g2_fill_1 FILLER_52_399 ();
 sg13g2_fill_1 FILLER_52_409 ();
 sg13g2_fill_1 FILLER_52_430 ();
 sg13g2_fill_1 FILLER_52_440 ();
 sg13g2_fill_2 FILLER_52_489 ();
 sg13g2_fill_1 FILLER_52_491 ();
 sg13g2_fill_1 FILLER_52_495 ();
 sg13g2_fill_1 FILLER_52_501 ();
 sg13g2_fill_1 FILLER_52_507 ();
 sg13g2_fill_1 FILLER_52_519 ();
 sg13g2_fill_1 FILLER_52_524 ();
 sg13g2_fill_1 FILLER_52_546 ();
 sg13g2_decap_4 FILLER_52_595 ();
 sg13g2_decap_8 FILLER_52_603 ();
 sg13g2_fill_1 FILLER_52_610 ();
 sg13g2_decap_4 FILLER_52_620 ();
 sg13g2_fill_1 FILLER_52_674 ();
 sg13g2_fill_1 FILLER_52_680 ();
 sg13g2_fill_1 FILLER_52_686 ();
 sg13g2_fill_2 FILLER_52_695 ();
 sg13g2_fill_2 FILLER_52_733 ();
 sg13g2_fill_1 FILLER_52_735 ();
 sg13g2_fill_1 FILLER_52_742 ();
 sg13g2_fill_1 FILLER_52_747 ();
 sg13g2_fill_1 FILLER_52_752 ();
 sg13g2_fill_1 FILLER_52_757 ();
 sg13g2_fill_2 FILLER_52_762 ();
 sg13g2_fill_2 FILLER_52_785 ();
 sg13g2_decap_8 FILLER_52_793 ();
 sg13g2_fill_1 FILLER_52_825 ();
 sg13g2_fill_1 FILLER_52_833 ();
 sg13g2_fill_1 FILLER_52_850 ();
 sg13g2_fill_1 FILLER_52_856 ();
 sg13g2_fill_1 FILLER_52_865 ();
 sg13g2_fill_1 FILLER_52_871 ();
 sg13g2_fill_2 FILLER_52_876 ();
 sg13g2_fill_1 FILLER_53_61 ();
 sg13g2_fill_2 FILLER_53_88 ();
 sg13g2_fill_1 FILLER_53_114 ();
 sg13g2_fill_2 FILLER_53_135 ();
 sg13g2_fill_1 FILLER_53_137 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_decap_8 FILLER_53_205 ();
 sg13g2_fill_1 FILLER_53_212 ();
 sg13g2_fill_2 FILLER_53_237 ();
 sg13g2_fill_1 FILLER_53_239 ();
 sg13g2_fill_2 FILLER_53_303 ();
 sg13g2_fill_2 FILLER_53_318 ();
 sg13g2_fill_1 FILLER_53_324 ();
 sg13g2_fill_2 FILLER_53_351 ();
 sg13g2_fill_2 FILLER_53_365 ();
 sg13g2_fill_1 FILLER_53_367 ();
 sg13g2_fill_1 FILLER_53_376 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_decap_4 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_410 ();
 sg13g2_fill_1 FILLER_53_415 ();
 sg13g2_fill_1 FILLER_53_420 ();
 sg13g2_fill_1 FILLER_53_458 ();
 sg13g2_fill_1 FILLER_53_492 ();
 sg13g2_fill_1 FILLER_53_497 ();
 sg13g2_fill_1 FILLER_53_502 ();
 sg13g2_fill_2 FILLER_53_507 ();
 sg13g2_fill_1 FILLER_53_529 ();
 sg13g2_decap_4 FILLER_53_538 ();
 sg13g2_fill_1 FILLER_53_542 ();
 sg13g2_fill_2 FILLER_53_547 ();
 sg13g2_fill_1 FILLER_53_566 ();
 sg13g2_fill_1 FILLER_53_570 ();
 sg13g2_fill_1 FILLER_53_575 ();
 sg13g2_fill_1 FILLER_53_580 ();
 sg13g2_fill_1 FILLER_53_585 ();
 sg13g2_fill_1 FILLER_53_590 ();
 sg13g2_fill_2 FILLER_53_594 ();
 sg13g2_fill_1 FILLER_53_596 ();
 sg13g2_fill_2 FILLER_53_601 ();
 sg13g2_fill_1 FILLER_53_650 ();
 sg13g2_fill_2 FILLER_53_698 ();
 sg13g2_fill_1 FILLER_53_704 ();
 sg13g2_decap_4 FILLER_53_739 ();
 sg13g2_fill_2 FILLER_53_743 ();
 sg13g2_fill_1 FILLER_53_782 ();
 sg13g2_fill_1 FILLER_53_787 ();
 sg13g2_decap_8 FILLER_53_814 ();
 sg13g2_decap_8 FILLER_53_821 ();
 sg13g2_fill_2 FILLER_53_828 ();
 sg13g2_fill_1 FILLER_53_834 ();
 sg13g2_fill_1 FILLER_53_873 ();
 sg13g2_fill_1 FILLER_54_30 ();
 sg13g2_fill_1 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_54 ();
 sg13g2_fill_1 FILLER_54_119 ();
 sg13g2_fill_2 FILLER_54_138 ();
 sg13g2_fill_1 FILLER_54_175 ();
 sg13g2_fill_1 FILLER_54_194 ();
 sg13g2_fill_1 FILLER_54_234 ();
 sg13g2_fill_1 FILLER_54_240 ();
 sg13g2_fill_1 FILLER_54_267 ();
 sg13g2_fill_1 FILLER_54_271 ();
 sg13g2_fill_1 FILLER_54_279 ();
 sg13g2_fill_2 FILLER_54_325 ();
 sg13g2_fill_1 FILLER_54_335 ();
 sg13g2_fill_2 FILLER_54_366 ();
 sg13g2_decap_4 FILLER_54_384 ();
 sg13g2_fill_2 FILLER_54_434 ();
 sg13g2_fill_1 FILLER_54_436 ();
 sg13g2_fill_1 FILLER_54_463 ();
 sg13g2_fill_2 FILLER_54_469 ();
 sg13g2_fill_1 FILLER_54_476 ();
 sg13g2_fill_2 FILLER_54_482 ();
 sg13g2_fill_1 FILLER_54_489 ();
 sg13g2_fill_1 FILLER_54_495 ();
 sg13g2_fill_2 FILLER_54_500 ();
 sg13g2_fill_2 FILLER_54_507 ();
 sg13g2_fill_2 FILLER_54_535 ();
 sg13g2_fill_1 FILLER_54_542 ();
 sg13g2_fill_1 FILLER_54_554 ();
 sg13g2_fill_1 FILLER_54_576 ();
 sg13g2_decap_4 FILLER_54_588 ();
 sg13g2_fill_1 FILLER_54_592 ();
 sg13g2_fill_1 FILLER_54_602 ();
 sg13g2_fill_2 FILLER_54_620 ();
 sg13g2_fill_1 FILLER_54_629 ();
 sg13g2_fill_2 FILLER_54_640 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_2 FILLER_54_676 ();
 sg13g2_fill_2 FILLER_54_683 ();
 sg13g2_fill_1 FILLER_54_750 ();
 sg13g2_fill_1 FILLER_54_759 ();
 sg13g2_fill_1 FILLER_54_768 ();
 sg13g2_fill_1 FILLER_54_777 ();
 sg13g2_fill_2 FILLER_54_796 ();
 sg13g2_fill_1 FILLER_54_798 ();
 sg13g2_fill_2 FILLER_54_819 ();
 sg13g2_fill_1 FILLER_54_821 ();
 sg13g2_fill_1 FILLER_54_835 ();
 sg13g2_fill_1 FILLER_54_840 ();
 sg13g2_fill_2 FILLER_54_865 ();
 sg13g2_fill_2 FILLER_54_872 ();
 sg13g2_fill_1 FILLER_54_877 ();
 sg13g2_fill_1 FILLER_55_17 ();
 sg13g2_fill_1 FILLER_55_47 ();
 sg13g2_fill_1 FILLER_55_83 ();
 sg13g2_fill_1 FILLER_55_89 ();
 sg13g2_fill_2 FILLER_55_123 ();
 sg13g2_fill_1 FILLER_55_132 ();
 sg13g2_fill_2 FILLER_55_169 ();
 sg13g2_fill_1 FILLER_55_176 ();
 sg13g2_fill_1 FILLER_55_185 ();
 sg13g2_fill_2 FILLER_55_189 ();
 sg13g2_fill_2 FILLER_55_212 ();
 sg13g2_fill_2 FILLER_55_245 ();
 sg13g2_fill_1 FILLER_55_247 ();
 sg13g2_fill_2 FILLER_55_256 ();
 sg13g2_decap_4 FILLER_55_263 ();
 sg13g2_fill_1 FILLER_55_289 ();
 sg13g2_fill_1 FILLER_55_293 ();
 sg13g2_fill_2 FILLER_55_308 ();
 sg13g2_fill_1 FILLER_55_310 ();
 sg13g2_fill_2 FILLER_55_341 ();
 sg13g2_fill_2 FILLER_55_347 ();
 sg13g2_fill_1 FILLER_55_369 ();
 sg13g2_fill_1 FILLER_55_374 ();
 sg13g2_fill_1 FILLER_55_380 ();
 sg13g2_fill_1 FILLER_55_384 ();
 sg13g2_fill_1 FILLER_55_389 ();
 sg13g2_fill_2 FILLER_55_446 ();
 sg13g2_fill_2 FILLER_55_469 ();
 sg13g2_decap_4 FILLER_55_483 ();
 sg13g2_fill_2 FILLER_55_487 ();
 sg13g2_fill_2 FILLER_55_494 ();
 sg13g2_fill_1 FILLER_55_500 ();
 sg13g2_fill_2 FILLER_55_505 ();
 sg13g2_fill_1 FILLER_55_511 ();
 sg13g2_fill_2 FILLER_55_517 ();
 sg13g2_fill_1 FILLER_55_519 ();
 sg13g2_fill_2 FILLER_55_528 ();
 sg13g2_fill_1 FILLER_55_530 ();
 sg13g2_decap_4 FILLER_55_553 ();
 sg13g2_fill_1 FILLER_55_561 ();
 sg13g2_decap_8 FILLER_55_578 ();
 sg13g2_fill_1 FILLER_55_585 ();
 sg13g2_fill_2 FILLER_55_639 ();
 sg13g2_fill_2 FILLER_55_678 ();
 sg13g2_fill_2 FILLER_55_691 ();
 sg13g2_fill_1 FILLER_55_697 ();
 sg13g2_fill_2 FILLER_55_718 ();
 sg13g2_fill_2 FILLER_55_724 ();
 sg13g2_fill_1 FILLER_55_756 ();
 sg13g2_fill_1 FILLER_55_762 ();
 sg13g2_fill_1 FILLER_55_788 ();
 sg13g2_fill_2 FILLER_55_793 ();
 sg13g2_fill_1 FILLER_55_795 ();
 sg13g2_fill_1 FILLER_55_827 ();
 sg13g2_fill_1 FILLER_55_845 ();
 sg13g2_fill_2 FILLER_55_876 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_31 ();
 sg13g2_fill_2 FILLER_56_112 ();
 sg13g2_fill_2 FILLER_56_140 ();
 sg13g2_fill_2 FILLER_56_184 ();
 sg13g2_fill_2 FILLER_56_223 ();
 sg13g2_fill_1 FILLER_56_229 ();
 sg13g2_fill_1 FILLER_56_233 ();
 sg13g2_decap_4 FILLER_56_250 ();
 sg13g2_fill_1 FILLER_56_267 ();
 sg13g2_fill_2 FILLER_56_285 ();
 sg13g2_decap_4 FILLER_56_308 ();
 sg13g2_fill_1 FILLER_56_312 ();
 sg13g2_fill_2 FILLER_56_321 ();
 sg13g2_fill_2 FILLER_56_331 ();
 sg13g2_fill_2 FILLER_56_337 ();
 sg13g2_fill_2 FILLER_56_343 ();
 sg13g2_fill_2 FILLER_56_349 ();
 sg13g2_fill_1 FILLER_56_351 ();
 sg13g2_fill_1 FILLER_56_385 ();
 sg13g2_fill_1 FILLER_56_391 ();
 sg13g2_fill_1 FILLER_56_396 ();
 sg13g2_decap_4 FILLER_56_415 ();
 sg13g2_fill_1 FILLER_56_424 ();
 sg13g2_fill_1 FILLER_56_430 ();
 sg13g2_fill_1 FILLER_56_435 ();
 sg13g2_fill_1 FILLER_56_440 ();
 sg13g2_decap_4 FILLER_56_475 ();
 sg13g2_fill_1 FILLER_56_488 ();
 sg13g2_fill_1 FILLER_56_493 ();
 sg13g2_fill_1 FILLER_56_499 ();
 sg13g2_fill_2 FILLER_56_527 ();
 sg13g2_fill_1 FILLER_56_541 ();
 sg13g2_fill_1 FILLER_56_546 ();
 sg13g2_fill_1 FILLER_56_555 ();
 sg13g2_fill_2 FILLER_56_560 ();
 sg13g2_fill_1 FILLER_56_566 ();
 sg13g2_fill_1 FILLER_56_571 ();
 sg13g2_decap_8 FILLER_56_584 ();
 sg13g2_decap_8 FILLER_56_591 ();
 sg13g2_fill_2 FILLER_56_598 ();
 sg13g2_fill_1 FILLER_56_626 ();
 sg13g2_fill_1 FILLER_56_635 ();
 sg13g2_fill_1 FILLER_56_649 ();
 sg13g2_fill_2 FILLER_56_672 ();
 sg13g2_fill_1 FILLER_56_678 ();
 sg13g2_fill_1 FILLER_56_691 ();
 sg13g2_fill_2 FILLER_56_705 ();
 sg13g2_decap_8 FILLER_56_716 ();
 sg13g2_fill_2 FILLER_56_726 ();
 sg13g2_fill_1 FILLER_56_728 ();
 sg13g2_fill_2 FILLER_56_736 ();
 sg13g2_fill_1 FILLER_56_738 ();
 sg13g2_decap_4 FILLER_56_747 ();
 sg13g2_fill_1 FILLER_56_755 ();
 sg13g2_fill_2 FILLER_56_765 ();
 sg13g2_fill_2 FILLER_56_771 ();
 sg13g2_fill_1 FILLER_56_785 ();
 sg13g2_fill_1 FILLER_56_844 ();
 sg13g2_fill_2 FILLER_56_875 ();
 sg13g2_fill_1 FILLER_56_877 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_45 ();
 sg13g2_fill_1 FILLER_57_61 ();
 sg13g2_fill_1 FILLER_57_86 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_fill_1 FILLER_57_162 ();
 sg13g2_fill_1 FILLER_57_172 ();
 sg13g2_fill_1 FILLER_57_177 ();
 sg13g2_fill_2 FILLER_57_183 ();
 sg13g2_fill_2 FILLER_57_198 ();
 sg13g2_fill_1 FILLER_57_200 ();
 sg13g2_fill_2 FILLER_57_220 ();
 sg13g2_fill_1 FILLER_57_280 ();
 sg13g2_decap_4 FILLER_57_297 ();
 sg13g2_fill_1 FILLER_57_309 ();
 sg13g2_fill_2 FILLER_57_343 ();
 sg13g2_fill_2 FILLER_57_362 ();
 sg13g2_fill_2 FILLER_57_386 ();
 sg13g2_fill_2 FILLER_57_413 ();
 sg13g2_fill_1 FILLER_57_426 ();
 sg13g2_fill_1 FILLER_57_432 ();
 sg13g2_decap_4 FILLER_57_438 ();
 sg13g2_fill_2 FILLER_57_463 ();
 sg13g2_fill_2 FILLER_57_469 ();
 sg13g2_fill_2 FILLER_57_476 ();
 sg13g2_fill_2 FILLER_57_494 ();
 sg13g2_fill_1 FILLER_57_496 ();
 sg13g2_fill_2 FILLER_57_502 ();
 sg13g2_fill_1 FILLER_57_504 ();
 sg13g2_fill_2 FILLER_57_532 ();
 sg13g2_fill_2 FILLER_57_579 ();
 sg13g2_fill_2 FILLER_57_590 ();
 sg13g2_fill_1 FILLER_57_600 ();
 sg13g2_fill_1 FILLER_57_606 ();
 sg13g2_fill_1 FILLER_57_611 ();
 sg13g2_decap_4 FILLER_57_616 ();
 sg13g2_fill_1 FILLER_57_624 ();
 sg13g2_fill_2 FILLER_57_664 ();
 sg13g2_fill_1 FILLER_57_682 ();
 sg13g2_fill_2 FILLER_57_695 ();
 sg13g2_fill_1 FILLER_57_697 ();
 sg13g2_fill_2 FILLER_57_743 ();
 sg13g2_fill_1 FILLER_57_749 ();
 sg13g2_fill_2 FILLER_57_777 ();
 sg13g2_fill_1 FILLER_57_819 ();
 sg13g2_decap_8 FILLER_57_870 ();
 sg13g2_fill_1 FILLER_57_877 ();
 sg13g2_fill_1 FILLER_58_26 ();
 sg13g2_fill_1 FILLER_58_40 ();
 sg13g2_fill_1 FILLER_58_84 ();
 sg13g2_fill_1 FILLER_58_124 ();
 sg13g2_fill_1 FILLER_58_129 ();
 sg13g2_fill_1 FILLER_58_143 ();
 sg13g2_fill_1 FILLER_58_156 ();
 sg13g2_fill_1 FILLER_58_196 ();
 sg13g2_fill_1 FILLER_58_233 ();
 sg13g2_fill_1 FILLER_58_237 ();
 sg13g2_fill_1 FILLER_58_243 ();
 sg13g2_fill_1 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_258 ();
 sg13g2_fill_1 FILLER_58_263 ();
 sg13g2_fill_1 FILLER_58_293 ();
 sg13g2_fill_2 FILLER_58_298 ();
 sg13g2_fill_1 FILLER_58_311 ();
 sg13g2_fill_2 FILLER_58_316 ();
 sg13g2_fill_1 FILLER_58_326 ();
 sg13g2_fill_2 FILLER_58_335 ();
 sg13g2_fill_1 FILLER_58_362 ();
 sg13g2_fill_1 FILLER_58_367 ();
 sg13g2_fill_1 FILLER_58_372 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_2 FILLER_58_410 ();
 sg13g2_fill_1 FILLER_58_421 ();
 sg13g2_fill_2 FILLER_58_441 ();
 sg13g2_fill_1 FILLER_58_451 ();
 sg13g2_fill_1 FILLER_58_455 ();
 sg13g2_fill_1 FILLER_58_460 ();
 sg13g2_fill_2 FILLER_58_509 ();
 sg13g2_fill_1 FILLER_58_529 ();
 sg13g2_decap_4 FILLER_58_534 ();
 sg13g2_fill_2 FILLER_58_567 ();
 sg13g2_fill_1 FILLER_58_574 ();
 sg13g2_fill_1 FILLER_58_579 ();
 sg13g2_fill_1 FILLER_58_584 ();
 sg13g2_fill_2 FILLER_58_590 ();
 sg13g2_fill_2 FILLER_58_604 ();
 sg13g2_fill_1 FILLER_58_606 ();
 sg13g2_fill_1 FILLER_58_616 ();
 sg13g2_fill_2 FILLER_58_620 ();
 sg13g2_fill_1 FILLER_58_622 ();
 sg13g2_fill_1 FILLER_58_647 ();
 sg13g2_fill_2 FILLER_58_662 ();
 sg13g2_fill_2 FILLER_58_697 ();
 sg13g2_fill_1 FILLER_58_699 ();
 sg13g2_fill_2 FILLER_58_721 ();
 sg13g2_fill_2 FILLER_58_850 ();
 sg13g2_fill_1 FILLER_59_70 ();
 sg13g2_fill_1 FILLER_59_122 ();
 sg13g2_fill_1 FILLER_59_126 ();
 sg13g2_fill_1 FILLER_59_178 ();
 sg13g2_fill_1 FILLER_59_186 ();
 sg13g2_fill_1 FILLER_59_196 ();
 sg13g2_fill_2 FILLER_59_244 ();
 sg13g2_fill_1 FILLER_59_250 ();
 sg13g2_fill_1 FILLER_59_309 ();
 sg13g2_fill_1 FILLER_59_318 ();
 sg13g2_fill_1 FILLER_59_327 ();
 sg13g2_fill_2 FILLER_59_334 ();
 sg13g2_fill_1 FILLER_59_362 ();
 sg13g2_fill_1 FILLER_59_375 ();
 sg13g2_decap_8 FILLER_59_391 ();
 sg13g2_fill_1 FILLER_59_398 ();
 sg13g2_fill_2 FILLER_59_412 ();
 sg13g2_fill_1 FILLER_59_419 ();
 sg13g2_fill_1 FILLER_59_424 ();
 sg13g2_fill_2 FILLER_59_449 ();
 sg13g2_fill_2 FILLER_59_482 ();
 sg13g2_fill_1 FILLER_59_488 ();
 sg13g2_fill_2 FILLER_59_493 ();
 sg13g2_fill_1 FILLER_59_549 ();
 sg13g2_fill_2 FILLER_59_563 ();
 sg13g2_fill_2 FILLER_59_573 ();
 sg13g2_fill_2 FILLER_59_583 ();
 sg13g2_fill_2 FILLER_59_589 ();
 sg13g2_decap_4 FILLER_59_594 ();
 sg13g2_fill_1 FILLER_59_598 ();
 sg13g2_decap_8 FILLER_59_628 ();
 sg13g2_decap_4 FILLER_59_635 ();
 sg13g2_fill_1 FILLER_59_643 ();
 sg13g2_decap_4 FILLER_59_739 ();
 sg13g2_fill_2 FILLER_59_743 ();
 sg13g2_fill_1 FILLER_59_750 ();
 sg13g2_fill_1 FILLER_59_755 ();
 sg13g2_fill_1 FILLER_59_760 ();
 sg13g2_fill_1 FILLER_59_765 ();
 sg13g2_fill_1 FILLER_59_770 ();
 sg13g2_fill_1 FILLER_59_797 ();
 sg13g2_fill_1 FILLER_59_802 ();
 sg13g2_fill_2 FILLER_59_820 ();
 sg13g2_fill_2 FILLER_59_868 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_126 ();
 sg13g2_fill_1 FILLER_60_154 ();
 sg13g2_fill_1 FILLER_60_188 ();
 sg13g2_decap_4 FILLER_60_210 ();
 sg13g2_fill_2 FILLER_60_244 ();
 sg13g2_fill_1 FILLER_60_257 ();
 sg13g2_decap_4 FILLER_60_266 ();
 sg13g2_fill_1 FILLER_60_270 ();
 sg13g2_fill_1 FILLER_60_304 ();
 sg13g2_fill_2 FILLER_60_334 ();
 sg13g2_fill_2 FILLER_60_355 ();
 sg13g2_decap_4 FILLER_60_405 ();
 sg13g2_fill_1 FILLER_60_426 ();
 sg13g2_fill_1 FILLER_60_431 ();
 sg13g2_decap_4 FILLER_60_441 ();
 sg13g2_fill_1 FILLER_60_458 ();
 sg13g2_fill_1 FILLER_60_464 ();
 sg13g2_fill_1 FILLER_60_475 ();
 sg13g2_fill_1 FILLER_60_483 ();
 sg13g2_fill_2 FILLER_60_493 ();
 sg13g2_fill_1 FILLER_60_495 ();
 sg13g2_fill_2 FILLER_60_520 ();
 sg13g2_fill_2 FILLER_60_544 ();
 sg13g2_fill_2 FILLER_60_564 ();
 sg13g2_fill_2 FILLER_60_571 ();
 sg13g2_fill_2 FILLER_60_603 ();
 sg13g2_fill_2 FILLER_60_609 ();
 sg13g2_fill_2 FILLER_60_628 ();
 sg13g2_fill_1 FILLER_60_630 ();
 sg13g2_fill_1 FILLER_60_640 ();
 sg13g2_fill_1 FILLER_60_646 ();
 sg13g2_fill_2 FILLER_60_659 ();
 sg13g2_fill_1 FILLER_60_666 ();
 sg13g2_decap_8 FILLER_60_685 ();
 sg13g2_fill_2 FILLER_60_705 ();
 sg13g2_fill_1 FILLER_60_707 ();
 sg13g2_fill_2 FILLER_60_716 ();
 sg13g2_fill_1 FILLER_60_718 ();
 sg13g2_fill_1 FILLER_60_779 ();
 sg13g2_fill_2 FILLER_60_802 ();
 sg13g2_fill_1 FILLER_60_847 ();
 sg13g2_fill_2 FILLER_61_54 ();
 sg13g2_fill_2 FILLER_61_66 ();
 sg13g2_fill_2 FILLER_61_177 ();
 sg13g2_decap_4 FILLER_61_191 ();
 sg13g2_fill_1 FILLER_61_195 ();
 sg13g2_fill_2 FILLER_61_228 ();
 sg13g2_fill_2 FILLER_61_264 ();
 sg13g2_fill_1 FILLER_61_277 ();
 sg13g2_fill_2 FILLER_61_353 ();
 sg13g2_fill_1 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_383 ();
 sg13g2_fill_2 FILLER_61_390 ();
 sg13g2_fill_1 FILLER_61_405 ();
 sg13g2_fill_1 FILLER_61_425 ();
 sg13g2_decap_4 FILLER_61_440 ();
 sg13g2_fill_1 FILLER_61_449 ();
 sg13g2_fill_1 FILLER_61_471 ();
 sg13g2_fill_1 FILLER_61_502 ();
 sg13g2_fill_2 FILLER_61_516 ();
 sg13g2_fill_1 FILLER_61_526 ();
 sg13g2_fill_1 FILLER_61_540 ();
 sg13g2_fill_2 FILLER_61_554 ();
 sg13g2_fill_1 FILLER_61_556 ();
 sg13g2_fill_2 FILLER_61_583 ();
 sg13g2_fill_2 FILLER_61_589 ();
 sg13g2_fill_2 FILLER_61_595 ();
 sg13g2_fill_1 FILLER_61_597 ();
 sg13g2_fill_1 FILLER_61_602 ();
 sg13g2_fill_2 FILLER_61_608 ();
 sg13g2_fill_1 FILLER_61_610 ();
 sg13g2_fill_2 FILLER_61_624 ();
 sg13g2_decap_8 FILLER_61_709 ();
 sg13g2_fill_1 FILLER_61_716 ();
 sg13g2_fill_1 FILLER_61_791 ();
 sg13g2_fill_1 FILLER_61_798 ();
 sg13g2_fill_2 FILLER_61_810 ();
 sg13g2_fill_2 FILLER_61_847 ();
 sg13g2_fill_2 FILLER_61_856 ();
 sg13g2_decap_4 FILLER_61_874 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_40 ();
 sg13g2_fill_2 FILLER_62_80 ();
 sg13g2_fill_1 FILLER_62_140 ();
 sg13g2_fill_1 FILLER_62_168 ();
 sg13g2_fill_1 FILLER_62_217 ();
 sg13g2_fill_1 FILLER_62_228 ();
 sg13g2_fill_2 FILLER_62_232 ();
 sg13g2_fill_1 FILLER_62_234 ();
 sg13g2_fill_2 FILLER_62_255 ();
 sg13g2_fill_1 FILLER_62_261 ();
 sg13g2_fill_2 FILLER_62_291 ();
 sg13g2_fill_2 FILLER_62_321 ();
 sg13g2_decap_8 FILLER_62_359 ();
 sg13g2_fill_2 FILLER_62_366 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_1 FILLER_62_376 ();
 sg13g2_decap_4 FILLER_62_399 ();
 sg13g2_fill_1 FILLER_62_403 ();
 sg13g2_fill_1 FILLER_62_416 ();
 sg13g2_fill_2 FILLER_62_425 ();
 sg13g2_fill_2 FILLER_62_432 ();
 sg13g2_fill_1 FILLER_62_439 ();
 sg13g2_fill_1 FILLER_62_444 ();
 sg13g2_fill_2 FILLER_62_449 ();
 sg13g2_decap_4 FILLER_62_469 ();
 sg13g2_fill_2 FILLER_62_473 ();
 sg13g2_fill_2 FILLER_62_493 ();
 sg13g2_fill_1 FILLER_62_628 ();
 sg13g2_fill_1 FILLER_62_640 ();
 sg13g2_fill_1 FILLER_62_645 ();
 sg13g2_decap_4 FILLER_62_652 ();
 sg13g2_fill_1 FILLER_62_660 ();
 sg13g2_decap_8 FILLER_62_678 ();
 sg13g2_fill_1 FILLER_62_685 ();
 sg13g2_fill_2 FILLER_62_690 ();
 sg13g2_fill_1 FILLER_62_700 ();
 sg13g2_fill_1 FILLER_62_720 ();
 sg13g2_fill_2 FILLER_62_731 ();
 sg13g2_fill_1 FILLER_62_746 ();
 sg13g2_fill_1 FILLER_62_781 ();
 sg13g2_fill_2 FILLER_62_818 ();
 sg13g2_fill_1 FILLER_62_829 ();
 sg13g2_fill_2 FILLER_62_856 ();
 sg13g2_decap_4 FILLER_62_874 ();
 sg13g2_fill_1 FILLER_63_44 ();
 sg13g2_fill_1 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_74 ();
 sg13g2_fill_2 FILLER_63_108 ();
 sg13g2_fill_1 FILLER_63_139 ();
 sg13g2_fill_1 FILLER_63_144 ();
 sg13g2_fill_1 FILLER_63_159 ();
 sg13g2_fill_1 FILLER_63_168 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_fill_1 FILLER_63_210 ();
 sg13g2_fill_1 FILLER_63_226 ();
 sg13g2_fill_2 FILLER_63_246 ();
 sg13g2_fill_1 FILLER_63_248 ();
 sg13g2_fill_2 FILLER_63_285 ();
 sg13g2_fill_1 FILLER_63_290 ();
 sg13g2_fill_2 FILLER_63_309 ();
 sg13g2_fill_2 FILLER_63_320 ();
 sg13g2_decap_4 FILLER_63_334 ();
 sg13g2_fill_1 FILLER_63_338 ();
 sg13g2_decap_8 FILLER_63_361 ();
 sg13g2_fill_2 FILLER_63_368 ();
 sg13g2_fill_1 FILLER_63_387 ();
 sg13g2_fill_2 FILLER_63_393 ();
 sg13g2_fill_1 FILLER_63_409 ();
 sg13g2_fill_2 FILLER_63_419 ();
 sg13g2_fill_2 FILLER_63_440 ();
 sg13g2_decap_4 FILLER_63_460 ();
 sg13g2_fill_2 FILLER_63_498 ();
 sg13g2_fill_1 FILLER_63_500 ();
 sg13g2_decap_4 FILLER_63_506 ();
 sg13g2_fill_2 FILLER_63_510 ();
 sg13g2_fill_2 FILLER_63_517 ();
 sg13g2_decap_8 FILLER_63_527 ();
 sg13g2_fill_2 FILLER_63_629 ();
 sg13g2_fill_1 FILLER_63_657 ();
 sg13g2_fill_2 FILLER_63_695 ();
 sg13g2_fill_1 FILLER_63_726 ();
 sg13g2_decap_8 FILLER_63_772 ();
 sg13g2_decap_8 FILLER_63_779 ();
 sg13g2_fill_1 FILLER_63_786 ();
 sg13g2_fill_2 FILLER_63_826 ();
 sg13g2_fill_2 FILLER_63_850 ();
 sg13g2_fill_1 FILLER_64_30 ();
 sg13g2_fill_2 FILLER_64_35 ();
 sg13g2_fill_1 FILLER_64_57 ();
 sg13g2_fill_1 FILLER_64_71 ();
 sg13g2_fill_1 FILLER_64_76 ();
 sg13g2_fill_1 FILLER_64_138 ();
 sg13g2_fill_2 FILLER_64_167 ();
 sg13g2_fill_2 FILLER_64_211 ();
 sg13g2_fill_2 FILLER_64_221 ();
 sg13g2_fill_1 FILLER_64_223 ();
 sg13g2_fill_1 FILLER_64_232 ();
 sg13g2_fill_2 FILLER_64_249 ();
 sg13g2_fill_1 FILLER_64_267 ();
 sg13g2_fill_2 FILLER_64_276 ();
 sg13g2_fill_2 FILLER_64_294 ();
 sg13g2_fill_1 FILLER_64_316 ();
 sg13g2_fill_1 FILLER_64_337 ();
 sg13g2_fill_1 FILLER_64_374 ();
 sg13g2_fill_1 FILLER_64_397 ();
 sg13g2_fill_1 FILLER_64_403 ();
 sg13g2_decap_4 FILLER_64_413 ();
 sg13g2_fill_2 FILLER_64_417 ();
 sg13g2_fill_1 FILLER_64_431 ();
 sg13g2_fill_1 FILLER_64_435 ();
 sg13g2_fill_1 FILLER_64_441 ();
 sg13g2_fill_1 FILLER_64_446 ();
 sg13g2_fill_1 FILLER_64_451 ();
 sg13g2_fill_1 FILLER_64_461 ();
 sg13g2_fill_2 FILLER_64_483 ();
 sg13g2_fill_1 FILLER_64_493 ();
 sg13g2_decap_8 FILLER_64_498 ();
 sg13g2_decap_4 FILLER_64_505 ();
 sg13g2_fill_1 FILLER_64_526 ();
 sg13g2_fill_2 FILLER_64_562 ();
 sg13g2_fill_1 FILLER_64_568 ();
 sg13g2_fill_1 FILLER_64_573 ();
 sg13g2_fill_1 FILLER_64_599 ();
 sg13g2_decap_4 FILLER_64_629 ();
 sg13g2_fill_1 FILLER_64_633 ();
 sg13g2_fill_1 FILLER_64_638 ();
 sg13g2_fill_2 FILLER_64_643 ();
 sg13g2_decap_4 FILLER_64_649 ();
 sg13g2_fill_2 FILLER_64_732 ();
 sg13g2_fill_2 FILLER_64_757 ();
 sg13g2_fill_2 FILLER_64_790 ();
 sg13g2_fill_2 FILLER_64_854 ();
 sg13g2_fill_2 FILLER_64_876 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_32 ();
 sg13g2_fill_1 FILLER_65_65 ();
 sg13g2_fill_1 FILLER_65_130 ();
 sg13g2_fill_1 FILLER_65_139 ();
 sg13g2_fill_1 FILLER_65_165 ();
 sg13g2_fill_2 FILLER_65_174 ();
 sg13g2_fill_1 FILLER_65_209 ();
 sg13g2_decap_4 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_232 ();
 sg13g2_fill_1 FILLER_65_247 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_fill_1 FILLER_65_265 ();
 sg13g2_fill_1 FILLER_65_279 ();
 sg13g2_fill_2 FILLER_65_284 ();
 sg13g2_fill_1 FILLER_65_286 ();
 sg13g2_fill_2 FILLER_65_361 ();
 sg13g2_fill_1 FILLER_65_363 ();
 sg13g2_fill_1 FILLER_65_373 ();
 sg13g2_fill_2 FILLER_65_401 ();
 sg13g2_fill_2 FILLER_65_412 ();
 sg13g2_fill_2 FILLER_65_419 ();
 sg13g2_fill_2 FILLER_65_437 ();
 sg13g2_fill_1 FILLER_65_489 ();
 sg13g2_fill_2 FILLER_65_498 ();
 sg13g2_fill_1 FILLER_65_599 ();
 sg13g2_fill_2 FILLER_65_641 ();
 sg13g2_fill_1 FILLER_65_651 ();
 sg13g2_fill_1 FILLER_65_688 ();
 sg13g2_fill_2 FILLER_65_702 ();
 sg13g2_fill_2 FILLER_65_730 ();
 sg13g2_fill_2 FILLER_65_780 ();
 sg13g2_fill_1 FILLER_65_829 ();
 sg13g2_fill_1 FILLER_66_69 ();
 sg13g2_fill_1 FILLER_66_90 ();
 sg13g2_fill_2 FILLER_66_105 ();
 sg13g2_fill_2 FILLER_66_180 ();
 sg13g2_fill_1 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_209 ();
 sg13g2_fill_1 FILLER_66_218 ();
 sg13g2_fill_1 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_236 ();
 sg13g2_fill_1 FILLER_66_272 ();
 sg13g2_decap_8 FILLER_66_277 ();
 sg13g2_fill_1 FILLER_66_284 ();
 sg13g2_fill_1 FILLER_66_301 ();
 sg13g2_fill_2 FILLER_66_316 ();
 sg13g2_decap_8 FILLER_66_322 ();
 sg13g2_fill_2 FILLER_66_329 ();
 sg13g2_fill_1 FILLER_66_340 ();
 sg13g2_fill_2 FILLER_66_355 ();
 sg13g2_fill_1 FILLER_66_368 ();
 sg13g2_fill_1 FILLER_66_417 ();
 sg13g2_fill_1 FILLER_66_422 ();
 sg13g2_fill_1 FILLER_66_427 ();
 sg13g2_fill_1 FILLER_66_433 ();
 sg13g2_fill_2 FILLER_66_437 ();
 sg13g2_fill_2 FILLER_66_447 ();
 sg13g2_fill_1 FILLER_66_453 ();
 sg13g2_fill_1 FILLER_66_462 ();
 sg13g2_decap_4 FILLER_66_482 ();
 sg13g2_decap_8 FILLER_66_495 ();
 sg13g2_fill_2 FILLER_66_519 ();
 sg13g2_fill_1 FILLER_66_596 ();
 sg13g2_fill_1 FILLER_66_605 ();
 sg13g2_fill_1 FILLER_66_612 ();
 sg13g2_fill_1 FILLER_66_622 ();
 sg13g2_decap_4 FILLER_66_647 ();
 sg13g2_fill_2 FILLER_66_651 ();
 sg13g2_fill_2 FILLER_66_763 ();
 sg13g2_fill_1 FILLER_66_785 ();
 sg13g2_fill_1 FILLER_66_790 ();
 sg13g2_fill_1 FILLER_66_800 ();
 sg13g2_fill_2 FILLER_66_819 ();
 sg13g2_fill_1 FILLER_66_826 ();
 sg13g2_fill_1 FILLER_66_831 ();
 sg13g2_fill_2 FILLER_66_845 ();
 sg13g2_fill_2 FILLER_66_863 ();
 sg13g2_fill_2 FILLER_66_876 ();
 sg13g2_fill_2 FILLER_67_65 ();
 sg13g2_fill_1 FILLER_67_109 ();
 sg13g2_fill_1 FILLER_67_114 ();
 sg13g2_fill_1 FILLER_67_152 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_fill_2 FILLER_67_166 ();
 sg13g2_fill_2 FILLER_67_201 ();
 sg13g2_fill_1 FILLER_67_237 ();
 sg13g2_fill_2 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_256 ();
 sg13g2_decap_8 FILLER_67_278 ();
 sg13g2_fill_2 FILLER_67_289 ();
 sg13g2_fill_2 FILLER_67_299 ();
 sg13g2_fill_1 FILLER_67_305 ();
 sg13g2_fill_2 FILLER_67_326 ();
 sg13g2_fill_1 FILLER_67_328 ();
 sg13g2_decap_4 FILLER_67_348 ();
 sg13g2_decap_4 FILLER_67_356 ();
 sg13g2_decap_8 FILLER_67_368 ();
 sg13g2_fill_2 FILLER_67_405 ();
 sg13g2_fill_1 FILLER_67_411 ();
 sg13g2_fill_1 FILLER_67_417 ();
 sg13g2_fill_2 FILLER_67_423 ();
 sg13g2_fill_2 FILLER_67_429 ();
 sg13g2_fill_2 FILLER_67_435 ();
 sg13g2_fill_2 FILLER_67_441 ();
 sg13g2_fill_1 FILLER_67_443 ();
 sg13g2_fill_1 FILLER_67_449 ();
 sg13g2_fill_1 FILLER_67_454 ();
 sg13g2_fill_1 FILLER_67_460 ();
 sg13g2_fill_2 FILLER_67_464 ();
 sg13g2_fill_2 FILLER_67_480 ();
 sg13g2_decap_4 FILLER_67_486 ();
 sg13g2_fill_1 FILLER_67_490 ();
 sg13g2_decap_4 FILLER_67_495 ();
 sg13g2_fill_2 FILLER_67_499 ();
 sg13g2_fill_1 FILLER_67_505 ();
 sg13g2_decap_8 FILLER_67_511 ();
 sg13g2_decap_8 FILLER_67_518 ();
 sg13g2_fill_1 FILLER_67_525 ();
 sg13g2_fill_2 FILLER_67_557 ();
 sg13g2_fill_1 FILLER_67_569 ();
 sg13g2_fill_1 FILLER_67_579 ();
 sg13g2_fill_1 FILLER_67_583 ();
 sg13g2_fill_1 FILLER_67_594 ();
 sg13g2_fill_2 FILLER_67_605 ();
 sg13g2_fill_2 FILLER_67_611 ();
 sg13g2_fill_1 FILLER_67_613 ();
 sg13g2_decap_8 FILLER_67_619 ();
 sg13g2_fill_1 FILLER_67_626 ();
 sg13g2_fill_1 FILLER_67_661 ();
 sg13g2_fill_1 FILLER_67_665 ();
 sg13g2_fill_1 FILLER_67_670 ();
 sg13g2_fill_2 FILLER_67_675 ();
 sg13g2_fill_2 FILLER_67_690 ();
 sg13g2_fill_2 FILLER_67_700 ();
 sg13g2_fill_2 FILLER_67_707 ();
 sg13g2_fill_1 FILLER_67_714 ();
 sg13g2_fill_1 FILLER_67_723 ();
 sg13g2_fill_1 FILLER_67_731 ();
 sg13g2_fill_2 FILLER_67_767 ();
 sg13g2_fill_2 FILLER_67_798 ();
 sg13g2_fill_1 FILLER_67_800 ();
 sg13g2_fill_1 FILLER_67_805 ();
 sg13g2_fill_1 FILLER_67_811 ();
 sg13g2_fill_2 FILLER_67_838 ();
 sg13g2_fill_1 FILLER_67_849 ();
 sg13g2_fill_2 FILLER_67_876 ();
 sg13g2_fill_2 FILLER_68_26 ();
 sg13g2_fill_1 FILLER_68_44 ();
 sg13g2_fill_1 FILLER_68_79 ();
 sg13g2_fill_2 FILLER_68_84 ();
 sg13g2_fill_2 FILLER_68_154 ();
 sg13g2_fill_1 FILLER_68_165 ();
 sg13g2_fill_1 FILLER_68_233 ();
 sg13g2_fill_1 FILLER_68_237 ();
 sg13g2_fill_1 FILLER_68_244 ();
 sg13g2_fill_1 FILLER_68_284 ();
 sg13g2_fill_2 FILLER_68_295 ();
 sg13g2_fill_1 FILLER_68_297 ();
 sg13g2_decap_8 FILLER_68_378 ();
 sg13g2_decap_4 FILLER_68_407 ();
 sg13g2_fill_2 FILLER_68_411 ();
 sg13g2_fill_1 FILLER_68_417 ();
 sg13g2_fill_2 FILLER_68_437 ();
 sg13g2_fill_2 FILLER_68_464 ();
 sg13g2_fill_2 FILLER_68_491 ();
 sg13g2_fill_2 FILLER_68_505 ();
 sg13g2_fill_1 FILLER_68_537 ();
 sg13g2_fill_1 FILLER_68_546 ();
 sg13g2_fill_2 FILLER_68_551 ();
 sg13g2_fill_1 FILLER_68_558 ();
 sg13g2_fill_2 FILLER_68_571 ();
 sg13g2_fill_1 FILLER_68_644 ();
 sg13g2_fill_1 FILLER_68_669 ();
 sg13g2_fill_1 FILLER_68_691 ();
 sg13g2_fill_1 FILLER_68_707 ();
 sg13g2_fill_2 FILLER_68_721 ();
 sg13g2_fill_1 FILLER_68_723 ();
 sg13g2_decap_8 FILLER_68_732 ();
 sg13g2_fill_1 FILLER_68_739 ();
 sg13g2_decap_8 FILLER_68_744 ();
 sg13g2_decap_4 FILLER_68_751 ();
 sg13g2_fill_1 FILLER_68_790 ();
 sg13g2_fill_1 FILLER_68_804 ();
 sg13g2_fill_1 FILLER_68_818 ();
 sg13g2_fill_1 FILLER_68_823 ();
 sg13g2_fill_1 FILLER_68_828 ();
 sg13g2_fill_1 FILLER_69_26 ();
 sg13g2_fill_1 FILLER_69_32 ();
 sg13g2_fill_1 FILLER_69_60 ();
 sg13g2_fill_1 FILLER_69_111 ();
 sg13g2_fill_1 FILLER_69_158 ();
 sg13g2_fill_2 FILLER_69_182 ();
 sg13g2_fill_1 FILLER_69_196 ();
 sg13g2_fill_1 FILLER_69_207 ();
 sg13g2_fill_1 FILLER_69_213 ();
 sg13g2_fill_1 FILLER_69_218 ();
 sg13g2_fill_1 FILLER_69_224 ();
 sg13g2_fill_2 FILLER_69_233 ();
 sg13g2_fill_1 FILLER_69_254 ();
 sg13g2_fill_1 FILLER_69_260 ();
 sg13g2_fill_1 FILLER_69_284 ();
 sg13g2_fill_2 FILLER_69_301 ();
 sg13g2_fill_1 FILLER_69_313 ();
 sg13g2_fill_2 FILLER_69_331 ();
 sg13g2_fill_1 FILLER_69_349 ();
 sg13g2_fill_1 FILLER_69_354 ();
 sg13g2_fill_1 FILLER_69_369 ();
 sg13g2_decap_4 FILLER_69_382 ();
 sg13g2_decap_4 FILLER_69_390 ();
 sg13g2_fill_2 FILLER_69_394 ();
 sg13g2_decap_8 FILLER_69_416 ();
 sg13g2_fill_2 FILLER_69_423 ();
 sg13g2_fill_2 FILLER_69_433 ();
 sg13g2_decap_8 FILLER_69_440 ();
 sg13g2_fill_2 FILLER_69_447 ();
 sg13g2_fill_1 FILLER_69_468 ();
 sg13g2_fill_1 FILLER_69_478 ();
 sg13g2_decap_8 FILLER_69_487 ();
 sg13g2_fill_1 FILLER_69_520 ();
 sg13g2_fill_2 FILLER_69_530 ();
 sg13g2_fill_1 FILLER_69_536 ();
 sg13g2_fill_2 FILLER_69_550 ();
 sg13g2_fill_1 FILLER_69_565 ();
 sg13g2_fill_1 FILLER_69_575 ();
 sg13g2_fill_1 FILLER_69_628 ();
 sg13g2_fill_2 FILLER_69_649 ();
 sg13g2_fill_1 FILLER_69_667 ();
 sg13g2_fill_2 FILLER_69_722 ();
 sg13g2_fill_1 FILLER_69_740 ();
 sg13g2_decap_4 FILLER_69_751 ();
 sg13g2_fill_2 FILLER_69_755 ();
 sg13g2_fill_1 FILLER_69_808 ();
 sg13g2_fill_1 FILLER_69_854 ();
 sg13g2_decap_8 FILLER_69_863 ();
 sg13g2_decap_4 FILLER_69_874 ();
 sg13g2_fill_2 FILLER_70_86 ();
 sg13g2_fill_1 FILLER_70_156 ();
 sg13g2_fill_2 FILLER_70_169 ();
 sg13g2_fill_1 FILLER_70_184 ();
 sg13g2_fill_1 FILLER_70_193 ();
 sg13g2_fill_2 FILLER_70_230 ();
 sg13g2_fill_2 FILLER_70_246 ();
 sg13g2_fill_1 FILLER_70_253 ();
 sg13g2_fill_2 FILLER_70_273 ();
 sg13g2_fill_1 FILLER_70_284 ();
 sg13g2_fill_1 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_70_302 ();
 sg13g2_fill_1 FILLER_70_330 ();
 sg13g2_fill_1 FILLER_70_335 ();
 sg13g2_fill_1 FILLER_70_341 ();
 sg13g2_fill_1 FILLER_70_359 ();
 sg13g2_decap_8 FILLER_70_365 ();
 sg13g2_fill_1 FILLER_70_372 ();
 sg13g2_decap_4 FILLER_70_386 ();
 sg13g2_fill_2 FILLER_70_390 ();
 sg13g2_fill_2 FILLER_70_419 ();
 sg13g2_fill_1 FILLER_70_437 ();
 sg13g2_fill_2 FILLER_70_442 ();
 sg13g2_fill_2 FILLER_70_448 ();
 sg13g2_fill_2 FILLER_70_472 ();
 sg13g2_fill_2 FILLER_70_479 ();
 sg13g2_decap_4 FILLER_70_485 ();
 sg13g2_decap_4 FILLER_70_503 ();
 sg13g2_decap_4 FILLER_70_514 ();
 sg13g2_fill_1 FILLER_70_518 ();
 sg13g2_fill_2 FILLER_70_577 ();
 sg13g2_decap_4 FILLER_70_583 ();
 sg13g2_fill_2 FILLER_70_591 ();
 sg13g2_fill_1 FILLER_70_593 ();
 sg13g2_decap_4 FILLER_70_602 ();
 sg13g2_fill_2 FILLER_70_606 ();
 sg13g2_decap_8 FILLER_70_619 ();
 sg13g2_decap_4 FILLER_70_626 ();
 sg13g2_fill_1 FILLER_70_663 ();
 sg13g2_fill_2 FILLER_70_687 ();
 sg13g2_fill_1 FILLER_70_728 ();
 sg13g2_fill_2 FILLER_70_762 ();
 sg13g2_fill_1 FILLER_70_764 ();
 sg13g2_fill_1 FILLER_70_773 ();
 sg13g2_fill_1 FILLER_70_778 ();
 sg13g2_fill_1 FILLER_70_783 ();
 sg13g2_fill_1 FILLER_70_789 ();
 sg13g2_fill_1 FILLER_70_802 ();
 sg13g2_fill_1 FILLER_70_808 ();
 sg13g2_fill_1 FILLER_70_813 ();
 sg13g2_decap_4 FILLER_70_817 ();
 sg13g2_fill_1 FILLER_70_832 ();
 sg13g2_fill_1 FILLER_70_841 ();
 sg13g2_fill_2 FILLER_70_846 ();
 sg13g2_fill_1 FILLER_70_852 ();
 sg13g2_fill_2 FILLER_70_857 ();
 sg13g2_fill_2 FILLER_70_864 ();
 sg13g2_decap_8 FILLER_70_870 ();
 sg13g2_fill_1 FILLER_70_877 ();
 sg13g2_fill_2 FILLER_71_30 ();
 sg13g2_fill_1 FILLER_71_45 ();
 sg13g2_fill_1 FILLER_71_112 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_fill_1 FILLER_71_145 ();
 sg13g2_fill_2 FILLER_71_163 ();
 sg13g2_fill_1 FILLER_71_187 ();
 sg13g2_fill_1 FILLER_71_208 ();
 sg13g2_fill_1 FILLER_71_273 ();
 sg13g2_fill_2 FILLER_71_289 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_fill_2 FILLER_71_327 ();
 sg13g2_fill_1 FILLER_71_329 ();
 sg13g2_fill_2 FILLER_71_341 ();
 sg13g2_fill_1 FILLER_71_351 ();
 sg13g2_fill_2 FILLER_71_355 ();
 sg13g2_fill_1 FILLER_71_383 ();
 sg13g2_fill_1 FILLER_71_389 ();
 sg13g2_fill_1 FILLER_71_420 ();
 sg13g2_fill_2 FILLER_71_434 ();
 sg13g2_fill_1 FILLER_71_444 ();
 sg13g2_fill_1 FILLER_71_449 ();
 sg13g2_fill_1 FILLER_71_472 ();
 sg13g2_fill_2 FILLER_71_487 ();
 sg13g2_fill_1 FILLER_71_489 ();
 sg13g2_fill_2 FILLER_71_498 ();
 sg13g2_decap_8 FILLER_71_504 ();
 sg13g2_fill_2 FILLER_71_547 ();
 sg13g2_fill_1 FILLER_71_557 ();
 sg13g2_fill_1 FILLER_71_562 ();
 sg13g2_fill_2 FILLER_71_566 ();
 sg13g2_fill_2 FILLER_71_576 ();
 sg13g2_fill_1 FILLER_71_586 ();
 sg13g2_fill_2 FILLER_71_597 ();
 sg13g2_fill_1 FILLER_71_602 ();
 sg13g2_fill_1 FILLER_71_607 ();
 sg13g2_fill_1 FILLER_71_631 ();
 sg13g2_fill_1 FILLER_71_636 ();
 sg13g2_fill_2 FILLER_71_664 ();
 sg13g2_fill_1 FILLER_71_679 ();
 sg13g2_fill_1 FILLER_71_697 ();
 sg13g2_fill_2 FILLER_71_724 ();
 sg13g2_fill_1 FILLER_71_730 ();
 sg13g2_fill_1 FILLER_71_736 ();
 sg13g2_fill_1 FILLER_71_755 ();
 sg13g2_decap_4 FILLER_71_761 ();
 sg13g2_fill_1 FILLER_71_775 ();
 sg13g2_fill_2 FILLER_71_784 ();
 sg13g2_fill_2 FILLER_71_790 ();
 sg13g2_fill_1 FILLER_71_798 ();
 sg13g2_fill_1 FILLER_71_823 ();
 sg13g2_decap_4 FILLER_71_874 ();
 sg13g2_fill_1 FILLER_72_40 ();
 sg13g2_fill_2 FILLER_72_45 ();
 sg13g2_fill_1 FILLER_72_101 ();
 sg13g2_fill_1 FILLER_72_162 ();
 sg13g2_fill_2 FILLER_72_168 ();
 sg13g2_fill_1 FILLER_72_277 ();
 sg13g2_fill_1 FILLER_72_301 ();
 sg13g2_fill_1 FILLER_72_309 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_8 FILLER_72_346 ();
 sg13g2_fill_1 FILLER_72_353 ();
 sg13g2_fill_1 FILLER_72_362 ();
 sg13g2_fill_2 FILLER_72_367 ();
 sg13g2_fill_1 FILLER_72_373 ();
 sg13g2_fill_1 FILLER_72_393 ();
 sg13g2_fill_2 FILLER_72_403 ();
 sg13g2_fill_2 FILLER_72_417 ();
 sg13g2_fill_1 FILLER_72_436 ();
 sg13g2_fill_1 FILLER_72_446 ();
 sg13g2_fill_2 FILLER_72_457 ();
 sg13g2_decap_4 FILLER_72_471 ();
 sg13g2_fill_2 FILLER_72_479 ();
 sg13g2_fill_1 FILLER_72_481 ();
 sg13g2_fill_2 FILLER_72_498 ();
 sg13g2_decap_4 FILLER_72_509 ();
 sg13g2_fill_2 FILLER_72_513 ();
 sg13g2_fill_2 FILLER_72_526 ();
 sg13g2_fill_1 FILLER_72_528 ();
 sg13g2_fill_1 FILLER_72_548 ();
 sg13g2_fill_2 FILLER_72_573 ();
 sg13g2_fill_1 FILLER_72_580 ();
 sg13g2_decap_4 FILLER_72_594 ();
 sg13g2_fill_2 FILLER_72_607 ();
 sg13g2_fill_1 FILLER_72_654 ();
 sg13g2_fill_2 FILLER_72_668 ();
 sg13g2_fill_2 FILLER_72_681 ();
 sg13g2_decap_8 FILLER_72_716 ();
 sg13g2_fill_2 FILLER_72_723 ();
 sg13g2_fill_1 FILLER_72_725 ();
 sg13g2_fill_1 FILLER_72_735 ();
 sg13g2_fill_1 FILLER_72_740 ();
 sg13g2_decap_8 FILLER_72_749 ();
 sg13g2_fill_1 FILLER_72_769 ();
 sg13g2_fill_2 FILLER_72_778 ();
 sg13g2_fill_1 FILLER_72_780 ();
 sg13g2_fill_1 FILLER_72_799 ();
 sg13g2_fill_1 FILLER_72_809 ();
 sg13g2_fill_1 FILLER_72_818 ();
 sg13g2_fill_1 FILLER_72_823 ();
 sg13g2_fill_2 FILLER_72_844 ();
 sg13g2_fill_2 FILLER_72_863 ();
 sg13g2_fill_1 FILLER_72_865 ();
 sg13g2_decap_4 FILLER_72_874 ();
 sg13g2_fill_1 FILLER_73_48 ();
 sg13g2_fill_2 FILLER_73_64 ();
 sg13g2_fill_2 FILLER_73_169 ();
 sg13g2_fill_2 FILLER_73_216 ();
 sg13g2_fill_1 FILLER_73_230 ();
 sg13g2_fill_1 FILLER_73_268 ();
 sg13g2_fill_1 FILLER_73_297 ();
 sg13g2_fill_2 FILLER_73_306 ();
 sg13g2_fill_1 FILLER_73_316 ();
 sg13g2_fill_2 FILLER_73_346 ();
 sg13g2_decap_4 FILLER_73_369 ();
 sg13g2_fill_1 FILLER_73_377 ();
 sg13g2_fill_2 FILLER_73_387 ();
 sg13g2_fill_1 FILLER_73_389 ();
 sg13g2_fill_1 FILLER_73_398 ();
 sg13g2_fill_1 FILLER_73_407 ();
 sg13g2_fill_1 FILLER_73_412 ();
 sg13g2_fill_1 FILLER_73_418 ();
 sg13g2_fill_1 FILLER_73_424 ();
 sg13g2_fill_2 FILLER_73_429 ();
 sg13g2_fill_2 FILLER_73_435 ();
 sg13g2_fill_1 FILLER_73_442 ();
 sg13g2_fill_1 FILLER_73_446 ();
 sg13g2_fill_1 FILLER_73_468 ();
 sg13g2_fill_2 FILLER_73_473 ();
 sg13g2_fill_1 FILLER_73_480 ();
 sg13g2_fill_2 FILLER_73_486 ();
 sg13g2_fill_1 FILLER_73_502 ();
 sg13g2_fill_1 FILLER_73_506 ();
 sg13g2_fill_2 FILLER_73_526 ();
 sg13g2_fill_1 FILLER_73_537 ();
 sg13g2_fill_1 FILLER_73_548 ();
 sg13g2_fill_2 FILLER_73_562 ();
 sg13g2_fill_1 FILLER_73_576 ();
 sg13g2_decap_4 FILLER_73_593 ();
 sg13g2_fill_1 FILLER_73_602 ();
 sg13g2_decap_8 FILLER_73_608 ();
 sg13g2_fill_2 FILLER_73_615 ();
 sg13g2_fill_1 FILLER_73_625 ();
 sg13g2_fill_2 FILLER_73_630 ();
 sg13g2_fill_2 FILLER_73_652 ();
 sg13g2_fill_1 FILLER_73_654 ();
 sg13g2_fill_1 FILLER_73_669 ();
 sg13g2_fill_1 FILLER_73_675 ();
 sg13g2_fill_1 FILLER_73_684 ();
 sg13g2_fill_2 FILLER_73_712 ();
 sg13g2_fill_2 FILLER_73_749 ();
 sg13g2_fill_2 FILLER_73_777 ();
 sg13g2_fill_1 FILLER_73_779 ();
 sg13g2_fill_1 FILLER_73_784 ();
 sg13g2_fill_2 FILLER_73_834 ();
 sg13g2_fill_2 FILLER_73_844 ();
 sg13g2_decap_4 FILLER_73_874 ();
 sg13g2_fill_1 FILLER_74_13 ();
 sg13g2_fill_1 FILLER_74_95 ();
 sg13g2_fill_1 FILLER_74_217 ();
 sg13g2_fill_1 FILLER_74_248 ();
 sg13g2_fill_1 FILLER_74_275 ();
 sg13g2_fill_1 FILLER_74_280 ();
 sg13g2_fill_2 FILLER_74_300 ();
 sg13g2_fill_2 FILLER_74_349 ();
 sg13g2_decap_8 FILLER_74_362 ();
 sg13g2_decap_4 FILLER_74_369 ();
 sg13g2_fill_2 FILLER_74_373 ();
 sg13g2_fill_1 FILLER_74_389 ();
 sg13g2_fill_1 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_422 ();
 sg13g2_fill_1 FILLER_74_428 ();
 sg13g2_fill_1 FILLER_74_433 ();
 sg13g2_fill_1 FILLER_74_439 ();
 sg13g2_fill_2 FILLER_74_448 ();
 sg13g2_decap_4 FILLER_74_458 ();
 sg13g2_fill_2 FILLER_74_462 ();
 sg13g2_fill_2 FILLER_74_476 ();
 sg13g2_fill_1 FILLER_74_478 ();
 sg13g2_decap_4 FILLER_74_506 ();
 sg13g2_fill_2 FILLER_74_510 ();
 sg13g2_fill_1 FILLER_74_520 ();
 sg13g2_decap_4 FILLER_74_525 ();
 sg13g2_fill_1 FILLER_74_529 ();
 sg13g2_fill_2 FILLER_74_537 ();
 sg13g2_fill_1 FILLER_74_539 ();
 sg13g2_fill_1 FILLER_74_548 ();
 sg13g2_fill_2 FILLER_74_563 ();
 sg13g2_fill_1 FILLER_74_571 ();
 sg13g2_fill_1 FILLER_74_577 ();
 sg13g2_fill_1 FILLER_74_590 ();
 sg13g2_fill_2 FILLER_74_609 ();
 sg13g2_fill_1 FILLER_74_614 ();
 sg13g2_decap_4 FILLER_74_619 ();
 sg13g2_fill_1 FILLER_74_688 ();
 sg13g2_fill_1 FILLER_74_745 ();
 sg13g2_fill_1 FILLER_74_759 ();
 sg13g2_fill_1 FILLER_74_772 ();
 sg13g2_fill_1 FILLER_74_786 ();
 sg13g2_fill_1 FILLER_74_806 ();
 sg13g2_fill_2 FILLER_74_862 ();
 sg13g2_fill_2 FILLER_74_876 ();
 sg13g2_fill_1 FILLER_75_60 ();
 sg13g2_fill_1 FILLER_75_102 ();
 sg13g2_fill_1 FILLER_75_107 ();
 sg13g2_fill_1 FILLER_75_116 ();
 sg13g2_fill_1 FILLER_75_121 ();
 sg13g2_fill_1 FILLER_75_153 ();
 sg13g2_fill_1 FILLER_75_159 ();
 sg13g2_fill_2 FILLER_75_218 ();
 sg13g2_fill_1 FILLER_75_274 ();
 sg13g2_fill_2 FILLER_75_300 ();
 sg13g2_fill_2 FILLER_75_323 ();
 sg13g2_fill_2 FILLER_75_350 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_fill_1 FILLER_75_370 ();
 sg13g2_fill_1 FILLER_75_379 ();
 sg13g2_fill_2 FILLER_75_384 ();
 sg13g2_fill_1 FILLER_75_391 ();
 sg13g2_fill_2 FILLER_75_396 ();
 sg13g2_fill_1 FILLER_75_401 ();
 sg13g2_fill_2 FILLER_75_406 ();
 sg13g2_fill_2 FILLER_75_416 ();
 sg13g2_fill_1 FILLER_75_422 ();
 sg13g2_fill_1 FILLER_75_432 ();
 sg13g2_fill_1 FILLER_75_440 ();
 sg13g2_fill_1 FILLER_75_444 ();
 sg13g2_fill_2 FILLER_75_448 ();
 sg13g2_decap_8 FILLER_75_454 ();
 sg13g2_fill_2 FILLER_75_461 ();
 sg13g2_fill_2 FILLER_75_475 ();
 sg13g2_fill_1 FILLER_75_504 ();
 sg13g2_decap_8 FILLER_75_513 ();
 sg13g2_fill_2 FILLER_75_520 ();
 sg13g2_fill_1 FILLER_75_522 ();
 sg13g2_fill_2 FILLER_75_527 ();
 sg13g2_fill_1 FILLER_75_543 ();
 sg13g2_fill_1 FILLER_75_552 ();
 sg13g2_fill_1 FILLER_75_558 ();
 sg13g2_fill_2 FILLER_75_564 ();
 sg13g2_fill_1 FILLER_75_574 ();
 sg13g2_fill_2 FILLER_75_579 ();
 sg13g2_fill_2 FILLER_75_617 ();
 sg13g2_fill_1 FILLER_75_674 ();
 sg13g2_fill_2 FILLER_75_679 ();
 sg13g2_fill_2 FILLER_75_694 ();
 sg13g2_fill_1 FILLER_75_702 ();
 sg13g2_fill_1 FILLER_75_711 ();
 sg13g2_fill_1 FILLER_75_720 ();
 sg13g2_fill_2 FILLER_75_754 ();
 sg13g2_fill_2 FILLER_75_773 ();
 sg13g2_fill_1 FILLER_75_775 ();
 sg13g2_decap_4 FILLER_75_780 ();
 sg13g2_decap_8 FILLER_75_793 ();
 sg13g2_fill_1 FILLER_75_813 ();
 sg13g2_fill_1 FILLER_75_820 ();
 sg13g2_fill_1 FILLER_75_833 ();
 sg13g2_fill_1 FILLER_75_871 ();
 sg13g2_fill_2 FILLER_75_876 ();
 sg13g2_fill_2 FILLER_76_10 ();
 sg13g2_fill_1 FILLER_76_79 ();
 sg13g2_fill_2 FILLER_76_148 ();
 sg13g2_fill_2 FILLER_76_192 ();
 sg13g2_fill_2 FILLER_76_216 ();
 sg13g2_fill_2 FILLER_76_283 ();
 sg13g2_fill_1 FILLER_76_309 ();
 sg13g2_fill_1 FILLER_76_340 ();
 sg13g2_fill_1 FILLER_76_350 ();
 sg13g2_fill_1 FILLER_76_356 ();
 sg13g2_fill_1 FILLER_76_361 ();
 sg13g2_fill_2 FILLER_76_367 ();
 sg13g2_fill_1 FILLER_76_377 ();
 sg13g2_fill_2 FILLER_76_382 ();
 sg13g2_fill_1 FILLER_76_392 ();
 sg13g2_fill_1 FILLER_76_406 ();
 sg13g2_fill_2 FILLER_76_411 ();
 sg13g2_fill_2 FILLER_76_421 ();
 sg13g2_fill_1 FILLER_76_423 ();
 sg13g2_decap_8 FILLER_76_428 ();
 sg13g2_decap_4 FILLER_76_438 ();
 sg13g2_fill_2 FILLER_76_442 ();
 sg13g2_fill_1 FILLER_76_456 ();
 sg13g2_fill_1 FILLER_76_476 ();
 sg13g2_fill_1 FILLER_76_504 ();
 sg13g2_fill_1 FILLER_76_517 ();
 sg13g2_fill_2 FILLER_76_526 ();
 sg13g2_fill_2 FILLER_76_536 ();
 sg13g2_fill_1 FILLER_76_542 ();
 sg13g2_decap_4 FILLER_76_547 ();
 sg13g2_fill_1 FILLER_76_555 ();
 sg13g2_fill_1 FILLER_76_564 ();
 sg13g2_fill_1 FILLER_76_570 ();
 sg13g2_fill_1 FILLER_76_574 ();
 sg13g2_fill_1 FILLER_76_579 ();
 sg13g2_decap_4 FILLER_76_600 ();
 sg13g2_fill_2 FILLER_76_604 ();
 sg13g2_fill_2 FILLER_76_633 ();
 sg13g2_fill_1 FILLER_76_635 ();
 sg13g2_fill_1 FILLER_76_644 ();
 sg13g2_fill_1 FILLER_76_649 ();
 sg13g2_fill_2 FILLER_76_668 ();
 sg13g2_fill_1 FILLER_76_684 ();
 sg13g2_fill_1 FILLER_76_693 ();
 sg13g2_fill_2 FILLER_76_702 ();
 sg13g2_fill_1 FILLER_76_728 ();
 sg13g2_decap_4 FILLER_76_733 ();
 sg13g2_fill_2 FILLER_76_737 ();
 sg13g2_decap_4 FILLER_76_743 ();
 sg13g2_fill_1 FILLER_76_747 ();
 sg13g2_fill_1 FILLER_76_751 ();
 sg13g2_fill_1 FILLER_76_776 ();
 sg13g2_fill_1 FILLER_76_801 ();
 sg13g2_decap_8 FILLER_76_840 ();
 sg13g2_decap_4 FILLER_76_850 ();
 sg13g2_fill_1 FILLER_76_854 ();
 sg13g2_fill_1 FILLER_76_877 ();
 sg13g2_fill_2 FILLER_77_25 ();
 sg13g2_fill_1 FILLER_77_41 ();
 sg13g2_fill_1 FILLER_77_68 ();
 sg13g2_fill_1 FILLER_77_79 ();
 sg13g2_fill_1 FILLER_77_89 ();
 sg13g2_fill_2 FILLER_77_110 ();
 sg13g2_fill_2 FILLER_77_234 ();
 sg13g2_fill_2 FILLER_77_293 ();
 sg13g2_fill_2 FILLER_77_307 ();
 sg13g2_fill_1 FILLER_77_314 ();
 sg13g2_fill_2 FILLER_77_335 ();
 sg13g2_fill_1 FILLER_77_341 ();
 sg13g2_fill_1 FILLER_77_346 ();
 sg13g2_fill_1 FILLER_77_352 ();
 sg13g2_fill_1 FILLER_77_357 ();
 sg13g2_fill_1 FILLER_77_363 ();
 sg13g2_fill_1 FILLER_77_377 ();
 sg13g2_fill_1 FILLER_77_382 ();
 sg13g2_fill_1 FILLER_77_388 ();
 sg13g2_fill_1 FILLER_77_392 ();
 sg13g2_fill_1 FILLER_77_401 ();
 sg13g2_fill_1 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_fill_2 FILLER_77_442 ();
 sg13g2_fill_2 FILLER_77_464 ();
 sg13g2_fill_1 FILLER_77_473 ();
 sg13g2_fill_2 FILLER_77_487 ();
 sg13g2_fill_1 FILLER_77_489 ();
 sg13g2_fill_2 FILLER_77_516 ();
 sg13g2_fill_1 FILLER_77_522 ();
 sg13g2_decap_4 FILLER_77_527 ();
 sg13g2_fill_2 FILLER_77_531 ();
 sg13g2_fill_1 FILLER_77_537 ();
 sg13g2_fill_1 FILLER_77_545 ();
 sg13g2_fill_2 FILLER_77_549 ();
 sg13g2_fill_1 FILLER_77_551 ();
 sg13g2_fill_2 FILLER_77_561 ();
 sg13g2_fill_1 FILLER_77_563 ();
 sg13g2_fill_2 FILLER_77_586 ();
 sg13g2_fill_1 FILLER_77_627 ();
 sg13g2_fill_2 FILLER_77_635 ();
 sg13g2_fill_1 FILLER_77_641 ();
 sg13g2_fill_2 FILLER_77_651 ();
 sg13g2_fill_2 FILLER_77_663 ();
 sg13g2_decap_8 FILLER_77_689 ();
 sg13g2_fill_1 FILLER_77_696 ();
 sg13g2_decap_8 FILLER_77_726 ();
 sg13g2_fill_2 FILLER_77_733 ();
 sg13g2_fill_2 FILLER_77_759 ();
 sg13g2_fill_1 FILLER_77_761 ();
 sg13g2_fill_2 FILLER_77_770 ();
 sg13g2_fill_1 FILLER_77_784 ();
 sg13g2_fill_1 FILLER_77_790 ();
 sg13g2_fill_2 FILLER_77_795 ();
 sg13g2_decap_8 FILLER_77_805 ();
 sg13g2_decap_4 FILLER_77_812 ();
 sg13g2_fill_1 FILLER_77_835 ();
 sg13g2_fill_1 FILLER_77_852 ();
 sg13g2_fill_1 FILLER_77_858 ();
 sg13g2_fill_1 FILLER_77_866 ();
 sg13g2_decap_8 FILLER_77_871 ();
 sg13g2_fill_1 FILLER_78_32 ();
 sg13g2_fill_1 FILLER_78_65 ();
 sg13g2_fill_1 FILLER_78_71 ();
 sg13g2_fill_1 FILLER_78_86 ();
 sg13g2_fill_1 FILLER_78_163 ();
 sg13g2_fill_1 FILLER_78_206 ();
 sg13g2_fill_1 FILLER_78_216 ();
 sg13g2_fill_2 FILLER_78_226 ();
 sg13g2_fill_2 FILLER_78_261 ();
 sg13g2_fill_1 FILLER_78_297 ();
 sg13g2_fill_1 FILLER_78_305 ();
 sg13g2_fill_1 FILLER_78_311 ();
 sg13g2_fill_2 FILLER_78_338 ();
 sg13g2_fill_1 FILLER_78_340 ();
 sg13g2_fill_2 FILLER_78_345 ();
 sg13g2_fill_1 FILLER_78_373 ();
 sg13g2_fill_1 FILLER_78_378 ();
 sg13g2_fill_2 FILLER_78_383 ();
 sg13g2_fill_1 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_401 ();
 sg13g2_fill_2 FILLER_78_408 ();
 sg13g2_fill_1 FILLER_78_410 ();
 sg13g2_fill_1 FILLER_78_420 ();
 sg13g2_fill_2 FILLER_78_426 ();
 sg13g2_fill_1 FILLER_78_428 ();
 sg13g2_decap_4 FILLER_78_461 ();
 sg13g2_fill_2 FILLER_78_465 ();
 sg13g2_fill_1 FILLER_78_489 ();
 sg13g2_decap_4 FILLER_78_494 ();
 sg13g2_fill_1 FILLER_78_506 ();
 sg13g2_decap_4 FILLER_78_520 ();
 sg13g2_fill_2 FILLER_78_528 ();
 sg13g2_fill_1 FILLER_78_530 ();
 sg13g2_fill_2 FILLER_78_540 ();
 sg13g2_fill_1 FILLER_78_547 ();
 sg13g2_fill_1 FILLER_78_561 ();
 sg13g2_fill_2 FILLER_78_570 ();
 sg13g2_fill_1 FILLER_78_594 ();
 sg13g2_fill_1 FILLER_78_607 ();
 sg13g2_fill_2 FILLER_78_652 ();
 sg13g2_fill_2 FILLER_78_659 ();
 sg13g2_fill_2 FILLER_78_670 ();
 sg13g2_decap_4 FILLER_78_711 ();
 sg13g2_fill_1 FILLER_78_741 ();
 sg13g2_fill_2 FILLER_78_781 ();
 sg13g2_fill_1 FILLER_78_783 ();
 sg13g2_fill_1 FILLER_78_796 ();
 sg13g2_decap_4 FILLER_78_809 ();
 sg13g2_fill_2 FILLER_78_813 ();
 sg13g2_fill_1 FILLER_78_845 ();
 sg13g2_fill_2 FILLER_78_851 ();
 sg13g2_decap_4 FILLER_78_874 ();
 sg13g2_fill_2 FILLER_79_28 ();
 sg13g2_fill_1 FILLER_79_42 ();
 sg13g2_fill_1 FILLER_79_67 ();
 sg13g2_fill_2 FILLER_79_132 ();
 sg13g2_fill_2 FILLER_79_160 ();
 sg13g2_fill_2 FILLER_79_180 ();
 sg13g2_fill_2 FILLER_79_258 ();
 sg13g2_fill_1 FILLER_79_294 ();
 sg13g2_fill_2 FILLER_79_300 ();
 sg13g2_fill_1 FILLER_79_306 ();
 sg13g2_fill_2 FILLER_79_311 ();
 sg13g2_fill_1 FILLER_79_317 ();
 sg13g2_fill_1 FILLER_79_322 ();
 sg13g2_fill_1 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_370 ();
 sg13g2_fill_1 FILLER_79_377 ();
 sg13g2_fill_1 FILLER_79_382 ();
 sg13g2_fill_1 FILLER_79_387 ();
 sg13g2_fill_1 FILLER_79_402 ();
 sg13g2_decap_4 FILLER_79_407 ();
 sg13g2_fill_1 FILLER_79_428 ();
 sg13g2_fill_2 FILLER_79_438 ();
 sg13g2_fill_1 FILLER_79_440 ();
 sg13g2_fill_1 FILLER_79_458 ();
 sg13g2_fill_2 FILLER_79_472 ();
 sg13g2_fill_1 FILLER_79_474 ();
 sg13g2_fill_1 FILLER_79_480 ();
 sg13g2_fill_1 FILLER_79_485 ();
 sg13g2_fill_2 FILLER_79_503 ();
 sg13g2_fill_1 FILLER_79_509 ();
 sg13g2_fill_2 FILLER_79_527 ();
 sg13g2_fill_1 FILLER_79_529 ();
 sg13g2_fill_1 FILLER_79_543 ();
 sg13g2_fill_1 FILLER_79_570 ();
 sg13g2_fill_1 FILLER_79_591 ();
 sg13g2_fill_1 FILLER_79_595 ();
 sg13g2_fill_1 FILLER_79_612 ();
 sg13g2_fill_1 FILLER_79_617 ();
 sg13g2_fill_1 FILLER_79_621 ();
 sg13g2_fill_2 FILLER_79_670 ();
 sg13g2_fill_1 FILLER_79_672 ();
 sg13g2_fill_1 FILLER_79_678 ();
 sg13g2_decap_4 FILLER_79_684 ();
 sg13g2_fill_2 FILLER_79_696 ();
 sg13g2_fill_1 FILLER_79_738 ();
 sg13g2_fill_1 FILLER_79_755 ();
 sg13g2_fill_2 FILLER_79_769 ();
 sg13g2_fill_1 FILLER_79_784 ();
 sg13g2_fill_1 FILLER_79_801 ();
 sg13g2_fill_1 FILLER_79_817 ();
 sg13g2_fill_2 FILLER_79_826 ();
 sg13g2_fill_1 FILLER_79_852 ();
 sg13g2_decap_4 FILLER_79_872 ();
 sg13g2_fill_2 FILLER_79_876 ();
 sg13g2_fill_2 FILLER_80_42 ();
 sg13g2_fill_1 FILLER_80_100 ();
 sg13g2_fill_1 FILLER_80_188 ();
 sg13g2_fill_1 FILLER_80_276 ();
 sg13g2_fill_1 FILLER_80_287 ();
 sg13g2_fill_2 FILLER_80_292 ();
 sg13g2_fill_2 FILLER_80_350 ();
 sg13g2_decap_8 FILLER_80_363 ();
 sg13g2_decap_8 FILLER_80_370 ();
 sg13g2_fill_2 FILLER_80_377 ();
 sg13g2_fill_2 FILLER_80_383 ();
 sg13g2_fill_1 FILLER_80_397 ();
 sg13g2_fill_2 FILLER_80_402 ();
 sg13g2_fill_2 FILLER_80_422 ();
 sg13g2_fill_1 FILLER_80_424 ();
 sg13g2_fill_2 FILLER_80_430 ();
 sg13g2_fill_1 FILLER_80_432 ();
 sg13g2_fill_2 FILLER_80_438 ();
 sg13g2_fill_1 FILLER_80_462 ();
 sg13g2_decap_8 FILLER_80_468 ();
 sg13g2_decap_8 FILLER_80_475 ();
 sg13g2_decap_4 FILLER_80_490 ();
 sg13g2_fill_1 FILLER_80_494 ();
 sg13g2_fill_1 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_531 ();
 sg13g2_decap_8 FILLER_80_538 ();
 sg13g2_fill_2 FILLER_80_545 ();
 sg13g2_fill_1 FILLER_80_547 ();
 sg13g2_decap_4 FILLER_80_565 ();
 sg13g2_fill_2 FILLER_80_569 ();
 sg13g2_fill_2 FILLER_80_575 ();
 sg13g2_fill_1 FILLER_80_598 ();
 sg13g2_fill_2 FILLER_80_619 ();
 sg13g2_decap_8 FILLER_80_632 ();
 sg13g2_decap_4 FILLER_80_639 ();
 sg13g2_fill_2 FILLER_80_643 ();
 sg13g2_fill_1 FILLER_80_690 ();
 sg13g2_decap_4 FILLER_80_699 ();
 sg13g2_fill_2 FILLER_80_703 ();
 sg13g2_fill_1 FILLER_80_713 ();
 sg13g2_decap_8 FILLER_80_746 ();
 sg13g2_decap_4 FILLER_80_757 ();
 sg13g2_fill_1 FILLER_80_761 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_fill_1 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_808 ();
 sg13g2_decap_4 FILLER_80_819 ();
 sg13g2_fill_1 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_fill_1 FILLER_80_835 ();
 sg13g2_fill_1 FILLER_80_843 ();
 sg13g2_decap_4 FILLER_80_872 ();
 sg13g2_fill_2 FILLER_80_876 ();
endmodule
