module tt_um_MichaelBell_tinyQV (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire clknet_leaf_0_clk;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire net1354;
 wire \addr[0] ;
 wire \addr[10] ;
 wire \addr[11] ;
 wire \addr[12] ;
 wire \addr[13] ;
 wire \addr[14] ;
 wire \addr[15] ;
 wire \addr[16] ;
 wire \addr[17] ;
 wire \addr[18] ;
 wire \addr[19] ;
 wire \addr[1] ;
 wire \addr[20] ;
 wire \addr[21] ;
 wire \addr[22] ;
 wire \addr[23] ;
 wire \addr[24] ;
 wire \addr[25] ;
 wire \addr[26] ;
 wire \addr[27] ;
 wire \addr[2] ;
 wire \addr[3] ;
 wire \addr[4] ;
 wire \addr[5] ;
 wire \addr[6] ;
 wire \addr[7] ;
 wire \addr[8] ;
 wire \addr[9] ;
 wire \data_to_write[0] ;
 wire \data_to_write[10] ;
 wire \data_to_write[11] ;
 wire \data_to_write[12] ;
 wire \data_to_write[13] ;
 wire \data_to_write[14] ;
 wire \data_to_write[15] ;
 wire \data_to_write[16] ;
 wire \data_to_write[17] ;
 wire \data_to_write[18] ;
 wire \data_to_write[19] ;
 wire \data_to_write[1] ;
 wire \data_to_write[20] ;
 wire \data_to_write[21] ;
 wire \data_to_write[22] ;
 wire \data_to_write[23] ;
 wire \data_to_write[24] ;
 wire \data_to_write[25] ;
 wire \data_to_write[26] ;
 wire \data_to_write[27] ;
 wire \data_to_write[28] ;
 wire \data_to_write[29] ;
 wire \data_to_write[2] ;
 wire \data_to_write[30] ;
 wire \data_to_write[31] ;
 wire \data_to_write[3] ;
 wire \data_to_write[4] ;
 wire \data_to_write[5] ;
 wire \data_to_write[6] ;
 wire \data_to_write[7] ;
 wire \data_to_write[8] ;
 wire \data_to_write[9] ;
 wire debug_data_continue;
 wire debug_instr_valid;
 wire \debug_rd[0] ;
 wire \debug_rd[1] ;
 wire \debug_rd[2] ;
 wire \debug_rd[3] ;
 wire \debug_rd_r[0] ;
 wire \debug_rd_r[1] ;
 wire \debug_rd_r[2] ;
 wire \debug_rd_r[3] ;
 wire debug_register_data;
 wire debug_uart_txd;
 wire \gpio_out[0] ;
 wire \gpio_out[1] ;
 wire \gpio_out[2] ;
 wire \gpio_out[3] ;
 wire \gpio_out[4] ;
 wire \gpio_out[5] ;
 wire \gpio_out[6] ;
 wire \gpio_out[7] ;
 wire \gpio_out_sel[0] ;
 wire \gpio_out_sel[1] ;
 wire \gpio_out_sel[2] ;
 wire \gpio_out_sel[3] ;
 wire \gpio_out_sel[4] ;
 wire \gpio_out_sel[5] ;
 wire \gpio_out_sel[6] ;
 wire \gpio_out_sel[7] ;
 wire \i_debug_uart_tx.cycle_counter[0] ;
 wire \i_debug_uart_tx.cycle_counter[1] ;
 wire \i_debug_uart_tx.cycle_counter[2] ;
 wire \i_debug_uart_tx.cycle_counter[3] ;
 wire \i_debug_uart_tx.cycle_counter[4] ;
 wire \i_debug_uart_tx.data_to_send[0] ;
 wire \i_debug_uart_tx.data_to_send[1] ;
 wire \i_debug_uart_tx.data_to_send[2] ;
 wire \i_debug_uart_tx.data_to_send[3] ;
 wire \i_debug_uart_tx.data_to_send[4] ;
 wire \i_debug_uart_tx.data_to_send[5] ;
 wire \i_debug_uart_tx.data_to_send[6] ;
 wire \i_debug_uart_tx.data_to_send[7] ;
 wire \i_debug_uart_tx.fsm_state[0] ;
 wire \i_debug_uart_tx.fsm_state[1] ;
 wire \i_debug_uart_tx.fsm_state[2] ;
 wire \i_debug_uart_tx.fsm_state[3] ;
 wire \i_debug_uart_tx.resetn ;
 wire \i_spi.bits_remaining[0] ;
 wire \i_spi.bits_remaining[1] ;
 wire \i_spi.bits_remaining[2] ;
 wire \i_spi.bits_remaining[3] ;
 wire \i_spi.busy ;
 wire \i_spi.clock_count[0] ;
 wire \i_spi.clock_count[1] ;
 wire \i_spi.clock_divider[0] ;
 wire \i_spi.clock_divider[1] ;
 wire \i_spi.data[0] ;
 wire \i_spi.data[1] ;
 wire \i_spi.data[2] ;
 wire \i_spi.data[3] ;
 wire \i_spi.data[4] ;
 wire \i_spi.data[5] ;
 wire \i_spi.data[6] ;
 wire \i_spi.data[7] ;
 wire \i_spi.end_txn_reg ;
 wire \i_spi.read_latency ;
 wire \i_spi.spi_clk_out ;
 wire \i_spi.spi_dc ;
 wire \i_spi.spi_select ;
 wire \i_tinyqv.cpu.additional_mem_ops[0] ;
 wire \i_tinyqv.cpu.additional_mem_ops[1] ;
 wire \i_tinyqv.cpu.additional_mem_ops[2] ;
 wire \i_tinyqv.cpu.alu_op[0] ;
 wire \i_tinyqv.cpu.alu_op[1] ;
 wire \i_tinyqv.cpu.alu_op[2] ;
 wire \i_tinyqv.cpu.alu_op[3] ;
 wire \i_tinyqv.cpu.counter[2] ;
 wire \i_tinyqv.cpu.counter[3] ;
 wire \i_tinyqv.cpu.counter[4] ;
 wire \i_tinyqv.cpu.data_read_n[0] ;
 wire \i_tinyqv.cpu.data_read_n[1] ;
 wire \i_tinyqv.cpu.data_ready_core ;
 wire \i_tinyqv.cpu.data_ready_latch ;
 wire \i_tinyqv.cpu.data_write_n[0] ;
 wire \i_tinyqv.cpu.data_write_n[1] ;
 wire \i_tinyqv.cpu.i_core.cmp ;
 wire \i_tinyqv.cpu.i_core.cmp_out ;
 wire \i_tinyqv.cpu.i_core.cy ;
 wire \i_tinyqv.cpu.i_core.cy_out ;
 wire \i_tinyqv.cpu.i_core.cycle[0] ;
 wire \i_tinyqv.cpu.i_core.cycle[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[0] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[2] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[3] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[4] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[5] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[6] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.cy ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.rstn ;
 wire \i_tinyqv.cpu.i_core.i_instrret.add ;
 wire \i_tinyqv.cpu.i_core.i_instrret.cy ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[0] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[1] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[2] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[3] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[10] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[11] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[12] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[13] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[14] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[15] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[16] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[17] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[18] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[19] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[20] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[21] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[22] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[23] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[24] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[25] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[26] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[27] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[28] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[29] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[30] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[31] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[4] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[5] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[6] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[7] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[8] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[9] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[0] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[10] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[11] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[1] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[2] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[3] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[5] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[6] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[7] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[8] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[9] ;
 wire \i_tinyqv.cpu.i_core.interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.is_double_fault_r ;
 wire \i_tinyqv.cpu.i_core.is_interrupt ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.load_done ;
 wire \i_tinyqv.cpu.i_core.load_top_bit ;
 wire \i_tinyqv.cpu.i_core.mcause[0] ;
 wire \i_tinyqv.cpu.i_core.mcause[1] ;
 wire \i_tinyqv.cpu.i_core.mcause[3] ;
 wire \i_tinyqv.cpu.i_core.mcause[4] ;
 wire \i_tinyqv.cpu.i_core.mem_op[0] ;
 wire \i_tinyqv.cpu.i_core.mem_op[1] ;
 wire \i_tinyqv.cpu.i_core.mem_op[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[0] ;
 wire \i_tinyqv.cpu.i_core.mepc[10] ;
 wire \i_tinyqv.cpu.i_core.mepc[11] ;
 wire \i_tinyqv.cpu.i_core.mepc[12] ;
 wire \i_tinyqv.cpu.i_core.mepc[13] ;
 wire \i_tinyqv.cpu.i_core.mepc[14] ;
 wire \i_tinyqv.cpu.i_core.mepc[15] ;
 wire \i_tinyqv.cpu.i_core.mepc[16] ;
 wire \i_tinyqv.cpu.i_core.mepc[17] ;
 wire \i_tinyqv.cpu.i_core.mepc[18] ;
 wire \i_tinyqv.cpu.i_core.mepc[19] ;
 wire \i_tinyqv.cpu.i_core.mepc[1] ;
 wire \i_tinyqv.cpu.i_core.mepc[20] ;
 wire \i_tinyqv.cpu.i_core.mepc[21] ;
 wire \i_tinyqv.cpu.i_core.mepc[22] ;
 wire \i_tinyqv.cpu.i_core.mepc[23] ;
 wire \i_tinyqv.cpu.i_core.mepc[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[3] ;
 wire \i_tinyqv.cpu.i_core.mepc[4] ;
 wire \i_tinyqv.cpu.i_core.mepc[5] ;
 wire \i_tinyqv.cpu.i_core.mepc[6] ;
 wire \i_tinyqv.cpu.i_core.mepc[7] ;
 wire \i_tinyqv.cpu.i_core.mepc[8] ;
 wire \i_tinyqv.cpu.i_core.mepc[9] ;
 wire \i_tinyqv.cpu.i_core.mie[16] ;
 wire \i_tinyqv.cpu.i_core.mie[17] ;
 wire \i_tinyqv.cpu.i_core.mie[18] ;
 wire \i_tinyqv.cpu.i_core.mie[19] ;
 wire \i_tinyqv.cpu.i_core.mip[16] ;
 wire \i_tinyqv.cpu.i_core.mip[17] ;
 wire \i_tinyqv.cpu.i_core.mstatus_mie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mpie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mte ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[0] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[10] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[11] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[12] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[13] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[14] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[15] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[1] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[2] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[3] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[4] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[5] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[6] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[7] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[8] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[9] ;
 wire \i_tinyqv.cpu.i_core.time_hi[0] ;
 wire \i_tinyqv.cpu.i_core.time_hi[1] ;
 wire \i_tinyqv.cpu.i_core.time_hi[2] ;
 wire \i_tinyqv.cpu.imm[12] ;
 wire \i_tinyqv.cpu.imm[13] ;
 wire \i_tinyqv.cpu.imm[14] ;
 wire \i_tinyqv.cpu.imm[15] ;
 wire \i_tinyqv.cpu.imm[16] ;
 wire \i_tinyqv.cpu.imm[17] ;
 wire \i_tinyqv.cpu.imm[18] ;
 wire \i_tinyqv.cpu.imm[19] ;
 wire \i_tinyqv.cpu.imm[20] ;
 wire \i_tinyqv.cpu.imm[21] ;
 wire \i_tinyqv.cpu.imm[22] ;
 wire \i_tinyqv.cpu.imm[23] ;
 wire \i_tinyqv.cpu.imm[24] ;
 wire \i_tinyqv.cpu.imm[25] ;
 wire \i_tinyqv.cpu.imm[26] ;
 wire \i_tinyqv.cpu.imm[27] ;
 wire \i_tinyqv.cpu.imm[28] ;
 wire \i_tinyqv.cpu.imm[29] ;
 wire \i_tinyqv.cpu.imm[30] ;
 wire \i_tinyqv.cpu.imm[31] ;
 wire \i_tinyqv.cpu.instr_data[0][0] ;
 wire \i_tinyqv.cpu.instr_data[0][10] ;
 wire \i_tinyqv.cpu.instr_data[0][11] ;
 wire \i_tinyqv.cpu.instr_data[0][12] ;
 wire \i_tinyqv.cpu.instr_data[0][13] ;
 wire \i_tinyqv.cpu.instr_data[0][14] ;
 wire \i_tinyqv.cpu.instr_data[0][15] ;
 wire \i_tinyqv.cpu.instr_data[0][1] ;
 wire \i_tinyqv.cpu.instr_data[0][2] ;
 wire \i_tinyqv.cpu.instr_data[0][3] ;
 wire \i_tinyqv.cpu.instr_data[0][4] ;
 wire \i_tinyqv.cpu.instr_data[0][5] ;
 wire \i_tinyqv.cpu.instr_data[0][6] ;
 wire \i_tinyqv.cpu.instr_data[0][7] ;
 wire \i_tinyqv.cpu.instr_data[0][8] ;
 wire \i_tinyqv.cpu.instr_data[0][9] ;
 wire \i_tinyqv.cpu.instr_data[1][0] ;
 wire \i_tinyqv.cpu.instr_data[1][10] ;
 wire \i_tinyqv.cpu.instr_data[1][11] ;
 wire \i_tinyqv.cpu.instr_data[1][12] ;
 wire \i_tinyqv.cpu.instr_data[1][13] ;
 wire \i_tinyqv.cpu.instr_data[1][14] ;
 wire \i_tinyqv.cpu.instr_data[1][15] ;
 wire \i_tinyqv.cpu.instr_data[1][1] ;
 wire \i_tinyqv.cpu.instr_data[1][2] ;
 wire \i_tinyqv.cpu.instr_data[1][3] ;
 wire \i_tinyqv.cpu.instr_data[1][4] ;
 wire \i_tinyqv.cpu.instr_data[1][5] ;
 wire \i_tinyqv.cpu.instr_data[1][6] ;
 wire \i_tinyqv.cpu.instr_data[1][7] ;
 wire \i_tinyqv.cpu.instr_data[1][8] ;
 wire \i_tinyqv.cpu.instr_data[1][9] ;
 wire \i_tinyqv.cpu.instr_data[2][0] ;
 wire \i_tinyqv.cpu.instr_data[2][10] ;
 wire \i_tinyqv.cpu.instr_data[2][11] ;
 wire \i_tinyqv.cpu.instr_data[2][12] ;
 wire \i_tinyqv.cpu.instr_data[2][13] ;
 wire \i_tinyqv.cpu.instr_data[2][14] ;
 wire \i_tinyqv.cpu.instr_data[2][15] ;
 wire \i_tinyqv.cpu.instr_data[2][1] ;
 wire \i_tinyqv.cpu.instr_data[2][2] ;
 wire \i_tinyqv.cpu.instr_data[2][3] ;
 wire \i_tinyqv.cpu.instr_data[2][4] ;
 wire \i_tinyqv.cpu.instr_data[2][5] ;
 wire \i_tinyqv.cpu.instr_data[2][6] ;
 wire \i_tinyqv.cpu.instr_data[2][7] ;
 wire \i_tinyqv.cpu.instr_data[2][8] ;
 wire \i_tinyqv.cpu.instr_data[2][9] ;
 wire \i_tinyqv.cpu.instr_data[3][0] ;
 wire \i_tinyqv.cpu.instr_data[3][10] ;
 wire \i_tinyqv.cpu.instr_data[3][11] ;
 wire \i_tinyqv.cpu.instr_data[3][12] ;
 wire \i_tinyqv.cpu.instr_data[3][13] ;
 wire \i_tinyqv.cpu.instr_data[3][14] ;
 wire \i_tinyqv.cpu.instr_data[3][15] ;
 wire \i_tinyqv.cpu.instr_data[3][1] ;
 wire \i_tinyqv.cpu.instr_data[3][2] ;
 wire \i_tinyqv.cpu.instr_data[3][3] ;
 wire \i_tinyqv.cpu.instr_data[3][4] ;
 wire \i_tinyqv.cpu.instr_data[3][5] ;
 wire \i_tinyqv.cpu.instr_data[3][6] ;
 wire \i_tinyqv.cpu.instr_data[3][7] ;
 wire \i_tinyqv.cpu.instr_data[3][8] ;
 wire \i_tinyqv.cpu.instr_data[3][9] ;
 wire \i_tinyqv.cpu.instr_data_in[0] ;
 wire \i_tinyqv.cpu.instr_data_in[10] ;
 wire \i_tinyqv.cpu.instr_data_in[11] ;
 wire \i_tinyqv.cpu.instr_data_in[12] ;
 wire \i_tinyqv.cpu.instr_data_in[13] ;
 wire \i_tinyqv.cpu.instr_data_in[14] ;
 wire \i_tinyqv.cpu.instr_data_in[15] ;
 wire \i_tinyqv.cpu.instr_data_in[1] ;
 wire \i_tinyqv.cpu.instr_data_in[2] ;
 wire \i_tinyqv.cpu.instr_data_in[3] ;
 wire \i_tinyqv.cpu.instr_data_in[4] ;
 wire \i_tinyqv.cpu.instr_data_in[5] ;
 wire \i_tinyqv.cpu.instr_data_in[6] ;
 wire \i_tinyqv.cpu.instr_data_in[7] ;
 wire \i_tinyqv.cpu.instr_data_in[8] ;
 wire \i_tinyqv.cpu.instr_data_in[9] ;
 wire \i_tinyqv.cpu.instr_data_start[10] ;
 wire \i_tinyqv.cpu.instr_data_start[11] ;
 wire \i_tinyqv.cpu.instr_data_start[12] ;
 wire \i_tinyqv.cpu.instr_data_start[13] ;
 wire \i_tinyqv.cpu.instr_data_start[14] ;
 wire \i_tinyqv.cpu.instr_data_start[15] ;
 wire \i_tinyqv.cpu.instr_data_start[16] ;
 wire \i_tinyqv.cpu.instr_data_start[17] ;
 wire \i_tinyqv.cpu.instr_data_start[18] ;
 wire \i_tinyqv.cpu.instr_data_start[19] ;
 wire \i_tinyqv.cpu.instr_data_start[20] ;
 wire \i_tinyqv.cpu.instr_data_start[21] ;
 wire \i_tinyqv.cpu.instr_data_start[22] ;
 wire \i_tinyqv.cpu.instr_data_start[23] ;
 wire \i_tinyqv.cpu.instr_data_start[3] ;
 wire \i_tinyqv.cpu.instr_data_start[4] ;
 wire \i_tinyqv.cpu.instr_data_start[5] ;
 wire \i_tinyqv.cpu.instr_data_start[6] ;
 wire \i_tinyqv.cpu.instr_data_start[7] ;
 wire \i_tinyqv.cpu.instr_data_start[8] ;
 wire \i_tinyqv.cpu.instr_data_start[9] ;
 wire \i_tinyqv.cpu.instr_fetch_running ;
 wire \i_tinyqv.cpu.instr_fetch_started ;
 wire \i_tinyqv.cpu.instr_fetch_stopped ;
 wire \i_tinyqv.cpu.instr_len[1] ;
 wire \i_tinyqv.cpu.instr_len[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[1] ;
 wire \i_tinyqv.cpu.instr_write_offset[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[3] ;
 wire \i_tinyqv.cpu.is_alu_imm ;
 wire \i_tinyqv.cpu.is_alu_reg ;
 wire \i_tinyqv.cpu.is_auipc ;
 wire \i_tinyqv.cpu.is_branch ;
 wire \i_tinyqv.cpu.is_jal ;
 wire \i_tinyqv.cpu.is_jalr ;
 wire \i_tinyqv.cpu.is_load ;
 wire \i_tinyqv.cpu.is_lui ;
 wire \i_tinyqv.cpu.is_store ;
 wire \i_tinyqv.cpu.is_system ;
 wire \i_tinyqv.cpu.load_started ;
 wire \i_tinyqv.cpu.mem_op_increment_reg ;
 wire \i_tinyqv.cpu.no_write_in_progress ;
 wire \i_tinyqv.cpu.pc[1] ;
 wire \i_tinyqv.cpu.pc[2] ;
 wire \i_tinyqv.cpu.was_early_branch ;
 wire \i_tinyqv.mem.data_from_read[16] ;
 wire \i_tinyqv.mem.data_from_read[17] ;
 wire \i_tinyqv.mem.data_from_read[18] ;
 wire \i_tinyqv.mem.data_from_read[19] ;
 wire \i_tinyqv.mem.data_from_read[20] ;
 wire \i_tinyqv.mem.data_from_read[21] ;
 wire \i_tinyqv.mem.data_from_read[22] ;
 wire \i_tinyqv.mem.data_from_read[23] ;
 wire \i_tinyqv.mem.data_stall ;
 wire \i_tinyqv.mem.instr_active ;
 wire \i_tinyqv.mem.q_ctrl.addr[0] ;
 wire \i_tinyqv.mem.q_ctrl.addr[10] ;
 wire \i_tinyqv.mem.q_ctrl.addr[11] ;
 wire \i_tinyqv.mem.q_ctrl.addr[12] ;
 wire \i_tinyqv.mem.q_ctrl.addr[13] ;
 wire \i_tinyqv.mem.q_ctrl.addr[14] ;
 wire \i_tinyqv.mem.q_ctrl.addr[15] ;
 wire \i_tinyqv.mem.q_ctrl.addr[16] ;
 wire \i_tinyqv.mem.q_ctrl.addr[17] ;
 wire \i_tinyqv.mem.q_ctrl.addr[18] ;
 wire \i_tinyqv.mem.q_ctrl.addr[19] ;
 wire \i_tinyqv.mem.q_ctrl.addr[1] ;
 wire \i_tinyqv.mem.q_ctrl.addr[20] ;
 wire \i_tinyqv.mem.q_ctrl.addr[21] ;
 wire \i_tinyqv.mem.q_ctrl.addr[22] ;
 wire \i_tinyqv.mem.q_ctrl.addr[23] ;
 wire \i_tinyqv.mem.q_ctrl.addr[2] ;
 wire \i_tinyqv.mem.q_ctrl.addr[3] ;
 wire \i_tinyqv.mem.q_ctrl.addr[4] ;
 wire \i_tinyqv.mem.q_ctrl.addr[5] ;
 wire \i_tinyqv.mem.q_ctrl.addr[6] ;
 wire \i_tinyqv.mem.q_ctrl.addr[7] ;
 wire \i_tinyqv.mem.q_ctrl.addr[8] ;
 wire \i_tinyqv.mem.q_ctrl.addr[9] ;
 wire \i_tinyqv.mem.q_ctrl.data_ready ;
 wire \i_tinyqv.mem.q_ctrl.data_req ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[0] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[1] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[2] ;
 wire \i_tinyqv.mem.q_ctrl.is_writing ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_a_sel ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_b_sel ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[0] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[1] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[2] ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_out ;
 wire \i_tinyqv.mem.q_ctrl.spi_data_oe[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_flash_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_a_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_b_select ;
 wire \i_tinyqv.mem.q_ctrl.stop_txn_reg ;
 wire \i_tinyqv.mem.qspi_data_buf[10] ;
 wire \i_tinyqv.mem.qspi_data_buf[11] ;
 wire \i_tinyqv.mem.qspi_data_buf[12] ;
 wire \i_tinyqv.mem.qspi_data_buf[13] ;
 wire \i_tinyqv.mem.qspi_data_buf[14] ;
 wire \i_tinyqv.mem.qspi_data_buf[15] ;
 wire \i_tinyqv.mem.qspi_data_buf[24] ;
 wire \i_tinyqv.mem.qspi_data_buf[25] ;
 wire \i_tinyqv.mem.qspi_data_buf[26] ;
 wire \i_tinyqv.mem.qspi_data_buf[27] ;
 wire \i_tinyqv.mem.qspi_data_buf[28] ;
 wire \i_tinyqv.mem.qspi_data_buf[29] ;
 wire \i_tinyqv.mem.qspi_data_buf[30] ;
 wire \i_tinyqv.mem.qspi_data_buf[31] ;
 wire \i_tinyqv.mem.qspi_data_buf[8] ;
 wire \i_tinyqv.mem.qspi_data_buf[9] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[0] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[1] ;
 wire \i_tinyqv.mem.qspi_write_done ;
 wire \i_uart_rx.bit_sample ;
 wire \i_uart_rx.cycle_counter[0] ;
 wire \i_uart_rx.cycle_counter[10] ;
 wire \i_uart_rx.cycle_counter[1] ;
 wire \i_uart_rx.cycle_counter[2] ;
 wire \i_uart_rx.cycle_counter[3] ;
 wire \i_uart_rx.cycle_counter[4] ;
 wire \i_uart_rx.cycle_counter[5] ;
 wire \i_uart_rx.cycle_counter[6] ;
 wire \i_uart_rx.cycle_counter[7] ;
 wire \i_uart_rx.cycle_counter[8] ;
 wire \i_uart_rx.cycle_counter[9] ;
 wire \i_uart_rx.fsm_state[0] ;
 wire \i_uart_rx.fsm_state[1] ;
 wire \i_uart_rx.fsm_state[2] ;
 wire \i_uart_rx.fsm_state[3] ;
 wire \i_uart_rx.recieved_data[0] ;
 wire \i_uart_rx.recieved_data[1] ;
 wire \i_uart_rx.recieved_data[2] ;
 wire \i_uart_rx.recieved_data[3] ;
 wire \i_uart_rx.recieved_data[4] ;
 wire \i_uart_rx.recieved_data[5] ;
 wire \i_uart_rx.recieved_data[6] ;
 wire \i_uart_rx.recieved_data[7] ;
 wire \i_uart_rx.rxd_reg[0] ;
 wire \i_uart_rx.rxd_reg[1] ;
 wire \i_uart_rx.uart_rts ;
 wire \i_uart_tx.cycle_counter[0] ;
 wire \i_uart_tx.cycle_counter[10] ;
 wire \i_uart_tx.cycle_counter[1] ;
 wire \i_uart_tx.cycle_counter[2] ;
 wire \i_uart_tx.cycle_counter[3] ;
 wire \i_uart_tx.cycle_counter[4] ;
 wire \i_uart_tx.cycle_counter[5] ;
 wire \i_uart_tx.cycle_counter[6] ;
 wire \i_uart_tx.cycle_counter[7] ;
 wire \i_uart_tx.cycle_counter[8] ;
 wire \i_uart_tx.cycle_counter[9] ;
 wire \i_uart_tx.data_to_send[0] ;
 wire \i_uart_tx.data_to_send[1] ;
 wire \i_uart_tx.data_to_send[2] ;
 wire \i_uart_tx.data_to_send[3] ;
 wire \i_uart_tx.data_to_send[4] ;
 wire \i_uart_tx.data_to_send[5] ;
 wire \i_uart_tx.data_to_send[6] ;
 wire \i_uart_tx.data_to_send[7] ;
 wire \i_uart_tx.fsm_state[0] ;
 wire \i_uart_tx.fsm_state[1] ;
 wire \i_uart_tx.fsm_state[2] ;
 wire \i_uart_tx.fsm_state[3] ;
 wire \i_uart_tx.txd_reg ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _06029_ (.A(\i_tinyqv.cpu.alu_op[1] ),
    .X(_00745_));
 sg13g2_buf_1 _06030_ (.A(\i_tinyqv.cpu.alu_op[2] ),
    .X(_00746_));
 sg13g2_and2_1 _06031_ (.A(_00745_),
    .B(net315),
    .X(_00747_));
 sg13g2_buf_1 _06032_ (.A(_00747_),
    .X(_00748_));
 sg13g2_nand2b_1 _06033_ (.Y(_00749_),
    .B(_00748_),
    .A_N(_00085_));
 sg13g2_buf_1 _06034_ (.A(_00749_),
    .X(_00750_));
 sg13g2_buf_2 _06035_ (.A(debug_instr_valid),
    .X(_00751_));
 sg13g2_o21ai_1 _06036_ (.B1(_00751_),
    .Y(_00752_),
    .A1(\i_tinyqv.cpu.is_auipc ),
    .A2(\i_tinyqv.cpu.is_jal ));
 sg13g2_buf_2 _06037_ (.A(_00752_),
    .X(_00753_));
 sg13g2_buf_1 _06038_ (.A(\i_tinyqv.cpu.counter[3] ),
    .X(_00754_));
 sg13g2_buf_1 _06039_ (.A(_00754_),
    .X(_00755_));
 sg13g2_inv_2 _06040_ (.Y(_00756_),
    .A(net277));
 sg13g2_buf_1 _06041_ (.A(_00756_),
    .X(_00757_));
 sg13g2_buf_2 _06042_ (.A(\i_tinyqv.cpu.pc[2] ),
    .X(_00758_));
 sg13g2_buf_1 _06043_ (.A(\i_tinyqv.cpu.instr_data_start[6] ),
    .X(_00759_));
 sg13g2_buf_1 _06044_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .X(_00760_));
 sg13g2_buf_2 _06045_ (.A(\i_tinyqv.cpu.counter[2] ),
    .X(_00761_));
 sg13g2_buf_8 _06046_ (.A(_00761_),
    .X(_00762_));
 sg13g2_buf_8 _06047_ (.A(net276),
    .X(_00763_));
 sg13g2_buf_1 _06048_ (.A(\i_tinyqv.cpu.counter[4] ),
    .X(_00764_));
 sg13g2_buf_1 _06049_ (.A(_00764_),
    .X(_00765_));
 sg13g2_buf_1 _06050_ (.A(net275),
    .X(_00766_));
 sg13g2_mux4_1 _06051_ (.S0(net228),
    .A0(_00758_),
    .A1(_00759_),
    .A2(\i_tinyqv.cpu.instr_data_start[18] ),
    .A3(_00760_),
    .S1(net227),
    .X(_00767_));
 sg13g2_buf_1 _06052_ (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .X(_00768_));
 sg13g2_buf_1 _06053_ (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .X(_00769_));
 sg13g2_buf_2 _06054_ (.A(net276),
    .X(_00770_));
 sg13g2_mux2_1 _06055_ (.A0(_00768_),
    .A1(_00769_),
    .S(net226),
    .X(_00771_));
 sg13g2_nor2_1 _06056_ (.A(_00756_),
    .B(_00765_),
    .Y(_00772_));
 sg13g2_a22oi_1 _06057_ (.Y(_00773_),
    .B1(_00771_),
    .B2(_00772_),
    .A2(_00767_),
    .A1(net211));
 sg13g2_nand2b_1 _06058_ (.Y(_00774_),
    .B(_00773_),
    .A_N(_00753_));
 sg13g2_buf_8 _06059_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .X(_00775_));
 sg13g2_buf_1 _06060_ (.A(net314),
    .X(_00776_));
 sg13g2_buf_8 _06061_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .X(_00777_));
 sg13g2_buf_1 _06062_ (.A(_00777_),
    .X(_00778_));
 sg13g2_buf_8 _06063_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .X(_00779_));
 sg13g2_buf_8 _06064_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .X(_00780_));
 sg13g2_and2_1 _06065_ (.A(_00779_),
    .B(_00780_),
    .X(_00781_));
 sg13g2_buf_1 _06066_ (.A(_00781_),
    .X(_00782_));
 sg13g2_buf_8 _06067_ (.A(_00779_),
    .X(_00783_));
 sg13g2_nor2_1 _06068_ (.A(net272),
    .B(_00780_),
    .Y(_00784_));
 sg13g2_a22oi_1 _06069_ (.Y(_00785_),
    .B1(_00784_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .A2(_00782_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ));
 sg13g2_buf_8 _06070_ (.A(_00780_),
    .X(_00786_));
 sg13g2_buf_8 _06071_ (.A(_00777_),
    .X(_00787_));
 sg13g2_nand3b_1 _06072_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .C(net270),
    .Y(_00788_),
    .A_N(net271));
 sg13g2_nand3b_1 _06073_ (.B(net271),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .Y(_00789_),
    .A_N(net270));
 sg13g2_buf_8 _06074_ (.A(net272),
    .X(_00790_));
 sg13g2_a21o_1 _06075_ (.A2(_00789_),
    .A1(_00788_),
    .B1(_00790_),
    .X(_00791_));
 sg13g2_o21ai_1 _06076_ (.B1(_00791_),
    .Y(_00792_),
    .A1(net273),
    .A2(_00785_));
 sg13g2_nand2_2 _06077_ (.Y(_00793_),
    .A(_00776_),
    .B(_00792_));
 sg13g2_inv_4 _06078_ (.A(_00786_),
    .Y(_00794_));
 sg13g2_and2_1 _06079_ (.A(_00779_),
    .B(net314),
    .X(_00795_));
 sg13g2_buf_8 _06080_ (.A(_00795_),
    .X(_00796_));
 sg13g2_mux2_1 _06081_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .S(_00777_),
    .X(_00797_));
 sg13g2_and3_1 _06082_ (.X(_00798_),
    .A(_00794_),
    .B(_00796_),
    .C(_00797_));
 sg13g2_inv_2 _06083_ (.Y(_00799_),
    .A(_00775_));
 sg13g2_mux2_1 _06084_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .S(_00780_),
    .X(_00800_));
 sg13g2_nor2b_1 _06085_ (.A(_00783_),
    .B_N(_00777_),
    .Y(_00801_));
 sg13g2_and3_1 _06086_ (.X(_00802_),
    .A(_00799_),
    .B(_00800_),
    .C(_00801_));
 sg13g2_nand2_1 _06087_ (.Y(_00803_),
    .A(_00779_),
    .B(_00777_));
 sg13g2_nor4_1 _06088_ (.A(_00799_),
    .B(_00794_),
    .C(_00090_),
    .D(_00803_),
    .Y(_00804_));
 sg13g2_nand2b_2 _06089_ (.Y(_00805_),
    .B(_00754_),
    .A_N(_00761_));
 sg13g2_or2_1 _06090_ (.X(_00806_),
    .B(_00780_),
    .A(_00775_));
 sg13g2_nor4_1 _06091_ (.A(_00764_),
    .B(_00805_),
    .C(_00803_),
    .D(_00806_),
    .Y(_00807_));
 sg13g2_nor4_1 _06092_ (.A(_00798_),
    .B(_00802_),
    .C(_00804_),
    .D(_00807_),
    .Y(_00808_));
 sg13g2_nor2b_1 _06093_ (.A(net270),
    .B_N(_00779_),
    .Y(_00809_));
 sg13g2_nand3_1 _06094_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .C(_00809_),
    .A(_00799_),
    .Y(_00810_));
 sg13g2_nand3_1 _06095_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .C(_00801_),
    .A(net274),
    .Y(_00811_));
 sg13g2_a21o_1 _06096_ (.A2(_00811_),
    .A1(_00810_),
    .B1(_00794_),
    .X(_00812_));
 sg13g2_inv_1 _06097_ (.Y(_00813_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ));
 sg13g2_or2_1 _06098_ (.X(_00814_),
    .B(net271),
    .A(net270));
 sg13g2_nand3_1 _06099_ (.B(net271),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .A(_00778_),
    .Y(_00815_));
 sg13g2_o21ai_1 _06100_ (.B1(_00815_),
    .Y(_00816_),
    .A1(_00813_),
    .A2(_00814_));
 sg13g2_nand3_1 _06101_ (.B(_00799_),
    .C(_00816_),
    .A(net225),
    .Y(_00817_));
 sg13g2_and3_1 _06102_ (.X(_00818_),
    .A(_00808_),
    .B(_00812_),
    .C(_00817_));
 sg13g2_buf_2 _06103_ (.A(_00818_),
    .X(_00819_));
 sg13g2_nand3_1 _06104_ (.B(_00793_),
    .C(_00819_),
    .A(_00753_),
    .Y(_00820_));
 sg13g2_nand3_1 _06105_ (.B(_00774_),
    .C(_00820_),
    .A(_00750_),
    .Y(_00821_));
 sg13g2_buf_2 _06106_ (.A(_00821_),
    .X(_00822_));
 sg13g2_buf_1 _06107_ (.A(\i_tinyqv.cpu.alu_op[3] ),
    .X(_00823_));
 sg13g2_buf_1 _06108_ (.A(_00089_),
    .X(_00824_));
 sg13g2_nor2b_1 _06109_ (.A(net313),
    .B_N(_00824_),
    .Y(_00825_));
 sg13g2_a21o_1 _06110_ (.A2(_00748_),
    .A1(net313),
    .B1(_00825_),
    .X(_00826_));
 sg13g2_buf_1 _06111_ (.A(_00826_),
    .X(_00827_));
 sg13g2_and2_1 _06112_ (.A(net314),
    .B(net271),
    .X(_00828_));
 sg13g2_buf_1 _06113_ (.A(_00780_),
    .X(_00829_));
 sg13g2_mux2_1 _06114_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .S(_00829_),
    .X(_00830_));
 sg13g2_a22oi_1 _06115_ (.Y(_00831_),
    .B1(_00830_),
    .B2(_00799_),
    .A2(_00828_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ));
 sg13g2_nand3b_1 _06116_ (.B(_00764_),
    .C(_00754_),
    .Y(_00832_),
    .A_N(_00761_));
 sg13g2_buf_1 _06117_ (.A(_00832_),
    .X(_00833_));
 sg13g2_nor2b_1 _06118_ (.A(net314),
    .B_N(_00780_),
    .Y(_00834_));
 sg13g2_buf_2 _06119_ (.A(_00834_),
    .X(_00835_));
 sg13g2_nand2b_1 _06120_ (.Y(_00836_),
    .B(_00835_),
    .A_N(_00833_));
 sg13g2_nor2b_1 _06121_ (.A(net271),
    .B_N(net314),
    .Y(_00837_));
 sg13g2_a21oi_1 _06122_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .A2(_00837_),
    .Y(_00838_),
    .B1(_00790_));
 sg13g2_a221oi_1 _06123_ (.B2(_00838_),
    .C1(net273),
    .B1(_00836_),
    .A1(net225),
    .Y(_00839_),
    .A2(_00831_));
 sg13g2_inv_2 _06124_ (.Y(_00840_),
    .A(_00777_));
 sg13g2_inv_1 _06125_ (.Y(_00841_),
    .A(_00087_));
 sg13g2_a22oi_1 _06126_ (.Y(_00842_),
    .B1(_00784_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .A2(_00782_),
    .A1(_00841_));
 sg13g2_nor3_1 _06127_ (.A(_00840_),
    .B(_00799_),
    .C(_00842_),
    .Y(_00843_));
 sg13g2_nor2_1 _06128_ (.A(net225),
    .B(net274),
    .Y(_00844_));
 sg13g2_a22oi_1 _06129_ (.Y(_00845_),
    .B1(_00844_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .A2(_00796_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ));
 sg13g2_nor3_1 _06130_ (.A(_00840_),
    .B(net269),
    .C(_00845_),
    .Y(_00846_));
 sg13g2_nand3b_1 _06131_ (.B(net269),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .Y(_00847_),
    .A_N(net225));
 sg13g2_nand3b_1 _06132_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .C(net225),
    .Y(_00848_),
    .A_N(net269));
 sg13g2_nand2b_1 _06133_ (.Y(_00849_),
    .B(net274),
    .A_N(net273));
 sg13g2_a21o_1 _06134_ (.A2(_00848_),
    .A1(_00847_),
    .B1(_00849_),
    .X(_00850_));
 sg13g2_mux2_1 _06135_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .S(net274),
    .X(_00851_));
 sg13g2_nand3_1 _06136_ (.B(_00801_),
    .C(_00851_),
    .A(net269),
    .Y(_00852_));
 sg13g2_nand4_1 _06137_ (.B(net273),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .A(net225),
    .Y(_00853_),
    .D(_00835_));
 sg13g2_nand3_1 _06138_ (.B(_00852_),
    .C(_00853_),
    .A(_00850_),
    .Y(_00854_));
 sg13g2_nor4_1 _06139_ (.A(_00839_),
    .B(_00843_),
    .C(_00846_),
    .D(_00854_),
    .Y(_00855_));
 sg13g2_buf_1 _06140_ (.A(_00855_),
    .X(_00856_));
 sg13g2_buf_1 _06141_ (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .X(_00857_));
 sg13g2_buf_1 _06142_ (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .X(_00858_));
 sg13g2_buf_2 _06143_ (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .X(_00859_));
 sg13g2_mux4_1 _06144_ (.S0(net228),
    .A0(_00857_),
    .A1(_00858_),
    .A2(_00859_),
    .A3(\i_tinyqv.cpu.instr_data_start[23] ),
    .S1(net275),
    .X(_00860_));
 sg13g2_buf_1 _06145_ (.A(\i_tinyqv.cpu.instr_data_start[15] ),
    .X(_00861_));
 sg13g2_mux2_1 _06146_ (.A0(\i_tinyqv.cpu.instr_data_start[11] ),
    .A1(_00861_),
    .S(net228),
    .X(_00862_));
 sg13g2_a22oi_1 _06147_ (.Y(_00863_),
    .B1(_00862_),
    .B2(_00772_),
    .A2(_00860_),
    .A1(_00756_));
 sg13g2_nor2b_1 _06148_ (.A(_00753_),
    .B_N(_00863_),
    .Y(_00864_));
 sg13g2_a21oi_1 _06149_ (.A1(_00753_),
    .A2(net154),
    .Y(_00865_),
    .B1(_00864_));
 sg13g2_nand2_1 _06150_ (.Y(_00866_),
    .A(_00750_),
    .B(_00865_));
 sg13g2_buf_2 _06151_ (.A(_00866_),
    .X(_00867_));
 sg13g2_buf_1 _06152_ (.A(\i_tinyqv.cpu.is_branch ),
    .X(_00868_));
 sg13g2_nor2_1 _06153_ (.A(\i_tinyqv.cpu.is_alu_reg ),
    .B(_00868_),
    .Y(_00869_));
 sg13g2_nor2b_1 _06154_ (.A(_00869_),
    .B_N(_00751_),
    .Y(_00870_));
 sg13g2_buf_1 _06155_ (.A(_00870_),
    .X(_00871_));
 sg13g2_buf_8 _06156_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .X(_00872_));
 sg13g2_buf_8 _06157_ (.A(_00872_),
    .X(_00873_));
 sg13g2_buf_8 _06158_ (.A(net268),
    .X(_00874_));
 sg13g2_inv_2 _06159_ (.Y(_00875_),
    .A(_00874_));
 sg13g2_buf_8 _06160_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .X(_00876_));
 sg13g2_buf_8 _06161_ (.A(_00876_),
    .X(_00877_));
 sg13g2_buf_8 _06162_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .X(_00878_));
 sg13g2_buf_8 _06163_ (.A(_00878_),
    .X(_00879_));
 sg13g2_nor2b_1 _06164_ (.A(_00877_),
    .B_N(_00879_),
    .Y(_00880_));
 sg13g2_mux2_1 _06165_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .S(_00879_),
    .X(_00881_));
 sg13g2_buf_8 _06166_ (.A(net267),
    .X(_00882_));
 sg13g2_buf_1 _06167_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .X(_00883_));
 sg13g2_buf_1 _06168_ (.A(_00883_),
    .X(_00884_));
 sg13g2_buf_1 _06169_ (.A(net265),
    .X(_00885_));
 sg13g2_a221oi_1 _06170_ (.B2(net223),
    .C1(net222),
    .B1(_00881_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .Y(_00886_),
    .A2(_00880_));
 sg13g2_buf_8 _06171_ (.A(net266),
    .X(_00887_));
 sg13g2_nor2b_1 _06172_ (.A(net221),
    .B_N(net267),
    .Y(_00888_));
 sg13g2_inv_1 _06173_ (.Y(_00889_),
    .A(_00883_));
 sg13g2_a221oi_1 _06174_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .C1(_00889_),
    .B1(_00888_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .Y(_00890_),
    .A2(_00880_));
 sg13g2_nor3_1 _06175_ (.A(_00875_),
    .B(_00886_),
    .C(_00890_),
    .Y(_00891_));
 sg13g2_inv_2 _06176_ (.Y(_00892_),
    .A(_00765_));
 sg13g2_nor2_1 _06177_ (.A(_00756_),
    .B(net228),
    .Y(_00893_));
 sg13g2_nor2_1 _06178_ (.A(net268),
    .B(net265),
    .Y(_00894_));
 sg13g2_nand3_1 _06179_ (.B(_00893_),
    .C(_00894_),
    .A(_00892_),
    .Y(_00895_));
 sg13g2_nor2_1 _06180_ (.A(_00875_),
    .B(_00090_),
    .Y(_00896_));
 sg13g2_nor2b_1 _06181_ (.A(net224),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .Y(_00897_));
 sg13g2_o21ai_1 _06182_ (.B1(_00885_),
    .Y(_00898_),
    .A1(_00896_),
    .A2(_00897_));
 sg13g2_nand2_1 _06183_ (.Y(_00899_),
    .A(_00876_),
    .B(_00878_));
 sg13g2_a21oi_1 _06184_ (.A1(_00895_),
    .A2(_00898_),
    .Y(_00900_),
    .B1(_00899_));
 sg13g2_nor2_1 _06185_ (.A(_00889_),
    .B(net267),
    .Y(_00901_));
 sg13g2_inv_2 _06186_ (.Y(_00902_),
    .A(net223));
 sg13g2_nor2_1 _06187_ (.A(net222),
    .B(_00902_),
    .Y(_00903_));
 sg13g2_a22oi_1 _06188_ (.Y(_00904_),
    .B1(_00903_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .A2(_00901_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ));
 sg13g2_nor2_1 _06189_ (.A(_00872_),
    .B(_00878_),
    .Y(_00905_));
 sg13g2_nor2b_1 _06190_ (.A(_00904_),
    .B_N(_00905_),
    .Y(_00906_));
 sg13g2_nand2_1 _06191_ (.Y(_00907_),
    .A(_00875_),
    .B(_00885_));
 sg13g2_a22oi_1 _06192_ (.Y(_00908_),
    .B1(_00888_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .A2(_00880_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ));
 sg13g2_nand3_1 _06193_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .C(_00894_),
    .A(net221),
    .Y(_00909_));
 sg13g2_inv_1 _06194_ (.Y(_00910_),
    .A(_00878_));
 sg13g2_and2_1 _06195_ (.A(net268),
    .B(net265),
    .X(_00911_));
 sg13g2_buf_1 _06196_ (.A(_00911_),
    .X(_00912_));
 sg13g2_nand3_1 _06197_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .C(_00912_),
    .A(_00910_),
    .Y(_00913_));
 sg13g2_a21o_1 _06198_ (.A2(_00913_),
    .A1(_00909_),
    .B1(net223),
    .X(_00914_));
 sg13g2_o21ai_1 _06199_ (.B1(_00914_),
    .Y(_00915_),
    .A1(_00907_),
    .A2(_00908_));
 sg13g2_nor4_2 _06200_ (.A(_00891_),
    .B(_00900_),
    .C(_00906_),
    .Y(_00916_),
    .D(_00915_));
 sg13g2_buf_2 _06201_ (.A(\i_tinyqv.cpu.imm[14] ),
    .X(_00917_));
 sg13g2_mux4_1 _06202_ (.S0(net228),
    .A0(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .A1(_00917_),
    .A2(\i_tinyqv.cpu.imm[26] ),
    .A3(\i_tinyqv.cpu.imm[30] ),
    .S1(net275),
    .X(_00918_));
 sg13g2_buf_1 _06203_ (.A(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .X(_00919_));
 sg13g2_buf_2 _06204_ (.A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .X(_00920_));
 sg13g2_buf_2 _06205_ (.A(\i_tinyqv.cpu.imm[18] ),
    .X(_00921_));
 sg13g2_mux4_1 _06206_ (.S0(net228),
    .A0(net311),
    .A1(_00920_),
    .A2(_00921_),
    .A3(\i_tinyqv.cpu.imm[22] ),
    .S1(net275),
    .X(_00922_));
 sg13g2_mux2_1 _06207_ (.A0(_00918_),
    .A1(_00922_),
    .S(_00756_),
    .X(_00923_));
 sg13g2_buf_1 _06208_ (.A(_00923_),
    .X(_00924_));
 sg13g2_nor2_1 _06209_ (.A(_00871_),
    .B(_00924_),
    .Y(_00925_));
 sg13g2_a21oi_1 _06210_ (.A1(_00871_),
    .A2(_00916_),
    .Y(_00926_),
    .B1(_00925_));
 sg13g2_buf_2 _06211_ (.A(_00926_),
    .X(_00927_));
 sg13g2_mux2_1 _06212_ (.A0(net193),
    .A1(_00867_),
    .S(_00927_),
    .X(_00928_));
 sg13g2_a21oi_1 _06213_ (.A1(net313),
    .A2(_00748_),
    .Y(_00929_),
    .B1(_00825_));
 sg13g2_buf_2 _06214_ (.A(_00929_),
    .X(_00930_));
 sg13g2_mux2_1 _06215_ (.A0(_00867_),
    .A1(_00930_),
    .S(_00927_),
    .X(_00931_));
 sg13g2_o21ai_1 _06216_ (.B1(_00751_),
    .Y(_00932_),
    .A1(\i_tinyqv.cpu.is_alu_reg ),
    .A2(_00868_));
 sg13g2_mux2_1 _06217_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .S(net221),
    .X(_00933_));
 sg13g2_nor3_1 _06218_ (.A(net223),
    .B(_00887_),
    .C(_00833_),
    .Y(_00934_));
 sg13g2_a21o_1 _06219_ (.A2(_00933_),
    .A1(net223),
    .B1(_00934_),
    .X(_00935_));
 sg13g2_nor2b_1 _06220_ (.A(_00883_),
    .B_N(_00872_),
    .Y(_00936_));
 sg13g2_and2_1 _06221_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .B(net223),
    .X(_00937_));
 sg13g2_a21oi_1 _06222_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .A2(_00902_),
    .Y(_00938_),
    .B1(_00937_));
 sg13g2_nor3_1 _06223_ (.A(_00889_),
    .B(net221),
    .C(_00938_),
    .Y(_00939_));
 sg13g2_and2_1 _06224_ (.A(net265),
    .B(_00878_),
    .X(_00940_));
 sg13g2_nor2_1 _06225_ (.A(net265),
    .B(net266),
    .Y(_00941_));
 sg13g2_a22oi_1 _06226_ (.Y(_00942_),
    .B1(_00941_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .A2(_00940_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ));
 sg13g2_nor2b_1 _06227_ (.A(_00087_),
    .B_N(net266),
    .Y(_00943_));
 sg13g2_nor2b_1 _06228_ (.A(net266),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .Y(_00944_));
 sg13g2_o21ai_1 _06229_ (.B1(_00912_),
    .Y(_00945_),
    .A1(_00943_),
    .A2(_00944_));
 sg13g2_o21ai_1 _06230_ (.B1(_00945_),
    .Y(_00946_),
    .A1(net224),
    .A2(_00942_));
 sg13g2_mux2_1 _06231_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .S(_00884_),
    .X(_00947_));
 sg13g2_a22oi_1 _06232_ (.Y(_00948_),
    .B1(_00947_),
    .B2(_00875_),
    .A2(_00936_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ));
 sg13g2_mux2_1 _06233_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .S(net266),
    .X(_00949_));
 sg13g2_nand2_1 _06234_ (.Y(_00950_),
    .A(_00912_),
    .B(_00949_));
 sg13g2_o21ai_1 _06235_ (.B1(_00950_),
    .Y(_00951_),
    .A1(_00910_),
    .A2(_00948_));
 sg13g2_mux2_1 _06236_ (.A0(_00946_),
    .A1(_00951_),
    .S(_00902_),
    .X(_00952_));
 sg13g2_a221oi_1 _06237_ (.B2(_00875_),
    .C1(_00952_),
    .B1(_00939_),
    .A1(_00935_),
    .Y(_00953_),
    .A2(_00936_));
 sg13g2_buf_1 _06238_ (.A(_00953_),
    .X(_00954_));
 sg13g2_buf_1 _06239_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .X(_00955_));
 sg13g2_buf_2 _06240_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .X(_00956_));
 sg13g2_mux2_1 _06241_ (.A0(_00955_),
    .A1(_00956_),
    .S(net276),
    .X(_00957_));
 sg13g2_nor2_1 _06242_ (.A(net277),
    .B(_00957_),
    .Y(_00958_));
 sg13g2_buf_2 _06243_ (.A(\i_tinyqv.cpu.imm[15] ),
    .X(_00959_));
 sg13g2_nand2_1 _06244_ (.Y(_00960_),
    .A(net277),
    .B(_00761_));
 sg13g2_buf_2 _06245_ (.A(_00960_),
    .X(_00961_));
 sg13g2_nor2_1 _06246_ (.A(_00959_),
    .B(_00961_),
    .Y(_00962_));
 sg13g2_o21ai_1 _06247_ (.B1(_00892_),
    .Y(_00963_),
    .A1(_00958_),
    .A2(_00962_));
 sg13g2_inv_1 _06248_ (.Y(_00964_),
    .A(net276));
 sg13g2_buf_2 _06249_ (.A(\i_tinyqv.cpu.imm[19] ),
    .X(_00965_));
 sg13g2_and2_1 _06250_ (.A(_00762_),
    .B(\i_tinyqv.cpu.imm[23] ),
    .X(_00966_));
 sg13g2_a21oi_1 _06251_ (.A1(_00964_),
    .A2(_00965_),
    .Y(_00967_),
    .B1(_00966_));
 sg13g2_nor2_1 _06252_ (.A(net277),
    .B(_00892_),
    .Y(_00968_));
 sg13g2_buf_1 _06253_ (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .X(_00969_));
 sg13g2_mux2_1 _06254_ (.A0(net310),
    .A1(\i_tinyqv.cpu.imm[27] ),
    .S(net275),
    .X(_00970_));
 sg13g2_nand3b_1 _06255_ (.B(net275),
    .C(net276),
    .Y(_00971_),
    .A_N(\i_tinyqv.cpu.imm[31] ));
 sg13g2_o21ai_1 _06256_ (.B1(_00971_),
    .Y(_00972_),
    .A1(net228),
    .A2(_00970_));
 sg13g2_a22oi_1 _06257_ (.Y(_00973_),
    .B1(_00972_),
    .B2(_00755_),
    .A2(_00968_),
    .A1(_00967_));
 sg13g2_and2_1 _06258_ (.A(_00963_),
    .B(_00973_),
    .X(_00974_));
 sg13g2_buf_1 _06259_ (.A(_00974_),
    .X(_00975_));
 sg13g2_nand2_1 _06260_ (.Y(_00976_),
    .A(_00932_),
    .B(_00975_));
 sg13g2_o21ai_1 _06261_ (.B1(_00976_),
    .Y(_00977_),
    .A1(_00932_),
    .A2(_00954_));
 sg13g2_buf_2 _06262_ (.A(_00977_),
    .X(_00978_));
 sg13g2_mux2_1 _06263_ (.A0(_00928_),
    .A1(_00931_),
    .S(_00978_),
    .X(_00979_));
 sg13g2_xnor2_1 _06264_ (.Y(_00980_),
    .A(_00930_),
    .B(_00978_));
 sg13g2_or2_1 _06265_ (.X(_00981_),
    .B(_00980_),
    .A(_00867_));
 sg13g2_o21ai_1 _06266_ (.B1(_00981_),
    .Y(_00982_),
    .A1(_00822_),
    .A2(_00979_));
 sg13g2_xnor2_1 _06267_ (.Y(_00983_),
    .A(_00927_),
    .B(_00822_));
 sg13g2_xnor2_1 _06268_ (.Y(_00984_),
    .A(_00978_),
    .B(_00867_));
 sg13g2_and3_1 _06269_ (.X(_00985_),
    .A(net193),
    .B(_00983_),
    .C(_00984_));
 sg13g2_nor3_1 _06270_ (.A(net193),
    .B(_00983_),
    .C(_00984_),
    .Y(_00986_));
 sg13g2_buf_1 _06271_ (.A(\i_tinyqv.cpu.pc[1] ),
    .X(_00987_));
 sg13g2_buf_1 _06272_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .X(_00988_));
 sg13g2_buf_1 _06273_ (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .X(_00989_));
 sg13g2_buf_1 _06274_ (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .X(_00990_));
 sg13g2_mux4_1 _06275_ (.S0(net228),
    .A0(_00987_),
    .A1(_00988_),
    .A2(net308),
    .A3(_00990_),
    .S1(_00766_),
    .X(_00991_));
 sg13g2_buf_1 _06276_ (.A(\i_tinyqv.cpu.instr_data_start[13] ),
    .X(_00992_));
 sg13g2_mux2_1 _06277_ (.A0(\i_tinyqv.cpu.instr_data_start[9] ),
    .A1(_00992_),
    .S(net226),
    .X(_00993_));
 sg13g2_a22oi_1 _06278_ (.Y(_00994_),
    .B1(_00993_),
    .B2(_00772_),
    .A2(_00991_),
    .A1(net211));
 sg13g2_nand2b_1 _06279_ (.Y(_00995_),
    .B(_00994_),
    .A_N(_00753_));
 sg13g2_nor2b_1 _06280_ (.A(net314),
    .B_N(net270),
    .Y(_00996_));
 sg13g2_nor2b_1 _06281_ (.A(net271),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .Y(_00997_));
 sg13g2_nor2b_1 _06282_ (.A(_00786_),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .Y(_00998_));
 sg13g2_nor2b_1 _06283_ (.A(_00787_),
    .B_N(net274),
    .Y(_00999_));
 sg13g2_a22oi_1 _06284_ (.Y(_01000_),
    .B1(_00998_),
    .B2(_00999_),
    .A2(_00997_),
    .A1(_00996_));
 sg13g2_and2_1 _06285_ (.A(net270),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .X(_01001_));
 sg13g2_and2_1 _06286_ (.A(_00787_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .X(_01002_));
 sg13g2_a22oi_1 _06287_ (.Y(_01003_),
    .B1(_01002_),
    .B2(_00837_),
    .A2(_01001_),
    .A1(_00835_));
 sg13g2_a21o_1 _06288_ (.A2(_01003_),
    .A1(_01000_),
    .B1(net225),
    .X(_01004_));
 sg13g2_inv_1 _06289_ (.Y(_01005_),
    .A(_00091_));
 sg13g2_mux4_1 _06290_ (.S0(_00840_),
    .A0(_01005_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .A2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A3(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .S1(_00794_),
    .X(_01006_));
 sg13g2_nand2_1 _06291_ (.Y(_01007_),
    .A(_00796_),
    .B(_01006_));
 sg13g2_mux2_1 _06292_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .S(_00780_),
    .X(_01008_));
 sg13g2_nand3_1 _06293_ (.B(_00809_),
    .C(_01008_),
    .A(_00799_),
    .Y(_01009_));
 sg13g2_nor2b_1 _06294_ (.A(net272),
    .B_N(net314),
    .Y(_01010_));
 sg13g2_mux2_1 _06295_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .S(_00777_),
    .X(_01011_));
 sg13g2_nand3_1 _06296_ (.B(_01010_),
    .C(_01011_),
    .A(net269),
    .Y(_01012_));
 sg13g2_nand4_1 _06297_ (.B(_00778_),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .A(net272),
    .Y(_01013_),
    .D(_00835_));
 sg13g2_and3_1 _06298_ (.X(_01014_),
    .A(_01009_),
    .B(_01012_),
    .C(_01013_));
 sg13g2_nand4_1 _06299_ (.B(_01004_),
    .C(_01007_),
    .A(_00753_),
    .Y(_01015_),
    .D(_01014_));
 sg13g2_nand3_1 _06300_ (.B(_00995_),
    .C(_01015_),
    .A(_00750_),
    .Y(_01016_));
 sg13g2_buf_2 _06301_ (.A(_01016_),
    .X(_01017_));
 sg13g2_nand2_1 _06302_ (.Y(_01018_),
    .A(_00878_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ));
 sg13g2_nand3b_1 _06303_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .C(_00872_),
    .Y(_01019_),
    .A_N(_00878_));
 sg13g2_o21ai_1 _06304_ (.B1(_01019_),
    .Y(_01020_),
    .A1(net268),
    .A2(_01018_));
 sg13g2_nand2_1 _06305_ (.Y(_01021_),
    .A(net267),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ));
 sg13g2_nand3b_1 _06306_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .C(net268),
    .Y(_01022_),
    .A_N(_00876_));
 sg13g2_o21ai_1 _06307_ (.B1(_01022_),
    .Y(_01023_),
    .A1(net268),
    .A2(_01021_));
 sg13g2_nor4_1 _06308_ (.A(net268),
    .B(net265),
    .C(_00899_),
    .D(_00833_),
    .Y(_01024_));
 sg13g2_a221oi_1 _06309_ (.B2(_00940_),
    .C1(_01024_),
    .B1(_01023_),
    .A1(_00901_),
    .Y(_01025_),
    .A2(_01020_));
 sg13g2_mux2_1 _06310_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .S(_00876_),
    .X(_01026_));
 sg13g2_nor2_1 _06311_ (.A(_00872_),
    .B(_00876_),
    .Y(_01027_));
 sg13g2_a22oi_1 _06312_ (.Y(_01028_),
    .B1(_01027_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .A2(_01026_),
    .A1(net268));
 sg13g2_or3_1 _06313_ (.A(_00884_),
    .B(_00910_),
    .C(_01028_),
    .X(_01029_));
 sg13g2_mux2_1 _06314_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .S(_00878_),
    .X(_01030_));
 sg13g2_a22oi_1 _06315_ (.Y(_01031_),
    .B1(_01030_),
    .B2(_00873_),
    .A2(_00905_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ));
 sg13g2_nand3b_1 _06316_ (.B(net223),
    .C(net222),
    .Y(_01032_),
    .A_N(_01031_));
 sg13g2_nand3b_1 _06317_ (.B(_00876_),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .Y(_01033_),
    .A_N(net265));
 sg13g2_nand3b_1 _06318_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .C(net265),
    .Y(_01034_),
    .A_N(_00876_));
 sg13g2_a21oi_1 _06319_ (.A1(_01033_),
    .A2(_01034_),
    .Y(_01035_),
    .B1(_00873_));
 sg13g2_and3_1 _06320_ (.X(_01036_),
    .A(net267),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .C(_00936_));
 sg13g2_o21ai_1 _06321_ (.B1(_00910_),
    .Y(_01037_),
    .A1(_01035_),
    .A2(_01036_));
 sg13g2_and4_1 _06322_ (.A(_01025_),
    .B(_01029_),
    .C(_01032_),
    .D(_01037_),
    .X(_01038_));
 sg13g2_buf_2 _06323_ (.A(_01038_),
    .X(_01039_));
 sg13g2_buf_1 _06324_ (.A(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .X(_01040_));
 sg13g2_buf_2 _06325_ (.A(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .X(_01041_));
 sg13g2_buf_1 _06326_ (.A(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .X(_01042_));
 sg13g2_buf_2 _06327_ (.A(\i_tinyqv.cpu.imm[12] ),
    .X(_01043_));
 sg13g2_mux4_1 _06328_ (.S0(net276),
    .A0(_01040_),
    .A1(_01041_),
    .A2(net306),
    .A3(_01043_),
    .S1(net277),
    .X(_01044_));
 sg13g2_buf_2 _06329_ (.A(\i_tinyqv.cpu.imm[16] ),
    .X(_01045_));
 sg13g2_buf_1 _06330_ (.A(\i_tinyqv.cpu.imm[20] ),
    .X(_01046_));
 sg13g2_mux4_1 _06331_ (.S0(_00761_),
    .A0(_01045_),
    .A1(_01046_),
    .A2(\i_tinyqv.cpu.imm[24] ),
    .A3(\i_tinyqv.cpu.imm[28] ),
    .S1(net277),
    .X(_01047_));
 sg13g2_and2_1 _06332_ (.A(net227),
    .B(_01047_),
    .X(_01048_));
 sg13g2_a21oi_1 _06333_ (.A1(_00892_),
    .A2(_01044_),
    .Y(_01049_),
    .B1(_01048_));
 sg13g2_mux2_1 _06334_ (.A0(_01039_),
    .A1(_01049_),
    .S(_00932_),
    .X(_01050_));
 sg13g2_buf_1 _06335_ (.A(_01050_),
    .X(_01051_));
 sg13g2_buf_1 _06336_ (.A(_01051_),
    .X(_01052_));
 sg13g2_buf_1 _06337_ (.A(_00084_),
    .X(_01053_));
 sg13g2_nor2_1 _06338_ (.A(net277),
    .B(_00761_),
    .Y(_01054_));
 sg13g2_buf_2 _06339_ (.A(_01054_),
    .X(_01055_));
 sg13g2_and2_1 _06340_ (.A(_01053_),
    .B(_01055_),
    .X(_01056_));
 sg13g2_buf_1 _06341_ (.A(_01056_),
    .X(_01057_));
 sg13g2_nand2_1 _06342_ (.Y(_01058_),
    .A(net193),
    .B(_01057_));
 sg13g2_nand2_1 _06343_ (.Y(_01059_),
    .A(_01053_),
    .B(_01055_));
 sg13g2_buf_1 _06344_ (.A(_01059_),
    .X(_01060_));
 sg13g2_nand2_1 _06345_ (.Y(_01061_),
    .A(_00092_),
    .B(net173));
 sg13g2_and2_1 _06346_ (.A(_01058_),
    .B(_01061_),
    .X(_01062_));
 sg13g2_buf_1 _06347_ (.A(_01062_),
    .X(_01063_));
 sg13g2_nand2_1 _06348_ (.Y(_01064_),
    .A(net125),
    .B(_01063_));
 sg13g2_nand3_1 _06349_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .C(_00880_),
    .A(_00889_),
    .Y(_01065_));
 sg13g2_nand3_1 _06350_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .C(_00888_),
    .A(net222),
    .Y(_01066_));
 sg13g2_a21oi_1 _06351_ (.A1(_01065_),
    .A2(_01066_),
    .Y(_01067_),
    .B1(_00875_));
 sg13g2_nor2b_1 _06352_ (.A(_00091_),
    .B_N(net266),
    .Y(_01068_));
 sg13g2_nor2b_1 _06353_ (.A(net221),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .Y(_01069_));
 sg13g2_a22oi_1 _06354_ (.Y(_01070_),
    .B1(_01069_),
    .B2(_00894_),
    .A2(_01068_),
    .A1(_00912_));
 sg13g2_nand3b_1 _06355_ (.B(net266),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .Y(_01071_),
    .A_N(net224));
 sg13g2_nand3b_1 _06356_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .C(net224),
    .Y(_01072_),
    .A_N(net266));
 sg13g2_nand2b_1 _06357_ (.Y(_01073_),
    .B(net222),
    .A_N(net267));
 sg13g2_a21o_1 _06358_ (.A2(_01072_),
    .A1(_01071_),
    .B1(_01073_),
    .X(_01074_));
 sg13g2_o21ai_1 _06359_ (.B1(_01074_),
    .Y(_01075_),
    .A1(_00902_),
    .A2(_01070_));
 sg13g2_and2_1 _06360_ (.A(net224),
    .B(_00877_),
    .X(_01076_));
 sg13g2_a221oi_1 _06361_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .C1(net222),
    .B1(_01076_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .Y(_01077_),
    .A2(_01027_));
 sg13g2_nor2b_1 _06362_ (.A(net224),
    .B_N(net267),
    .Y(_01078_));
 sg13g2_nor2b_1 _06363_ (.A(_00882_),
    .B_N(_00874_),
    .Y(_01079_));
 sg13g2_a221oi_1 _06364_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .C1(_00889_),
    .B1(_01079_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .Y(_01080_),
    .A2(_01078_));
 sg13g2_nor3_1 _06365_ (.A(_00910_),
    .B(_01077_),
    .C(_01080_),
    .Y(_01081_));
 sg13g2_nand3_1 _06366_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .C(_00936_),
    .A(net223),
    .Y(_01082_));
 sg13g2_nor2b_1 _06367_ (.A(net224),
    .B_N(net222),
    .Y(_01083_));
 sg13g2_mux2_1 _06368_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .S(net267),
    .X(_01084_));
 sg13g2_nand2_1 _06369_ (.Y(_01085_),
    .A(_01083_),
    .B(_01084_));
 sg13g2_a21oi_1 _06370_ (.A1(_01082_),
    .A2(_01085_),
    .Y(_01086_),
    .B1(_00887_));
 sg13g2_nor4_2 _06371_ (.A(_01067_),
    .B(_01075_),
    .C(_01081_),
    .Y(_01087_),
    .D(_01086_));
 sg13g2_buf_2 _06372_ (.A(\i_tinyqv.cpu.imm[13] ),
    .X(_01088_));
 sg13g2_mux4_1 _06373_ (.S0(net276),
    .A0(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .A1(_01088_),
    .A2(\i_tinyqv.cpu.imm[25] ),
    .A3(\i_tinyqv.cpu.imm[29] ),
    .S1(net275),
    .X(_01089_));
 sg13g2_buf_2 _06374_ (.A(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .X(_01090_));
 sg13g2_buf_2 _06375_ (.A(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .X(_01091_));
 sg13g2_buf_1 _06376_ (.A(\i_tinyqv.cpu.imm[17] ),
    .X(_01092_));
 sg13g2_buf_1 _06377_ (.A(\i_tinyqv.cpu.imm[21] ),
    .X(_01093_));
 sg13g2_mux4_1 _06378_ (.S0(net276),
    .A0(_01090_),
    .A1(_01091_),
    .A2(_01092_),
    .A3(_01093_),
    .S1(net275),
    .X(_01094_));
 sg13g2_mux2_1 _06379_ (.A0(_01089_),
    .A1(_01094_),
    .S(_00756_),
    .X(_01095_));
 sg13g2_buf_1 _06380_ (.A(_01095_),
    .X(_01096_));
 sg13g2_nor2_1 _06381_ (.A(_00871_),
    .B(_01096_),
    .Y(_01097_));
 sg13g2_a21oi_1 _06382_ (.A1(_00871_),
    .A2(_01087_),
    .Y(_01098_),
    .B1(_01097_));
 sg13g2_a21oi_1 _06383_ (.A1(_01017_),
    .A2(_01064_),
    .Y(_01099_),
    .B1(_01098_));
 sg13g2_nor2_1 _06384_ (.A(_01017_),
    .B(_01064_),
    .Y(_01100_));
 sg13g2_nor3_1 _06385_ (.A(net193),
    .B(_01099_),
    .C(_01100_),
    .Y(_01101_));
 sg13g2_nand2b_1 _06386_ (.Y(_01102_),
    .B(_01063_),
    .A_N(_01051_));
 sg13g2_a21o_1 _06387_ (.A2(_01087_),
    .A1(_00871_),
    .B1(_01097_),
    .X(_01103_));
 sg13g2_buf_2 _06388_ (.A(_01103_),
    .X(_01104_));
 sg13g2_a21oi_1 _06389_ (.A1(_01017_),
    .A2(_01102_),
    .Y(_01105_),
    .B1(_01104_));
 sg13g2_nor2_1 _06390_ (.A(_01017_),
    .B(_01102_),
    .Y(_01106_));
 sg13g2_nor3_1 _06391_ (.A(_00930_),
    .B(_01105_),
    .C(_01106_),
    .Y(_01107_));
 sg13g2_nor2b_1 _06392_ (.A(_00085_),
    .B_N(_00748_),
    .Y(_01108_));
 sg13g2_buf_1 _06393_ (.A(_01108_),
    .X(_01109_));
 sg13g2_nand3_1 _06394_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .C(_00796_),
    .A(_00794_),
    .Y(_01110_));
 sg13g2_nor2b_1 _06395_ (.A(net272),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .Y(_01111_));
 sg13g2_a21oi_1 _06396_ (.A1(_00835_),
    .A2(_01111_),
    .Y(_01112_),
    .B1(_00840_));
 sg13g2_nand3_1 _06397_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .C(_01010_),
    .A(net269),
    .Y(_01113_));
 sg13g2_nor2_1 _06398_ (.A(net274),
    .B(_00829_),
    .Y(_01114_));
 sg13g2_and2_1 _06399_ (.A(_00783_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .X(_01115_));
 sg13g2_a21oi_1 _06400_ (.A1(_01114_),
    .A2(_01115_),
    .Y(_01116_),
    .B1(net273));
 sg13g2_a22oi_1 _06401_ (.Y(_01117_),
    .B1(_01113_),
    .B2(_01116_),
    .A2(_01112_),
    .A1(_01110_));
 sg13g2_and2_1 _06402_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .B(_00828_),
    .X(_01118_));
 sg13g2_and3_1 _06403_ (.X(_01119_),
    .A(net272),
    .B(net271),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_a21o_1 _06404_ (.A2(_00784_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .B1(_01119_),
    .X(_01120_));
 sg13g2_nor3_1 _06405_ (.A(_00833_),
    .B(_00803_),
    .C(_00806_),
    .Y(_01121_));
 sg13g2_a221oi_1 _06406_ (.B2(_00996_),
    .C1(_01121_),
    .B1(_01120_),
    .A1(_00809_),
    .Y(_01122_),
    .A2(_01118_));
 sg13g2_nand2b_1 _06407_ (.Y(_01123_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .A_N(net314));
 sg13g2_nand3_1 _06408_ (.B(net274),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .A(net270),
    .Y(_01124_));
 sg13g2_o21ai_1 _06409_ (.B1(_01124_),
    .Y(_01125_),
    .A1(net273),
    .A2(_01123_));
 sg13g2_inv_1 _06410_ (.Y(_01126_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ));
 sg13g2_nand3_1 _06411_ (.B(net269),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .A(net273),
    .Y(_01127_));
 sg13g2_o21ai_1 _06412_ (.B1(_01127_),
    .Y(_01128_),
    .A1(_01126_),
    .A2(_00814_));
 sg13g2_nand3b_1 _06413_ (.B(net273),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .Y(_01129_),
    .A_N(net272));
 sg13g2_nand3b_1 _06414_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .C(net272),
    .Y(_01130_),
    .A_N(net270));
 sg13g2_nand2b_1 _06415_ (.Y(_01131_),
    .B(net274),
    .A_N(net269));
 sg13g2_a21oi_1 _06416_ (.A1(_01129_),
    .A2(_01130_),
    .Y(_01132_),
    .B1(_01131_));
 sg13g2_a221oi_1 _06417_ (.B2(_01010_),
    .C1(_01132_),
    .B1(_01128_),
    .A1(_00782_),
    .Y(_01133_),
    .A2(_01125_));
 sg13g2_nand3b_1 _06418_ (.B(_01122_),
    .C(_01133_),
    .Y(_01134_),
    .A_N(_01117_));
 sg13g2_buf_2 _06419_ (.A(_01134_),
    .X(_01135_));
 sg13g2_buf_8 _06420_ (.A(_01135_),
    .X(_01136_));
 sg13g2_buf_1 _06421_ (.A(\i_tinyqv.cpu.instr_data_start[16] ),
    .X(_01137_));
 sg13g2_buf_2 _06422_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .X(_01138_));
 sg13g2_mux2_1 _06423_ (.A0(net305),
    .A1(_01138_),
    .S(_00763_),
    .X(_01139_));
 sg13g2_nand2_1 _06424_ (.Y(_01140_),
    .A(_00756_),
    .B(_01139_));
 sg13g2_buf_2 _06425_ (.A(net277),
    .X(_01141_));
 sg13g2_buf_1 _06426_ (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .X(_01142_));
 sg13g2_mux2_1 _06427_ (.A0(net304),
    .A1(\i_tinyqv.cpu.instr_data_start[12] ),
    .S(_00763_),
    .X(_01143_));
 sg13g2_nor2b_1 _06428_ (.A(_00755_),
    .B_N(_00762_),
    .Y(_01144_));
 sg13g2_buf_1 _06429_ (.A(_01144_),
    .X(_01145_));
 sg13g2_buf_1 _06430_ (.A(\i_tinyqv.cpu.instr_data_start[4] ),
    .X(_01146_));
 sg13g2_a22oi_1 _06431_ (.Y(_01147_),
    .B1(_01145_),
    .B2(net303),
    .A2(_01143_),
    .A1(net220));
 sg13g2_mux2_1 _06432_ (.A0(_01140_),
    .A1(_01147_),
    .S(_00892_),
    .X(_01148_));
 sg13g2_nor2_1 _06433_ (.A(_00753_),
    .B(_01148_),
    .Y(_01149_));
 sg13g2_a21oi_1 _06434_ (.A1(_00753_),
    .A2(net153),
    .Y(_01150_),
    .B1(_01149_));
 sg13g2_nor2_1 _06435_ (.A(_01109_),
    .B(_01150_),
    .Y(_01151_));
 sg13g2_buf_2 _06436_ (.A(_01151_),
    .X(_01152_));
 sg13g2_nor2_1 _06437_ (.A(_00930_),
    .B(_01063_),
    .Y(_01153_));
 sg13g2_nor3_1 _06438_ (.A(net193),
    .B(net125),
    .C(_01063_),
    .Y(_01154_));
 sg13g2_a21oi_1 _06439_ (.A1(net125),
    .A2(_01153_),
    .Y(_01155_),
    .B1(_01154_));
 sg13g2_and2_1 _06440_ (.A(_01104_),
    .B(_01017_),
    .X(_01156_));
 sg13g2_nand2_1 _06441_ (.Y(_01157_),
    .A(_00827_),
    .B(_01156_));
 sg13g2_nand3_1 _06442_ (.B(_01098_),
    .C(_01017_),
    .A(_00930_),
    .Y(_01158_));
 sg13g2_nand4_1 _06443_ (.B(_01155_),
    .C(_01157_),
    .A(_01152_),
    .Y(_01159_),
    .D(_01158_));
 sg13g2_o21ai_1 _06444_ (.B1(_01159_),
    .Y(_01160_),
    .A1(_01101_),
    .A2(_01107_));
 sg13g2_buf_1 _06445_ (.A(_01160_),
    .X(_01161_));
 sg13g2_o21ai_1 _06446_ (.B1(_01161_),
    .Y(_01162_),
    .A1(_00985_),
    .A2(_00986_));
 sg13g2_nand2b_1 _06447_ (.Y(\i_tinyqv.cpu.i_core.cy_out ),
    .B(_01162_),
    .A_N(_00982_));
 sg13g2_buf_1 _06448_ (.A(_01053_),
    .X(_01163_));
 sg13g2_nor2_1 _06449_ (.A(net264),
    .B(_00961_),
    .Y(_01164_));
 sg13g2_buf_1 _06450_ (.A(_01164_),
    .X(_01165_));
 sg13g2_buf_1 _06451_ (.A(net172),
    .X(_01166_));
 sg13g2_buf_1 _06452_ (.A(_00750_),
    .X(_01167_));
 sg13g2_or2_1 _06453_ (.X(_01168_),
    .B(\i_tinyqv.cpu.is_alu_imm ),
    .A(\i_tinyqv.cpu.is_alu_reg ));
 sg13g2_buf_1 _06454_ (.A(_01168_),
    .X(_01169_));
 sg13g2_buf_1 _06455_ (.A(\i_tinyqv.cpu.is_load ),
    .X(_01170_));
 sg13g2_nand2b_1 _06456_ (.Y(_01171_),
    .B(_01170_),
    .A_N(_00083_));
 sg13g2_nor2_1 _06457_ (.A(_01169_),
    .B(_01171_),
    .Y(_01172_));
 sg13g2_buf_2 _06458_ (.A(_00086_),
    .X(_01173_));
 sg13g2_buf_1 _06459_ (.A(_01173_),
    .X(_01174_));
 sg13g2_nor2b_1 _06460_ (.A(net315),
    .B_N(_00745_),
    .Y(_01175_));
 sg13g2_buf_1 _06461_ (.A(_01175_),
    .X(_01176_));
 sg13g2_buf_2 _06462_ (.A(\i_tinyqv.cpu.alu_op[0] ),
    .X(_01177_));
 sg13g2_nand2b_1 _06463_ (.Y(_01178_),
    .B(_01177_),
    .A_N(_00745_));
 sg13g2_buf_2 _06464_ (.A(_01178_),
    .X(_01179_));
 sg13g2_nor2b_1 _06465_ (.A(_01176_),
    .B_N(_01179_),
    .Y(_01180_));
 sg13g2_xnor2_1 _06466_ (.Y(_01181_),
    .A(net263),
    .B(_01180_));
 sg13g2_a22oi_1 _06467_ (.Y(_01182_),
    .B1(_01181_),
    .B2(_01169_),
    .A2(_01172_),
    .A1(\i_tinyqv.cpu.i_core.load_done ));
 sg13g2_buf_1 _06468_ (.A(_00751_),
    .X(_01183_));
 sg13g2_nor2b_1 _06469_ (.A(_01182_),
    .B_N(net262),
    .Y(_01184_));
 sg13g2_buf_1 _06470_ (.A(_00093_),
    .X(_01185_));
 sg13g2_buf_2 _06471_ (.A(_00094_),
    .X(_01186_));
 sg13g2_and2_1 _06472_ (.A(net262),
    .B(\i_tinyqv.cpu.is_system ),
    .X(_01187_));
 sg13g2_nor2_1 _06473_ (.A(_00745_),
    .B(_01177_),
    .Y(_01188_));
 sg13g2_and2_1 _06474_ (.A(_01187_),
    .B(_01188_),
    .X(_01189_));
 sg13g2_buf_1 _06475_ (.A(_01189_),
    .X(_01190_));
 sg13g2_buf_1 _06476_ (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .X(_01191_));
 sg13g2_nor2_1 _06477_ (.A(_01191_),
    .B(net306),
    .Y(_01192_));
 sg13g2_nand3_1 _06478_ (.B(_01190_),
    .C(_01192_),
    .A(_01186_),
    .Y(_01193_));
 sg13g2_buf_1 _06479_ (.A(_01193_),
    .X(_01194_));
 sg13g2_nand2_1 _06480_ (.Y(_01195_),
    .A(_01185_),
    .B(_01194_));
 sg13g2_buf_2 _06481_ (.A(\i_tinyqv.cpu.is_store ),
    .X(_01196_));
 sg13g2_and2_1 _06482_ (.A(_01196_),
    .B(\i_tinyqv.cpu.no_write_in_progress ),
    .X(_01197_));
 sg13g2_buf_2 _06483_ (.A(_01197_),
    .X(_01198_));
 sg13g2_and2_1 _06484_ (.A(net262),
    .B(_00868_),
    .X(_01199_));
 sg13g2_buf_1 _06485_ (.A(_01199_),
    .X(_01200_));
 sg13g2_nor4_1 _06486_ (.A(\i_tinyqv.cpu.is_auipc ),
    .B(\i_tinyqv.cpu.is_system ),
    .C(_01198_),
    .D(_01200_),
    .Y(_01201_));
 sg13g2_o21ai_1 _06487_ (.B1(_00083_),
    .Y(_01202_),
    .A1(_01170_),
    .A2(_01196_));
 sg13g2_and2_1 _06488_ (.A(_01183_),
    .B(_01202_),
    .X(_01203_));
 sg13g2_buf_1 _06489_ (.A(_01203_),
    .X(_01204_));
 sg13g2_or2_1 _06490_ (.X(_01205_),
    .B(\i_tinyqv.cpu.is_jalr ),
    .A(\i_tinyqv.cpu.is_jal ));
 sg13g2_buf_1 _06491_ (.A(_01205_),
    .X(_01206_));
 sg13g2_o21ai_1 _06492_ (.B1(net262),
    .Y(_01207_),
    .A1(\i_tinyqv.cpu.is_lui ),
    .A2(_01206_));
 sg13g2_nand3_1 _06493_ (.B(_01204_),
    .C(_01207_),
    .A(_01201_),
    .Y(_01208_));
 sg13g2_nor3_1 _06494_ (.A(_01184_),
    .B(_01195_),
    .C(_01208_),
    .Y(_01209_));
 sg13g2_nand2_1 _06495_ (.Y(_01210_),
    .A(net171),
    .B(_01209_));
 sg13g2_xnor2_1 _06496_ (.Y(_01211_),
    .A(_01152_),
    .B(net125));
 sg13g2_inv_1 _06497_ (.Y(_01212_),
    .A(\i_tinyqv.cpu.i_core.cmp ));
 sg13g2_nor2_1 _06498_ (.A(_00824_),
    .B(_01109_),
    .Y(_01213_));
 sg13g2_a21oi_1 _06499_ (.A1(_01212_),
    .A2(net173),
    .Y(_01214_),
    .B1(_01213_));
 sg13g2_xnor2_1 _06500_ (.Y(_01215_),
    .A(_01104_),
    .B(_01017_));
 sg13g2_nand2_1 _06501_ (.Y(_01216_),
    .A(_01214_),
    .B(_01215_));
 sg13g2_nor4_2 _06502_ (.A(_00983_),
    .B(_00984_),
    .C(_01211_),
    .Y(_01217_),
    .D(_01216_));
 sg13g2_xnor2_1 _06503_ (.Y(_01218_),
    .A(_01177_),
    .B(_01217_));
 sg13g2_inv_1 _06504_ (.Y(_01219_),
    .A(_01173_));
 sg13g2_buf_1 _06505_ (.A(_01219_),
    .X(_01220_));
 sg13g2_buf_1 _06506_ (.A(_01195_),
    .X(_01221_));
 sg13g2_nor4_2 _06507_ (.A(net219),
    .B(net171),
    .C(net137),
    .Y(_01222_),
    .D(_01208_));
 sg13g2_nand2_1 _06508_ (.Y(_01223_),
    .A(_01218_),
    .B(_01222_));
 sg13g2_nand3_1 _06509_ (.B(_01210_),
    .C(_01223_),
    .A(net160),
    .Y(_01224_));
 sg13g2_nor2b_1 _06510_ (.A(_01204_),
    .B_N(_01185_),
    .Y(_01225_));
 sg13g2_nor2_1 _06511_ (.A(_01224_),
    .B(_01225_),
    .Y(_00029_));
 sg13g2_or3_1 _06512_ (.A(\addr[26] ),
    .B(\addr[25] ),
    .C(\addr[27] ),
    .X(_01226_));
 sg13g2_buf_2 _06513_ (.A(_01226_),
    .X(_01227_));
 sg13g2_a21oi_1 _06514_ (.A1(\i_tinyqv.cpu.data_write_n[1] ),
    .A2(\i_tinyqv.cpu.data_read_n[1] ),
    .Y(_01228_),
    .B1(_01227_));
 sg13g2_buf_1 _06515_ (.A(_01228_),
    .X(_01229_));
 sg13g2_buf_1 _06516_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .X(_01230_));
 sg13g2_buf_1 _06517_ (.A(_00157_),
    .X(_01231_));
 sg13g2_buf_1 _06518_ (.A(\i_tinyqv.cpu.data_write_n[0] ),
    .X(_01232_));
 sg13g2_buf_1 _06519_ (.A(\i_tinyqv.cpu.data_read_n[0] ),
    .X(_01233_));
 sg13g2_and2_1 _06520_ (.A(_01232_),
    .B(_01233_),
    .X(_01234_));
 sg13g2_buf_2 _06521_ (.A(_01234_),
    .X(_01235_));
 sg13g2_xnor2_1 _06522_ (.Y(_01236_),
    .A(_01231_),
    .B(_01235_));
 sg13g2_nor2_1 _06523_ (.A(_01230_),
    .B(_01236_),
    .Y(_01237_));
 sg13g2_nor2_1 _06524_ (.A(_01231_),
    .B(net210),
    .Y(_01238_));
 sg13g2_a22oi_1 _06525_ (.Y(_01239_),
    .B1(_01238_),
    .B2(_01230_),
    .A2(_01237_),
    .A1(_01229_));
 sg13g2_buf_1 _06526_ (.A(\i_tinyqv.mem.q_ctrl.data_req ),
    .X(_01240_));
 sg13g2_nor2b_1 _06527_ (.A(_01239_),
    .B_N(_01240_),
    .Y(_00082_));
 sg13g2_mux2_1 _06528_ (.A0(\i_uart_tx.txd_reg ),
    .A1(\gpio_out[0] ),
    .S(\gpio_out_sel[0] ),
    .X(net28));
 sg13g2_buf_1 _06529_ (.A(debug_register_data),
    .X(_01241_));
 sg13g2_nor2b_1 _06530_ (.A(net301),
    .B_N(\i_spi.spi_select ),
    .Y(_01242_));
 sg13g2_a21oi_1 _06531_ (.A1(\debug_rd_r[2] ),
    .A2(net301),
    .Y(_01243_),
    .B1(_01242_));
 sg13g2_nand2_1 _06532_ (.Y(_01244_),
    .A(\gpio_out_sel[4] ),
    .B(\gpio_out[4] ));
 sg13g2_o21ai_1 _06533_ (.B1(_01244_),
    .Y(net32),
    .A1(\gpio_out_sel[4] ),
    .A2(_01243_));
 sg13g2_mux2_1 _06534_ (.A0(\i_uart_rx.uart_rts ),
    .A1(\gpio_out[1] ),
    .S(\gpio_out_sel[1] ),
    .X(net29));
 sg13g2_buf_1 _06535_ (.A(\i_spi.spi_clk_out ),
    .X(_01245_));
 sg13g2_inv_1 _06536_ (.Y(_01246_),
    .A(_01245_));
 sg13g2_nor2_1 _06537_ (.A(_01246_),
    .B(net301),
    .Y(_01247_));
 sg13g2_a21oi_1 _06538_ (.A1(net301),
    .A2(\debug_rd_r[3] ),
    .Y(_01248_),
    .B1(_01247_));
 sg13g2_nand2_1 _06539_ (.Y(_01249_),
    .A(\gpio_out_sel[5] ),
    .B(\gpio_out[5] ));
 sg13g2_o21ai_1 _06540_ (.B1(_01249_),
    .Y(net33),
    .A1(\gpio_out_sel[5] ),
    .A2(_01248_));
 sg13g2_nor2b_1 _06541_ (.A(net301),
    .B_N(\i_spi.spi_dc ),
    .Y(_01250_));
 sg13g2_a21oi_1 _06542_ (.A1(net301),
    .A2(\debug_rd_r[0] ),
    .Y(_01251_),
    .B1(_01250_));
 sg13g2_nand2_1 _06543_ (.Y(_01252_),
    .A(\gpio_out_sel[2] ),
    .B(\gpio_out[2] ));
 sg13g2_o21ai_1 _06544_ (.B1(_01252_),
    .Y(net30),
    .A1(\gpio_out_sel[2] ),
    .A2(_01251_));
 sg13g2_mux2_1 _06545_ (.A0(debug_uart_txd),
    .A1(\gpio_out[6] ),
    .S(\gpio_out_sel[6] ),
    .X(net34));
 sg13g2_nor2b_1 _06546_ (.A(net301),
    .B_N(\i_spi.data[7] ),
    .Y(_01253_));
 sg13g2_a21oi_1 _06547_ (.A1(net301),
    .A2(\debug_rd_r[1] ),
    .Y(_01254_),
    .B1(_01253_));
 sg13g2_nand2_1 _06548_ (.Y(_01255_),
    .A(\gpio_out_sel[3] ),
    .B(\gpio_out[3] ));
 sg13g2_o21ai_1 _06549_ (.B1(_01255_),
    .Y(net31),
    .A1(\gpio_out_sel[3] ),
    .A2(_01254_));
 sg13g2_buf_1 _06550_ (.A(\gpio_out_sel[7] ),
    .X(_01256_));
 sg13g2_buf_1 _06551_ (.A(net5),
    .X(_01257_));
 sg13g2_buf_2 _06552_ (.A(ui_in[5]),
    .X(_01258_));
 sg13g2_and2_1 _06553_ (.A(net317),
    .B(_01258_),
    .X(_01259_));
 sg13g2_buf_1 _06554_ (.A(ui_in[3]),
    .X(_01260_));
 sg13g2_nand2_1 _06555_ (.Y(_01261_),
    .A(net262),
    .B(_00868_));
 sg13g2_buf_2 _06556_ (.A(_01261_),
    .X(_01262_));
 sg13g2_buf_2 _06557_ (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .X(_01263_));
 sg13g2_xnor2_1 _06558_ (.Y(_01264_),
    .A(_00867_),
    .B(_00980_));
 sg13g2_nand2_1 _06559_ (.Y(_01265_),
    .A(_01177_),
    .B(_00750_));
 sg13g2_o21ai_1 _06560_ (.B1(_01265_),
    .Y(_01266_),
    .A1(_01217_),
    .A2(_01264_));
 sg13g2_xor2_1 _06561_ (.B(net125),
    .A(_01152_),
    .X(_01267_));
 sg13g2_nand4_1 _06562_ (.B(_01214_),
    .C(_01215_),
    .A(_01267_),
    .Y(_01268_),
    .D(_01265_));
 sg13g2_a21o_1 _06563_ (.A2(_01268_),
    .A1(_00986_),
    .B1(_00985_),
    .X(_01269_));
 sg13g2_nand2_1 _06564_ (.Y(_01270_),
    .A(_00867_),
    .B(_00980_));
 sg13g2_a221oi_1 _06565_ (.B2(_01270_),
    .C1(_01217_),
    .B1(_01213_),
    .A1(_01177_),
    .Y(_01271_),
    .A2(net171));
 sg13g2_a221oi_1 _06566_ (.B2(_01161_),
    .C1(_01271_),
    .B1(_01269_),
    .A1(_00982_),
    .Y(\i_tinyqv.cpu.i_core.cmp_out ),
    .A2(_01266_));
 sg13g2_xnor2_1 _06567_ (.Y(_01272_),
    .A(_01263_),
    .B(\i_tinyqv.cpu.i_core.cmp_out ));
 sg13g2_and2_1 _06568_ (.A(net262),
    .B(_01206_),
    .X(_01273_));
 sg13g2_buf_1 _06569_ (.A(_01273_),
    .X(_01274_));
 sg13g2_and4_1 _06570_ (.A(net302),
    .B(net306),
    .C(_01186_),
    .D(_01190_),
    .X(_01275_));
 sg13g2_buf_1 _06571_ (.A(_01275_),
    .X(_01276_));
 sg13g2_nor3_1 _06572_ (.A(net137),
    .B(_01274_),
    .C(_01276_),
    .Y(_01277_));
 sg13g2_o21ai_1 _06573_ (.B1(_01277_),
    .Y(_01278_),
    .A1(_01262_),
    .A2(_01272_));
 sg13g2_buf_2 _06574_ (.A(_01278_),
    .X(_01279_));
 sg13g2_and2_1 _06575_ (.A(net172),
    .B(_01279_),
    .X(_01280_));
 sg13g2_buf_1 _06576_ (.A(_01280_),
    .X(_01281_));
 sg13g2_buf_2 _06577_ (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .X(_01282_));
 sg13g2_buf_1 _06578_ (.A(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .X(_01283_));
 sg13g2_buf_1 _06579_ (.A(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .X(_01284_));
 sg13g2_nor3_1 _06580_ (.A(_01283_),
    .B(_01284_),
    .C(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .Y(_01285_));
 sg13g2_buf_2 _06581_ (.A(_01285_),
    .X(_01286_));
 sg13g2_nand3_1 _06582_ (.B(_01210_),
    .C(_01286_),
    .A(_01202_),
    .Y(_01287_));
 sg13g2_buf_1 _06583_ (.A(net262),
    .X(_01288_));
 sg13g2_a22oi_1 _06584_ (.Y(_01289_),
    .B1(_01287_),
    .B2(net218),
    .A2(_01222_),
    .A1(_01218_));
 sg13g2_buf_2 _06585_ (.A(\i_tinyqv.cpu.instr_len[1] ),
    .X(_01290_));
 sg13g2_xnor2_1 _06586_ (.Y(_01291_),
    .A(_01290_),
    .B(net309));
 sg13g2_buf_1 _06587_ (.A(_00100_),
    .X(_01292_));
 sg13g2_nor2b_1 _06588_ (.A(_00751_),
    .B_N(_01292_),
    .Y(_01293_));
 sg13g2_a21o_1 _06589_ (.A2(_01291_),
    .A1(_00751_),
    .B1(_01293_),
    .X(_01294_));
 sg13g2_buf_1 _06590_ (.A(_01294_),
    .X(_01295_));
 sg13g2_buf_1 _06591_ (.A(_01295_),
    .X(_01296_));
 sg13g2_buf_1 _06592_ (.A(net192),
    .X(_01297_));
 sg13g2_nand2_2 _06593_ (.Y(_01298_),
    .A(_01290_),
    .B(net309));
 sg13g2_xor2_1 _06594_ (.B(_00758_),
    .A(\i_tinyqv.cpu.instr_len[2] ),
    .X(_01299_));
 sg13g2_xnor2_1 _06595_ (.Y(_01300_),
    .A(_01298_),
    .B(_01299_));
 sg13g2_nor2_1 _06596_ (.A(_00751_),
    .B(_00101_),
    .Y(_01301_));
 sg13g2_a21oi_2 _06597_ (.B1(_01301_),
    .Y(_01302_),
    .A2(_01300_),
    .A1(_00751_));
 sg13g2_buf_8 _06598_ (.A(_01302_),
    .X(_01303_));
 sg13g2_buf_8 _06599_ (.A(net191),
    .X(_01304_));
 sg13g2_mux2_1 _06600_ (.A0(\i_tinyqv.cpu.instr_data[3][0] ),
    .A1(\i_tinyqv.cpu.instr_data[1][0] ),
    .S(net169),
    .X(_01305_));
 sg13g2_nor2_1 _06601_ (.A(net170),
    .B(_01305_),
    .Y(_01306_));
 sg13g2_mux2_1 _06602_ (.A0(\i_tinyqv.cpu.instr_data[2][0] ),
    .A1(\i_tinyqv.cpu.instr_data[0][0] ),
    .S(net169),
    .X(_01307_));
 sg13g2_nand2b_1 _06603_ (.Y(_01308_),
    .B(_01297_),
    .A_N(_01307_));
 sg13g2_nor2b_1 _06604_ (.A(_01306_),
    .B_N(_01308_),
    .Y(_01309_));
 sg13g2_buf_1 _06605_ (.A(_01309_),
    .X(_01310_));
 sg13g2_mux2_1 _06606_ (.A0(_00121_),
    .A1(_00118_),
    .S(net191),
    .X(_01311_));
 sg13g2_nor2_1 _06607_ (.A(net170),
    .B(_01311_),
    .Y(_01312_));
 sg13g2_mux2_1 _06608_ (.A0(_00120_),
    .A1(_00119_),
    .S(net169),
    .X(_01313_));
 sg13g2_nand2b_1 _06609_ (.Y(_01314_),
    .B(net170),
    .A_N(_01313_));
 sg13g2_nor2b_1 _06610_ (.A(_01312_),
    .B_N(_01314_),
    .Y(_01315_));
 sg13g2_buf_1 _06611_ (.A(_01315_),
    .X(_01316_));
 sg13g2_mux2_1 _06612_ (.A0(_00125_),
    .A1(_00122_),
    .S(net191),
    .X(_01317_));
 sg13g2_nor2_1 _06613_ (.A(_01296_),
    .B(_01317_),
    .Y(_01318_));
 sg13g2_mux2_1 _06614_ (.A0(_00124_),
    .A1(_00123_),
    .S(net191),
    .X(_01319_));
 sg13g2_nand2b_1 _06615_ (.Y(_01320_),
    .B(net192),
    .A_N(_01319_));
 sg13g2_nand2b_1 _06616_ (.Y(_01321_),
    .B(_01320_),
    .A_N(_01318_));
 sg13g2_buf_2 _06617_ (.A(_01321_),
    .X(_01322_));
 sg13g2_nor2_1 _06618_ (.A(_01316_),
    .B(_01322_),
    .Y(_01323_));
 sg13g2_buf_1 _06619_ (.A(_01323_),
    .X(_01324_));
 sg13g2_mux2_1 _06620_ (.A0(\i_tinyqv.cpu.instr_data[3][2] ),
    .A1(\i_tinyqv.cpu.instr_data[1][2] ),
    .S(_01302_),
    .X(_01325_));
 sg13g2_mux2_1 _06621_ (.A0(\i_tinyqv.cpu.instr_data[2][2] ),
    .A1(\i_tinyqv.cpu.instr_data[0][2] ),
    .S(net191),
    .X(_01326_));
 sg13g2_mux2_1 _06622_ (.A0(_01325_),
    .A1(_01326_),
    .S(net192),
    .X(_01327_));
 sg13g2_buf_1 _06623_ (.A(_01327_),
    .X(_01328_));
 sg13g2_mux2_1 _06624_ (.A0(\i_tinyqv.cpu.instr_data[3][3] ),
    .A1(\i_tinyqv.cpu.instr_data[1][3] ),
    .S(_01302_),
    .X(_01329_));
 sg13g2_mux2_1 _06625_ (.A0(\i_tinyqv.cpu.instr_data[2][3] ),
    .A1(\i_tinyqv.cpu.instr_data[0][3] ),
    .S(net191),
    .X(_01330_));
 sg13g2_mux2_1 _06626_ (.A0(_01329_),
    .A1(_01330_),
    .S(_01295_),
    .X(_01331_));
 sg13g2_buf_2 _06627_ (.A(_01331_),
    .X(_01332_));
 sg13g2_a21oi_1 _06628_ (.A1(_01183_),
    .A2(_01291_),
    .Y(_01333_),
    .B1(_01293_));
 sg13g2_buf_2 _06629_ (.A(_01333_),
    .X(_01334_));
 sg13g2_mux2_1 _06630_ (.A0(_00109_),
    .A1(_00106_),
    .S(net169),
    .X(_01335_));
 sg13g2_mux2_1 _06631_ (.A0(_00108_),
    .A1(_00107_),
    .S(_01304_),
    .X(_01336_));
 sg13g2_and2_1 _06632_ (.A(net170),
    .B(_01336_),
    .X(_01337_));
 sg13g2_a21oi_1 _06633_ (.A1(_01334_),
    .A2(_01335_),
    .Y(_01338_),
    .B1(_01337_));
 sg13g2_buf_1 _06634_ (.A(_01338_),
    .X(_01339_));
 sg13g2_mux2_1 _06635_ (.A0(_00113_),
    .A1(_00110_),
    .S(net191),
    .X(_01340_));
 sg13g2_nor2_1 _06636_ (.A(net192),
    .B(_01340_),
    .Y(_01341_));
 sg13g2_mux2_1 _06637_ (.A0(_00112_),
    .A1(_00111_),
    .S(_01303_),
    .X(_01342_));
 sg13g2_nand2b_1 _06638_ (.Y(_01343_),
    .B(net192),
    .A_N(_01342_));
 sg13g2_nand2b_1 _06639_ (.Y(_01344_),
    .B(_01343_),
    .A_N(_01341_));
 sg13g2_buf_2 _06640_ (.A(_01344_),
    .X(_01345_));
 sg13g2_mux2_1 _06641_ (.A0(_00117_),
    .A1(_00114_),
    .S(net191),
    .X(_01346_));
 sg13g2_nor2_1 _06642_ (.A(net192),
    .B(_01346_),
    .Y(_01347_));
 sg13g2_mux2_1 _06643_ (.A0(_00116_),
    .A1(_00115_),
    .S(_01303_),
    .X(_01348_));
 sg13g2_nand2b_1 _06644_ (.Y(_01349_),
    .B(net192),
    .A_N(_01348_));
 sg13g2_nand2b_1 _06645_ (.Y(_01350_),
    .B(_01349_),
    .A_N(_01347_));
 sg13g2_buf_2 _06646_ (.A(_01350_),
    .X(_01351_));
 sg13g2_nand2_2 _06647_ (.Y(_01352_),
    .A(_01345_),
    .B(_01351_));
 sg13g2_nor2_1 _06648_ (.A(net123),
    .B(_01352_),
    .Y(_01353_));
 sg13g2_and3_1 _06649_ (.X(_01354_),
    .A(_01328_),
    .B(_01332_),
    .C(_01353_));
 sg13g2_buf_2 _06650_ (.A(_01354_),
    .X(_01355_));
 sg13g2_mux2_1 _06651_ (.A0(_00105_),
    .A1(_00104_),
    .S(net192),
    .X(_01356_));
 sg13g2_nor2_1 _06652_ (.A(net169),
    .B(_01356_),
    .Y(_01357_));
 sg13g2_nand2_1 _06653_ (.Y(_01358_),
    .A(_00103_),
    .B(_01296_));
 sg13g2_nand2_1 _06654_ (.Y(_01359_),
    .A(_00102_),
    .B(_01334_));
 sg13g2_nand3_1 _06655_ (.B(_01358_),
    .C(_01359_),
    .A(net169),
    .Y(_01360_));
 sg13g2_nand2b_1 _06656_ (.Y(_01361_),
    .B(_01360_),
    .A_N(_01357_));
 sg13g2_buf_2 _06657_ (.A(_01361_),
    .X(_01362_));
 sg13g2_mux2_1 _06658_ (.A0(_01324_),
    .A1(_01355_),
    .S(_01362_),
    .X(_01363_));
 sg13g2_and2_1 _06659_ (.A(net124),
    .B(_01363_),
    .X(_01364_));
 sg13g2_nand4_1 _06660_ (.B(net172),
    .C(_01289_),
    .A(_01282_),
    .Y(_01365_),
    .D(_01364_));
 sg13g2_or2_1 _06661_ (.X(_01366_),
    .B(_00961_),
    .A(net264));
 sg13g2_buf_1 _06662_ (.A(_01366_),
    .X(_01367_));
 sg13g2_a221oi_1 _06663_ (.B2(_01222_),
    .C1(net168),
    .B1(_01218_),
    .A1(net171),
    .Y(_01368_),
    .A2(_01209_));
 sg13g2_buf_1 _06664_ (.A(_01368_),
    .X(_01369_));
 sg13g2_buf_1 _06665_ (.A(\i_tinyqv.cpu.i_core.mip[17] ),
    .X(_01370_));
 sg13g2_nand2_1 _06666_ (.Y(_01371_),
    .A(\i_tinyqv.cpu.i_core.mie[17] ),
    .B(_01370_));
 sg13g2_nand2_1 _06667_ (.Y(_01372_),
    .A(\i_tinyqv.cpu.i_core.mie[16] ),
    .B(\i_tinyqv.cpu.i_core.mip[16] ));
 sg13g2_nand2_1 _06668_ (.Y(_01373_),
    .A(_01371_),
    .B(_01372_));
 sg13g2_buf_1 _06669_ (.A(\i_tinyqv.cpu.i_core.mie[18] ),
    .X(_01374_));
 sg13g2_buf_1 _06670_ (.A(\i_uart_rx.fsm_state[0] ),
    .X(_01375_));
 sg13g2_buf_1 _06671_ (.A(\i_uart_rx.fsm_state[2] ),
    .X(_01376_));
 sg13g2_buf_2 _06672_ (.A(\i_uart_rx.fsm_state[1] ),
    .X(_01377_));
 sg13g2_nand2_1 _06673_ (.Y(_01378_),
    .A(_01377_),
    .B(\i_uart_rx.fsm_state[3] ));
 sg13g2_nor2_1 _06674_ (.A(net299),
    .B(_01378_),
    .Y(_01379_));
 sg13g2_and2_1 _06675_ (.A(net300),
    .B(_01379_),
    .X(_01380_));
 sg13g2_buf_1 _06676_ (.A(_01380_),
    .X(_01381_));
 sg13g2_buf_2 _06677_ (.A(\i_uart_tx.fsm_state[1] ),
    .X(_01382_));
 sg13g2_buf_1 _06678_ (.A(\i_uart_tx.fsm_state[2] ),
    .X(_01383_));
 sg13g2_nor2_1 _06679_ (.A(_01382_),
    .B(_01383_),
    .Y(_01384_));
 sg13g2_buf_2 _06680_ (.A(\i_uart_tx.fsm_state[0] ),
    .X(_01385_));
 sg13g2_buf_2 _06681_ (.A(\i_uart_tx.fsm_state[3] ),
    .X(_01386_));
 sg13g2_nor2_1 _06682_ (.A(_01385_),
    .B(_01386_),
    .Y(_01387_));
 sg13g2_and2_1 _06683_ (.A(_01384_),
    .B(_01387_),
    .X(_01388_));
 sg13g2_buf_1 _06684_ (.A(_01388_),
    .X(_01389_));
 sg13g2_buf_1 _06685_ (.A(\i_tinyqv.cpu.i_core.mie[19] ),
    .X(_01390_));
 sg13g2_a22oi_1 _06686_ (.Y(_01391_),
    .B1(net209),
    .B2(_01390_),
    .A2(_01381_),
    .A1(_01374_));
 sg13g2_inv_1 _06687_ (.Y(_01392_),
    .A(_01391_));
 sg13g2_o21ai_1 _06688_ (.B1(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .Y(_01393_),
    .A1(_01373_),
    .A2(_01392_));
 sg13g2_inv_1 _06689_ (.Y(_01394_),
    .A(_01393_));
 sg13g2_nand2_1 _06690_ (.Y(_01395_),
    .A(_01310_),
    .B(_01362_));
 sg13g2_buf_2 _06691_ (.A(\i_tinyqv.cpu.instr_write_offset[1] ),
    .X(_01396_));
 sg13g2_buf_1 _06692_ (.A(_01297_),
    .X(_01397_));
 sg13g2_xnor2_1 _06693_ (.Y(_01398_),
    .A(_01396_),
    .B(_01397_));
 sg13g2_buf_2 _06694_ (.A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .X(_01399_));
 sg13g2_inv_1 _06695_ (.Y(_01400_),
    .A(_00758_));
 sg13g2_nand3_1 _06696_ (.B(_01290_),
    .C(net309),
    .A(_00758_),
    .Y(_01401_));
 sg13g2_nor2b_1 _06697_ (.A(\i_tinyqv.cpu.instr_len[2] ),
    .B_N(_01401_),
    .Y(_01402_));
 sg13g2_a21oi_2 _06698_ (.B1(_01402_),
    .Y(_01403_),
    .A2(_01298_),
    .A1(_01400_));
 sg13g2_nor2b_1 _06699_ (.A(_00099_),
    .B_N(_01403_),
    .Y(_01404_));
 sg13g2_xnor2_1 _06700_ (.Y(_01405_),
    .A(_01399_),
    .B(_01404_));
 sg13g2_buf_1 _06701_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .X(_01406_));
 sg13g2_buf_1 _06702_ (.A(net169),
    .X(_01407_));
 sg13g2_buf_1 _06703_ (.A(_00095_),
    .X(_01408_));
 sg13g2_nand2_1 _06704_ (.Y(_01409_),
    .A(_01408_),
    .B(_01334_));
 sg13g2_xor2_1 _06705_ (.B(_01409_),
    .A(_01407_),
    .X(_01410_));
 sg13g2_nand2_1 _06706_ (.Y(_01411_),
    .A(_01407_),
    .B(_01409_));
 sg13g2_nor2_1 _06707_ (.A(net298),
    .B(_01411_),
    .Y(_01412_));
 sg13g2_a21oi_1 _06708_ (.A1(net298),
    .A2(_01410_),
    .Y(_01413_),
    .B1(_01412_));
 sg13g2_nor3_1 _06709_ (.A(net298),
    .B(net158),
    .C(_01409_),
    .Y(_01414_));
 sg13g2_nor2_1 _06710_ (.A(_01405_),
    .B(_01414_),
    .Y(_01415_));
 sg13g2_a221oi_1 _06711_ (.B2(_01413_),
    .C1(_01415_),
    .B1(_01405_),
    .A1(_01395_),
    .Y(_01416_),
    .A2(_01398_));
 sg13g2_nand2b_1 _06712_ (.Y(_01417_),
    .B(_00098_),
    .A_N(_01416_));
 sg13g2_a21o_1 _06713_ (.A2(_01394_),
    .A1(_01369_),
    .B1(_01417_),
    .X(_01418_));
 sg13g2_buf_1 _06714_ (.A(_01418_),
    .X(_01419_));
 sg13g2_nor4_1 _06715_ (.A(net316),
    .B(_01279_),
    .C(_01365_),
    .D(_01419_),
    .Y(_01420_));
 sg13g2_a21oi_1 _06716_ (.A1(net316),
    .A2(net83),
    .Y(_01421_),
    .B1(_01420_));
 sg13g2_inv_2 _06717_ (.Y(_01422_),
    .A(net316));
 sg13g2_inv_1 _06718_ (.Y(_01423_),
    .A(_00097_));
 sg13g2_buf_1 _06719_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .X(_01424_));
 sg13g2_nor2b_1 _06720_ (.A(_01230_),
    .B_N(_01424_),
    .Y(_01425_));
 sg13g2_buf_1 _06721_ (.A(_01425_),
    .X(_01426_));
 sg13g2_buf_1 _06722_ (.A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .X(_01427_));
 sg13g2_buf_1 _06723_ (.A(\i_tinyqv.mem.instr_active ),
    .X(_01428_));
 sg13g2_nand2_1 _06724_ (.Y(_01429_),
    .A(_01427_),
    .B(_01428_));
 sg13g2_nand3_1 _06725_ (.B(_01426_),
    .C(_01429_),
    .A(_01423_),
    .Y(_01430_));
 sg13g2_buf_2 _06726_ (.A(_00096_),
    .X(_01431_));
 sg13g2_nand3_1 _06727_ (.B(_01428_),
    .C(_01426_),
    .A(net297),
    .Y(_01432_));
 sg13g2_buf_1 _06728_ (.A(_01432_),
    .X(_01433_));
 sg13g2_nor3_2 _06729_ (.A(_01431_),
    .B(_01408_),
    .C(_01433_),
    .Y(_01434_));
 sg13g2_nand2_1 _06730_ (.Y(_01435_),
    .A(net298),
    .B(_01434_));
 sg13g2_xor2_1 _06731_ (.B(_01435_),
    .A(_01399_),
    .X(_01436_));
 sg13g2_nand4_1 _06732_ (.B(_01369_),
    .C(_01286_),
    .A(_01204_),
    .Y(_01437_),
    .D(_01403_));
 sg13g2_xnor2_1 _06733_ (.Y(_01438_),
    .A(_01436_),
    .B(_01437_));
 sg13g2_nor2_1 _06734_ (.A(_01431_),
    .B(_01433_),
    .Y(_01439_));
 sg13g2_xor2_1 _06735_ (.B(_01439_),
    .A(_01292_),
    .X(_01440_));
 sg13g2_nor3_1 _06736_ (.A(_01408_),
    .B(_01292_),
    .C(_01439_),
    .Y(_01441_));
 sg13g2_a21oi_1 _06737_ (.A1(_01408_),
    .A2(_01440_),
    .Y(_01442_),
    .B1(_01441_));
 sg13g2_nand2_1 _06738_ (.Y(_01443_),
    .A(_01292_),
    .B(_01434_));
 sg13g2_xor2_1 _06739_ (.B(_00158_),
    .A(_00101_),
    .X(_01444_));
 sg13g2_mux2_1 _06740_ (.A0(_01442_),
    .A1(_01443_),
    .S(_01444_),
    .X(_01445_));
 sg13g2_nor3_2 _06741_ (.A(_01430_),
    .B(_01438_),
    .C(_01445_),
    .Y(_01446_));
 sg13g2_nor4_1 _06742_ (.A(net317),
    .B(_01258_),
    .C(_01422_),
    .D(_01446_),
    .Y(_01447_));
 sg13g2_a21oi_1 _06743_ (.A1(_01259_),
    .A2(_01421_),
    .Y(_01448_),
    .B1(_01447_));
 sg13g2_nor2b_1 _06744_ (.A(_01341_),
    .B_N(_01343_),
    .Y(_01449_));
 sg13g2_buf_1 _06745_ (.A(_01449_),
    .X(_01450_));
 sg13g2_nor2_1 _06746_ (.A(_01328_),
    .B(_01332_),
    .Y(_01451_));
 sg13g2_nand2b_1 _06747_ (.Y(_01452_),
    .B(_01451_),
    .A_N(_01338_));
 sg13g2_buf_2 _06748_ (.A(_01452_),
    .X(_01453_));
 sg13g2_nor2_1 _06749_ (.A(_01453_),
    .B(_01351_),
    .Y(_01454_));
 sg13g2_nand2_2 _06750_ (.Y(_01455_),
    .A(_01450_),
    .B(_01454_));
 sg13g2_nand2b_1 _06751_ (.Y(_01456_),
    .B(_01308_),
    .A_N(_01306_));
 sg13g2_buf_2 _06752_ (.A(_01456_),
    .X(_01457_));
 sg13g2_nand2_2 _06753_ (.Y(_01458_),
    .A(_01457_),
    .B(_01362_));
 sg13g2_mux2_1 _06754_ (.A0(_00129_),
    .A1(_00126_),
    .S(net169),
    .X(_01459_));
 sg13g2_nor2_1 _06755_ (.A(net170),
    .B(_01459_),
    .Y(_01460_));
 sg13g2_mux2_1 _06756_ (.A0(_00128_),
    .A1(_00127_),
    .S(_01304_),
    .X(_01461_));
 sg13g2_nand2b_1 _06757_ (.Y(_01462_),
    .B(net170),
    .A_N(_01461_));
 sg13g2_nand2b_1 _06758_ (.Y(_01463_),
    .B(_01462_),
    .A_N(_01460_));
 sg13g2_buf_1 _06759_ (.A(_01463_),
    .X(_01464_));
 sg13g2_nand2b_1 _06760_ (.Y(_01465_),
    .B(_01314_),
    .A_N(_01312_));
 sg13g2_nor2_2 _06761_ (.A(_01465_),
    .B(_01322_),
    .Y(_01466_));
 sg13g2_nand2_2 _06762_ (.Y(_01467_),
    .A(_01464_),
    .B(_01466_));
 sg13g2_nor2_1 _06763_ (.A(_01458_),
    .B(_01467_),
    .Y(_01468_));
 sg13g2_nor2b_1 _06764_ (.A(_01455_),
    .B_N(_01468_),
    .Y(_01469_));
 sg13g2_mux2_1 _06765_ (.A0(_00145_),
    .A1(_00142_),
    .S(net158),
    .X(_01470_));
 sg13g2_mux2_1 _06766_ (.A0(_00144_),
    .A1(_00143_),
    .S(net158),
    .X(_01471_));
 sg13g2_mux2_1 _06767_ (.A0(_01470_),
    .A1(_01471_),
    .S(net170),
    .X(_01472_));
 sg13g2_buf_2 _06768_ (.A(_01472_),
    .X(_01473_));
 sg13g2_inv_2 _06769_ (.Y(_01474_),
    .A(_01473_));
 sg13g2_mux2_1 _06770_ (.A0(_00141_),
    .A1(_00138_),
    .S(net158),
    .X(_01475_));
 sg13g2_mux2_1 _06771_ (.A0(_00140_),
    .A1(_00139_),
    .S(net158),
    .X(_01476_));
 sg13g2_mux2_1 _06772_ (.A0(_01475_),
    .A1(_01476_),
    .S(net170),
    .X(_01477_));
 sg13g2_buf_1 _06773_ (.A(_01477_),
    .X(_01478_));
 sg13g2_inv_1 _06774_ (.Y(_01479_),
    .A(_01478_));
 sg13g2_nor2_1 _06775_ (.A(_01474_),
    .B(_01479_),
    .Y(_01480_));
 sg13g2_buf_1 _06776_ (.A(net158),
    .X(_01481_));
 sg13g2_mux4_1 _06777_ (.S0(net159),
    .A0(_00137_),
    .A1(_00136_),
    .A2(_00134_),
    .A3(_00135_),
    .S1(_01481_),
    .X(_01482_));
 sg13g2_buf_1 _06778_ (.A(_01482_),
    .X(_01483_));
 sg13g2_mux2_1 _06779_ (.A0(_00149_),
    .A1(_00146_),
    .S(net158),
    .X(_01484_));
 sg13g2_nor2_1 _06780_ (.A(net159),
    .B(_01484_),
    .Y(_01485_));
 sg13g2_mux2_1 _06781_ (.A0(_00148_),
    .A1(_00147_),
    .S(net158),
    .X(_01486_));
 sg13g2_nand2b_1 _06782_ (.Y(_01487_),
    .B(net159),
    .A_N(_01486_));
 sg13g2_nand2b_1 _06783_ (.Y(_01488_),
    .B(_01487_),
    .A_N(_01485_));
 sg13g2_buf_2 _06784_ (.A(_01488_),
    .X(_01489_));
 sg13g2_mux4_1 _06785_ (.S0(net159),
    .A0(_00133_),
    .A1(_00132_),
    .A2(_00130_),
    .A3(_00131_),
    .S1(net152),
    .X(_01490_));
 sg13g2_buf_2 _06786_ (.A(_01490_),
    .X(_01491_));
 sg13g2_nor2_1 _06787_ (.A(_01489_),
    .B(_01491_),
    .Y(_01492_));
 sg13g2_nand4_1 _06788_ (.B(_01480_),
    .C(net122),
    .A(_01469_),
    .Y(_01493_),
    .D(_01492_));
 sg13g2_buf_1 _06789_ (.A(_01493_),
    .X(_01494_));
 sg13g2_nand2_1 _06790_ (.Y(_01495_),
    .A(net124),
    .B(_01363_));
 sg13g2_a21oi_1 _06791_ (.A1(_01210_),
    .A2(_01394_),
    .Y(_01496_),
    .B1(_01417_));
 sg13g2_nand4_1 _06792_ (.B(_01164_),
    .C(_01289_),
    .A(_01282_),
    .Y(_01497_),
    .D(_01496_));
 sg13g2_a21o_1 _06793_ (.A2(_01495_),
    .A1(_01494_),
    .B1(_01497_),
    .X(_01498_));
 sg13g2_nand2_1 _06794_ (.Y(_01499_),
    .A(_00098_),
    .B(_01165_));
 sg13g2_mux2_1 _06795_ (.A0(_01498_),
    .A1(_01499_),
    .S(_01279_),
    .X(_01500_));
 sg13g2_nand2_1 _06796_ (.Y(_01501_),
    .A(_01431_),
    .B(_01500_));
 sg13g2_nor2b_1 _06797_ (.A(_01446_),
    .B_N(\i_tinyqv.cpu.instr_fetch_started ),
    .Y(_01502_));
 sg13g2_nor3_1 _06798_ (.A(net317),
    .B(_01258_),
    .C(net316),
    .Y(_01503_));
 sg13g2_xor2_1 _06799_ (.B(_01437_),
    .A(_01436_),
    .X(_01504_));
 sg13g2_nor3_1 _06800_ (.A(\addr[26] ),
    .B(\addr[25] ),
    .C(\addr[27] ),
    .Y(_01505_));
 sg13g2_buf_2 _06801_ (.A(_01505_),
    .X(_01506_));
 sg13g2_nand2_1 _06802_ (.Y(_01507_),
    .A(_01232_),
    .B(_01233_));
 sg13g2_buf_2 _06803_ (.A(_01507_),
    .X(_01508_));
 sg13g2_a21oi_2 _06804_ (.B1(_01229_),
    .Y(_01509_),
    .A2(_01508_),
    .A1(_01506_));
 sg13g2_nor2_1 _06805_ (.A(_01445_),
    .B(_01509_),
    .Y(_01510_));
 sg13g2_nand2_1 _06806_ (.Y(_01511_),
    .A(net297),
    .B(_01426_));
 sg13g2_buf_1 _06807_ (.A(_01511_),
    .X(_01512_));
 sg13g2_o21ai_1 _06808_ (.B1(_01428_),
    .Y(_01513_),
    .A1(net190),
    .A2(_01509_));
 sg13g2_a21oi_1 _06809_ (.A1(_01504_),
    .A2(_01510_),
    .Y(_01514_),
    .B1(_01513_));
 sg13g2_and2_1 _06810_ (.A(_01503_),
    .B(_01514_),
    .X(_01515_));
 sg13g2_o21ai_1 _06811_ (.B1(_01515_),
    .Y(_01516_),
    .A1(_01501_),
    .A2(_01502_));
 sg13g2_buf_1 _06812_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .X(_01517_));
 sg13g2_buf_1 _06813_ (.A(_00155_),
    .X(_01518_));
 sg13g2_inv_2 _06814_ (.Y(_01519_),
    .A(_01518_));
 sg13g2_nor3_2 _06815_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .B(_01517_),
    .C(_01519_),
    .Y(_01520_));
 sg13g2_and2_1 _06816_ (.A(_00154_),
    .B(_01520_),
    .X(_01521_));
 sg13g2_buf_1 _06817_ (.A(_01521_),
    .X(_01522_));
 sg13g2_nor2_1 _06818_ (.A(net297),
    .B(_01240_),
    .Y(_01523_));
 sg13g2_nor3_1 _06819_ (.A(debug_data_continue),
    .B(_01239_),
    .C(_01523_),
    .Y(_01524_));
 sg13g2_nor2_1 _06820_ (.A(_01428_),
    .B(_01524_),
    .Y(_01525_));
 sg13g2_nor2_1 _06821_ (.A(_01522_),
    .B(_01525_),
    .Y(_01526_));
 sg13g2_inv_1 _06822_ (.Y(_01527_),
    .A(_01526_));
 sg13g2_nor2b_1 _06823_ (.A(net317),
    .B_N(_01258_),
    .Y(_01528_));
 sg13g2_nor3_1 _06824_ (.A(_01279_),
    .B(_01497_),
    .C(_01494_),
    .Y(_01529_));
 sg13g2_nor2_1 _06825_ (.A(\i_tinyqv.cpu.is_auipc ),
    .B(_01169_),
    .Y(_01530_));
 sg13g2_nor2b_1 _06826_ (.A(_01530_),
    .B_N(net218),
    .Y(_01531_));
 sg13g2_buf_1 _06827_ (.A(_01531_),
    .X(_01532_));
 sg13g2_nand2_1 _06828_ (.Y(_01533_),
    .A(net262),
    .B(\i_tinyqv.cpu.data_ready_core ));
 sg13g2_or2_1 _06829_ (.X(_01534_),
    .B(_01533_),
    .A(_01171_));
 sg13g2_buf_2 _06830_ (.A(_01534_),
    .X(_01535_));
 sg13g2_nand2b_1 _06831_ (.Y(_01536_),
    .B(_01187_),
    .A_N(_01188_));
 sg13g2_buf_1 _06832_ (.A(_01536_),
    .X(_01537_));
 sg13g2_nand3_1 _06833_ (.B(_01535_),
    .C(_01537_),
    .A(_01207_),
    .Y(_01538_));
 sg13g2_nand4_1 _06834_ (.B(net263),
    .C(_01176_),
    .A(net313),
    .Y(_01539_),
    .D(_01532_));
 sg13g2_o21ai_1 _06835_ (.B1(_01539_),
    .Y(_01540_),
    .A1(net189),
    .A2(_01538_));
 sg13g2_buf_1 _06836_ (.A(_01540_),
    .X(_01541_));
 sg13g2_nand2_1 _06837_ (.Y(_01542_),
    .A(_01422_),
    .B(_01541_));
 sg13g2_o21ai_1 _06838_ (.B1(_01542_),
    .Y(_01543_),
    .A1(_01422_),
    .A2(_01529_));
 sg13g2_nor2b_1 _06839_ (.A(_01258_),
    .B_N(net317),
    .Y(_01544_));
 sg13g2_nand2_1 _06840_ (.Y(_01545_),
    .A(net316),
    .B(_01060_));
 sg13g2_o21ai_1 _06841_ (.B1(_01545_),
    .Y(_01546_),
    .A1(debug_data_continue),
    .A2(net316));
 sg13g2_a21o_1 _06842_ (.A2(_01546_),
    .A1(_01544_),
    .B1(net6),
    .X(_01547_));
 sg13g2_a221oi_1 _06843_ (.B2(_01543_),
    .C1(_01547_),
    .B1(_01528_),
    .A1(_01503_),
    .Y(_01548_),
    .A2(_01527_));
 sg13g2_nand3_1 _06844_ (.B(_01516_),
    .C(_01548_),
    .A(_01448_),
    .Y(_01549_));
 sg13g2_nor2_1 _06845_ (.A(net317),
    .B(net316),
    .Y(_01550_));
 sg13g2_nand3_1 _06846_ (.B(_01500_),
    .C(_01550_),
    .A(_01431_),
    .Y(_01551_));
 sg13g2_and2_1 _06847_ (.A(_01204_),
    .B(_01369_),
    .X(_01552_));
 sg13g2_buf_2 _06848_ (.A(_01552_),
    .X(_01553_));
 sg13g2_nand2_1 _06849_ (.Y(_01554_),
    .A(_01286_),
    .B(_01553_));
 sg13g2_nand2b_1 _06850_ (.Y(_01555_),
    .B(_01422_),
    .A_N(_01433_));
 sg13g2_o21ai_1 _06851_ (.B1(_01555_),
    .Y(_01556_),
    .A1(_01422_),
    .A2(_01554_));
 sg13g2_nand2b_1 _06852_ (.Y(_01557_),
    .B(_01288_),
    .A_N(net5));
 sg13g2_o21ai_1 _06853_ (.B1(_01258_),
    .Y(_01558_),
    .A1(_01422_),
    .A2(_01557_));
 sg13g2_a21oi_1 _06854_ (.A1(net317),
    .A2(_01556_),
    .Y(_01559_),
    .B1(_01558_));
 sg13g2_nor2b_1 _06855_ (.A(_01239_),
    .B_N(_01427_),
    .Y(_01560_));
 sg13g2_nor2b_1 _06856_ (.A(_01560_),
    .B_N(_00154_),
    .Y(_01561_));
 sg13g2_nor2_1 _06857_ (.A(_01423_),
    .B(_01561_),
    .Y(_01562_));
 sg13g2_buf_2 _06858_ (.A(_01562_),
    .X(_01563_));
 sg13g2_nand2b_1 _06859_ (.Y(_01564_),
    .B(_01506_),
    .A_N(_01563_));
 sg13g2_buf_1 _06860_ (.A(_01564_),
    .X(_01565_));
 sg13g2_a21oi_1 _06861_ (.A1(_01232_),
    .A2(\i_tinyqv.cpu.data_write_n[1] ),
    .Y(_01566_),
    .B1(_01506_));
 sg13g2_buf_1 _06862_ (.A(_01566_),
    .X(_01567_));
 sg13g2_a21oi_1 _06863_ (.A1(_01233_),
    .A2(\i_tinyqv.cpu.data_read_n[1] ),
    .Y(_01568_),
    .B1(_01506_));
 sg13g2_mux4_1 _06864_ (.S0(_01260_),
    .A0(_01394_),
    .A1(_01565_),
    .A2(net208),
    .A3(_01568_),
    .S1(net317),
    .X(_01569_));
 sg13g2_o21ai_1 _06865_ (.B1(net6),
    .Y(_01570_),
    .A1(_01258_),
    .A2(_01569_));
 sg13g2_a21o_1 _06866_ (.A2(_01559_),
    .A1(_01551_),
    .B1(_01570_),
    .X(_01571_));
 sg13g2_a21oi_1 _06867_ (.A1(_01549_),
    .A2(_01571_),
    .Y(_01572_),
    .B1(_01256_));
 sg13g2_a21o_1 _06868_ (.A2(\gpio_out[7] ),
    .A1(_01256_),
    .B1(_01572_),
    .X(net35));
 sg13g2_buf_2 _06869_ (.A(\data_to_write[0] ),
    .X(_01573_));
 sg13g2_inv_1 _06870_ (.Y(_01574_),
    .A(_01573_));
 sg13g2_buf_1 _06871_ (.A(\addr[4] ),
    .X(_01575_));
 sg13g2_buf_1 _06872_ (.A(\addr[5] ),
    .X(_01576_));
 sg13g2_nor2_1 _06873_ (.A(_01575_),
    .B(net296),
    .Y(_01577_));
 sg13g2_buf_2 _06874_ (.A(\addr[2] ),
    .X(_01578_));
 sg13g2_buf_1 _06875_ (.A(\addr[3] ),
    .X(_01579_));
 sg13g2_nor4_1 _06876_ (.A(\addr[16] ),
    .B(\addr[19] ),
    .C(\addr[18] ),
    .D(\addr[21] ),
    .Y(_01580_));
 sg13g2_nor4_1 _06877_ (.A(\addr[20] ),
    .B(\addr[23] ),
    .C(\addr[22] ),
    .D(\addr[24] ),
    .Y(_01581_));
 sg13g2_nor4_1 _06878_ (.A(\addr[0] ),
    .B(\addr[7] ),
    .C(\addr[6] ),
    .D(\addr[9] ),
    .Y(_01582_));
 sg13g2_inv_1 _06879_ (.Y(_01583_),
    .A(\addr[27] ));
 sg13g2_nor4_1 _06880_ (.A(_01583_),
    .B(\addr[1] ),
    .C(\addr[14] ),
    .D(\addr[17] ),
    .Y(_01584_));
 sg13g2_nand4_1 _06881_ (.B(_01581_),
    .C(_01582_),
    .A(_01580_),
    .Y(_01585_),
    .D(_01584_));
 sg13g2_nor4_1 _06882_ (.A(\addr[11] ),
    .B(\addr[10] ),
    .C(\addr[13] ),
    .D(\addr[15] ),
    .Y(_01586_));
 sg13g2_nor4_1 _06883_ (.A(\addr[26] ),
    .B(\addr[25] ),
    .C(\addr[8] ),
    .D(\addr[12] ),
    .Y(_01587_));
 sg13g2_nand2_1 _06884_ (.Y(_01588_),
    .A(_01586_),
    .B(_01587_));
 sg13g2_nor2_2 _06885_ (.A(_01585_),
    .B(_01588_),
    .Y(_01589_));
 sg13g2_inv_1 _06886_ (.Y(_01590_),
    .A(_01589_));
 sg13g2_nor3_2 _06887_ (.A(_01578_),
    .B(net295),
    .C(_01590_),
    .Y(_01591_));
 sg13g2_and2_1 _06888_ (.A(_01577_),
    .B(_01591_),
    .X(_01592_));
 sg13g2_buf_2 _06889_ (.A(_01592_),
    .X(_01593_));
 sg13g2_nand2_1 _06890_ (.Y(_01594_),
    .A(net208),
    .B(_01593_));
 sg13g2_buf_2 _06891_ (.A(_01594_),
    .X(_01595_));
 sg13g2_buf_1 _06892_ (.A(_01595_),
    .X(_01596_));
 sg13g2_buf_1 _06893_ (.A(\i_debug_uart_tx.resetn ),
    .X(_01597_));
 sg13g2_buf_1 _06894_ (.A(net261),
    .X(_01598_));
 sg13g2_nand3_1 _06895_ (.B(\gpio_out[0] ),
    .C(net110),
    .A(net217),
    .Y(_01599_));
 sg13g2_o21ai_1 _06896_ (.B1(_01599_),
    .Y(_00000_),
    .A1(_01574_),
    .A2(net110));
 sg13g2_buf_2 _06897_ (.A(\data_to_write[1] ),
    .X(_01600_));
 sg13g2_inv_1 _06898_ (.Y(_01601_),
    .A(_01600_));
 sg13g2_nand3_1 _06899_ (.B(\gpio_out[1] ),
    .C(net110),
    .A(net217),
    .Y(_01602_));
 sg13g2_o21ai_1 _06900_ (.B1(_01602_),
    .Y(_00001_),
    .A1(_01601_),
    .A2(_01596_));
 sg13g2_buf_2 _06901_ (.A(\data_to_write[2] ),
    .X(_01603_));
 sg13g2_inv_1 _06902_ (.Y(_01604_),
    .A(_01603_));
 sg13g2_nand3_1 _06903_ (.B(\gpio_out[2] ),
    .C(_01595_),
    .A(net217),
    .Y(_01605_));
 sg13g2_o21ai_1 _06904_ (.B1(_01605_),
    .Y(_00002_),
    .A1(_01604_),
    .A2(net110));
 sg13g2_buf_2 _06905_ (.A(\data_to_write[3] ),
    .X(_01606_));
 sg13g2_inv_1 _06906_ (.Y(_01607_),
    .A(_01606_));
 sg13g2_nand3_1 _06907_ (.B(\gpio_out[3] ),
    .C(_01595_),
    .A(net217),
    .Y(_01608_));
 sg13g2_o21ai_1 _06908_ (.B1(_01608_),
    .Y(_00003_),
    .A1(_01607_),
    .A2(net110));
 sg13g2_buf_1 _06909_ (.A(\data_to_write[4] ),
    .X(_01609_));
 sg13g2_inv_1 _06910_ (.Y(_01610_),
    .A(_01609_));
 sg13g2_nand3_1 _06911_ (.B(\gpio_out[4] ),
    .C(_01595_),
    .A(net217),
    .Y(_01611_));
 sg13g2_o21ai_1 _06912_ (.B1(_01611_),
    .Y(_00004_),
    .A1(_01610_),
    .A2(net110));
 sg13g2_buf_1 _06913_ (.A(\data_to_write[5] ),
    .X(_01612_));
 sg13g2_inv_1 _06914_ (.Y(_01613_),
    .A(_01612_));
 sg13g2_buf_1 _06915_ (.A(net261),
    .X(_01614_));
 sg13g2_nand3_1 _06916_ (.B(\gpio_out[5] ),
    .C(_01595_),
    .A(net216),
    .Y(_01615_));
 sg13g2_o21ai_1 _06917_ (.B1(_01615_),
    .Y(_00005_),
    .A1(_01613_),
    .A2(net110));
 sg13g2_buf_1 _06918_ (.A(\data_to_write[6] ),
    .X(_01616_));
 sg13g2_inv_1 _06919_ (.Y(_01617_),
    .A(_01616_));
 sg13g2_nand3_1 _06920_ (.B(\gpio_out[6] ),
    .C(_01595_),
    .A(_01614_),
    .Y(_01618_));
 sg13g2_o21ai_1 _06921_ (.B1(_01618_),
    .Y(_00006_),
    .A1(_01617_),
    .A2(_01596_));
 sg13g2_inv_1 _06922_ (.Y(_01619_),
    .A(\data_to_write[7] ));
 sg13g2_nand3_1 _06923_ (.B(\gpio_out[7] ),
    .C(_01595_),
    .A(net216),
    .Y(_01620_));
 sg13g2_o21ai_1 _06924_ (.B1(_01620_),
    .Y(_00007_),
    .A1(_01619_),
    .A2(net110));
 sg13g2_and4_1 _06925_ (.A(_01578_),
    .B(net295),
    .C(_01577_),
    .D(_01589_),
    .X(_01621_));
 sg13g2_buf_1 _06926_ (.A(_01621_),
    .X(_01622_));
 sg13g2_and2_1 _06927_ (.A(net208),
    .B(net167),
    .X(_01623_));
 sg13g2_buf_1 _06928_ (.A(_01623_),
    .X(_01624_));
 sg13g2_buf_1 _06929_ (.A(_01624_),
    .X(_01625_));
 sg13g2_nand2_1 _06930_ (.Y(_01626_),
    .A(net216),
    .B(\gpio_out_sel[0] ));
 sg13g2_nand2_1 _06931_ (.Y(_01627_),
    .A(_01573_),
    .B(net135));
 sg13g2_o21ai_1 _06932_ (.B1(_01627_),
    .Y(_00008_),
    .A1(net135),
    .A2(_01626_));
 sg13g2_nand2_1 _06933_ (.Y(_01628_),
    .A(net216),
    .B(\gpio_out_sel[1] ));
 sg13g2_nand2_1 _06934_ (.Y(_01629_),
    .A(_01600_),
    .B(net135));
 sg13g2_o21ai_1 _06935_ (.B1(_01629_),
    .Y(_00009_),
    .A1(net135),
    .A2(_01628_));
 sg13g2_nand2_1 _06936_ (.Y(_01630_),
    .A(net216),
    .B(\gpio_out_sel[2] ));
 sg13g2_nand2_1 _06937_ (.Y(_01631_),
    .A(_01603_),
    .B(_01624_));
 sg13g2_o21ai_1 _06938_ (.B1(_01631_),
    .Y(_00010_),
    .A1(_01625_),
    .A2(_01630_));
 sg13g2_nand2_1 _06939_ (.Y(_01632_),
    .A(net216),
    .B(\gpio_out_sel[3] ));
 sg13g2_nand2_1 _06940_ (.Y(_01633_),
    .A(_01606_),
    .B(_01624_));
 sg13g2_o21ai_1 _06941_ (.B1(_01633_),
    .Y(_00011_),
    .A1(net135),
    .A2(_01632_));
 sg13g2_nand2_1 _06942_ (.Y(_01634_),
    .A(net216),
    .B(\gpio_out_sel[4] ));
 sg13g2_nand2_1 _06943_ (.Y(_01635_),
    .A(_01609_),
    .B(_01624_));
 sg13g2_o21ai_1 _06944_ (.B1(_01635_),
    .Y(_00012_),
    .A1(_01625_),
    .A2(_01634_));
 sg13g2_nand2_1 _06945_ (.Y(_01636_),
    .A(net216),
    .B(\gpio_out_sel[5] ));
 sg13g2_nand2_1 _06946_ (.Y(_01637_),
    .A(_01612_),
    .B(_01624_));
 sg13g2_o21ai_1 _06947_ (.B1(_01637_),
    .Y(_00013_),
    .A1(net135),
    .A2(_01636_));
 sg13g2_nand2_1 _06948_ (.Y(_01638_),
    .A(net261),
    .B(\gpio_out_sel[6] ));
 sg13g2_nand2_1 _06949_ (.Y(_01639_),
    .A(_01616_),
    .B(_01624_));
 sg13g2_o21ai_1 _06950_ (.B1(_01639_),
    .Y(_00014_),
    .A1(net135),
    .A2(_01638_));
 sg13g2_nor2_1 _06951_ (.A(net261),
    .B(_01257_),
    .Y(_01640_));
 sg13g2_a221oi_1 _06952_ (.B2(net167),
    .C1(_01640_),
    .B1(net208),
    .A1(net261),
    .Y(_01641_),
    .A2(_01256_));
 sg13g2_a21oi_1 _06953_ (.A1(_01619_),
    .A2(net135),
    .Y(_00015_),
    .B1(_01641_));
 sg13g2_buf_1 _06954_ (.A(_00164_),
    .X(_01642_));
 sg13g2_buf_1 _06955_ (.A(_01642_),
    .X(_01643_));
 sg13g2_buf_1 _06956_ (.A(_01554_),
    .X(_01644_));
 sg13g2_a21oi_1 _06957_ (.A1(_01170_),
    .A2(net85),
    .Y(_01645_),
    .B1(_01196_));
 sg13g2_buf_1 _06958_ (.A(\i_tinyqv.cpu.i_core.cycle[0] ),
    .X(_01646_));
 sg13g2_buf_1 _06959_ (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .X(_01647_));
 sg13g2_nor2_2 _06960_ (.A(_01646_),
    .B(_01647_),
    .Y(_01648_));
 sg13g2_nand2_1 _06961_ (.Y(_01649_),
    .A(_01196_),
    .B(\i_tinyqv.cpu.no_write_in_progress ));
 sg13g2_nand2_1 _06962_ (.Y(_01650_),
    .A(_01171_),
    .B(_01649_));
 sg13g2_and4_1 _06963_ (.A(net218),
    .B(net160),
    .C(_01648_),
    .D(_01650_),
    .X(_01651_));
 sg13g2_buf_1 _06964_ (.A(_01651_),
    .X(_01652_));
 sg13g2_nand2b_1 _06965_ (.Y(_01653_),
    .B(_01652_),
    .A_N(_01645_));
 sg13g2_nand4_1 _06966_ (.B(net160),
    .C(_01648_),
    .A(net218),
    .Y(_01654_),
    .D(_01650_));
 sg13g2_buf_1 _06967_ (.A(_01654_),
    .X(_01655_));
 sg13g2_nor2_1 _06968_ (.A(_01286_),
    .B(net134),
    .Y(_01656_));
 sg13g2_a22oi_1 _06969_ (.Y(_01657_),
    .B1(_01656_),
    .B2(_01196_),
    .A2(_01653_),
    .A1(debug_data_continue));
 sg13g2_buf_1 _06970_ (.A(net85),
    .X(_01658_));
 sg13g2_nand3_1 _06971_ (.B(net82),
    .C(_01656_),
    .A(_01170_),
    .Y(_01659_));
 sg13g2_o21ai_1 _06972_ (.B1(_01659_),
    .Y(_00028_),
    .A1(net260),
    .A2(_01657_));
 sg13g2_buf_1 _06973_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .X(_01660_));
 sg13g2_buf_1 _06974_ (.A(_01660_),
    .X(_01661_));
 sg13g2_buf_1 _06975_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .X(_01662_));
 sg13g2_and2_1 _06976_ (.A(net259),
    .B(_01662_),
    .X(_01663_));
 sg13g2_buf_2 _06977_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .X(_01664_));
 sg13g2_a21oi_1 _06978_ (.A1(_00793_),
    .A2(_00819_),
    .Y(_01665_),
    .B1(_01173_));
 sg13g2_buf_2 _06979_ (.A(_01665_),
    .X(_01666_));
 sg13g2_or2_1 _06980_ (.X(_01667_),
    .B(_01666_),
    .A(_01664_));
 sg13g2_and2_1 _06981_ (.A(_00776_),
    .B(_00792_),
    .X(_01668_));
 sg13g2_buf_2 _06982_ (.A(_01668_),
    .X(_01669_));
 sg13g2_nand3_1 _06983_ (.B(_00812_),
    .C(_00817_),
    .A(_00808_),
    .Y(_01670_));
 sg13g2_buf_2 _06984_ (.A(_01670_),
    .X(_01671_));
 sg13g2_inv_1 _06985_ (.Y(_01672_),
    .A(_01664_));
 sg13g2_nor2_1 _06986_ (.A(_01173_),
    .B(_01672_),
    .Y(_01673_));
 sg13g2_o21ai_1 _06987_ (.B1(_01673_),
    .Y(_01674_),
    .A1(_01669_),
    .A2(_01671_));
 sg13g2_buf_2 _06988_ (.A(_01674_),
    .X(_01675_));
 sg13g2_and2_1 _06989_ (.A(net219),
    .B(_01135_),
    .X(_01676_));
 sg13g2_buf_1 _06990_ (.A(_01676_),
    .X(_01677_));
 sg13g2_nand3_1 _06991_ (.B(_01007_),
    .C(_01014_),
    .A(_01004_),
    .Y(_01678_));
 sg13g2_buf_1 _06992_ (.A(_01678_),
    .X(_01679_));
 sg13g2_and2_1 _06993_ (.A(net219),
    .B(_01679_),
    .X(_01680_));
 sg13g2_buf_2 _06994_ (.A(_01680_),
    .X(_01681_));
 sg13g2_nand2_1 _06995_ (.Y(_01682_),
    .A(_01677_),
    .B(_01681_));
 sg13g2_a21oi_1 _06996_ (.A1(_01667_),
    .A2(_01675_),
    .Y(_01683_),
    .B1(_01682_));
 sg13g2_and2_1 _06997_ (.A(_01663_),
    .B(_01683_),
    .X(_01684_));
 sg13g2_inv_1 _06998_ (.Y(_01685_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[2] ));
 sg13g2_nor2_1 _06999_ (.A(_01669_),
    .B(_01671_),
    .Y(_01686_));
 sg13g2_nor2b_1 _07000_ (.A(_01173_),
    .B_N(_01660_),
    .Y(_01687_));
 sg13g2_and4_1 _07001_ (.A(_01672_),
    .B(_01686_),
    .C(net153),
    .D(_01687_),
    .X(_01688_));
 sg13g2_inv_1 _07002_ (.Y(_01689_),
    .A(_01662_));
 sg13g2_nor2_2 _07003_ (.A(_01173_),
    .B(_01689_),
    .Y(_01690_));
 sg13g2_and3_1 _07004_ (.X(_01691_),
    .A(_01135_),
    .B(_01679_),
    .C(_01690_));
 sg13g2_nor3_1 _07005_ (.A(net263),
    .B(_01660_),
    .C(_01672_),
    .Y(_01692_));
 sg13g2_a21oi_1 _07006_ (.A1(_00793_),
    .A2(_00819_),
    .Y(_01693_),
    .B1(net153));
 sg13g2_and3_1 _07007_ (.X(_01694_),
    .A(_01679_),
    .B(_01690_),
    .C(_01687_));
 sg13g2_a22oi_1 _07008_ (.Y(_01695_),
    .B1(_01693_),
    .B2(_01694_),
    .A2(_01692_),
    .A1(_01691_));
 sg13g2_nand2_2 _07009_ (.Y(_01696_),
    .A(_00793_),
    .B(_00819_));
 sg13g2_nand4_1 _07010_ (.B(_01696_),
    .C(net153),
    .A(_01664_),
    .Y(_01697_),
    .D(_01687_));
 sg13g2_nand3b_1 _07011_ (.B(_01695_),
    .C(_01697_),
    .Y(_01698_),
    .A_N(_01688_));
 sg13g2_buf_1 _07012_ (.A(_01679_),
    .X(_01699_));
 sg13g2_and2_1 _07013_ (.A(net151),
    .B(_01690_),
    .X(_01700_));
 sg13g2_a21oi_1 _07014_ (.A1(_01664_),
    .A2(_01135_),
    .Y(_01701_),
    .B1(_01660_));
 sg13g2_nor3_1 _07015_ (.A(_01669_),
    .B(_01671_),
    .C(net153),
    .Y(_01702_));
 sg13g2_nor3_1 _07016_ (.A(net263),
    .B(_01701_),
    .C(_01702_),
    .Y(_01703_));
 sg13g2_nor2_1 _07017_ (.A(_01700_),
    .B(_01703_),
    .Y(_01704_));
 sg13g2_nor3_1 _07018_ (.A(_01685_),
    .B(_01698_),
    .C(_01704_),
    .Y(_01705_));
 sg13g2_nor2_1 _07019_ (.A(_01684_),
    .B(_01705_),
    .Y(_01706_));
 sg13g2_buf_2 _07020_ (.A(_01706_),
    .X(_01707_));
 sg13g2_nand2_1 _07021_ (.Y(_01708_),
    .A(net151),
    .B(_01690_));
 sg13g2_buf_1 _07022_ (.A(net153),
    .X(_01709_));
 sg13g2_a22oi_1 _07023_ (.Y(_01710_),
    .B1(net133),
    .B2(_01664_),
    .A2(_01696_),
    .A1(net259));
 sg13g2_o21ai_1 _07024_ (.B1(_01697_),
    .Y(_01711_),
    .A1(_01708_),
    .A2(_01710_));
 sg13g2_inv_1 _07025_ (.Y(_01712_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[3] ));
 sg13g2_o21ai_1 _07026_ (.B1(_01690_),
    .Y(_01713_),
    .A1(_01669_),
    .A2(_01671_));
 sg13g2_buf_2 _07027_ (.A(_01713_),
    .X(_01714_));
 sg13g2_inv_1 _07028_ (.Y(_01715_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ));
 sg13g2_nor2_1 _07029_ (.A(_01173_),
    .B(_01715_),
    .Y(_01716_));
 sg13g2_nand2_1 _07030_ (.Y(_01717_),
    .A(_01135_),
    .B(_01716_));
 sg13g2_buf_2 _07031_ (.A(_01717_),
    .X(_01718_));
 sg13g2_nand3_1 _07032_ (.B(_01012_),
    .C(_01013_),
    .A(_01009_),
    .Y(_01719_));
 sg13g2_and2_1 _07033_ (.A(_01219_),
    .B(_00796_),
    .X(_01720_));
 sg13g2_inv_1 _07034_ (.Y(_01721_),
    .A(net225));
 sg13g2_nand2_1 _07035_ (.Y(_01722_),
    .A(_01721_),
    .B(_01219_));
 sg13g2_a21oi_1 _07036_ (.A1(_01000_),
    .A2(_01003_),
    .Y(_01723_),
    .B1(_01722_));
 sg13g2_a221oi_1 _07037_ (.B2(_01006_),
    .C1(_01723_),
    .B1(_01720_),
    .A1(net219),
    .Y(_01724_),
    .A2(_01719_));
 sg13g2_buf_2 _07038_ (.A(_01724_),
    .X(_01725_));
 sg13g2_or2_1 _07039_ (.X(_01726_),
    .B(_01725_),
    .A(_01672_));
 sg13g2_buf_1 _07040_ (.A(_01726_),
    .X(_01727_));
 sg13g2_xor2_1 _07041_ (.B(_01727_),
    .A(_01718_),
    .X(_01728_));
 sg13g2_xnor2_1 _07042_ (.Y(_01729_),
    .A(_01714_),
    .B(_01728_));
 sg13g2_xnor2_1 _07043_ (.Y(_01730_),
    .A(_01712_),
    .B(_01729_));
 sg13g2_xnor2_1 _07044_ (.Y(_01731_),
    .A(_01711_),
    .B(_01730_));
 sg13g2_buf_2 _07045_ (.A(_01731_),
    .X(_01732_));
 sg13g2_or3_1 _07046_ (.A(_01685_),
    .B(_01698_),
    .C(_01704_),
    .X(_01733_));
 sg13g2_buf_1 _07047_ (.A(_01733_),
    .X(_01734_));
 sg13g2_buf_1 _07048_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .X(_01735_));
 sg13g2_nand2_2 _07049_ (.Y(_01736_),
    .A(net219),
    .B(_01135_));
 sg13g2_nor2_1 _07050_ (.A(_01689_),
    .B(_01736_),
    .Y(_01737_));
 sg13g2_nand2_1 _07051_ (.Y(_01738_),
    .A(net259),
    .B(_01681_));
 sg13g2_nand3_1 _07052_ (.B(_01737_),
    .C(_01738_),
    .A(_01735_),
    .Y(_01739_));
 sg13g2_buf_1 _07053_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .X(_01740_));
 sg13g2_or2_1 _07054_ (.X(_01741_),
    .B(_01735_),
    .A(_01740_));
 sg13g2_mux2_1 _07055_ (.A0(_01689_),
    .A1(_01735_),
    .S(_01736_),
    .X(_01742_));
 sg13g2_nand4_1 _07056_ (.B(_01681_),
    .C(_01741_),
    .A(_01661_),
    .Y(_01743_),
    .D(_01742_));
 sg13g2_a21o_1 _07057_ (.A2(_01725_),
    .A1(_01662_),
    .B1(_01735_),
    .X(_01744_));
 sg13g2_nand4_1 _07058_ (.B(_01740_),
    .C(_01677_),
    .A(_01661_),
    .Y(_01745_),
    .D(_01744_));
 sg13g2_nand3_1 _07059_ (.B(_01743_),
    .C(_01745_),
    .A(_01739_),
    .Y(_01746_));
 sg13g2_buf_1 _07060_ (.A(_01746_),
    .X(_01747_));
 sg13g2_o21ai_1 _07061_ (.B1(_01685_),
    .Y(_01748_),
    .A1(_01698_),
    .A2(_01704_));
 sg13g2_buf_1 _07062_ (.A(_01748_),
    .X(_01749_));
 sg13g2_nand3_1 _07063_ (.B(_01747_),
    .C(_01749_),
    .A(_01734_),
    .Y(_01750_));
 sg13g2_buf_2 _07064_ (.A(_01750_),
    .X(_01751_));
 sg13g2_and2_1 _07065_ (.A(_01732_),
    .B(_01751_),
    .X(_01752_));
 sg13g2_o21ai_1 _07066_ (.B1(_01707_),
    .Y(_01753_),
    .A1(_01732_),
    .A2(_01751_));
 sg13g2_nand2b_1 _07067_ (.Y(_01754_),
    .B(_01753_),
    .A_N(_01752_));
 sg13g2_nor2_1 _07068_ (.A(net263),
    .B(net154),
    .Y(_01755_));
 sg13g2_buf_1 _07069_ (.A(_01755_),
    .X(_01756_));
 sg13g2_nand2_1 _07070_ (.Y(_01757_),
    .A(net259),
    .B(net121));
 sg13g2_buf_1 _07071_ (.A(_01757_),
    .X(_01758_));
 sg13g2_nor4_1 _07072_ (.A(_01707_),
    .B(_01732_),
    .C(net98),
    .D(_01751_),
    .Y(_01759_));
 sg13g2_a221oi_1 _07073_ (.B2(net98),
    .C1(_01759_),
    .B1(_01754_),
    .A1(_01707_),
    .Y(_01760_),
    .A2(_01752_));
 sg13g2_nand2_1 _07074_ (.Y(_01761_),
    .A(_01711_),
    .B(_01729_));
 sg13g2_nor2_1 _07075_ (.A(_01711_),
    .B(_01729_),
    .Y(_01762_));
 sg13g2_a21oi_2 _07076_ (.B1(_01762_),
    .Y(_01763_),
    .A2(_01761_),
    .A1(_01712_));
 sg13g2_nor3_2 _07077_ (.A(net263),
    .B(_01689_),
    .C(net154),
    .Y(_01764_));
 sg13g2_buf_1 _07078_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .X(_01765_));
 sg13g2_nor2b_1 _07079_ (.A(_01173_),
    .B_N(_01765_),
    .Y(_01766_));
 sg13g2_buf_1 _07080_ (.A(_01766_),
    .X(_01767_));
 sg13g2_nand2_1 _07081_ (.Y(_01768_),
    .A(_01135_),
    .B(_01767_));
 sg13g2_buf_2 _07082_ (.A(_01768_),
    .X(_01769_));
 sg13g2_nor2_1 _07083_ (.A(_01715_),
    .B(_01725_),
    .Y(_01770_));
 sg13g2_xnor2_1 _07084_ (.Y(_01771_),
    .A(_01769_),
    .B(_01770_));
 sg13g2_xnor2_1 _07085_ (.Y(_01772_),
    .A(_01675_),
    .B(_01771_));
 sg13g2_o21ai_1 _07086_ (.B1(_01727_),
    .Y(_01773_),
    .A1(_01718_),
    .A2(_01714_));
 sg13g2_a21oi_1 _07087_ (.A1(_01718_),
    .A2(_01714_),
    .Y(_01774_),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[4] ));
 sg13g2_and2_1 _07088_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .B(_01727_),
    .X(_01775_));
 sg13g2_or2_1 _07089_ (.X(_01776_),
    .B(_01714_),
    .A(_01718_));
 sg13g2_and3_1 _07090_ (.X(_01777_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .B(_01718_),
    .C(_01714_));
 sg13g2_a221oi_1 _07091_ (.B2(_01776_),
    .C1(_01777_),
    .B1(_01775_),
    .A1(_01773_),
    .Y(_01778_),
    .A2(_01774_));
 sg13g2_xnor2_1 _07092_ (.Y(_01779_),
    .A(_01772_),
    .B(_01778_));
 sg13g2_xnor2_1 _07093_ (.Y(_01780_),
    .A(_01764_),
    .B(_01779_));
 sg13g2_xnor2_1 _07094_ (.Y(_01781_),
    .A(_01763_),
    .B(_01780_));
 sg13g2_xor2_1 _07095_ (.B(_01781_),
    .A(_01760_),
    .X(_00016_));
 sg13g2_nor4_1 _07096_ (.A(_01732_),
    .B(net98),
    .C(_01763_),
    .D(_01780_),
    .Y(_01782_));
 sg13g2_a21o_1 _07097_ (.A2(_01761_),
    .A1(_01712_),
    .B1(_01762_),
    .X(_01783_));
 sg13g2_buf_1 _07098_ (.A(_01783_),
    .X(_01784_));
 sg13g2_xor2_1 _07099_ (.B(_01779_),
    .A(_01764_),
    .X(_01785_));
 sg13g2_nor4_1 _07100_ (.A(_01732_),
    .B(net98),
    .C(_01784_),
    .D(_01785_),
    .Y(_01786_));
 sg13g2_nor4_1 _07101_ (.A(net98),
    .B(_01751_),
    .C(_01763_),
    .D(_01780_),
    .Y(_01787_));
 sg13g2_nor4_1 _07102_ (.A(_01759_),
    .B(_01782_),
    .C(_01786_),
    .D(_01787_),
    .Y(_01788_));
 sg13g2_nor4_1 _07103_ (.A(net98),
    .B(_01751_),
    .C(_01784_),
    .D(_01785_),
    .Y(_01789_));
 sg13g2_nor4_1 _07104_ (.A(_01707_),
    .B(net98),
    .C(_01763_),
    .D(_01780_),
    .Y(_01790_));
 sg13g2_nor4_1 _07105_ (.A(_01707_),
    .B(net98),
    .C(_01784_),
    .D(_01785_),
    .Y(_01791_));
 sg13g2_nor3_1 _07106_ (.A(_01789_),
    .B(_01790_),
    .C(_01791_),
    .Y(_01792_));
 sg13g2_a221oi_1 _07107_ (.B2(_01749_),
    .C1(_01705_),
    .B1(_01747_),
    .A1(_01663_),
    .Y(_01793_),
    .A2(_01683_));
 sg13g2_nand4_1 _07108_ (.B(_01734_),
    .C(_01747_),
    .A(_01684_),
    .Y(_01794_),
    .D(_01749_));
 sg13g2_o21ai_1 _07109_ (.B1(_01794_),
    .Y(_01795_),
    .A1(_01732_),
    .A2(_01793_));
 sg13g2_nand2_1 _07110_ (.Y(_01796_),
    .A(_01795_),
    .B(_01781_));
 sg13g2_nand3_1 _07111_ (.B(_01792_),
    .C(_01796_),
    .A(_01788_),
    .Y(_01797_));
 sg13g2_nor2_1 _07112_ (.A(_01764_),
    .B(_01779_),
    .Y(_01798_));
 sg13g2_nand2_1 _07113_ (.Y(_01799_),
    .A(_01764_),
    .B(_01779_));
 sg13g2_o21ai_1 _07114_ (.B1(_01799_),
    .Y(_01800_),
    .A1(_01784_),
    .A2(_01798_));
 sg13g2_nand2_1 _07115_ (.Y(_01801_),
    .A(_01718_),
    .B(_01714_));
 sg13g2_and2_1 _07116_ (.A(_01773_),
    .B(_01801_),
    .X(_01802_));
 sg13g2_nand2_1 _07117_ (.Y(_01803_),
    .A(_01802_),
    .B(_01772_));
 sg13g2_o21ai_1 _07118_ (.B1(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .Y(_01804_),
    .A1(_01802_),
    .A2(_01772_));
 sg13g2_nand2_1 _07119_ (.Y(_01805_),
    .A(_01803_),
    .B(_01804_));
 sg13g2_nand2_1 _07120_ (.Y(_01806_),
    .A(net151),
    .B(_01767_));
 sg13g2_o21ai_1 _07121_ (.B1(_01716_),
    .Y(_01807_),
    .A1(_01669_),
    .A2(_01671_));
 sg13g2_buf_1 _07122_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .X(_01808_));
 sg13g2_inv_1 _07123_ (.Y(_01809_),
    .A(_01808_));
 sg13g2_nor2_2 _07124_ (.A(net263),
    .B(_01809_),
    .Y(_01810_));
 sg13g2_nand2_1 _07125_ (.Y(_01811_),
    .A(net153),
    .B(_01810_));
 sg13g2_xnor2_1 _07126_ (.Y(_01812_),
    .A(_01807_),
    .B(_01811_));
 sg13g2_xnor2_1 _07127_ (.Y(_01813_),
    .A(_01806_),
    .B(_01812_));
 sg13g2_buf_8 _07128_ (.A(_01725_),
    .X(_01814_));
 sg13g2_or2_1 _07129_ (.X(_01815_),
    .B(net132),
    .A(_01715_));
 sg13g2_o21ai_1 _07130_ (.B1(_01815_),
    .Y(_01816_),
    .A1(_01675_),
    .A2(_01769_));
 sg13g2_a21oi_1 _07131_ (.A1(_01675_),
    .A2(_01769_),
    .Y(_01817_),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[5] ));
 sg13g2_inv_1 _07132_ (.Y(_01818_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ));
 sg13g2_nor2_1 _07133_ (.A(_01818_),
    .B(_01770_),
    .Y(_01819_));
 sg13g2_or2_1 _07134_ (.X(_01820_),
    .B(_01769_),
    .A(_01675_));
 sg13g2_and3_1 _07135_ (.X(_01821_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .B(_01675_),
    .C(_01769_));
 sg13g2_a221oi_1 _07136_ (.B2(_01820_),
    .C1(_01821_),
    .B1(_01819_),
    .A1(_01816_),
    .Y(_01822_),
    .A2(_01817_));
 sg13g2_xnor2_1 _07137_ (.Y(_01823_),
    .A(_01813_),
    .B(_01822_));
 sg13g2_nand2_1 _07138_ (.Y(_01824_),
    .A(_01664_),
    .B(net121));
 sg13g2_xnor2_1 _07139_ (.Y(_01825_),
    .A(_01823_),
    .B(_01824_));
 sg13g2_xnor2_1 _07140_ (.Y(_01826_),
    .A(_01805_),
    .B(_01825_));
 sg13g2_xnor2_1 _07141_ (.Y(_01827_),
    .A(_01800_),
    .B(_01826_));
 sg13g2_xnor2_1 _07142_ (.Y(_00019_),
    .A(_01797_),
    .B(_01827_));
 sg13g2_or2_1 _07143_ (.X(_01828_),
    .B(_01826_),
    .A(_01800_));
 sg13g2_inv_1 _07144_ (.Y(_01829_),
    .A(_01828_));
 sg13g2_a22oi_1 _07145_ (.Y(_01830_),
    .B1(_01800_),
    .B2(_01826_),
    .A2(_01781_),
    .A1(_01795_));
 sg13g2_and3_1 _07146_ (.X(_01831_),
    .A(_01788_),
    .B(_01792_),
    .C(_01830_));
 sg13g2_buf_1 _07147_ (.A(_01831_),
    .X(_01832_));
 sg13g2_or2_1 _07148_ (.X(_01833_),
    .B(_01832_),
    .A(_01829_));
 sg13g2_nand2_1 _07149_ (.Y(_01834_),
    .A(_01823_),
    .B(_01824_));
 sg13g2_nor2_1 _07150_ (.A(_01823_),
    .B(_01824_),
    .Y(_01835_));
 sg13g2_a21oi_1 _07151_ (.A1(_01805_),
    .A2(_01834_),
    .Y(_01836_),
    .B1(_01835_));
 sg13g2_nand2_1 _07152_ (.Y(_01837_),
    .A(_01675_),
    .B(_01769_));
 sg13g2_nand2_1 _07153_ (.Y(_01838_),
    .A(_01816_),
    .B(_01837_));
 sg13g2_o21ai_1 _07154_ (.B1(_01818_),
    .Y(_01839_),
    .A1(_01813_),
    .A2(_01838_));
 sg13g2_nand2_1 _07155_ (.Y(_01840_),
    .A(_01813_),
    .B(_01838_));
 sg13g2_and2_1 _07156_ (.A(_01839_),
    .B(_01840_),
    .X(_01841_));
 sg13g2_nand2_1 _07157_ (.Y(_01842_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net121));
 sg13g2_nand2_1 _07158_ (.Y(_01843_),
    .A(net219),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[6] ));
 sg13g2_nand2b_1 _07159_ (.Y(_01844_),
    .B(net133),
    .A_N(_01843_));
 sg13g2_or2_1 _07160_ (.X(_01845_),
    .B(_01725_),
    .A(_01809_));
 sg13g2_buf_1 _07161_ (.A(_01845_),
    .X(_01846_));
 sg13g2_o21ai_1 _07162_ (.B1(_01767_),
    .Y(_01847_),
    .A1(_01669_),
    .A2(_01671_));
 sg13g2_buf_1 _07163_ (.A(_01847_),
    .X(_01848_));
 sg13g2_xor2_1 _07164_ (.B(_01848_),
    .A(_01846_),
    .X(_01849_));
 sg13g2_xnor2_1 _07165_ (.Y(_01850_),
    .A(_01844_),
    .B(_01849_));
 sg13g2_nand4_1 _07166_ (.B(net151),
    .C(_01767_),
    .A(net133),
    .Y(_01851_),
    .D(_01810_));
 sg13g2_a22oi_1 _07167_ (.Y(_01852_),
    .B1(_01810_),
    .B2(net133),
    .A2(_01767_),
    .A1(net151));
 sg13g2_a21oi_2 _07168_ (.B1(_01852_),
    .Y(_01853_),
    .A2(_01851_),
    .A1(_01807_));
 sg13g2_xnor2_1 _07169_ (.Y(_01854_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .B(_01853_));
 sg13g2_xnor2_1 _07170_ (.Y(_01855_),
    .A(_01850_),
    .B(_01854_));
 sg13g2_xnor2_1 _07171_ (.Y(_01856_),
    .A(_01842_),
    .B(_01855_));
 sg13g2_xnor2_1 _07172_ (.Y(_01857_),
    .A(_01841_),
    .B(_01856_));
 sg13g2_and2_1 _07173_ (.A(_01836_),
    .B(_01857_),
    .X(_01858_));
 sg13g2_nor2_1 _07174_ (.A(_01836_),
    .B(_01857_),
    .Y(_01859_));
 sg13g2_nor2_1 _07175_ (.A(_01858_),
    .B(_01859_),
    .Y(_01860_));
 sg13g2_xnor2_1 _07176_ (.Y(_00020_),
    .A(_01833_),
    .B(_01860_));
 sg13g2_inv_1 _07177_ (.Y(_01861_),
    .A(_01859_));
 sg13g2_a21oi_1 _07178_ (.A1(_01833_),
    .A2(_01861_),
    .Y(_01862_),
    .B1(_01858_));
 sg13g2_a21oi_1 _07179_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A2(net121),
    .Y(_01863_),
    .B1(_01855_));
 sg13g2_nand2_1 _07180_ (.Y(_01864_),
    .A(_01853_),
    .B(_01850_));
 sg13g2_o21ai_1 _07181_ (.B1(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .Y(_01865_),
    .A1(_01853_),
    .A2(_01850_));
 sg13g2_and2_1 _07182_ (.A(_01864_),
    .B(_01865_),
    .X(_01866_));
 sg13g2_nand2_1 _07183_ (.Y(_01867_),
    .A(_01765_),
    .B(net121));
 sg13g2_inv_1 _07184_ (.Y(_01868_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[6] ));
 sg13g2_or2_1 _07185_ (.X(_01869_),
    .B(net132),
    .A(_01868_));
 sg13g2_buf_2 _07186_ (.A(_01869_),
    .X(_01870_));
 sg13g2_o21ai_1 _07187_ (.B1(_01810_),
    .Y(_01871_),
    .A1(_01669_),
    .A2(_01671_));
 sg13g2_buf_1 _07188_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .X(_01872_));
 sg13g2_nand3_1 _07189_ (.B(_01872_),
    .C(net153),
    .A(net219),
    .Y(_01873_));
 sg13g2_buf_2 _07190_ (.A(_01873_),
    .X(_01874_));
 sg13g2_xnor2_1 _07191_ (.Y(_01875_),
    .A(_01871_),
    .B(_01874_));
 sg13g2_xnor2_1 _07192_ (.Y(_01876_),
    .A(_01870_),
    .B(_01875_));
 sg13g2_o21ai_1 _07193_ (.B1(_01844_),
    .Y(_01877_),
    .A1(_01846_),
    .A2(_01848_));
 sg13g2_buf_1 _07194_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[7] ),
    .X(_01878_));
 sg13g2_a21oi_1 _07195_ (.A1(_01846_),
    .A2(_01848_),
    .Y(_01879_),
    .B1(_01878_));
 sg13g2_and2_1 _07196_ (.A(_01878_),
    .B(_01844_),
    .X(_01880_));
 sg13g2_or2_1 _07197_ (.X(_01881_),
    .B(_01848_),
    .A(_01846_));
 sg13g2_and3_1 _07198_ (.X(_01882_),
    .A(_01878_),
    .B(_01846_),
    .C(_01848_));
 sg13g2_a221oi_1 _07199_ (.B2(_01881_),
    .C1(_01882_),
    .B1(_01880_),
    .A1(_01877_),
    .Y(_01883_),
    .A2(_01879_));
 sg13g2_xor2_1 _07200_ (.B(_01883_),
    .A(_01876_),
    .X(_01884_));
 sg13g2_xor2_1 _07201_ (.B(_01884_),
    .A(_01867_),
    .X(_01885_));
 sg13g2_xnor2_1 _07202_ (.Y(_01886_),
    .A(_01866_),
    .B(_01885_));
 sg13g2_nor2b_1 _07203_ (.A(_01842_),
    .B_N(_01855_),
    .Y(_01887_));
 sg13g2_nor2_1 _07204_ (.A(_01841_),
    .B(_01887_),
    .Y(_01888_));
 sg13g2_nor3_1 _07205_ (.A(_01863_),
    .B(_01886_),
    .C(_01888_),
    .Y(_01889_));
 sg13g2_o21ai_1 _07206_ (.B1(_01886_),
    .Y(_01890_),
    .A1(_01863_),
    .A2(_01888_));
 sg13g2_nand2b_1 _07207_ (.Y(_01891_),
    .B(_01890_),
    .A_N(_01889_));
 sg13g2_xnor2_1 _07208_ (.Y(_00021_),
    .A(_01862_),
    .B(_01891_));
 sg13g2_nand2_1 _07209_ (.Y(_01892_),
    .A(_01836_),
    .B(_01857_));
 sg13g2_nand3_1 _07210_ (.B(_01892_),
    .C(_01890_),
    .A(_01828_),
    .Y(_01893_));
 sg13g2_a21oi_1 _07211_ (.A1(_01859_),
    .A2(_01890_),
    .Y(_01894_),
    .B1(_01889_));
 sg13g2_o21ai_1 _07212_ (.B1(_01894_),
    .Y(_01895_),
    .A1(_01832_),
    .A2(_01893_));
 sg13g2_nor2b_1 _07213_ (.A(_01884_),
    .B_N(_01867_),
    .Y(_01896_));
 sg13g2_nand2b_1 _07214_ (.Y(_01897_),
    .B(_01884_),
    .A_N(_01867_));
 sg13g2_o21ai_1 _07215_ (.B1(_01897_),
    .Y(_01898_),
    .A1(_01866_),
    .A2(_01896_));
 sg13g2_buf_2 _07216_ (.A(_01898_),
    .X(_01899_));
 sg13g2_nand2_1 _07217_ (.Y(_01900_),
    .A(_01846_),
    .B(_01848_));
 sg13g2_nand2_1 _07218_ (.Y(_01901_),
    .A(_01877_),
    .B(_01900_));
 sg13g2_nand2_1 _07219_ (.Y(_01902_),
    .A(_01876_),
    .B(_01901_));
 sg13g2_nor2_1 _07220_ (.A(_01876_),
    .B(_01901_),
    .Y(_01903_));
 sg13g2_a21oi_2 _07221_ (.B1(_01903_),
    .Y(_01904_),
    .A2(_01902_),
    .A1(_01878_));
 sg13g2_inv_1 _07222_ (.Y(_01905_),
    .A(_01872_));
 sg13g2_nor2_1 _07223_ (.A(_01905_),
    .B(_01725_),
    .Y(_01906_));
 sg13g2_buf_1 _07224_ (.A(_01906_),
    .X(_01907_));
 sg13g2_a21oi_1 _07225_ (.A1(_00793_),
    .A2(_00819_),
    .Y(_01908_),
    .B1(_01843_));
 sg13g2_buf_2 _07226_ (.A(_01908_),
    .X(_01909_));
 sg13g2_buf_1 _07227_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .X(_01910_));
 sg13g2_and3_1 _07228_ (.X(_01911_),
    .A(net219),
    .B(_01910_),
    .C(_01136_));
 sg13g2_buf_1 _07229_ (.A(_01911_),
    .X(_01912_));
 sg13g2_xnor2_1 _07230_ (.Y(_01913_),
    .A(_01909_),
    .B(_01912_));
 sg13g2_xnor2_1 _07231_ (.Y(_01914_),
    .A(_01907_),
    .B(_01913_));
 sg13g2_or2_1 _07232_ (.X(_01915_),
    .B(_01874_),
    .A(_01870_));
 sg13g2_buf_1 _07233_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .X(_01916_));
 sg13g2_and2_1 _07234_ (.A(_01916_),
    .B(_01871_),
    .X(_01917_));
 sg13g2_a21oi_1 _07235_ (.A1(_01870_),
    .A2(_01874_),
    .Y(_01918_),
    .B1(_01916_));
 sg13g2_o21ai_1 _07236_ (.B1(_01871_),
    .Y(_01919_),
    .A1(_01870_),
    .A2(_01874_));
 sg13g2_and3_1 _07237_ (.X(_01920_),
    .A(_01916_),
    .B(_01870_),
    .C(_01874_));
 sg13g2_a221oi_1 _07238_ (.B2(_01919_),
    .C1(_01920_),
    .B1(_01918_),
    .A1(_01915_),
    .Y(_01921_),
    .A2(_01917_));
 sg13g2_xnor2_1 _07239_ (.Y(_01922_),
    .A(_01914_),
    .B(_01921_));
 sg13g2_nand2_1 _07240_ (.Y(_01923_),
    .A(_01808_),
    .B(net121));
 sg13g2_xnor2_1 _07241_ (.Y(_01924_),
    .A(_01922_),
    .B(_01923_));
 sg13g2_xnor2_1 _07242_ (.Y(_01925_),
    .A(_01904_),
    .B(_01924_));
 sg13g2_xnor2_1 _07243_ (.Y(_01926_),
    .A(_01899_),
    .B(_01925_));
 sg13g2_xnor2_1 _07244_ (.Y(_00022_),
    .A(_01895_),
    .B(_01926_));
 sg13g2_nand2_1 _07245_ (.Y(_01927_),
    .A(_01870_),
    .B(_01874_));
 sg13g2_a22oi_1 _07246_ (.Y(_01928_),
    .B1(_01914_),
    .B2(_01916_),
    .A2(_01919_),
    .A1(_01927_));
 sg13g2_nor2_1 _07247_ (.A(_01916_),
    .B(_01914_),
    .Y(_01929_));
 sg13g2_nor2_1 _07248_ (.A(_01928_),
    .B(_01929_),
    .Y(_01930_));
 sg13g2_nand2_1 _07249_ (.Y(_01931_),
    .A(_01872_),
    .B(_01666_));
 sg13g2_inv_1 _07250_ (.Y(_01932_),
    .A(_01910_));
 sg13g2_nor2_1 _07251_ (.A(_01932_),
    .B(_01814_),
    .Y(_01933_));
 sg13g2_buf_1 _07252_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .X(_01934_));
 sg13g2_and3_1 _07253_ (.X(_01935_),
    .A(_01220_),
    .B(_01934_),
    .C(_01136_));
 sg13g2_buf_1 _07254_ (.A(_01935_),
    .X(_01936_));
 sg13g2_xnor2_1 _07255_ (.Y(_01937_),
    .A(_01933_),
    .B(_01936_));
 sg13g2_xor2_1 _07256_ (.B(_01937_),
    .A(_01931_),
    .X(_01938_));
 sg13g2_o21ai_1 _07257_ (.B1(_01912_),
    .Y(_01939_),
    .A1(_01907_),
    .A2(_01909_));
 sg13g2_buf_1 _07258_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .X(_01940_));
 sg13g2_a21oi_1 _07259_ (.A1(_01907_),
    .A2(_01909_),
    .Y(_01941_),
    .B1(_01940_));
 sg13g2_and2_1 _07260_ (.A(_01940_),
    .B(_01912_),
    .X(_01942_));
 sg13g2_or2_1 _07261_ (.X(_01943_),
    .B(_01909_),
    .A(_01907_));
 sg13g2_and3_1 _07262_ (.X(_01944_),
    .A(_01940_),
    .B(_01907_),
    .C(_01909_));
 sg13g2_a221oi_1 _07263_ (.B2(_01943_),
    .C1(_01944_),
    .B1(_01942_),
    .A1(_01939_),
    .Y(_01945_),
    .A2(_01941_));
 sg13g2_xnor2_1 _07264_ (.Y(_01946_),
    .A(_01938_),
    .B(_01945_));
 sg13g2_nor3_1 _07265_ (.A(net263),
    .B(_01868_),
    .C(net154),
    .Y(_01947_));
 sg13g2_xor2_1 _07266_ (.B(_01947_),
    .A(_01946_),
    .X(_01948_));
 sg13g2_xor2_1 _07267_ (.B(_01948_),
    .A(_01930_),
    .X(_01949_));
 sg13g2_nor2_1 _07268_ (.A(_01832_),
    .B(_01893_),
    .Y(_01950_));
 sg13g2_nor2b_1 _07269_ (.A(_01950_),
    .B_N(_01894_),
    .Y(_01951_));
 sg13g2_nand3_1 _07270_ (.B(net121),
    .C(_01922_),
    .A(_01808_),
    .Y(_01952_));
 sg13g2_nor2b_2 _07271_ (.A(_01922_),
    .B_N(_01923_),
    .Y(_01953_));
 sg13g2_a21oi_2 _07272_ (.B1(_01953_),
    .Y(_01954_),
    .A2(_01952_),
    .A1(_01904_));
 sg13g2_nand2_1 _07273_ (.Y(_01955_),
    .A(_01904_),
    .B(_01953_));
 sg13g2_o21ai_1 _07274_ (.B1(_01955_),
    .Y(_01956_),
    .A1(_01899_),
    .A2(_01954_));
 sg13g2_a21o_1 _07275_ (.A2(_01902_),
    .A1(_01878_),
    .B1(_01903_),
    .X(_01957_));
 sg13g2_buf_1 _07276_ (.A(net121),
    .X(_01958_));
 sg13g2_and3_1 _07277_ (.X(_01959_),
    .A(_01808_),
    .B(_01958_),
    .C(_01922_));
 sg13g2_buf_1 _07278_ (.A(_01959_),
    .X(_01960_));
 sg13g2_a22oi_1 _07279_ (.Y(_01961_),
    .B1(_01954_),
    .B2(_01899_),
    .A2(_01960_),
    .A1(_01957_));
 sg13g2_nand2_1 _07280_ (.Y(_01962_),
    .A(_01899_),
    .B(_01957_));
 sg13g2_inv_1 _07281_ (.Y(_01963_),
    .A(_01962_));
 sg13g2_nor2_1 _07282_ (.A(_01899_),
    .B(_01957_),
    .Y(_01964_));
 sg13g2_a22oi_1 _07283_ (.Y(_01965_),
    .B1(_01964_),
    .B2(_01953_),
    .A2(_01963_),
    .A1(_01960_));
 sg13g2_o21ai_1 _07284_ (.B1(_01965_),
    .Y(_01966_),
    .A1(_01951_),
    .A2(_01961_));
 sg13g2_a21oi_1 _07285_ (.A1(_01951_),
    .A2(_01956_),
    .Y(_01967_),
    .B1(_01966_));
 sg13g2_xnor2_1 _07286_ (.Y(_00023_),
    .A(_01949_),
    .B(_01967_));
 sg13g2_xnor2_1 _07287_ (.Y(_01968_),
    .A(_01930_),
    .B(_01948_));
 sg13g2_nand2_1 _07288_ (.Y(_01969_),
    .A(_01949_),
    .B(_01962_));
 sg13g2_nor2_1 _07289_ (.A(_01949_),
    .B(_01964_),
    .Y(_01970_));
 sg13g2_a21oi_1 _07290_ (.A1(_01895_),
    .A2(_01969_),
    .Y(_01971_),
    .B1(_01970_));
 sg13g2_o21ai_1 _07291_ (.B1(_01962_),
    .Y(_01972_),
    .A1(_01951_),
    .A2(_01964_));
 sg13g2_o21ai_1 _07292_ (.B1(_01972_),
    .Y(_01973_),
    .A1(_01960_),
    .A2(_01968_));
 sg13g2_o21ai_1 _07293_ (.B1(_01973_),
    .Y(_01974_),
    .A1(_01953_),
    .A2(_01971_));
 sg13g2_a21o_1 _07294_ (.A2(_01968_),
    .A1(_01960_),
    .B1(_01974_),
    .X(_01975_));
 sg13g2_nor2_1 _07295_ (.A(_01933_),
    .B(_01936_),
    .Y(_01976_));
 sg13g2_a22oi_1 _07296_ (.Y(_01977_),
    .B1(_01933_),
    .B2(_01936_),
    .A2(_01666_),
    .A1(_01872_));
 sg13g2_or3_1 _07297_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .B(_01976_),
    .C(_01977_),
    .X(_01978_));
 sg13g2_o21ai_1 _07298_ (.B1(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .Y(_01979_),
    .A1(_01976_),
    .A2(_01977_));
 sg13g2_nand2_1 _07299_ (.Y(_01980_),
    .A(_01910_),
    .B(_01666_));
 sg13g2_inv_1 _07300_ (.Y(_01981_),
    .A(_01934_));
 sg13g2_nor2_1 _07301_ (.A(_01981_),
    .B(net132),
    .Y(_01982_));
 sg13g2_buf_1 _07302_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .X(_01983_));
 sg13g2_nand3_1 _07303_ (.B(net294),
    .C(net133),
    .A(_01220_),
    .Y(_01984_));
 sg13g2_xor2_1 _07304_ (.B(_01984_),
    .A(_01982_),
    .X(_01985_));
 sg13g2_xnor2_1 _07305_ (.Y(_01986_),
    .A(_01980_),
    .B(_01985_));
 sg13g2_a21oi_1 _07306_ (.A1(_01978_),
    .A2(_01979_),
    .Y(_01987_),
    .B1(_01986_));
 sg13g2_and3_1 _07307_ (.X(_01988_),
    .A(_01986_),
    .B(_01978_),
    .C(_01979_));
 sg13g2_buf_1 _07308_ (.A(_01988_),
    .X(_01989_));
 sg13g2_nand2_1 _07309_ (.Y(_01990_),
    .A(_01872_),
    .B(_01756_));
 sg13g2_o21ai_1 _07310_ (.B1(_01990_),
    .Y(_01991_),
    .A1(_01987_),
    .A2(_01989_));
 sg13g2_or3_1 _07311_ (.A(_01990_),
    .B(_01987_),
    .C(_01989_),
    .X(_01992_));
 sg13g2_nand2_1 _07312_ (.Y(_01993_),
    .A(_01940_),
    .B(_01938_));
 sg13g2_nand2_1 _07313_ (.Y(_01994_),
    .A(_01907_),
    .B(_01909_));
 sg13g2_nand2_1 _07314_ (.Y(_01995_),
    .A(_01939_),
    .B(_01994_));
 sg13g2_o21ai_1 _07315_ (.B1(_01995_),
    .Y(_01996_),
    .A1(_01940_),
    .A2(_01938_));
 sg13g2_nand2_1 _07316_ (.Y(_01997_),
    .A(_01993_),
    .B(_01996_));
 sg13g2_a21o_1 _07317_ (.A2(_01992_),
    .A1(_01991_),
    .B1(_01997_),
    .X(_01998_));
 sg13g2_nand3_1 _07318_ (.B(_01991_),
    .C(_01992_),
    .A(_01997_),
    .Y(_01999_));
 sg13g2_and2_1 _07319_ (.A(_01998_),
    .B(_01999_),
    .X(_02000_));
 sg13g2_o21ai_1 _07320_ (.B1(_01946_),
    .Y(_02001_),
    .A1(_01928_),
    .A2(_01929_));
 sg13g2_nor3_1 _07321_ (.A(_01928_),
    .B(_01929_),
    .C(_01946_),
    .Y(_02002_));
 sg13g2_a21o_1 _07322_ (.A2(_02001_),
    .A1(_01947_),
    .B1(_02002_),
    .X(_02003_));
 sg13g2_buf_1 _07323_ (.A(_02003_),
    .X(_02004_));
 sg13g2_xnor2_1 _07324_ (.Y(_02005_),
    .A(_02000_),
    .B(_02004_));
 sg13g2_xnor2_1 _07325_ (.Y(_00024_),
    .A(_01975_),
    .B(_02005_));
 sg13g2_nor2_1 _07326_ (.A(_01968_),
    .B(_01954_),
    .Y(_02006_));
 sg13g2_nor2_1 _07327_ (.A(_01899_),
    .B(_01925_),
    .Y(_02007_));
 sg13g2_a21oi_1 _07328_ (.A1(_01998_),
    .A2(_01999_),
    .Y(_02008_),
    .B1(_02004_));
 sg13g2_or2_1 _07329_ (.X(_02009_),
    .B(_02008_),
    .A(_02007_));
 sg13g2_nor3_1 _07330_ (.A(_01951_),
    .B(_02006_),
    .C(_02009_),
    .Y(_02010_));
 sg13g2_nand2_1 _07331_ (.Y(_02011_),
    .A(_02000_),
    .B(_02004_));
 sg13g2_a22oi_1 _07332_ (.Y(_02012_),
    .B1(_01968_),
    .B2(_01954_),
    .A2(_01925_),
    .A1(_01899_));
 sg13g2_or3_1 _07333_ (.A(_02006_),
    .B(_02008_),
    .C(_02012_),
    .X(_02013_));
 sg13g2_nand3b_1 _07334_ (.B(_02011_),
    .C(_02013_),
    .Y(_02014_),
    .A_N(_02010_));
 sg13g2_nor3_1 _07335_ (.A(_01990_),
    .B(_01987_),
    .C(_01989_),
    .Y(_02015_));
 sg13g2_o21ai_1 _07336_ (.B1(_01991_),
    .Y(_02016_),
    .A1(_01997_),
    .A2(_02015_));
 sg13g2_buf_1 _07337_ (.A(_02016_),
    .X(_02017_));
 sg13g2_or2_1 _07338_ (.X(_02018_),
    .B(_01977_),
    .A(_01976_));
 sg13g2_nand2b_1 _07339_ (.Y(_02019_),
    .B(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .A_N(_01986_));
 sg13g2_nor2b_1 _07340_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .B_N(_01986_),
    .Y(_02020_));
 sg13g2_a21oi_2 _07341_ (.B1(_02020_),
    .Y(_02021_),
    .A2(_02019_),
    .A1(_02018_));
 sg13g2_nand2_1 _07342_ (.Y(_02022_),
    .A(net294),
    .B(_01681_));
 sg13g2_nand2_1 _07343_ (.Y(_02023_),
    .A(_01934_),
    .B(_01666_));
 sg13g2_buf_1 _07344_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .X(_02024_));
 sg13g2_nand2_1 _07345_ (.Y(_02025_),
    .A(net293),
    .B(_01677_));
 sg13g2_xnor2_1 _07346_ (.Y(_02026_),
    .A(_02023_),
    .B(_02025_));
 sg13g2_xnor2_1 _07347_ (.Y(_02027_),
    .A(_02022_),
    .B(_02026_));
 sg13g2_nand3_1 _07348_ (.B(_01677_),
    .C(_01982_),
    .A(net294),
    .Y(_02028_));
 sg13g2_nor2b_1 _07349_ (.A(_01982_),
    .B_N(_01984_),
    .Y(_02029_));
 sg13g2_a21o_1 _07350_ (.A2(_02028_),
    .A1(_01980_),
    .B1(_02029_),
    .X(_02030_));
 sg13g2_buf_1 _07351_ (.A(_02030_),
    .X(_02031_));
 sg13g2_xor2_1 _07352_ (.B(_02031_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .X(_02032_));
 sg13g2_xnor2_1 _07353_ (.Y(_02033_),
    .A(_02027_),
    .B(_02032_));
 sg13g2_nand2_1 _07354_ (.Y(_02034_),
    .A(_01910_),
    .B(_01756_));
 sg13g2_xor2_1 _07355_ (.B(_02034_),
    .A(_02033_),
    .X(_02035_));
 sg13g2_xnor2_1 _07356_ (.Y(_02036_),
    .A(_02021_),
    .B(_02035_));
 sg13g2_xnor2_1 _07357_ (.Y(_02037_),
    .A(_02017_),
    .B(_02036_));
 sg13g2_xnor2_1 _07358_ (.Y(_00025_),
    .A(_02014_),
    .B(_02037_));
 sg13g2_nand2_1 _07359_ (.Y(_02038_),
    .A(_02031_),
    .B(_02027_));
 sg13g2_nor2_1 _07360_ (.A(_02031_),
    .B(_02027_),
    .Y(_02039_));
 sg13g2_a21o_1 _07361_ (.A2(_02038_),
    .A1(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .B1(_02039_),
    .X(_02040_));
 sg13g2_buf_1 _07362_ (.A(_02040_),
    .X(_02041_));
 sg13g2_nor3_1 _07363_ (.A(_01174_),
    .B(_01981_),
    .C(_00856_),
    .Y(_02042_));
 sg13g2_nand2_1 _07364_ (.Y(_02043_),
    .A(net293),
    .B(_01681_));
 sg13g2_nand2_1 _07365_ (.Y(_02044_),
    .A(net294),
    .B(_01666_));
 sg13g2_buf_2 _07366_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .X(_02045_));
 sg13g2_buf_1 _07367_ (.A(_01677_),
    .X(_02046_));
 sg13g2_nand2_1 _07368_ (.Y(_02047_),
    .A(_02045_),
    .B(net120));
 sg13g2_xnor2_1 _07369_ (.Y(_02048_),
    .A(_02044_),
    .B(_02047_));
 sg13g2_xnor2_1 _07370_ (.Y(_02049_),
    .A(_02043_),
    .B(_02048_));
 sg13g2_a22oi_1 _07371_ (.Y(_02050_),
    .B1(_01681_),
    .B2(net294),
    .A2(net120),
    .A1(net293));
 sg13g2_nand4_1 _07372_ (.B(net293),
    .C(net120),
    .A(net294),
    .Y(_02051_),
    .D(_01681_));
 sg13g2_o21ai_1 _07373_ (.B1(_02051_),
    .Y(_02052_),
    .A1(_02023_),
    .A2(_02050_));
 sg13g2_xnor2_1 _07374_ (.Y(_02053_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[12] ),
    .B(_02052_));
 sg13g2_xnor2_1 _07375_ (.Y(_02054_),
    .A(_02049_),
    .B(_02053_));
 sg13g2_xor2_1 _07376_ (.B(_02054_),
    .A(_02042_),
    .X(_02055_));
 sg13g2_xnor2_1 _07377_ (.Y(_02056_),
    .A(_02041_),
    .B(_02055_));
 sg13g2_nor2b_1 _07378_ (.A(_02021_),
    .B_N(_02033_),
    .Y(_02057_));
 sg13g2_nand2b_1 _07379_ (.Y(_02058_),
    .B(_02021_),
    .A_N(_02033_));
 sg13g2_o21ai_1 _07380_ (.B1(_02058_),
    .Y(_02059_),
    .A1(_02034_),
    .A2(_02057_));
 sg13g2_nor2_1 _07381_ (.A(_02056_),
    .B(_02059_),
    .Y(_02060_));
 sg13g2_nand2_1 _07382_ (.Y(_02061_),
    .A(_02056_),
    .B(_02059_));
 sg13g2_buf_1 _07383_ (.A(_02061_),
    .X(_02062_));
 sg13g2_nor2b_1 _07384_ (.A(_02060_),
    .B_N(_02062_),
    .Y(_02063_));
 sg13g2_nand2_1 _07385_ (.Y(_02064_),
    .A(_02017_),
    .B(_02036_));
 sg13g2_nor2_1 _07386_ (.A(_02017_),
    .B(_02036_),
    .Y(_02065_));
 sg13g2_a21oi_1 _07387_ (.A1(_02014_),
    .A2(_02064_),
    .Y(_02066_),
    .B1(_02065_));
 sg13g2_xnor2_1 _07388_ (.Y(_00026_),
    .A(_02063_),
    .B(_02066_));
 sg13g2_inv_1 _07389_ (.Y(_02067_),
    .A(_02060_));
 sg13g2_and2_1 _07390_ (.A(_02017_),
    .B(_02036_),
    .X(_02068_));
 sg13g2_nor4_1 _07391_ (.A(_02006_),
    .B(_02009_),
    .C(_02060_),
    .D(_02068_),
    .Y(_02069_));
 sg13g2_a221oi_1 _07392_ (.B2(_02036_),
    .C1(_02060_),
    .B1(_02017_),
    .A1(_02011_),
    .Y(_02070_),
    .A2(_02013_));
 sg13g2_a221oi_1 _07393_ (.B2(_01895_),
    .C1(_02070_),
    .B1(_02069_),
    .A1(_02067_),
    .Y(_02071_),
    .A2(_02065_));
 sg13g2_buf_1 _07394_ (.A(_02071_),
    .X(_02072_));
 sg13g2_nand2_1 _07395_ (.Y(_02073_),
    .A(_02062_),
    .B(_02072_));
 sg13g2_nand2b_1 _07396_ (.Y(_02074_),
    .B(_02054_),
    .A_N(_02041_));
 sg13g2_nor2b_1 _07397_ (.A(_02054_),
    .B_N(_02041_),
    .Y(_02075_));
 sg13g2_a21oi_1 _07398_ (.A1(_02042_),
    .A2(_02074_),
    .Y(_02076_),
    .B1(_02075_));
 sg13g2_buf_1 _07399_ (.A(_02076_),
    .X(_02077_));
 sg13g2_nand2_1 _07400_ (.Y(_02078_),
    .A(_02043_),
    .B(_02047_));
 sg13g2_o21ai_1 _07401_ (.B1(_02044_),
    .Y(_02079_),
    .A1(_02043_),
    .A2(_02047_));
 sg13g2_nand2_1 _07402_ (.Y(_02080_),
    .A(_02078_),
    .B(_02079_));
 sg13g2_buf_1 _07403_ (.A(_01666_),
    .X(_02081_));
 sg13g2_and2_1 _07404_ (.A(net293),
    .B(net119),
    .X(_02082_));
 sg13g2_buf_1 _07405_ (.A(_01681_),
    .X(_02083_));
 sg13g2_nand2_1 _07406_ (.Y(_02084_),
    .A(_02045_),
    .B(net118));
 sg13g2_buf_1 _07407_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .X(_02085_));
 sg13g2_nand2_1 _07408_ (.Y(_02086_),
    .A(net292),
    .B(net120));
 sg13g2_xor2_1 _07409_ (.B(_02086_),
    .A(_02084_),
    .X(_02087_));
 sg13g2_xnor2_1 _07410_ (.Y(_02088_),
    .A(_02082_),
    .B(_02087_));
 sg13g2_xnor2_1 _07411_ (.Y(_02089_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[13] ),
    .B(_02088_));
 sg13g2_xnor2_1 _07412_ (.Y(_02090_),
    .A(_02080_),
    .B(_02089_));
 sg13g2_buf_2 _07413_ (.A(_02090_),
    .X(_02091_));
 sg13g2_nand2_1 _07414_ (.Y(_02092_),
    .A(_02023_),
    .B(_02051_));
 sg13g2_nand2b_1 _07415_ (.Y(_02093_),
    .B(_02092_),
    .A_N(_02050_));
 sg13g2_nand2_1 _07416_ (.Y(_02094_),
    .A(_02093_),
    .B(_02049_));
 sg13g2_nor2_1 _07417_ (.A(_02093_),
    .B(_02049_),
    .Y(_02095_));
 sg13g2_a21oi_1 _07418_ (.A1(\i_tinyqv.cpu.i_core.multiplier.accum[12] ),
    .A2(_02094_),
    .Y(_02096_),
    .B1(_02095_));
 sg13g2_buf_2 _07419_ (.A(_02096_),
    .X(_02097_));
 sg13g2_nand2_2 _07420_ (.Y(_02098_),
    .A(net294),
    .B(net109));
 sg13g2_xor2_1 _07421_ (.B(_02098_),
    .A(_02097_),
    .X(_02099_));
 sg13g2_xnor2_1 _07422_ (.Y(_02100_),
    .A(_02091_),
    .B(_02099_));
 sg13g2_xnor2_1 _07423_ (.Y(_02101_),
    .A(_02077_),
    .B(_02100_));
 sg13g2_xnor2_1 _07424_ (.Y(_00027_),
    .A(_02073_),
    .B(_02101_));
 sg13g2_inv_1 _07425_ (.Y(_02102_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[13] ));
 sg13g2_a21o_1 _07426_ (.A2(_02088_),
    .A1(_02080_),
    .B1(_02102_),
    .X(_02103_));
 sg13g2_o21ai_1 _07427_ (.B1(_02103_),
    .Y(_02104_),
    .A1(_02080_),
    .A2(_02088_));
 sg13g2_buf_1 _07428_ (.A(_02104_),
    .X(_02105_));
 sg13g2_nand2_2 _07429_ (.Y(_02106_),
    .A(net292),
    .B(net118));
 sg13g2_nand2_1 _07430_ (.Y(_02107_),
    .A(_02045_),
    .B(_01666_));
 sg13g2_buf_1 _07431_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .X(_02108_));
 sg13g2_nand2_1 _07432_ (.Y(_02109_),
    .A(_02108_),
    .B(net120));
 sg13g2_xnor2_1 _07433_ (.Y(_02110_),
    .A(_02107_),
    .B(_02109_));
 sg13g2_xnor2_1 _07434_ (.Y(_02111_),
    .A(_02106_),
    .B(_02110_));
 sg13g2_nand2_1 _07435_ (.Y(_02112_),
    .A(_02084_),
    .B(_02086_));
 sg13g2_nor2_1 _07436_ (.A(_02084_),
    .B(_02086_),
    .Y(_02113_));
 sg13g2_a21oi_1 _07437_ (.A1(_02082_),
    .A2(_02112_),
    .Y(_02114_),
    .B1(_02113_));
 sg13g2_xor2_1 _07438_ (.B(_02114_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[14] ),
    .X(_02115_));
 sg13g2_xnor2_1 _07439_ (.Y(_02116_),
    .A(_02111_),
    .B(_02115_));
 sg13g2_nand2_1 _07440_ (.Y(_02117_),
    .A(net293),
    .B(_01958_));
 sg13g2_xor2_1 _07441_ (.B(_02117_),
    .A(_02116_),
    .X(_02118_));
 sg13g2_xnor2_1 _07442_ (.Y(_02119_),
    .A(_02105_),
    .B(_02118_));
 sg13g2_a21oi_1 _07443_ (.A1(_02062_),
    .A2(_02072_),
    .Y(_02120_),
    .B1(_02098_));
 sg13g2_nor2b_1 _07444_ (.A(_02097_),
    .B_N(_02091_),
    .Y(_02121_));
 sg13g2_nand3_1 _07445_ (.B(_02072_),
    .C(_02098_),
    .A(_02062_),
    .Y(_02122_));
 sg13g2_o21ai_1 _07446_ (.B1(_02122_),
    .Y(_02123_),
    .A1(_02091_),
    .A2(_02120_));
 sg13g2_nand2_1 _07447_ (.Y(_02124_),
    .A(_02091_),
    .B(_02120_));
 sg13g2_o21ai_1 _07448_ (.B1(_02124_),
    .Y(_02125_),
    .A1(_02097_),
    .A2(_02123_));
 sg13g2_or2_1 _07449_ (.X(_02126_),
    .B(_02125_),
    .A(_02077_));
 sg13g2_nor2_1 _07450_ (.A(_02091_),
    .B(_02122_),
    .Y(_02127_));
 sg13g2_a21oi_1 _07451_ (.A1(_02097_),
    .A2(_02123_),
    .Y(_02128_),
    .B1(_02127_));
 sg13g2_nand2_1 _07452_ (.Y(_02129_),
    .A(_02077_),
    .B(_02128_));
 sg13g2_nor2b_1 _07453_ (.A(_02091_),
    .B_N(_02097_),
    .Y(_02130_));
 sg13g2_nor2b_1 _07454_ (.A(_02122_),
    .B_N(_02130_),
    .Y(_02131_));
 sg13g2_a221oi_1 _07455_ (.B2(_02129_),
    .C1(_02131_),
    .B1(_02126_),
    .A1(_02120_),
    .Y(_02132_),
    .A2(_02121_));
 sg13g2_xnor2_1 _07456_ (.Y(_00017_),
    .A(_02119_),
    .B(_02132_));
 sg13g2_and2_1 _07457_ (.A(_02062_),
    .B(_02119_),
    .X(_02133_));
 sg13g2_nand2_1 _07458_ (.Y(_02134_),
    .A(_02077_),
    .B(_02097_));
 sg13g2_nor2b_1 _07459_ (.A(_02134_),
    .B_N(_02062_),
    .Y(_02135_));
 sg13g2_o21ai_1 _07460_ (.B1(_02072_),
    .Y(_02136_),
    .A1(_02133_),
    .A2(_02135_));
 sg13g2_nand2b_1 _07461_ (.Y(_02137_),
    .B(_02098_),
    .A_N(_02091_));
 sg13g2_o21ai_1 _07462_ (.B1(_02119_),
    .Y(_02138_),
    .A1(_02077_),
    .A2(_02097_));
 sg13g2_and2_1 _07463_ (.A(_02137_),
    .B(_02138_),
    .X(_02139_));
 sg13g2_nand2b_1 _07464_ (.Y(_02140_),
    .B(_02091_),
    .A_N(_02098_));
 sg13g2_o21ai_1 _07465_ (.B1(_02062_),
    .Y(_02141_),
    .A1(_02119_),
    .A2(_02140_));
 sg13g2_nor2b_1 _07466_ (.A(_02141_),
    .B_N(_02097_),
    .Y(_02142_));
 sg13g2_nor2b_1 _07467_ (.A(_02141_),
    .B_N(_02077_),
    .Y(_02143_));
 sg13g2_o21ai_1 _07468_ (.B1(_02072_),
    .Y(_02144_),
    .A1(_02142_),
    .A2(_02143_));
 sg13g2_xor2_1 _07469_ (.B(_02118_),
    .A(_02105_),
    .X(_02145_));
 sg13g2_inv_1 _07470_ (.Y(_02146_),
    .A(_02140_));
 sg13g2_a21oi_1 _07471_ (.A1(_02145_),
    .A2(_02146_),
    .Y(_02147_),
    .B1(_02134_));
 sg13g2_a21oi_1 _07472_ (.A1(_02119_),
    .A2(_02140_),
    .Y(_02148_),
    .B1(_02147_));
 sg13g2_a22oi_1 _07473_ (.Y(_02149_),
    .B1(_02144_),
    .B2(_02148_),
    .A2(_02139_),
    .A1(_02136_));
 sg13g2_buf_1 _07474_ (.A(_02149_),
    .X(_02150_));
 sg13g2_inv_1 _07475_ (.Y(_02151_),
    .A(_02116_));
 sg13g2_nor2_1 _07476_ (.A(_02105_),
    .B(_02151_),
    .Y(_02152_));
 sg13g2_nor2_1 _07477_ (.A(_02117_),
    .B(_02152_),
    .Y(_02153_));
 sg13g2_a21oi_1 _07478_ (.A1(_02105_),
    .A2(_02151_),
    .Y(_02154_),
    .B1(_02153_));
 sg13g2_buf_1 _07479_ (.A(_02154_),
    .X(_02155_));
 sg13g2_nor2_1 _07480_ (.A(_02114_),
    .B(_02111_),
    .Y(_02156_));
 sg13g2_nor2_1 _07481_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[14] ),
    .B(_02156_),
    .Y(_02157_));
 sg13g2_a21oi_1 _07482_ (.A1(_02114_),
    .A2(_02111_),
    .Y(_02158_),
    .B1(_02157_));
 sg13g2_buf_2 _07483_ (.A(_02158_),
    .X(_02159_));
 sg13g2_nand2_1 _07484_ (.Y(_02160_),
    .A(_02108_),
    .B(net118));
 sg13g2_nand2_1 _07485_ (.Y(_02161_),
    .A(net292),
    .B(net119));
 sg13g2_buf_1 _07486_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .X(_02162_));
 sg13g2_nand2_1 _07487_ (.Y(_02163_),
    .A(net291),
    .B(net120));
 sg13g2_xnor2_1 _07488_ (.Y(_02164_),
    .A(_02161_),
    .B(_02163_));
 sg13g2_xnor2_1 _07489_ (.Y(_02165_),
    .A(_02160_),
    .B(_02164_));
 sg13g2_nand2_1 _07490_ (.Y(_02166_),
    .A(_02106_),
    .B(_02109_));
 sg13g2_o21ai_1 _07491_ (.B1(_02107_),
    .Y(_02167_),
    .A1(_02106_),
    .A2(_02109_));
 sg13g2_nand2_1 _07492_ (.Y(_02168_),
    .A(_02166_),
    .B(_02167_));
 sg13g2_xnor2_1 _07493_ (.Y(_02169_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .B(_02168_));
 sg13g2_xnor2_1 _07494_ (.Y(_02170_),
    .A(_02165_),
    .B(_02169_));
 sg13g2_and3_1 _07495_ (.X(_02171_),
    .A(_02045_),
    .B(net109),
    .C(_02170_));
 sg13g2_buf_1 _07496_ (.A(_02171_),
    .X(_02172_));
 sg13g2_a21o_1 _07497_ (.A2(net109),
    .A1(_02045_),
    .B1(_02170_),
    .X(_02173_));
 sg13g2_buf_1 _07498_ (.A(_02173_),
    .X(_02174_));
 sg13g2_nand2b_1 _07499_ (.Y(_02175_),
    .B(_02174_),
    .A_N(_02172_));
 sg13g2_xnor2_1 _07500_ (.Y(_02176_),
    .A(_02159_),
    .B(_02175_));
 sg13g2_xnor2_1 _07501_ (.Y(_02177_),
    .A(_02155_),
    .B(_02176_));
 sg13g2_xnor2_1 _07502_ (.Y(_00018_),
    .A(_02150_),
    .B(_02177_));
 sg13g2_buf_1 _07503_ (.A(net211),
    .X(_02178_));
 sg13g2_inv_1 _07504_ (.Y(_02179_),
    .A(_01575_));
 sg13g2_nor3_2 _07505_ (.A(_02179_),
    .B(net296),
    .C(_01590_),
    .Y(_02180_));
 sg13g2_and2_1 _07506_ (.A(_01591_),
    .B(_02180_),
    .X(_02181_));
 sg13g2_buf_1 _07507_ (.A(_02181_),
    .X(_02182_));
 sg13g2_nor2b_1 _07508_ (.A(_01575_),
    .B_N(net296),
    .Y(_02183_));
 sg13g2_and2_1 _07509_ (.A(_01591_),
    .B(_02183_),
    .X(_02184_));
 sg13g2_buf_1 _07510_ (.A(_02184_),
    .X(_02185_));
 sg13g2_buf_1 _07511_ (.A(_02185_),
    .X(_02186_));
 sg13g2_and2_1 _07512_ (.A(\gpio_out_sel[4] ),
    .B(net167),
    .X(_02187_));
 sg13g2_a221oi_1 _07513_ (.B2(\i_spi.data[4] ),
    .C1(_02187_),
    .B1(net131),
    .A1(\i_uart_rx.recieved_data[4] ),
    .Y(_02188_),
    .A2(net150));
 sg13g2_nand2_1 _07514_ (.Y(_02189_),
    .A(_01578_),
    .B(_01589_));
 sg13g2_nor2_1 _07515_ (.A(net295),
    .B(_02189_),
    .Y(_02190_));
 sg13g2_and2_1 _07516_ (.A(_01577_),
    .B(_02190_),
    .X(_02191_));
 sg13g2_buf_1 _07517_ (.A(_02191_),
    .X(_02192_));
 sg13g2_buf_1 _07518_ (.A(_00964_),
    .X(_02193_));
 sg13g2_a221oi_1 _07519_ (.B2(_01257_),
    .C1(net207),
    .B1(_02192_),
    .A1(net32),
    .Y(_02194_),
    .A2(_01593_));
 sg13g2_buf_1 _07520_ (.A(\i_debug_uart_tx.fsm_state[1] ),
    .X(_02195_));
 sg13g2_buf_2 _07521_ (.A(\i_debug_uart_tx.fsm_state[2] ),
    .X(_02196_));
 sg13g2_nor2_1 _07522_ (.A(net290),
    .B(_02196_),
    .Y(_02197_));
 sg13g2_buf_2 _07523_ (.A(\i_debug_uart_tx.fsm_state[0] ),
    .X(_02198_));
 sg13g2_buf_2 _07524_ (.A(\i_debug_uart_tx.fsm_state[3] ),
    .X(_02199_));
 sg13g2_nor2_1 _07525_ (.A(_02198_),
    .B(_02199_),
    .Y(_02200_));
 sg13g2_nand2_1 _07526_ (.Y(_02201_),
    .A(_02197_),
    .B(_02200_));
 sg13g2_buf_1 _07527_ (.A(_02201_),
    .X(_02202_));
 sg13g2_nor2_1 _07528_ (.A(net295),
    .B(net209),
    .Y(_02203_));
 sg13g2_a21oi_1 _07529_ (.A1(net295),
    .A2(net206),
    .Y(_02204_),
    .B1(_02203_));
 sg13g2_or4_1 _07530_ (.A(_02179_),
    .B(net296),
    .C(_02189_),
    .D(_02204_),
    .X(_02205_));
 sg13g2_nand2_1 _07531_ (.Y(_02206_),
    .A(\gpio_out_sel[0] ),
    .B(_01622_));
 sg13g2_buf_1 _07532_ (.A(_00167_),
    .X(_02207_));
 sg13g2_nand2b_1 _07533_ (.Y(_02208_),
    .B(net296),
    .A_N(_02207_));
 sg13g2_nand2b_1 _07534_ (.Y(_02209_),
    .B(net2),
    .A_N(net296));
 sg13g2_a21oi_1 _07535_ (.A1(_02208_),
    .A2(_02209_),
    .Y(_02210_),
    .B1(_01575_));
 sg13g2_a22oi_1 _07536_ (.Y(_02211_),
    .B1(_02190_),
    .B2(_02210_),
    .A2(_02186_),
    .A1(\i_spi.data[0] ));
 sg13g2_and4_1 _07537_ (.A(net207),
    .B(_02205_),
    .C(_02206_),
    .D(_02211_),
    .X(_02212_));
 sg13g2_a22oi_1 _07538_ (.Y(_02213_),
    .B1(_02180_),
    .B2(\i_uart_rx.recieved_data[0] ),
    .A2(_01577_),
    .A1(net28));
 sg13g2_nand2b_1 _07539_ (.Y(_02214_),
    .B(_01591_),
    .A_N(_02213_));
 sg13g2_a22oi_1 _07540_ (.Y(_02215_),
    .B1(_02212_),
    .B2(_02214_),
    .A2(_02194_),
    .A1(_02188_));
 sg13g2_and2_1 _07541_ (.A(_01575_),
    .B(net296),
    .X(_02216_));
 sg13g2_nor2_1 _07542_ (.A(net295),
    .B(_02216_),
    .Y(_02217_));
 sg13g2_nor2b_1 _07543_ (.A(net296),
    .B_N(_01578_),
    .Y(_02218_));
 sg13g2_o21ai_1 _07544_ (.B1(_01589_),
    .Y(_02219_),
    .A1(_02217_),
    .A2(_02218_));
 sg13g2_buf_1 _07545_ (.A(_02219_),
    .X(_02220_));
 sg13g2_a21oi_1 _07546_ (.A1(net188),
    .A2(_02215_),
    .Y(_02221_),
    .B1(net166));
 sg13g2_buf_1 _07547_ (.A(net226),
    .X(_02222_));
 sg13g2_buf_1 _07548_ (.A(_02222_),
    .X(_02223_));
 sg13g2_nand2_1 _07549_ (.Y(_02224_),
    .A(net187),
    .B(\i_tinyqv.cpu.instr_data_in[12] ));
 sg13g2_buf_1 _07550_ (.A(_00964_),
    .X(_02225_));
 sg13g2_buf_1 _07551_ (.A(\i_tinyqv.cpu.instr_data_in[8] ),
    .X(_02226_));
 sg13g2_nand2_1 _07552_ (.Y(_02227_),
    .A(net204),
    .B(_02226_));
 sg13g2_nand2_1 _07553_ (.Y(_02228_),
    .A(net210),
    .B(_01563_));
 sg13g2_a21oi_1 _07554_ (.A1(_02224_),
    .A2(_02227_),
    .Y(_02229_),
    .B1(_02228_));
 sg13g2_nor2_1 _07555_ (.A(net188),
    .B(_02229_),
    .Y(_02230_));
 sg13g2_buf_1 _07556_ (.A(net220),
    .X(_02231_));
 sg13g2_buf_1 _07557_ (.A(net203),
    .X(_02232_));
 sg13g2_buf_1 _07558_ (.A(net205),
    .X(_02233_));
 sg13g2_inv_1 _07559_ (.Y(_02234_),
    .A(\i_tinyqv.cpu.instr_data_in[0] ));
 sg13g2_buf_1 _07560_ (.A(\i_tinyqv.cpu.instr_data_in[4] ),
    .X(_02235_));
 sg13g2_nand2_1 _07561_ (.Y(_02236_),
    .A(net187),
    .B(_02235_));
 sg13g2_o21ai_1 _07562_ (.B1(_02236_),
    .Y(_02237_),
    .A1(net185),
    .A2(_02234_));
 sg13g2_nor2_1 _07563_ (.A(net186),
    .B(_02237_),
    .Y(_02238_));
 sg13g2_nor3_1 _07564_ (.A(_01508_),
    .B(_02230_),
    .C(_02238_),
    .Y(_02239_));
 sg13g2_a22oi_1 _07565_ (.Y(_02240_),
    .B1(_02237_),
    .B2(_02228_),
    .A2(_02229_),
    .A1(_01508_));
 sg13g2_and2_1 _07566_ (.A(net210),
    .B(_01563_),
    .X(_02241_));
 sg13g2_buf_2 _07567_ (.A(_02241_),
    .X(_02242_));
 sg13g2_nand2_1 _07568_ (.Y(_02243_),
    .A(_01235_),
    .B(_02242_));
 sg13g2_mux2_1 _07569_ (.A0(\i_tinyqv.mem.qspi_data_buf[8] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[12] ),
    .S(net185),
    .X(_02244_));
 sg13g2_nand3_1 _07570_ (.B(_02243_),
    .C(_02244_),
    .A(net186),
    .Y(_02245_));
 sg13g2_o21ai_1 _07571_ (.B1(_02245_),
    .Y(_02246_),
    .A1(net186),
    .A2(_02240_));
 sg13g2_buf_1 _07572_ (.A(_00892_),
    .X(_02247_));
 sg13g2_nand2_1 _07573_ (.Y(_02248_),
    .A(net202),
    .B(_01506_));
 sg13g2_nor3_1 _07574_ (.A(_02239_),
    .B(_02246_),
    .C(_02248_),
    .Y(_02249_));
 sg13g2_buf_1 _07575_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .X(_02250_));
 sg13g2_nor2_1 _07576_ (.A(net211),
    .B(_01263_),
    .Y(_02251_));
 sg13g2_nor2_1 _07577_ (.A(net227),
    .B(_02251_),
    .Y(_02252_));
 sg13g2_nor2_1 _07578_ (.A(_02250_),
    .B(_02252_),
    .Y(_02253_));
 sg13g2_buf_2 _07579_ (.A(_02253_),
    .X(_02254_));
 sg13g2_mux4_1 _07580_ (.S0(net185),
    .A0(\i_tinyqv.mem.qspi_data_buf[24] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[28] ),
    .A2(_02226_),
    .A3(\i_tinyqv.cpu.instr_data_in[12] ),
    .S1(_01563_),
    .X(_02255_));
 sg13g2_nor2_1 _07581_ (.A(_02178_),
    .B(_02255_),
    .Y(_02256_));
 sg13g2_mux2_1 _07582_ (.A0(\i_tinyqv.mem.data_from_read[16] ),
    .A1(\i_tinyqv.mem.data_from_read[20] ),
    .S(net185),
    .X(_02257_));
 sg13g2_nor2_1 _07583_ (.A(net186),
    .B(_02257_),
    .Y(_02258_));
 sg13g2_o21ai_1 _07584_ (.B1(_01506_),
    .Y(_02259_),
    .A1(_02256_),
    .A2(_02258_));
 sg13g2_a21oi_1 _07585_ (.A1(net166),
    .A2(_02259_),
    .Y(_02260_),
    .B1(net202));
 sg13g2_nor4_1 _07586_ (.A(_02221_),
    .B(_02249_),
    .C(_02254_),
    .D(_02260_),
    .Y(_02261_));
 sg13g2_nand2_1 _07587_ (.Y(_02262_),
    .A(\i_tinyqv.cpu.i_core.load_top_bit ),
    .B(_02254_));
 sg13g2_nand2b_1 _07588_ (.Y(_02263_),
    .B(_02262_),
    .A_N(_01535_));
 sg13g2_buf_1 _07589_ (.A(net227),
    .X(_02264_));
 sg13g2_buf_1 _07590_ (.A(\i_tinyqv.cpu.instr_data_start[12] ),
    .X(_02265_));
 sg13g2_buf_1 _07591_ (.A(_00759_),
    .X(_02266_));
 sg13g2_nand2_1 _07592_ (.Y(_02267_),
    .A(_00858_),
    .B(net258));
 sg13g2_nand2_1 _07593_ (.Y(_02268_),
    .A(net312),
    .B(_01403_));
 sg13g2_buf_2 _07594_ (.A(_02268_),
    .X(_02269_));
 sg13g2_nand2_1 _07595_ (.Y(_02270_),
    .A(_00988_),
    .B(net303));
 sg13g2_nor2_2 _07596_ (.A(_02269_),
    .B(_02270_),
    .Y(_02271_));
 sg13g2_nand2b_1 _07597_ (.Y(_02272_),
    .B(_02271_),
    .A_N(_02267_));
 sg13g2_buf_1 _07598_ (.A(_02272_),
    .X(_02273_));
 sg13g2_buf_1 _07599_ (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .X(_02274_));
 sg13g2_buf_1 _07600_ (.A(_00768_),
    .X(_02275_));
 sg13g2_buf_1 _07601_ (.A(\i_tinyqv.cpu.instr_data_start[9] ),
    .X(_02276_));
 sg13g2_and3_1 _07602_ (.X(_02277_),
    .A(_02275_),
    .B(net287),
    .C(net304));
 sg13g2_buf_1 _07603_ (.A(_02277_),
    .X(_02278_));
 sg13g2_nand2_1 _07604_ (.Y(_02279_),
    .A(net288),
    .B(_02278_));
 sg13g2_nor2_1 _07605_ (.A(_02273_),
    .B(_02279_),
    .Y(_02280_));
 sg13g2_xor2_1 _07606_ (.B(_02280_),
    .A(net289),
    .X(_02281_));
 sg13g2_xnor2_1 _07607_ (.Y(_02282_),
    .A(_01142_),
    .B(_02273_));
 sg13g2_mux2_1 _07608_ (.A0(_02281_),
    .A1(_02282_),
    .S(net204),
    .X(_02283_));
 sg13g2_buf_1 _07609_ (.A(_00161_),
    .X(_02284_));
 sg13g2_nor2_1 _07610_ (.A(_02284_),
    .B(_02269_),
    .Y(_02285_));
 sg13g2_buf_2 _07611_ (.A(_02285_),
    .X(_02286_));
 sg13g2_and2_1 _07612_ (.A(_02284_),
    .B(_02269_),
    .X(_02287_));
 sg13g2_nor2_1 _07613_ (.A(_02286_),
    .B(_02287_),
    .Y(_02288_));
 sg13g2_a22oi_1 _07614_ (.Y(_02289_),
    .B1(_02288_),
    .B2(_01145_),
    .A2(_02283_),
    .A1(net203));
 sg13g2_buf_1 _07615_ (.A(_00988_),
    .X(_02290_));
 sg13g2_buf_1 _07616_ (.A(_00858_),
    .X(_02291_));
 sg13g2_buf_1 _07617_ (.A(_00769_),
    .X(_02292_));
 sg13g2_and4_1 _07618_ (.A(net288),
    .B(_00992_),
    .C(net289),
    .D(_02278_),
    .X(_02293_));
 sg13g2_buf_1 _07619_ (.A(_02293_),
    .X(_02294_));
 sg13g2_and4_1 _07620_ (.A(net255),
    .B(net258),
    .C(net254),
    .D(_02294_),
    .X(_02295_));
 sg13g2_buf_1 _07621_ (.A(_02295_),
    .X(_02296_));
 sg13g2_buf_1 _07622_ (.A(\i_tinyqv.cpu.instr_data_start[18] ),
    .X(_02297_));
 sg13g2_and2_1 _07623_ (.A(_00861_),
    .B(net305),
    .X(_02298_));
 sg13g2_buf_1 _07624_ (.A(_02298_),
    .X(_02299_));
 sg13g2_and3_1 _07625_ (.X(_02300_),
    .A(_02297_),
    .B(net308),
    .C(_02299_));
 sg13g2_buf_1 _07626_ (.A(_02300_),
    .X(_02301_));
 sg13g2_and2_1 _07627_ (.A(_00859_),
    .B(_02301_),
    .X(_02302_));
 sg13g2_nand4_1 _07628_ (.B(net303),
    .C(_02296_),
    .A(net256),
    .Y(_02303_),
    .D(_02302_));
 sg13g2_nor2_1 _07629_ (.A(_02269_),
    .B(_02303_),
    .Y(_02304_));
 sg13g2_xnor2_1 _07630_ (.Y(_02305_),
    .A(_01138_),
    .B(_02304_));
 sg13g2_buf_1 _07631_ (.A(_00861_),
    .X(_02306_));
 sg13g2_inv_1 _07632_ (.Y(_02307_),
    .A(_02273_));
 sg13g2_buf_1 _07633_ (.A(_00992_),
    .X(_02308_));
 sg13g2_and4_1 _07634_ (.A(net288),
    .B(net254),
    .C(net252),
    .D(net289),
    .X(_02309_));
 sg13g2_buf_1 _07635_ (.A(_02309_),
    .X(_02310_));
 sg13g2_nand4_1 _07636_ (.B(_02278_),
    .C(_02307_),
    .A(net253),
    .Y(_02311_),
    .D(_02310_));
 sg13g2_xnor2_1 _07637_ (.Y(_02312_),
    .A(net305),
    .B(_02311_));
 sg13g2_nand2_1 _07638_ (.Y(_02313_),
    .A(net204),
    .B(_02312_));
 sg13g2_o21ai_1 _07639_ (.B1(_02313_),
    .Y(_02314_),
    .A1(net207),
    .A2(_02305_));
 sg13g2_nand3_1 _07640_ (.B(_00088_),
    .C(_02314_),
    .A(net201),
    .Y(_02315_));
 sg13g2_o21ai_1 _07641_ (.B1(_02315_),
    .Y(_02316_),
    .A1(net201),
    .A2(_02289_));
 sg13g2_inv_1 _07642_ (.Y(_02317_),
    .A(net311));
 sg13g2_buf_1 _07643_ (.A(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .X(_02318_));
 sg13g2_nand2_1 _07644_ (.Y(_02319_),
    .A(net302),
    .B(net306));
 sg13g2_nor3_1 _07645_ (.A(net310),
    .B(net285),
    .C(_02319_),
    .Y(_02320_));
 sg13g2_nor3_1 _07646_ (.A(_00956_),
    .B(_01091_),
    .C(_01041_),
    .Y(_02321_));
 sg13g2_nor2b_1 _07647_ (.A(_00920_),
    .B_N(_02321_),
    .Y(_02322_));
 sg13g2_nand2_2 _07648_ (.Y(_02323_),
    .A(_02320_),
    .B(_02322_));
 sg13g2_nor3_1 _07649_ (.A(_02317_),
    .B(_01040_),
    .C(_02323_),
    .Y(_02324_));
 sg13g2_inv_1 _07650_ (.Y(_02325_),
    .A(_01040_));
 sg13g2_nand3_1 _07651_ (.B(_02320_),
    .C(_02321_),
    .A(_00920_),
    .Y(_02326_));
 sg13g2_buf_1 _07652_ (.A(_02326_),
    .X(_02327_));
 sg13g2_nor3_1 _07653_ (.A(net311),
    .B(_02325_),
    .C(_02327_),
    .Y(_02328_));
 sg13g2_nor2_1 _07654_ (.A(_00955_),
    .B(_01090_),
    .Y(_02329_));
 sg13g2_o21ai_1 _07655_ (.B1(_02329_),
    .Y(_02330_),
    .A1(_02324_),
    .A2(_02328_));
 sg13g2_nand3_1 _07656_ (.B(_01040_),
    .C(_02329_),
    .A(_02317_),
    .Y(_02331_));
 sg13g2_or2_1 _07657_ (.X(_02332_),
    .B(_02331_),
    .A(_02323_));
 sg13g2_inv_1 _07658_ (.Y(_02333_),
    .A(_02332_));
 sg13g2_nand4_1 _07659_ (.B(net285),
    .C(_01192_),
    .A(net310),
    .Y(_02334_),
    .D(_02322_));
 sg13g2_buf_1 _07660_ (.A(_02334_),
    .X(_02335_));
 sg13g2_nand2_1 _07661_ (.Y(_02336_),
    .A(_02325_),
    .B(_02329_));
 sg13g2_nor3_2 _07662_ (.A(net311),
    .B(_02335_),
    .C(_02336_),
    .Y(_02337_));
 sg13g2_inv_1 _07663_ (.Y(_02338_),
    .A(_00955_));
 sg13g2_nand4_1 _07664_ (.B(_02317_),
    .C(_01090_),
    .A(_02338_),
    .Y(_02339_),
    .D(_02325_));
 sg13g2_nor2_2 _07665_ (.A(_02327_),
    .B(_02339_),
    .Y(_02340_));
 sg13g2_nor2_2 _07666_ (.A(_02335_),
    .B(_02339_),
    .Y(_02341_));
 sg13g2_nor4_1 _07667_ (.A(_02333_),
    .B(_02337_),
    .C(_02340_),
    .D(_02341_),
    .Y(_02342_));
 sg13g2_nand2_1 _07668_ (.Y(_02343_),
    .A(_02330_),
    .B(_02342_));
 sg13g2_nor3_2 _07669_ (.A(net311),
    .B(_02323_),
    .C(_02336_),
    .Y(_02344_));
 sg13g2_nor2_1 _07670_ (.A(_02331_),
    .B(_02335_),
    .Y(_02345_));
 sg13g2_buf_2 _07671_ (.A(_02345_),
    .X(_02346_));
 sg13g2_nand3_1 _07672_ (.B(_02325_),
    .C(_02329_),
    .A(net311),
    .Y(_02347_));
 sg13g2_or2_1 _07673_ (.X(_02348_),
    .B(_02347_),
    .A(_02327_));
 sg13g2_buf_1 _07674_ (.A(_02348_),
    .X(_02349_));
 sg13g2_inv_1 _07675_ (.Y(_02350_),
    .A(_02349_));
 sg13g2_nor4_1 _07676_ (.A(_02343_),
    .B(_02344_),
    .C(_02346_),
    .D(_02350_),
    .Y(_02351_));
 sg13g2_or3_1 _07677_ (.A(_01206_),
    .B(_01537_),
    .C(_02351_),
    .X(_02352_));
 sg13g2_inv_1 _07678_ (.Y(_02353_),
    .A(_02352_));
 sg13g2_nor2_2 _07679_ (.A(net211),
    .B(_00892_),
    .Y(_02354_));
 sg13g2_or2_1 _07680_ (.X(_02355_),
    .B(_02331_),
    .A(_02327_));
 sg13g2_nor2_1 _07681_ (.A(_02354_),
    .B(_02355_),
    .Y(_02356_));
 sg13g2_nand2_1 _07682_ (.Y(_02357_),
    .A(net227),
    .B(_01055_));
 sg13g2_buf_2 _07683_ (.A(_02357_),
    .X(_02358_));
 sg13g2_nor2_2 _07684_ (.A(_02349_),
    .B(_02358_),
    .Y(_02359_));
 sg13g2_and3_1 _07685_ (.X(_02360_),
    .A(\i_tinyqv.cpu.i_core.mcause[0] ),
    .B(_01057_),
    .C(_02340_));
 sg13g2_a221oi_1 _07686_ (.B2(\i_tinyqv.cpu.i_core.mip[16] ),
    .C1(_02360_),
    .B1(_02359_),
    .A1(\i_tinyqv.cpu.i_core.mepc[0] ),
    .Y(_02361_),
    .A2(_02356_));
 sg13g2_and2_1 _07687_ (.A(\i_tinyqv.cpu.i_core.mcause[4] ),
    .B(_02340_),
    .X(_02362_));
 sg13g2_nand2_1 _07688_ (.Y(_02363_),
    .A(net264),
    .B(_01145_));
 sg13g2_inv_1 _07689_ (.Y(_02364_),
    .A(_02363_));
 sg13g2_o21ai_1 _07690_ (.B1(_02364_),
    .Y(_02365_),
    .A1(_02333_),
    .A2(_02362_));
 sg13g2_buf_1 _07691_ (.A(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .X(_02366_));
 sg13g2_a22oi_1 _07692_ (.Y(_02367_),
    .B1(_02346_),
    .B2(_02366_),
    .A2(_02337_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[0] ));
 sg13g2_inv_1 _07693_ (.Y(_02368_),
    .A(_00168_));
 sg13g2_nor3_2 _07694_ (.A(_02323_),
    .B(_02347_),
    .C(_02358_),
    .Y(_02369_));
 sg13g2_a22oi_1 _07695_ (.Y(_02370_),
    .B1(_02369_),
    .B2(\i_tinyqv.cpu.i_core.mie[16] ),
    .A2(_02341_),
    .A1(_02368_));
 sg13g2_nand4_1 _07696_ (.B(_02365_),
    .C(_02367_),
    .A(_02361_),
    .Y(_02371_),
    .D(_02370_));
 sg13g2_a22oi_1 _07697_ (.Y(_02372_),
    .B1(_02353_),
    .B2(_02371_),
    .A2(_02316_),
    .A1(_01274_));
 sg13g2_nand2_1 _07698_ (.Y(_02373_),
    .A(net218),
    .B(\i_tinyqv.cpu.is_lui ));
 sg13g2_buf_2 _07699_ (.A(_02373_),
    .X(_02374_));
 sg13g2_mux2_1 _07700_ (.A0(_01049_),
    .A1(_02372_),
    .S(_02374_),
    .X(_02375_));
 sg13g2_nand2_1 _07701_ (.Y(_02376_),
    .A(_01535_),
    .B(_02375_));
 sg13g2_o21ai_1 _07702_ (.B1(_02376_),
    .Y(_02377_),
    .A1(_02261_),
    .A2(_02263_));
 sg13g2_nand2b_1 _07703_ (.Y(_02378_),
    .B(_01646_),
    .A_N(_01647_));
 sg13g2_buf_1 _07704_ (.A(_02378_),
    .X(_02379_));
 sg13g2_o21ai_1 _07705_ (.B1(_01109_),
    .Y(_02380_),
    .A1(_00169_),
    .A2(_02379_));
 sg13g2_buf_1 _07706_ (.A(_01057_),
    .X(_02381_));
 sg13g2_nor2_1 _07707_ (.A(net313),
    .B(_02379_),
    .Y(_02382_));
 sg13g2_and3_1 _07708_ (.X(_02383_),
    .A(net157),
    .B(_01176_),
    .C(_02382_));
 sg13g2_buf_1 _07709_ (.A(_02383_),
    .X(_02384_));
 sg13g2_nand2_1 _07710_ (.Y(_02385_),
    .A(net313),
    .B(_01176_));
 sg13g2_buf_1 _07711_ (.A(_02385_),
    .X(_02386_));
 sg13g2_nand2_1 _07712_ (.Y(_02387_),
    .A(net259),
    .B(net120));
 sg13g2_xor2_1 _07713_ (.B(_02387_),
    .A(_01740_),
    .X(_02388_));
 sg13g2_nor2b_1 _07714_ (.A(_01152_),
    .B_N(_01052_),
    .Y(_02389_));
 sg13g2_inv_1 _07715_ (.Y(_02390_),
    .A(_01177_));
 sg13g2_and4_1 _07716_ (.A(_00824_),
    .B(_02390_),
    .C(_01186_),
    .D(net171),
    .X(_02391_));
 sg13g2_buf_1 _07717_ (.A(_02391_),
    .X(_02392_));
 sg13g2_xnor2_1 _07718_ (.Y(_02393_),
    .A(net193),
    .B(_01063_));
 sg13g2_and2_1 _07719_ (.A(_02392_),
    .B(_02393_),
    .X(_02394_));
 sg13g2_nor3_1 _07720_ (.A(_00824_),
    .B(_01186_),
    .C(_01109_),
    .Y(_02395_));
 sg13g2_nor2_1 _07721_ (.A(_02394_),
    .B(_02395_),
    .Y(_02396_));
 sg13g2_nor2_1 _07722_ (.A(_01052_),
    .B(_02396_),
    .Y(_02397_));
 sg13g2_a22oi_1 _07723_ (.Y(_02398_),
    .B1(_02397_),
    .B2(_01152_),
    .A2(_02394_),
    .A1(_02389_));
 sg13g2_o21ai_1 _07724_ (.B1(net171),
    .Y(_02399_),
    .A1(_01177_),
    .A2(_01186_));
 sg13g2_buf_1 _07725_ (.A(_02399_),
    .X(_02400_));
 sg13g2_nand4_1 _07726_ (.B(_02390_),
    .C(_01186_),
    .A(_00824_),
    .Y(_02401_),
    .D(net171));
 sg13g2_nor2_1 _07727_ (.A(_02401_),
    .B(_02393_),
    .Y(_02402_));
 sg13g2_o21ai_1 _07728_ (.B1(_01211_),
    .Y(_02403_),
    .A1(_02400_),
    .A2(_02402_));
 sg13g2_nand2_1 _07729_ (.Y(_02404_),
    .A(_02398_),
    .B(_02403_));
 sg13g2_nand2_1 _07730_ (.Y(_02405_),
    .A(net184),
    .B(_02404_));
 sg13g2_o21ai_1 _07731_ (.B1(_02405_),
    .Y(_02406_),
    .A1(net184),
    .A2(_02388_));
 sg13g2_nor2_1 _07732_ (.A(_01179_),
    .B(_02379_),
    .Y(_02407_));
 sg13g2_buf_2 _07733_ (.A(_02407_),
    .X(_02408_));
 sg13g2_buf_2 _07734_ (.A(net315),
    .X(_02409_));
 sg13g2_buf_2 _07735_ (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .X(_02410_));
 sg13g2_xor2_1 _07736_ (.B(_02410_),
    .A(net251),
    .X(_02411_));
 sg13g2_mux2_1 _07737_ (.A0(_00195_),
    .A1(_00194_),
    .S(_02411_),
    .X(_02412_));
 sg13g2_buf_1 _07738_ (.A(net315),
    .X(_02413_));
 sg13g2_buf_1 _07739_ (.A(_02410_),
    .X(_02414_));
 sg13g2_mux4_1 _07740_ (.S0(net250),
    .A0(_00187_),
    .A1(_00186_),
    .A2(_00189_),
    .A3(_00188_),
    .S1(net249),
    .X(_02415_));
 sg13g2_buf_1 _07741_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .X(_02416_));
 sg13g2_xnor2_1 _07742_ (.Y(_02417_),
    .A(net315),
    .B(_02416_));
 sg13g2_xnor2_1 _07743_ (.Y(_02418_),
    .A(net226),
    .B(_02417_));
 sg13g2_buf_2 _07744_ (.A(_02418_),
    .X(_02419_));
 sg13g2_buf_1 _07745_ (.A(_02419_),
    .X(_02420_));
 sg13g2_mux2_1 _07746_ (.A0(_02412_),
    .A1(_02415_),
    .S(net165),
    .X(_02421_));
 sg13g2_mux4_1 _07747_ (.S0(net250),
    .A0(_00192_),
    .A1(_00193_),
    .A2(_00190_),
    .A3(_00191_),
    .S1(net249),
    .X(_02422_));
 sg13g2_buf_2 _07748_ (.A(net315),
    .X(_02423_));
 sg13g2_mux4_1 _07749_ (.S0(net248),
    .A0(_00191_),
    .A1(_00190_),
    .A2(_00193_),
    .A3(_00192_),
    .S1(net249),
    .X(_02424_));
 sg13g2_buf_1 _07750_ (.A(_02419_),
    .X(_02425_));
 sg13g2_mux2_1 _07751_ (.A0(_02422_),
    .A1(_02424_),
    .S(net164),
    .X(_02426_));
 sg13g2_buf_1 _07752_ (.A(_02410_),
    .X(_02427_));
 sg13g2_mux4_1 _07753_ (.S0(net248),
    .A0(_00179_),
    .A1(_00178_),
    .A2(_00181_),
    .A3(_00180_),
    .S1(net247),
    .X(_02428_));
 sg13g2_buf_1 _07754_ (.A(_00170_),
    .X(_02429_));
 sg13g2_buf_2 _07755_ (.A(net315),
    .X(_02430_));
 sg13g2_buf_1 _07756_ (.A(_02410_),
    .X(_02431_));
 sg13g2_mux4_1 _07757_ (.S0(net246),
    .A0(_00171_),
    .A1(_02429_),
    .A2(_00173_),
    .A3(_00172_),
    .S1(net245),
    .X(_02432_));
 sg13g2_mux2_1 _07758_ (.A0(_02428_),
    .A1(_02432_),
    .S(net165),
    .X(_02433_));
 sg13g2_mux4_1 _07759_ (.S0(net248),
    .A0(_00183_),
    .A1(_00182_),
    .A2(_00185_),
    .A3(_00184_),
    .S1(net247),
    .X(_02434_));
 sg13g2_mux4_1 _07760_ (.S0(_02430_),
    .A0(_00175_),
    .A1(_00174_),
    .A2(_00177_),
    .A3(_00176_),
    .S1(net247),
    .X(_02435_));
 sg13g2_mux2_1 _07761_ (.A0(_02434_),
    .A1(_02435_),
    .S(net165),
    .X(_02436_));
 sg13g2_buf_1 _07762_ (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .X(_02437_));
 sg13g2_buf_1 _07763_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .X(_02438_));
 sg13g2_xor2_1 _07764_ (.B(_02438_),
    .A(net220),
    .X(_02439_));
 sg13g2_nor2b_1 _07765_ (.A(_02416_),
    .B_N(net251),
    .Y(_02440_));
 sg13g2_a21oi_1 _07766_ (.A1(_00964_),
    .A2(_02416_),
    .Y(_02441_),
    .B1(_02440_));
 sg13g2_xnor2_1 _07767_ (.Y(_02442_),
    .A(_02439_),
    .B(_02441_));
 sg13g2_buf_4 _07768_ (.X(_02443_),
    .A(_02442_));
 sg13g2_mux4_1 _07769_ (.S0(net284),
    .A0(_02421_),
    .A1(_02426_),
    .A2(_02433_),
    .A3(_02436_),
    .S1(_02443_),
    .X(_02444_));
 sg13g2_buf_1 _07770_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .X(_02445_));
 sg13g2_nand2_2 _07771_ (.Y(_02446_),
    .A(net313),
    .B(_02445_));
 sg13g2_nand2_1 _07772_ (.Y(_02447_),
    .A(net251),
    .B(_00200_));
 sg13g2_nand2b_1 _07773_ (.Y(_02448_),
    .B(_00169_),
    .A_N(net251));
 sg13g2_a21oi_1 _07774_ (.A1(_02447_),
    .A2(_02448_),
    .Y(_02449_),
    .B1(net245));
 sg13g2_a21oi_1 _07775_ (.A1(_02414_),
    .A2(_02446_),
    .Y(_02450_),
    .B1(_02449_));
 sg13g2_mux4_1 _07776_ (.S0(net251),
    .A0(_00172_),
    .A1(_00173_),
    .A2(_02429_),
    .A3(_00171_),
    .S1(_02410_),
    .X(_02451_));
 sg13g2_nand2_1 _07777_ (.Y(_02452_),
    .A(_02419_),
    .B(_02451_));
 sg13g2_o21ai_1 _07778_ (.B1(_02452_),
    .Y(_02453_),
    .A1(_02425_),
    .A2(_02450_));
 sg13g2_buf_1 _07779_ (.A(_00196_),
    .X(_02454_));
 sg13g2_buf_1 _07780_ (.A(_00198_),
    .X(_02455_));
 sg13g2_mux4_1 _07781_ (.S0(net246),
    .A0(_02454_),
    .A1(_00197_),
    .A2(_02455_),
    .A3(_00199_),
    .S1(net245),
    .X(_02456_));
 sg13g2_nor2b_1 _07782_ (.A(_02419_),
    .B_N(_02446_),
    .Y(_02457_));
 sg13g2_a21o_1 _07783_ (.A2(_02456_),
    .A1(net164),
    .B1(_02457_),
    .X(_02458_));
 sg13g2_mux4_1 _07784_ (.S0(net246),
    .A0(_00180_),
    .A1(_00181_),
    .A2(_00178_),
    .A3(_00179_),
    .S1(net247),
    .X(_02459_));
 sg13g2_mux4_1 _07785_ (.S0(net251),
    .A0(_00188_),
    .A1(_00189_),
    .A2(_00186_),
    .A3(_00187_),
    .S1(net245),
    .X(_02460_));
 sg13g2_mux2_1 _07786_ (.A0(_02459_),
    .A1(_02460_),
    .S(_02419_),
    .X(_02461_));
 sg13g2_mux4_1 _07787_ (.S0(net246),
    .A0(_00176_),
    .A1(_00177_),
    .A2(_00174_),
    .A3(_00175_),
    .S1(net247),
    .X(_02462_));
 sg13g2_mux4_1 _07788_ (.S0(net246),
    .A0(_00184_),
    .A1(_00185_),
    .A2(_00182_),
    .A3(_00183_),
    .S1(_02427_),
    .X(_02463_));
 sg13g2_mux2_1 _07789_ (.A0(_02462_),
    .A1(_02463_),
    .S(net165),
    .X(_02464_));
 sg13g2_mux4_1 _07790_ (.S0(net284),
    .A0(_02453_),
    .A1(_02458_),
    .A2(_02461_),
    .A3(_02464_),
    .S1(_02443_),
    .X(_02465_));
 sg13g2_buf_1 _07791_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .X(_02466_));
 sg13g2_xor2_1 _07792_ (.B(net227),
    .A(_00746_),
    .X(_02467_));
 sg13g2_xnor2_1 _07793_ (.Y(_02468_),
    .A(_02466_),
    .B(_02467_));
 sg13g2_nor2_1 _07794_ (.A(net226),
    .B(_00746_),
    .Y(_02469_));
 sg13g2_a21oi_1 _07795_ (.A1(_00770_),
    .A2(_02438_),
    .Y(_02470_),
    .B1(_02469_));
 sg13g2_mux2_1 _07796_ (.A0(_02438_),
    .A1(net315),
    .S(_00770_),
    .X(_02471_));
 sg13g2_nand2_1 _07797_ (.Y(_02472_),
    .A(net220),
    .B(_02471_));
 sg13g2_o21ai_1 _07798_ (.B1(_02472_),
    .Y(_02473_),
    .A1(_01141_),
    .A2(_02470_));
 sg13g2_xnor2_1 _07799_ (.Y(_02474_),
    .A(_01141_),
    .B(net251));
 sg13g2_a22oi_1 _07800_ (.Y(_02475_),
    .B1(_02474_),
    .B2(_02438_),
    .A2(_02473_),
    .A1(_02416_));
 sg13g2_nand2b_1 _07801_ (.Y(_02476_),
    .B(_02475_),
    .A_N(_02468_));
 sg13g2_buf_4 _07802_ (.X(_02477_),
    .A(_02476_));
 sg13g2_mux2_1 _07803_ (.A0(_02444_),
    .A1(_02465_),
    .S(_02477_),
    .X(_02478_));
 sg13g2_nand2b_1 _07804_ (.Y(_02479_),
    .B(_02466_),
    .A_N(_02475_));
 sg13g2_nor2b_1 _07805_ (.A(_02466_),
    .B_N(_02475_),
    .Y(_02480_));
 sg13g2_a21oi_2 _07806_ (.B1(_02480_),
    .Y(_02481_),
    .A2(_02467_),
    .A1(_02479_));
 sg13g2_mux2_1 _07807_ (.A0(_02478_),
    .A1(_02446_),
    .S(_02481_),
    .X(_02482_));
 sg13g2_mux4_1 _07808_ (.S0(net248),
    .A0(_00189_),
    .A1(_00188_),
    .A2(_00191_),
    .A3(_00190_),
    .S1(net249),
    .X(_02483_));
 sg13g2_mux4_1 _07809_ (.S0(net248),
    .A0(_00181_),
    .A1(_00180_),
    .A2(_00183_),
    .A3(_00182_),
    .S1(net249),
    .X(_02484_));
 sg13g2_mux2_1 _07810_ (.A0(_02483_),
    .A1(_02484_),
    .S(net165),
    .X(_02485_));
 sg13g2_mux4_1 _07811_ (.S0(_02423_),
    .A0(_00193_),
    .A1(_00192_),
    .A2(_00195_),
    .A3(_00194_),
    .S1(_02414_),
    .X(_02486_));
 sg13g2_mux4_1 _07812_ (.S0(_02423_),
    .A0(_00185_),
    .A1(_00184_),
    .A2(_00187_),
    .A3(_00186_),
    .S1(_02427_),
    .X(_02487_));
 sg13g2_mux2_1 _07813_ (.A0(_02486_),
    .A1(_02487_),
    .S(_02420_),
    .X(_02488_));
 sg13g2_mux4_1 _07814_ (.S0(_02410_),
    .A0(_02429_),
    .A1(_02454_),
    .A2(_00171_),
    .A3(_00197_),
    .S1(net250),
    .X(_02489_));
 sg13g2_mux4_1 _07815_ (.S0(net246),
    .A0(_00178_),
    .A1(_00179_),
    .A2(_00176_),
    .A3(_00177_),
    .S1(net245),
    .X(_02490_));
 sg13g2_mux2_1 _07816_ (.A0(_02489_),
    .A1(_02490_),
    .S(net165),
    .X(_02491_));
 sg13g2_mux4_1 _07817_ (.S0(net246),
    .A0(_02455_),
    .A1(_00199_),
    .A2(_00169_),
    .A3(_00200_),
    .S1(net247),
    .X(_02492_));
 sg13g2_mux4_1 _07818_ (.S0(net251),
    .A0(_00174_),
    .A1(_00175_),
    .A2(_00172_),
    .A3(_00173_),
    .S1(net245),
    .X(_02493_));
 sg13g2_mux2_1 _07819_ (.A0(_02492_),
    .A1(_02493_),
    .S(_02419_),
    .X(_02494_));
 sg13g2_mux4_1 _07820_ (.S0(net284),
    .A0(_02485_),
    .A1(_02488_),
    .A2(_02491_),
    .A3(_02494_),
    .S1(_02477_),
    .X(_02495_));
 sg13g2_mux4_1 _07821_ (.S0(net248),
    .A0(_00173_),
    .A1(_00172_),
    .A2(_00175_),
    .A3(_00174_),
    .S1(net249),
    .X(_02496_));
 sg13g2_mux4_1 _07822_ (.S0(_02410_),
    .A0(_00200_),
    .A1(_00199_),
    .A2(_00169_),
    .A3(_02455_),
    .S1(net250),
    .X(_02497_));
 sg13g2_mux2_1 _07823_ (.A0(_02496_),
    .A1(_02497_),
    .S(_02420_),
    .X(_02498_));
 sg13g2_mux4_1 _07824_ (.S0(net248),
    .A0(_00177_),
    .A1(_00176_),
    .A2(_00179_),
    .A3(_00178_),
    .S1(net247),
    .X(_02499_));
 sg13g2_mux4_1 _07825_ (.S0(net248),
    .A0(_00197_),
    .A1(_02454_),
    .A2(_00171_),
    .A3(_02429_),
    .S1(net247),
    .X(_02500_));
 sg13g2_mux2_1 _07826_ (.A0(_02499_),
    .A1(_02500_),
    .S(net165),
    .X(_02501_));
 sg13g2_mux4_1 _07827_ (.S0(_02430_),
    .A0(_00186_),
    .A1(_00187_),
    .A2(_00184_),
    .A3(_00185_),
    .S1(net245),
    .X(_02502_));
 sg13g2_mux4_1 _07828_ (.S0(_02409_),
    .A0(_00194_),
    .A1(_00195_),
    .A2(_00192_),
    .A3(_00193_),
    .S1(net245),
    .X(_02503_));
 sg13g2_mux2_1 _07829_ (.A0(_02502_),
    .A1(_02503_),
    .S(net165),
    .X(_02504_));
 sg13g2_mux4_1 _07830_ (.S0(net246),
    .A0(_00182_),
    .A1(_00183_),
    .A2(_00180_),
    .A3(_00181_),
    .S1(_02431_),
    .X(_02505_));
 sg13g2_mux4_1 _07831_ (.S0(_02409_),
    .A0(_00190_),
    .A1(_00191_),
    .A2(_00188_),
    .A3(_00189_),
    .S1(_02431_),
    .X(_02506_));
 sg13g2_mux2_1 _07832_ (.A0(_02505_),
    .A1(_02506_),
    .S(_02419_),
    .X(_02507_));
 sg13g2_mux4_1 _07833_ (.S0(net284),
    .A0(_02498_),
    .A1(_02501_),
    .A2(_02504_),
    .A3(_02507_),
    .S1(_02477_),
    .X(_02508_));
 sg13g2_mux2_1 _07834_ (.A0(_02495_),
    .A1(_02508_),
    .S(_02443_),
    .X(_02509_));
 sg13g2_mux2_1 _07835_ (.A0(_02509_),
    .A1(_02446_),
    .S(_02481_),
    .X(_02510_));
 sg13g2_mux2_1 _07836_ (.A0(_02482_),
    .A1(_02510_),
    .S(net250),
    .X(_02511_));
 sg13g2_nand2_1 _07837_ (.Y(_02512_),
    .A(_02408_),
    .B(_02511_));
 sg13g2_o21ai_1 _07838_ (.B1(_02512_),
    .Y(_02513_),
    .A1(_02406_),
    .A2(_02408_));
 sg13g2_nor2_1 _07839_ (.A(_02513_),
    .B(_02384_),
    .Y(_02514_));
 sg13g2_a21oi_1 _07840_ (.A1(\i_tinyqv.cpu.i_core.cmp ),
    .A2(_02384_),
    .Y(_02515_),
    .B1(_02514_));
 sg13g2_nand2_1 _07841_ (.Y(_02516_),
    .A(net171),
    .B(_02515_));
 sg13g2_nand3_1 _07842_ (.B(_02380_),
    .C(_02516_),
    .A(_01532_),
    .Y(_02517_));
 sg13g2_o21ai_1 _07843_ (.B1(_02517_),
    .Y(_02518_),
    .A1(net189),
    .A2(_02377_));
 sg13g2_buf_1 _07844_ (.A(_02518_),
    .X(_02519_));
 sg13g2_buf_1 _07845_ (.A(_02519_),
    .X(\debug_rd[0] ));
 sg13g2_buf_2 _07846_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .X(_02520_));
 sg13g2_buf_2 _07847_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .X(_02521_));
 sg13g2_nand2_2 _07848_ (.Y(_02522_),
    .A(_02520_),
    .B(_02521_));
 sg13g2_inv_1 _07849_ (.Y(_02523_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ));
 sg13g2_buf_1 _07850_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .X(_02524_));
 sg13g2_inv_1 _07851_ (.Y(_02525_),
    .A(_02524_));
 sg13g2_or3_1 _07852_ (.A(_02523_),
    .B(_02525_),
    .C(_01541_),
    .X(_02526_));
 sg13g2_buf_2 _07853_ (.A(_02526_),
    .X(_02527_));
 sg13g2_nor2_2 _07854_ (.A(_02522_),
    .B(_02527_),
    .Y(_02528_));
 sg13g2_mux2_1 _07855_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .A1(net64),
    .S(_02528_),
    .X(_00050_));
 sg13g2_nor2_1 _07856_ (.A(_01109_),
    .B(_02384_),
    .Y(_02529_));
 sg13g2_nand2_1 _07857_ (.Y(_02530_),
    .A(_01152_),
    .B(net125));
 sg13g2_o21ai_1 _07858_ (.B1(_01063_),
    .Y(_02531_),
    .A1(_01152_),
    .A2(net125));
 sg13g2_nand3_1 _07859_ (.B(_02530_),
    .C(_02531_),
    .A(_00930_),
    .Y(_02532_));
 sg13g2_nand2_1 _07860_ (.Y(_02533_),
    .A(_01058_),
    .B(_01061_));
 sg13g2_nand2_1 _07861_ (.Y(_02534_),
    .A(net125),
    .B(_02533_));
 sg13g2_nand2b_1 _07862_ (.Y(_02535_),
    .B(_01102_),
    .A_N(_01152_));
 sg13g2_nand3_1 _07863_ (.B(_02534_),
    .C(_02535_),
    .A(net193),
    .Y(_02536_));
 sg13g2_and2_1 _07864_ (.A(_02532_),
    .B(_02536_),
    .X(_02537_));
 sg13g2_a21oi_1 _07865_ (.A1(_02392_),
    .A2(_02537_),
    .Y(_02538_),
    .B1(_02400_));
 sg13g2_nor2_1 _07866_ (.A(_02401_),
    .B(_02537_),
    .Y(_02539_));
 sg13g2_or2_1 _07867_ (.X(_02540_),
    .B(_02539_),
    .A(_02395_));
 sg13g2_nor2_1 _07868_ (.A(_01104_),
    .B(_01017_),
    .Y(_02541_));
 sg13g2_a22oi_1 _07869_ (.Y(_02542_),
    .B1(_02540_),
    .B2(_02541_),
    .A2(_02539_),
    .A1(_01156_));
 sg13g2_o21ai_1 _07870_ (.B1(_02542_),
    .Y(_02543_),
    .A1(_01215_),
    .A2(_02538_));
 sg13g2_nor2_1 _07871_ (.A(_01740_),
    .B(_01662_),
    .Y(_02544_));
 sg13g2_o21ai_1 _07872_ (.B1(net118),
    .Y(_02545_),
    .A1(_01736_),
    .A2(_02544_));
 sg13g2_nor3_1 _07873_ (.A(_01662_),
    .B(_01736_),
    .C(net118),
    .Y(_02546_));
 sg13g2_o21ai_1 _07874_ (.B1(_01740_),
    .Y(_02547_),
    .A1(_01700_),
    .A2(_02546_));
 sg13g2_nand2_1 _07875_ (.Y(_02548_),
    .A(_02545_),
    .B(_02547_));
 sg13g2_o21ai_1 _07876_ (.B1(net259),
    .Y(_02549_),
    .A1(_01740_),
    .A2(net118));
 sg13g2_a22oi_1 _07877_ (.Y(_02550_),
    .B1(_02549_),
    .B2(_01737_),
    .A2(_02548_),
    .A1(net259));
 sg13g2_xor2_1 _07878_ (.B(_02550_),
    .A(_01735_),
    .X(_02551_));
 sg13g2_nor2_1 _07879_ (.A(net184),
    .B(_02551_),
    .Y(_02552_));
 sg13g2_a21oi_1 _07880_ (.A1(net184),
    .A2(_02543_),
    .Y(_02553_),
    .B1(_02552_));
 sg13g2_mux2_1 _07881_ (.A0(_02503_),
    .A1(_02483_),
    .S(net164),
    .X(_02554_));
 sg13g2_mux2_1 _07882_ (.A0(_02484_),
    .A1(_02496_),
    .S(net164),
    .X(_02555_));
 sg13g2_mux4_1 _07883_ (.S0(_02443_),
    .A0(_02488_),
    .A1(_02501_),
    .A2(_02554_),
    .A3(_02555_),
    .S1(net284),
    .X(_02556_));
 sg13g2_a21o_1 _07884_ (.A2(_02489_),
    .A1(net164),
    .B1(_02457_),
    .X(_02557_));
 sg13g2_mux2_1 _07885_ (.A0(_02490_),
    .A1(_02502_),
    .S(_02425_),
    .X(_02558_));
 sg13g2_mux4_1 _07886_ (.S0(_02443_),
    .A0(_02494_),
    .A1(_02507_),
    .A2(_02557_),
    .A3(_02558_),
    .S1(_02437_),
    .X(_02559_));
 sg13g2_mux2_1 _07887_ (.A0(_02556_),
    .A1(_02559_),
    .S(_02477_),
    .X(_02560_));
 sg13g2_mux2_1 _07888_ (.A0(_02560_),
    .A1(_02446_),
    .S(_02481_),
    .X(_02561_));
 sg13g2_mux2_1 _07889_ (.A0(_02421_),
    .A1(_02453_),
    .S(_02477_),
    .X(_02562_));
 sg13g2_mux4_1 _07890_ (.S0(net164),
    .A0(_02424_),
    .A1(_02434_),
    .A2(_02456_),
    .A3(_02462_),
    .S1(_02477_),
    .X(_02563_));
 sg13g2_nor2b_1 _07891_ (.A(net284),
    .B_N(_02563_),
    .Y(_02564_));
 sg13g2_a21oi_1 _07892_ (.A1(net284),
    .A2(_02562_),
    .Y(_02565_),
    .B1(_02564_));
 sg13g2_mux4_1 _07893_ (.S0(net250),
    .A0(_00199_),
    .A1(_02455_),
    .A2(_00197_),
    .A3(_02454_),
    .S1(net249),
    .X(_02566_));
 sg13g2_mux2_1 _07894_ (.A0(_02435_),
    .A1(_02566_),
    .S(net164),
    .X(_02567_));
 sg13g2_mux2_1 _07895_ (.A0(_02463_),
    .A1(_02422_),
    .S(net164),
    .X(_02568_));
 sg13g2_mux4_1 _07896_ (.S0(_02477_),
    .A0(_02567_),
    .A1(_02568_),
    .A2(_02433_),
    .A3(_02461_),
    .S1(net284),
    .X(_02569_));
 sg13g2_nand2_1 _07897_ (.Y(_02570_),
    .A(_02443_),
    .B(_02569_));
 sg13g2_o21ai_1 _07898_ (.B1(_02570_),
    .Y(_02571_),
    .A1(_02443_),
    .A2(_02565_));
 sg13g2_mux2_1 _07899_ (.A0(_02571_),
    .A1(_02446_),
    .S(_02481_),
    .X(_02572_));
 sg13g2_mux2_1 _07900_ (.A0(_02561_),
    .A1(_02572_),
    .S(_02413_),
    .X(_02573_));
 sg13g2_nand2b_1 _07901_ (.Y(_02574_),
    .B(_02408_),
    .A_N(_02573_));
 sg13g2_o21ai_1 _07902_ (.B1(_02574_),
    .Y(_02575_),
    .A1(_02408_),
    .A2(_02553_));
 sg13g2_or2_1 _07903_ (.X(_02576_),
    .B(_02379_),
    .A(_01167_));
 sg13g2_buf_1 _07904_ (.A(_02576_),
    .X(_02577_));
 sg13g2_nor2_1 _07905_ (.A(_02455_),
    .B(_02577_),
    .Y(_02578_));
 sg13g2_a21oi_1 _07906_ (.A1(_02529_),
    .A2(_02575_),
    .Y(_02579_),
    .B1(_02578_));
 sg13g2_and2_1 _07907_ (.A(net205),
    .B(\i_tinyqv.mem.data_from_read[21] ),
    .X(_02580_));
 sg13g2_a21oi_1 _07908_ (.A1(net204),
    .A2(\i_tinyqv.mem.data_from_read[17] ),
    .Y(_02581_),
    .B1(_02580_));
 sg13g2_buf_1 _07909_ (.A(\i_tinyqv.cpu.instr_data_in[9] ),
    .X(_02582_));
 sg13g2_mux4_1 _07910_ (.S0(net205),
    .A0(\i_tinyqv.mem.qspi_data_buf[25] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[29] ),
    .A2(_02582_),
    .A3(\i_tinyqv.cpu.instr_data_in[13] ),
    .S1(_01563_),
    .X(_02583_));
 sg13g2_nand2_1 _07911_ (.Y(_02584_),
    .A(net220),
    .B(_02583_));
 sg13g2_o21ai_1 _07912_ (.B1(_02584_),
    .Y(_02585_),
    .A1(net203),
    .A2(_02581_));
 sg13g2_mux2_1 _07913_ (.A0(\i_tinyqv.mem.qspi_data_buf[9] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[13] ),
    .S(net205),
    .X(_02586_));
 sg13g2_nand3_1 _07914_ (.B(_02243_),
    .C(_02586_),
    .A(net220),
    .Y(_02587_));
 sg13g2_mux2_1 _07915_ (.A0(_02582_),
    .A1(\i_tinyqv.cpu.instr_data_in[13] ),
    .S(net226),
    .X(_02588_));
 sg13g2_nand3_1 _07916_ (.B(_02242_),
    .C(_02588_),
    .A(_01508_),
    .Y(_02589_));
 sg13g2_inv_1 _07917_ (.Y(_02590_),
    .A(\i_tinyqv.cpu.instr_data_in[1] ));
 sg13g2_buf_1 _07918_ (.A(\i_tinyqv.cpu.instr_data_in[5] ),
    .X(_02591_));
 sg13g2_nand2_1 _07919_ (.Y(_02592_),
    .A(net226),
    .B(_02591_));
 sg13g2_o21ai_1 _07920_ (.B1(_02592_),
    .Y(_02593_),
    .A1(net226),
    .A2(_02590_));
 sg13g2_nand2_1 _07921_ (.Y(_02594_),
    .A(_02228_),
    .B(_02593_));
 sg13g2_nand2_1 _07922_ (.Y(_02595_),
    .A(_02589_),
    .B(_02594_));
 sg13g2_nor2_1 _07923_ (.A(net220),
    .B(_02593_),
    .Y(_02596_));
 sg13g2_a21oi_1 _07924_ (.A1(_02242_),
    .A2(_02588_),
    .Y(_02597_),
    .B1(net211));
 sg13g2_nor2_1 _07925_ (.A(_02596_),
    .B(_02597_),
    .Y(_02598_));
 sg13g2_a22oi_1 _07926_ (.Y(_02599_),
    .B1(_02598_),
    .B2(_01235_),
    .A2(_02595_),
    .A1(net211));
 sg13g2_a21oi_1 _07927_ (.A1(_02587_),
    .A2(_02599_),
    .Y(_02600_),
    .B1(net227));
 sg13g2_a21oi_1 _07928_ (.A1(net201),
    .A2(_02585_),
    .Y(_02601_),
    .B1(_02600_));
 sg13g2_nand2_1 _07929_ (.Y(_02602_),
    .A(_01506_),
    .B(_02601_));
 sg13g2_buf_1 _07930_ (.A(net185),
    .X(_02603_));
 sg13g2_a221oi_1 _07931_ (.B2(net3),
    .C1(_02603_),
    .B1(_02192_),
    .A1(\gpio_out_sel[1] ),
    .Y(_02604_),
    .A2(_01622_));
 sg13g2_nand2_1 _07932_ (.Y(_02605_),
    .A(\i_spi.data[1] ),
    .B(net131));
 sg13g2_nand3_1 _07933_ (.B(_02180_),
    .C(_02190_),
    .A(_01381_),
    .Y(_02606_));
 sg13g2_a22oi_1 _07934_ (.Y(_02607_),
    .B1(net150),
    .B2(\i_uart_rx.recieved_data[1] ),
    .A2(_01593_),
    .A1(net29));
 sg13g2_nand4_1 _07935_ (.B(_02605_),
    .C(_02606_),
    .A(_02604_),
    .Y(_02608_),
    .D(_02607_));
 sg13g2_nand2_1 _07936_ (.Y(_02609_),
    .A(\i_uart_rx.recieved_data[5] ),
    .B(net150));
 sg13g2_a22oi_1 _07937_ (.Y(_02610_),
    .B1(net131),
    .B2(\i_spi.data[5] ),
    .A2(_01593_),
    .A1(net33));
 sg13g2_a221oi_1 _07938_ (.B2(_01258_),
    .C1(net207),
    .B1(_02192_),
    .A1(\gpio_out_sel[5] ),
    .Y(_02611_),
    .A2(net167));
 sg13g2_and3_1 _07939_ (.X(_02612_),
    .A(_02609_),
    .B(_02610_),
    .C(_02611_));
 sg13g2_nor3_1 _07940_ (.A(net186),
    .B(net201),
    .C(_02612_),
    .Y(_02613_));
 sg13g2_a22oi_1 _07941_ (.Y(_02614_),
    .B1(_02608_),
    .B2(_02613_),
    .A2(_02602_),
    .A1(net166));
 sg13g2_o21ai_1 _07942_ (.B1(_02262_),
    .Y(_02615_),
    .A1(_02254_),
    .A2(_02614_));
 sg13g2_nand2_1 _07943_ (.Y(_02616_),
    .A(net288),
    .B(_02265_));
 sg13g2_and4_1 _07944_ (.A(net255),
    .B(net258),
    .C(net256),
    .D(_02278_),
    .X(_02617_));
 sg13g2_buf_1 _07945_ (.A(_02617_),
    .X(_02618_));
 sg13g2_nand2_1 _07946_ (.Y(_02619_),
    .A(_02286_),
    .B(_02618_));
 sg13g2_nor2_1 _07947_ (.A(_02616_),
    .B(_02619_),
    .Y(_02620_));
 sg13g2_xor2_1 _07948_ (.B(_02620_),
    .A(net252),
    .X(_02621_));
 sg13g2_nand4_1 _07949_ (.B(net258),
    .C(net256),
    .A(_02291_),
    .Y(_02622_),
    .D(net304));
 sg13g2_nor3_1 _07950_ (.A(_02284_),
    .B(_02269_),
    .C(_02622_),
    .Y(_02623_));
 sg13g2_xor2_1 _07951_ (.B(_02623_),
    .A(_02276_),
    .X(_02624_));
 sg13g2_mux2_1 _07952_ (.A0(_02621_),
    .A1(_02624_),
    .S(net204),
    .X(_02625_));
 sg13g2_xnor2_1 _07953_ (.Y(_02626_),
    .A(net256),
    .B(_02286_));
 sg13g2_mux2_1 _07954_ (.A0(_01291_),
    .A1(_02626_),
    .S(net187),
    .X(_02627_));
 sg13g2_nand2_1 _07955_ (.Y(_02628_),
    .A(_00757_),
    .B(_02627_));
 sg13g2_o21ai_1 _07956_ (.B1(_02628_),
    .Y(_02629_),
    .A1(_00757_),
    .A2(_02625_));
 sg13g2_and2_1 _07957_ (.A(_01138_),
    .B(_02302_),
    .X(_02630_));
 sg13g2_buf_1 _07958_ (.A(_02630_),
    .X(_02631_));
 sg13g2_nand3_1 _07959_ (.B(_02618_),
    .C(_02631_),
    .A(_02310_),
    .Y(_02632_));
 sg13g2_nor3_1 _07960_ (.A(_02284_),
    .B(_02269_),
    .C(_02632_),
    .Y(_02633_));
 sg13g2_xnor2_1 _07961_ (.Y(_02634_),
    .A(net307),
    .B(_02633_));
 sg13g2_nand2_1 _07962_ (.Y(_02635_),
    .A(net253),
    .B(_01137_));
 sg13g2_nand3_1 _07963_ (.B(_02286_),
    .C(_02618_),
    .A(_02310_),
    .Y(_02636_));
 sg13g2_buf_1 _07964_ (.A(_02636_),
    .X(_02637_));
 sg13g2_nor2_1 _07965_ (.A(_02635_),
    .B(_02637_),
    .Y(_02638_));
 sg13g2_xor2_1 _07966_ (.B(_02638_),
    .A(net308),
    .X(_02639_));
 sg13g2_nor2_1 _07967_ (.A(net187),
    .B(_02639_),
    .Y(_02640_));
 sg13g2_a21oi_1 _07968_ (.A1(net185),
    .A2(_02634_),
    .Y(_02641_),
    .B1(_02640_));
 sg13g2_a21oi_1 _07969_ (.A1(_00088_),
    .A2(_02641_),
    .Y(_02642_),
    .B1(net202));
 sg13g2_a21oi_1 _07970_ (.A1(net202),
    .A2(_02629_),
    .Y(_02643_),
    .B1(_02642_));
 sg13g2_buf_1 _07971_ (.A(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .X(_02644_));
 sg13g2_mux2_1 _07972_ (.A0(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .A1(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .S(net172),
    .X(_02645_));
 sg13g2_a22oi_1 _07973_ (.Y(_02646_),
    .B1(_02346_),
    .B2(_02645_),
    .A2(_02337_),
    .A1(_02644_));
 sg13g2_a22oi_1 _07974_ (.Y(_02647_),
    .B1(_02369_),
    .B2(\i_tinyqv.cpu.i_core.mie[17] ),
    .A2(_02341_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[1] ));
 sg13g2_nand3_1 _07975_ (.B(net157),
    .C(_02340_),
    .A(\i_tinyqv.cpu.i_core.mcause[1] ),
    .Y(_02648_));
 sg13g2_a22oi_1 _07976_ (.Y(_02649_),
    .B1(_02359_),
    .B2(_01370_),
    .A2(_02356_),
    .A1(\i_tinyqv.cpu.i_core.mepc[1] ));
 sg13g2_nand4_1 _07977_ (.B(_02647_),
    .C(_02648_),
    .A(_02646_),
    .Y(_02650_),
    .D(_02649_));
 sg13g2_a22oi_1 _07978_ (.Y(_02651_),
    .B1(_02650_),
    .B2(_02353_),
    .A2(_02643_),
    .A1(_01274_));
 sg13g2_nor2_1 _07979_ (.A(_01096_),
    .B(_02374_),
    .Y(_02652_));
 sg13g2_a21oi_1 _07980_ (.A1(_02374_),
    .A2(_02651_),
    .Y(_02653_),
    .B1(_02652_));
 sg13g2_mux2_1 _07981_ (.A0(_02615_),
    .A1(_02653_),
    .S(_01535_),
    .X(_02654_));
 sg13g2_nor2_1 _07982_ (.A(net189),
    .B(_02654_),
    .Y(_02655_));
 sg13g2_a21oi_1 _07983_ (.A1(net189),
    .A2(_02579_),
    .Y(_02656_),
    .B1(_02655_));
 sg13g2_buf_1 _07984_ (.A(_02656_),
    .X(_02657_));
 sg13g2_buf_1 _07985_ (.A(_02657_),
    .X(\debug_rd[1] ));
 sg13g2_mux2_1 _07986_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .A1(net63),
    .S(_02528_),
    .X(_00051_));
 sg13g2_mux2_1 _07987_ (.A0(_02572_),
    .A1(_02561_),
    .S(_02413_),
    .X(_02658_));
 sg13g2_a21o_1 _07988_ (.A2(_01749_),
    .A1(_01734_),
    .B1(_01747_),
    .X(_02659_));
 sg13g2_nand2_1 _07989_ (.Y(_02660_),
    .A(_01751_),
    .B(_02659_));
 sg13g2_xnor2_1 _07990_ (.Y(_02661_),
    .A(_00827_),
    .B(_00927_));
 sg13g2_xor2_1 _07991_ (.B(_02661_),
    .A(_00822_),
    .X(_02662_));
 sg13g2_xnor2_1 _07992_ (.Y(_02663_),
    .A(_01161_),
    .B(_02662_));
 sg13g2_nand2_1 _07993_ (.Y(_02664_),
    .A(_02392_),
    .B(_02663_));
 sg13g2_mux2_1 _07994_ (.A0(_02400_),
    .A1(_02395_),
    .S(_00927_),
    .X(_02665_));
 sg13g2_nand2b_1 _07995_ (.Y(_02666_),
    .B(_02665_),
    .A_N(_00822_));
 sg13g2_nand3_1 _07996_ (.B(_00822_),
    .C(_02400_),
    .A(_00927_),
    .Y(_02667_));
 sg13g2_nand3_1 _07997_ (.B(_02666_),
    .C(_02667_),
    .A(_02664_),
    .Y(_02668_));
 sg13g2_nand2_1 _07998_ (.Y(_02669_),
    .A(net184),
    .B(_02668_));
 sg13g2_o21ai_1 _07999_ (.B1(_02669_),
    .Y(_02670_),
    .A1(net184),
    .A2(_02660_));
 sg13g2_nor2_1 _08000_ (.A(_02408_),
    .B(_02670_),
    .Y(_02671_));
 sg13g2_a21oi_1 _08001_ (.A1(_02408_),
    .A2(_02658_),
    .Y(_02672_),
    .B1(_02671_));
 sg13g2_nor2_1 _08002_ (.A(_02454_),
    .B(_02577_),
    .Y(_02673_));
 sg13g2_a21oi_1 _08003_ (.A1(_02529_),
    .A2(_02672_),
    .Y(_02674_),
    .B1(_02673_));
 sg13g2_buf_1 _08004_ (.A(\i_tinyqv.cpu.instr_data_in[10] ),
    .X(_02675_));
 sg13g2_buf_1 _08005_ (.A(\i_tinyqv.cpu.instr_data_in[14] ),
    .X(_02676_));
 sg13g2_mux4_1 _08006_ (.S0(net205),
    .A0(\i_tinyqv.mem.qspi_data_buf[26] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[30] ),
    .A2(_02675_),
    .A3(_02676_),
    .S1(_01563_),
    .X(_02677_));
 sg13g2_mux2_1 _08007_ (.A0(\i_tinyqv.mem.data_from_read[18] ),
    .A1(\i_tinyqv.mem.data_from_read[22] ),
    .S(net187),
    .X(_02678_));
 sg13g2_mux2_1 _08008_ (.A0(_02677_),
    .A1(_02678_),
    .S(net211),
    .X(_02679_));
 sg13g2_o21ai_1 _08009_ (.B1(net166),
    .Y(_02680_),
    .A1(_01227_),
    .A2(_02679_));
 sg13g2_buf_1 _08010_ (.A(\i_tinyqv.cpu.instr_data_in[2] ),
    .X(_02681_));
 sg13g2_buf_1 _08011_ (.A(\i_tinyqv.cpu.instr_data_in[6] ),
    .X(_02682_));
 sg13g2_and2_1 _08012_ (.A(net205),
    .B(_02682_),
    .X(_02683_));
 sg13g2_a21oi_1 _08013_ (.A1(net204),
    .A2(_02681_),
    .Y(_02684_),
    .B1(_02683_));
 sg13g2_mux2_1 _08014_ (.A0(_02675_),
    .A1(_02676_),
    .S(net205),
    .X(_02685_));
 sg13g2_nand2_1 _08015_ (.Y(_02686_),
    .A(_02242_),
    .B(_02685_));
 sg13g2_o21ai_1 _08016_ (.B1(_02686_),
    .Y(_02687_),
    .A1(_02242_),
    .A2(_02684_));
 sg13g2_and2_1 _08017_ (.A(net187),
    .B(\i_tinyqv.mem.qspi_data_buf[14] ),
    .X(_02688_));
 sg13g2_a21oi_1 _08018_ (.A1(net207),
    .A2(\i_tinyqv.mem.qspi_data_buf[10] ),
    .Y(_02689_),
    .B1(_02688_));
 sg13g2_a22oi_1 _08019_ (.Y(_02690_),
    .B1(_02689_),
    .B2(net186),
    .A2(_02242_),
    .A1(_01235_));
 sg13g2_o21ai_1 _08020_ (.B1(_02690_),
    .Y(_02691_),
    .A1(net186),
    .A2(_02687_));
 sg13g2_nand3_1 _08021_ (.B(_02242_),
    .C(_02685_),
    .A(net203),
    .Y(_02692_));
 sg13g2_o21ai_1 _08022_ (.B1(_02692_),
    .Y(_02693_),
    .A1(net203),
    .A2(_02684_));
 sg13g2_a21oi_1 _08023_ (.A1(_01235_),
    .A2(_02693_),
    .Y(_02694_),
    .B1(_02248_));
 sg13g2_a221oi_1 _08024_ (.B2(net4),
    .C1(_02233_),
    .B1(_02192_),
    .A1(\i_uart_rx.recieved_data[2] ),
    .Y(_02695_),
    .A2(net150));
 sg13g2_and2_1 _08025_ (.A(\gpio_out_sel[2] ),
    .B(net167),
    .X(_02696_));
 sg13g2_a221oi_1 _08026_ (.B2(\i_spi.data[2] ),
    .C1(_02696_),
    .B1(net131),
    .A1(net30),
    .Y(_02697_),
    .A2(_01593_));
 sg13g2_and2_1 _08027_ (.A(\gpio_out_sel[6] ),
    .B(net167),
    .X(_02698_));
 sg13g2_a221oi_1 _08028_ (.B2(\i_spi.data[6] ),
    .C1(_02698_),
    .B1(net131),
    .A1(net34),
    .Y(_02699_),
    .A2(_01593_));
 sg13g2_a221oi_1 _08029_ (.B2(net6),
    .C1(net207),
    .B1(_02192_),
    .A1(\i_uart_rx.recieved_data[6] ),
    .Y(_02700_),
    .A2(net150));
 sg13g2_a221oi_1 _08030_ (.B2(_02700_),
    .C1(net203),
    .B1(_02699_),
    .A1(_02695_),
    .Y(_02701_),
    .A2(_02697_));
 sg13g2_inv_1 _08031_ (.Y(_02702_),
    .A(_02250_));
 sg13g2_o21ai_1 _08032_ (.B1(_02702_),
    .Y(_02703_),
    .A1(net227),
    .A2(_02251_));
 sg13g2_o21ai_1 _08033_ (.B1(_02703_),
    .Y(_02704_),
    .A1(_02220_),
    .A2(_02701_));
 sg13g2_a221oi_1 _08034_ (.B2(_02694_),
    .C1(_02704_),
    .B1(_02691_),
    .A1(net201),
    .Y(_02705_),
    .A2(_02680_));
 sg13g2_a21oi_1 _08035_ (.A1(\i_tinyqv.cpu.i_core.load_top_bit ),
    .A2(_02254_),
    .Y(_02706_),
    .B1(_02705_));
 sg13g2_nand2_1 _08036_ (.Y(_02707_),
    .A(_02276_),
    .B(net304));
 sg13g2_nor2_1 _08037_ (.A(_02707_),
    .B(_02273_),
    .Y(_02708_));
 sg13g2_xnor2_1 _08038_ (.Y(_02709_),
    .A(net257),
    .B(_02708_));
 sg13g2_and2_1 _08039_ (.A(_02294_),
    .B(_02307_),
    .X(_02710_));
 sg13g2_xor2_1 _08040_ (.B(_02710_),
    .A(net254),
    .X(_02711_));
 sg13g2_nand2_1 _08041_ (.Y(_02712_),
    .A(net187),
    .B(_02711_));
 sg13g2_o21ai_1 _08042_ (.B1(_02712_),
    .Y(_02713_),
    .A1(net187),
    .A2(_02709_));
 sg13g2_xnor2_1 _08043_ (.Y(_02714_),
    .A(net258),
    .B(_02271_));
 sg13g2_nand2_1 _08044_ (.Y(_02715_),
    .A(_02222_),
    .B(_02714_));
 sg13g2_o21ai_1 _08045_ (.B1(_02715_),
    .Y(_02716_),
    .A1(_02223_),
    .A2(_01300_));
 sg13g2_nor2_1 _08046_ (.A(net203),
    .B(_02716_),
    .Y(_02717_));
 sg13g2_a21oi_1 _08047_ (.A1(net203),
    .A2(_02713_),
    .Y(_02718_),
    .B1(_02717_));
 sg13g2_inv_2 _08048_ (.Y(_02719_),
    .A(_00760_));
 sg13g2_nand4_1 _08049_ (.B(_02296_),
    .C(_02271_),
    .A(net307),
    .Y(_02720_),
    .D(_02631_));
 sg13g2_xnor2_1 _08050_ (.Y(_02721_),
    .A(_02719_),
    .B(_02720_));
 sg13g2_nand4_1 _08051_ (.B(_02296_),
    .C(_02299_),
    .A(net308),
    .Y(_02722_),
    .D(_02271_));
 sg13g2_xnor2_1 _08052_ (.Y(_02723_),
    .A(net286),
    .B(_02722_));
 sg13g2_nand2_1 _08053_ (.Y(_02724_),
    .A(net204),
    .B(_02723_));
 sg13g2_o21ai_1 _08054_ (.B1(_02724_),
    .Y(_02725_),
    .A1(net207),
    .A2(_02721_));
 sg13g2_a21oi_1 _08055_ (.A1(_00088_),
    .A2(_02725_),
    .Y(_02726_),
    .B1(net202));
 sg13g2_a21oi_1 _08056_ (.A1(_02247_),
    .A2(_02718_),
    .Y(_02727_),
    .B1(_02726_));
 sg13g2_buf_1 _08057_ (.A(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .X(_02728_));
 sg13g2_a21o_1 _08058_ (.A2(_02344_),
    .A1(_02728_),
    .B1(_02333_),
    .X(_02729_));
 sg13g2_a21o_1 _08059_ (.A2(_02346_),
    .A1(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .B1(_02333_),
    .X(_02730_));
 sg13g2_a22oi_1 _08060_ (.Y(_02731_),
    .B1(_02730_),
    .B2(net172),
    .A2(_02729_),
    .A1(_01057_));
 sg13g2_a22oi_1 _08061_ (.Y(_02732_),
    .B1(_02359_),
    .B2(_01381_),
    .A2(_02356_),
    .A1(\i_tinyqv.cpu.i_core.mepc[2] ));
 sg13g2_buf_1 _08062_ (.A(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .X(_02733_));
 sg13g2_and2_1 _08063_ (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .B(net168),
    .X(_02734_));
 sg13g2_a22oi_1 _08064_ (.Y(_02735_),
    .B1(_02346_),
    .B2(_02734_),
    .A2(_02337_),
    .A1(_02733_));
 sg13g2_a22oi_1 _08065_ (.Y(_02736_),
    .B1(_02369_),
    .B2(_01374_),
    .A2(_02341_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[2] ));
 sg13g2_nand4_1 _08066_ (.B(_02732_),
    .C(_02735_),
    .A(_02731_),
    .Y(_02737_),
    .D(_02736_));
 sg13g2_a22oi_1 _08067_ (.Y(_02738_),
    .B1(_02737_),
    .B2(_02353_),
    .A2(_02727_),
    .A1(_01274_));
 sg13g2_nor2_1 _08068_ (.A(_00924_),
    .B(_02374_),
    .Y(_02739_));
 sg13g2_a21oi_1 _08069_ (.A1(_02374_),
    .A2(_02738_),
    .Y(_02740_),
    .B1(_02739_));
 sg13g2_nand2_1 _08070_ (.Y(_02741_),
    .A(_01535_),
    .B(_02740_));
 sg13g2_o21ai_1 _08071_ (.B1(_02741_),
    .Y(_02742_),
    .A1(_01535_),
    .A2(_02706_));
 sg13g2_nor2_1 _08072_ (.A(net189),
    .B(_02742_),
    .Y(_02743_));
 sg13g2_a21oi_1 _08073_ (.A1(net189),
    .A2(_02674_),
    .Y(_02744_),
    .B1(_02743_));
 sg13g2_buf_1 _08074_ (.A(_02744_),
    .X(_02745_));
 sg13g2_buf_1 _08075_ (.A(_02745_),
    .X(\debug_rd[2] ));
 sg13g2_mux2_1 _08076_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .A1(net57),
    .S(_02528_),
    .X(_00052_));
 sg13g2_xor2_1 _08077_ (.B(_02637_),
    .A(net253),
    .X(_02746_));
 sg13g2_xnor2_1 _08078_ (.Y(_02747_),
    .A(net288),
    .B(_02619_));
 sg13g2_nand2_1 _08079_ (.Y(_02748_),
    .A(net204),
    .B(_02747_));
 sg13g2_o21ai_1 _08080_ (.B1(_02748_),
    .Y(_02749_),
    .A1(_02225_),
    .A2(_02746_));
 sg13g2_xnor2_1 _08081_ (.Y(_02750_),
    .A(net312),
    .B(_01403_));
 sg13g2_and2_1 _08082_ (.A(_02225_),
    .B(_02750_),
    .X(_02751_));
 sg13g2_nor2_1 _08083_ (.A(_00964_),
    .B(net255),
    .Y(_02752_));
 sg13g2_nand3_1 _08084_ (.B(net256),
    .C(_02286_),
    .A(net258),
    .Y(_02753_));
 sg13g2_mux2_1 _08085_ (.A0(net255),
    .A1(_02752_),
    .S(_02753_),
    .X(_02754_));
 sg13g2_nor3_1 _08086_ (.A(_02231_),
    .B(_02751_),
    .C(_02754_),
    .Y(_02755_));
 sg13g2_a21oi_1 _08087_ (.A1(_02231_),
    .A2(_02749_),
    .Y(_02756_),
    .B1(_02755_));
 sg13g2_nand4_1 _08088_ (.B(_02310_),
    .C(_02286_),
    .A(_02301_),
    .Y(_02757_),
    .D(_02618_));
 sg13g2_xor2_1 _08089_ (.B(_02757_),
    .A(_00859_),
    .X(_02758_));
 sg13g2_nand3_1 _08090_ (.B(net307),
    .C(_02631_),
    .A(_00760_),
    .Y(_02759_));
 sg13g2_nor2_1 _08091_ (.A(_02637_),
    .B(_02759_),
    .Y(_02760_));
 sg13g2_xnor2_1 _08092_ (.Y(_02761_),
    .A(_00160_),
    .B(_02760_));
 sg13g2_nand2_1 _08093_ (.Y(_02762_),
    .A(_02223_),
    .B(_02761_));
 sg13g2_o21ai_1 _08094_ (.B1(_02762_),
    .Y(_02763_),
    .A1(_02233_),
    .A2(_02758_));
 sg13g2_nand3_1 _08095_ (.B(_00088_),
    .C(_02763_),
    .A(_00766_),
    .Y(_02764_));
 sg13g2_o21ai_1 _08096_ (.B1(_02764_),
    .Y(_02765_),
    .A1(_02264_),
    .A2(_02756_));
 sg13g2_mux2_1 _08097_ (.A0(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .A1(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .S(net172),
    .X(_02766_));
 sg13g2_a22oi_1 _08098_ (.Y(_02767_),
    .B1(_02346_),
    .B2(_02766_),
    .A2(_02341_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[3] ));
 sg13g2_a22oi_1 _08099_ (.Y(_02768_),
    .B1(_02369_),
    .B2(_01390_),
    .A2(_02337_),
    .A1(_02366_));
 sg13g2_nand2_1 _08100_ (.Y(_02769_),
    .A(net209),
    .B(_02359_));
 sg13g2_a22oi_1 _08101_ (.Y(_02770_),
    .B1(net172),
    .B2(\i_tinyqv.cpu.i_core.mcause[4] ),
    .A2(_01057_),
    .A1(\i_tinyqv.cpu.i_core.mcause[3] ));
 sg13g2_inv_1 _08102_ (.Y(_02771_),
    .A(_02770_));
 sg13g2_a22oi_1 _08103_ (.Y(_02772_),
    .B1(_02364_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .A2(_01057_),
    .A1(\i_tinyqv.cpu.i_core.mstatus_mie ));
 sg13g2_nor2b_1 _08104_ (.A(_02772_),
    .B_N(_02344_),
    .Y(_02773_));
 sg13g2_a221oi_1 _08105_ (.B2(_02340_),
    .C1(_02773_),
    .B1(_02771_),
    .A1(\i_tinyqv.cpu.i_core.mepc[3] ),
    .Y(_02774_),
    .A2(_02356_));
 sg13g2_nand4_1 _08106_ (.B(_02768_),
    .C(_02769_),
    .A(_02767_),
    .Y(_02775_),
    .D(_02774_));
 sg13g2_a22oi_1 _08107_ (.Y(_02776_),
    .B1(_02775_),
    .B2(_02353_),
    .A2(_02765_),
    .A1(_01274_));
 sg13g2_nand2_1 _08108_ (.Y(_02777_),
    .A(_02374_),
    .B(_02776_));
 sg13g2_o21ai_1 _08109_ (.B1(_02777_),
    .Y(_02778_),
    .A1(_00975_),
    .A2(_02374_));
 sg13g2_a21o_1 _08110_ (.A2(_02778_),
    .A1(_01535_),
    .B1(net189),
    .X(_02779_));
 sg13g2_buf_1 _08111_ (.A(\i_tinyqv.cpu.instr_data_in[15] ),
    .X(_02780_));
 sg13g2_buf_1 _08112_ (.A(\i_tinyqv.cpu.instr_data_in[7] ),
    .X(_02781_));
 sg13g2_nand2_1 _08113_ (.Y(_02782_),
    .A(_01508_),
    .B(_02242_));
 sg13g2_mux2_1 _08114_ (.A0(_02780_),
    .A1(_02781_),
    .S(_02782_),
    .X(_02783_));
 sg13g2_o21ai_1 _08115_ (.B1(_01145_),
    .Y(_02784_),
    .A1(_01227_),
    .A2(_02783_));
 sg13g2_a21oi_1 _08116_ (.A1(_01256_),
    .A2(net167),
    .Y(_02785_),
    .B1(net166));
 sg13g2_nand2_1 _08117_ (.Y(_02786_),
    .A(net7),
    .B(_02192_));
 sg13g2_a22oi_1 _08118_ (.Y(_02787_),
    .B1(net131),
    .B2(\i_spi.data[7] ),
    .A2(net150),
    .A1(\i_uart_rx.recieved_data[7] ));
 sg13g2_nand3_1 _08119_ (.B(_02786_),
    .C(_02787_),
    .A(_02785_),
    .Y(_02788_));
 sg13g2_nand2b_1 _08120_ (.Y(_02789_),
    .B(_02788_),
    .A_N(_02784_));
 sg13g2_buf_1 _08121_ (.A(\i_tinyqv.cpu.instr_data_in[11] ),
    .X(_02790_));
 sg13g2_buf_1 _08122_ (.A(\i_tinyqv.cpu.instr_data_in[3] ),
    .X(_02791_));
 sg13g2_mux2_1 _08123_ (.A0(_02790_),
    .A1(_02791_),
    .S(_02782_),
    .X(_02792_));
 sg13g2_nand2_1 _08124_ (.Y(_02793_),
    .A(\i_uart_rx.recieved_data[3] ),
    .B(net150));
 sg13g2_a22oi_1 _08125_ (.Y(_02794_),
    .B1(_02185_),
    .B2(\i_spi.data[3] ),
    .A2(_01593_),
    .A1(net31));
 sg13g2_a221oi_1 _08126_ (.B2(net316),
    .C1(net166),
    .B1(_02192_),
    .A1(\gpio_out_sel[3] ),
    .Y(_02795_),
    .A2(net167));
 sg13g2_nand3_1 _08127_ (.B(_02794_),
    .C(_02795_),
    .A(_02793_),
    .Y(_02796_));
 sg13g2_and2_1 _08128_ (.A(_01055_),
    .B(_02796_),
    .X(_02797_));
 sg13g2_o21ai_1 _08129_ (.B1(_02797_),
    .Y(_02798_),
    .A1(_01227_),
    .A2(_02792_));
 sg13g2_mux4_1 _08130_ (.S0(net205),
    .A0(_02790_),
    .A1(_02780_),
    .A2(\i_tinyqv.mem.qspi_data_buf[11] ),
    .A3(\i_tinyqv.mem.qspi_data_buf[15] ),
    .S1(_02243_),
    .X(_02799_));
 sg13g2_and2_1 _08131_ (.A(net220),
    .B(net166),
    .X(_02800_));
 sg13g2_o21ai_1 _08132_ (.B1(_02800_),
    .Y(_02801_),
    .A1(_01227_),
    .A2(_02799_));
 sg13g2_nand4_1 _08133_ (.B(_02789_),
    .C(_02798_),
    .A(net202),
    .Y(_02802_),
    .D(_02801_));
 sg13g2_nor2_1 _08134_ (.A(_01256_),
    .B(_02802_),
    .Y(_02803_));
 sg13g2_and2_1 _08135_ (.A(_01571_),
    .B(_02803_),
    .X(_02804_));
 sg13g2_mux4_1 _08136_ (.S0(net185),
    .A0(\i_tinyqv.mem.qspi_data_buf[27] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[31] ),
    .A2(_02790_),
    .A3(_02780_),
    .S1(_01563_),
    .X(_02805_));
 sg13g2_mux2_1 _08137_ (.A0(\i_tinyqv.mem.data_from_read[19] ),
    .A1(\i_tinyqv.mem.data_from_read[23] ),
    .S(net185),
    .X(_02806_));
 sg13g2_mux2_1 _08138_ (.A0(_02805_),
    .A1(_02806_),
    .S(net188),
    .X(_02807_));
 sg13g2_o21ai_1 _08139_ (.B1(net166),
    .Y(_02808_),
    .A1(_01227_),
    .A2(_02807_));
 sg13g2_nand2b_1 _08140_ (.Y(_02809_),
    .B(_01256_),
    .A_N(\gpio_out[7] ));
 sg13g2_inv_1 _08141_ (.Y(_02810_),
    .A(_01593_));
 sg13g2_nor2_1 _08142_ (.A(_02810_),
    .B(_02784_),
    .Y(_02811_));
 sg13g2_a21oi_1 _08143_ (.A1(_02809_),
    .A2(_02811_),
    .Y(_02812_),
    .B1(_02802_));
 sg13g2_a221oi_1 _08144_ (.B2(net201),
    .C1(_02812_),
    .B1(_02808_),
    .A1(_01549_),
    .Y(_02813_),
    .A2(_02804_));
 sg13g2_a21oi_1 _08145_ (.A1(_02703_),
    .A2(_02813_),
    .Y(_02814_),
    .B1(_02263_));
 sg13g2_mux2_1 _08146_ (.A0(_02395_),
    .A1(_02400_),
    .S(_00867_),
    .X(_02815_));
 sg13g2_nor2_1 _08147_ (.A(_00978_),
    .B(_00867_),
    .Y(_02816_));
 sg13g2_nor2_1 _08148_ (.A(_01161_),
    .B(_02661_),
    .Y(_02817_));
 sg13g2_nor2_1 _08149_ (.A(_00822_),
    .B(_02817_),
    .Y(_02818_));
 sg13g2_a21oi_1 _08150_ (.A1(_01161_),
    .A2(_02661_),
    .Y(_02819_),
    .B1(_02818_));
 sg13g2_xnor2_1 _08151_ (.Y(_02820_),
    .A(_01264_),
    .B(_02819_));
 sg13g2_nor2_1 _08152_ (.A(_02401_),
    .B(_02820_),
    .Y(_02821_));
 sg13g2_a221oi_1 _08153_ (.B2(_02400_),
    .C1(_02821_),
    .B1(_02816_),
    .A1(_00978_),
    .Y(_02822_),
    .A2(_02815_));
 sg13g2_a21oi_1 _08154_ (.A1(_00823_),
    .A2(_01176_),
    .Y(_02823_),
    .B1(_02408_));
 sg13g2_mux2_1 _08155_ (.A0(_02510_),
    .A1(_02482_),
    .S(net250),
    .X(_02824_));
 sg13g2_xnor2_1 _08156_ (.Y(_02825_),
    .A(_01732_),
    .B(_01758_));
 sg13g2_xor2_1 _08157_ (.B(_01751_),
    .A(_01707_),
    .X(_02826_));
 sg13g2_xnor2_1 _08158_ (.Y(_02827_),
    .A(_02825_),
    .B(_02826_));
 sg13g2_nor2_1 _08159_ (.A(net184),
    .B(_02827_),
    .Y(_02828_));
 sg13g2_a221oi_1 _08160_ (.B2(_02408_),
    .C1(_02828_),
    .B1(_02824_),
    .A1(_02822_),
    .Y(_02829_),
    .A2(_02823_));
 sg13g2_and2_1 _08161_ (.A(_02529_),
    .B(_02829_),
    .X(_02830_));
 sg13g2_nor2_1 _08162_ (.A(_02429_),
    .B(_02577_),
    .Y(_02831_));
 sg13g2_o21ai_1 _08163_ (.B1(net189),
    .Y(_02832_),
    .A1(_02830_),
    .A2(_02831_));
 sg13g2_o21ai_1 _08164_ (.B1(_02832_),
    .Y(_02833_),
    .A1(_02779_),
    .A2(_02814_));
 sg13g2_buf_2 _08165_ (.A(_02833_),
    .X(_02834_));
 sg13g2_buf_8 _08166_ (.A(_02834_),
    .X(\debug_rd[3] ));
 sg13g2_mux2_1 _08167_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .A1(net44),
    .S(_02528_),
    .X(_00053_));
 sg13g2_nand2b_1 _08168_ (.Y(_02835_),
    .B(_02520_),
    .A_N(_02521_));
 sg13g2_buf_1 _08169_ (.A(_02835_),
    .X(_02836_));
 sg13g2_nor2_2 _08170_ (.A(_02527_),
    .B(_02836_),
    .Y(_02837_));
 sg13g2_mux2_1 _08171_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .A1(net64),
    .S(_02837_),
    .X(_00046_));
 sg13g2_mux2_1 _08172_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .A1(net63),
    .S(_02837_),
    .X(_00047_));
 sg13g2_mux2_1 _08173_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .A1(net57),
    .S(_02837_),
    .X(_00048_));
 sg13g2_mux2_1 _08174_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .A1(net44),
    .S(_02837_),
    .X(_00049_));
 sg13g2_inv_1 _08175_ (.Y(_02838_),
    .A(_02520_));
 sg13g2_nand2_2 _08176_ (.Y(_02839_),
    .A(_02838_),
    .B(_02521_));
 sg13g2_nor2_2 _08177_ (.A(_02527_),
    .B(_02839_),
    .Y(_02840_));
 sg13g2_mux2_1 _08178_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .A1(net64),
    .S(_02840_),
    .X(_00042_));
 sg13g2_mux2_1 _08179_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .A1(net63),
    .S(_02840_),
    .X(_00043_));
 sg13g2_mux2_1 _08180_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .A1(net57),
    .S(_02840_),
    .X(_00044_));
 sg13g2_mux2_1 _08181_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .A1(net44),
    .S(_02840_),
    .X(_00045_));
 sg13g2_nor3_2 _08182_ (.A(_02520_),
    .B(_02521_),
    .C(_02527_),
    .Y(_02841_));
 sg13g2_mux2_1 _08183_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .A1(net64),
    .S(_02841_),
    .X(_00038_));
 sg13g2_mux2_1 _08184_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .A1(net63),
    .S(_02841_),
    .X(_00039_));
 sg13g2_mux2_1 _08185_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .A1(net57),
    .S(_02841_),
    .X(_00040_));
 sg13g2_mux2_1 _08186_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .A1(net44),
    .S(_02841_),
    .X(_00041_));
 sg13g2_nand3b_1 _08187_ (.B(_02523_),
    .C(_02524_),
    .Y(_02842_),
    .A_N(_01541_));
 sg13g2_buf_1 _08188_ (.A(_02842_),
    .X(_02843_));
 sg13g2_nor2_2 _08189_ (.A(_02522_),
    .B(_02843_),
    .Y(_02844_));
 sg13g2_mux2_1 _08190_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .A1(net64),
    .S(_02844_),
    .X(_00034_));
 sg13g2_mux2_1 _08191_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A1(net63),
    .S(_02844_),
    .X(_00035_));
 sg13g2_mux2_1 _08192_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .A1(net57),
    .S(_02844_),
    .X(_00036_));
 sg13g2_mux2_1 _08193_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .A1(net44),
    .S(_02844_),
    .X(_00037_));
 sg13g2_nor2_2 _08194_ (.A(_02836_),
    .B(_02843_),
    .Y(_02845_));
 sg13g2_mux2_1 _08195_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .A1(net64),
    .S(_02845_),
    .X(_00030_));
 sg13g2_mux2_1 _08196_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .A1(net63),
    .S(_02845_),
    .X(_00031_));
 sg13g2_mux2_1 _08197_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .A1(net57),
    .S(_02845_),
    .X(_00032_));
 sg13g2_mux2_1 _08198_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .A1(net44),
    .S(_02845_),
    .X(_00033_));
 sg13g2_nor2_2 _08199_ (.A(_02839_),
    .B(_02843_),
    .Y(_02846_));
 sg13g2_mux2_1 _08200_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .A1(_02519_),
    .S(_02846_),
    .X(_00078_));
 sg13g2_mux2_1 _08201_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .A1(_02657_),
    .S(_02846_),
    .X(_00079_));
 sg13g2_mux2_1 _08202_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .A1(_02745_),
    .S(_02846_),
    .X(_00080_));
 sg13g2_mux2_1 _08203_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .A1(_02834_),
    .S(_02846_),
    .X(_00081_));
 sg13g2_or3_1 _08204_ (.A(_02520_),
    .B(_02521_),
    .C(_02843_),
    .X(_02847_));
 sg13g2_buf_1 _08205_ (.A(_02847_),
    .X(_02848_));
 sg13g2_mux2_1 _08206_ (.A0(net64),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .S(_02848_),
    .X(_00074_));
 sg13g2_mux2_1 _08207_ (.A0(net63),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .S(_02848_),
    .X(_00075_));
 sg13g2_mux2_1 _08208_ (.A0(net57),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .S(_02848_),
    .X(_00076_));
 sg13g2_mux2_1 _08209_ (.A0(net44),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .S(_02848_),
    .X(_00077_));
 sg13g2_nor3_1 _08210_ (.A(_02523_),
    .B(_02524_),
    .C(_01541_),
    .Y(_02849_));
 sg13g2_nor2b_1 _08211_ (.A(_02522_),
    .B_N(_02849_),
    .Y(_02850_));
 sg13g2_buf_1 _08212_ (.A(_02850_),
    .X(_02851_));
 sg13g2_mux2_1 _08213_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .A1(_02519_),
    .S(_02851_),
    .X(_00070_));
 sg13g2_mux2_1 _08214_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .A1(_02657_),
    .S(_02851_),
    .X(_00071_));
 sg13g2_mux2_1 _08215_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .A1(_02745_),
    .S(_02851_),
    .X(_00072_));
 sg13g2_mux2_1 _08216_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .A1(_02834_),
    .S(_02851_),
    .X(_00073_));
 sg13g2_nor2b_1 _08217_ (.A(_02836_),
    .B_N(_02849_),
    .Y(_02852_));
 sg13g2_buf_1 _08218_ (.A(_02852_),
    .X(_02853_));
 sg13g2_mux2_1 _08219_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .A1(_02519_),
    .S(_02853_),
    .X(_00066_));
 sg13g2_mux2_1 _08220_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .A1(_02657_),
    .S(_02853_),
    .X(_00067_));
 sg13g2_mux2_1 _08221_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .A1(_02745_),
    .S(_02853_),
    .X(_00068_));
 sg13g2_mux2_1 _08222_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .A1(_02834_),
    .S(_02853_),
    .X(_00069_));
 sg13g2_nor2b_1 _08223_ (.A(_02839_),
    .B_N(_02849_),
    .Y(_02854_));
 sg13g2_buf_1 _08224_ (.A(_02854_),
    .X(_02855_));
 sg13g2_mux2_1 _08225_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .A1(_02519_),
    .S(_02855_),
    .X(_00062_));
 sg13g2_mux2_1 _08226_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .A1(_02657_),
    .S(_02855_),
    .X(_00063_));
 sg13g2_mux2_1 _08227_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .A1(_02745_),
    .S(_02855_),
    .X(_00064_));
 sg13g2_mux2_1 _08228_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .A1(_02834_),
    .S(_02855_),
    .X(_00065_));
 sg13g2_nor3_1 _08229_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .B(_02524_),
    .C(_01541_),
    .Y(_02856_));
 sg13g2_nand2b_1 _08230_ (.Y(_02857_),
    .B(_02856_),
    .A_N(_02836_));
 sg13g2_buf_1 _08231_ (.A(_02857_),
    .X(_02858_));
 sg13g2_mux2_1 _08232_ (.A0(net64),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .S(_02858_),
    .X(_00058_));
 sg13g2_mux2_1 _08233_ (.A0(net63),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .S(_02858_),
    .X(_00059_));
 sg13g2_mux2_1 _08234_ (.A0(net57),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .S(_02858_),
    .X(_00060_));
 sg13g2_mux2_1 _08235_ (.A0(net44),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .S(_02858_),
    .X(_00061_));
 sg13g2_nand2b_1 _08236_ (.Y(_02859_),
    .B(_02856_),
    .A_N(_02839_));
 sg13g2_buf_1 _08237_ (.A(_02859_),
    .X(_02860_));
 sg13g2_mux2_1 _08238_ (.A0(\debug_rd[0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .S(_02860_),
    .X(_00054_));
 sg13g2_mux2_1 _08239_ (.A0(\debug_rd[1] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .S(_02860_),
    .X(_00055_));
 sg13g2_mux2_1 _08240_ (.A0(\debug_rd[2] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .S(_02860_),
    .X(_00056_));
 sg13g2_mux2_1 _08241_ (.A0(\debug_rd[3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .S(_02860_),
    .X(_00057_));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_1 _08243_ (.A(_00156_),
    .X(_02861_));
 sg13g2_buf_1 _08244_ (.A(_02861_),
    .X(_02862_));
 sg13g2_a21oi_1 _08245_ (.A1(_01591_),
    .A2(_02216_),
    .Y(_02863_),
    .B1(_02862_));
 sg13g2_mux2_1 _08246_ (.A0(_01422_),
    .A1(_01574_),
    .S(_01597_),
    .X(_02864_));
 sg13g2_nand2_1 _08247_ (.Y(_02865_),
    .A(_01241_),
    .B(_02863_));
 sg13g2_o21ai_1 _08248_ (.B1(_02865_),
    .Y(_00228_),
    .A1(_02863_),
    .A2(_02864_));
 sg13g2_buf_1 _08249_ (.A(\i_spi.busy ),
    .X(_02866_));
 sg13g2_buf_1 _08250_ (.A(net283),
    .X(_02867_));
 sg13g2_nand2_1 _08251_ (.Y(_02868_),
    .A(net208),
    .B(net131));
 sg13g2_buf_1 _08252_ (.A(_02868_),
    .X(_02869_));
 sg13g2_buf_1 _08253_ (.A(\i_spi.bits_remaining[3] ),
    .X(_02870_));
 sg13g2_nor2b_1 _08254_ (.A(_02870_),
    .B_N(\i_spi.read_latency ),
    .Y(_02871_));
 sg13g2_xor2_1 _08255_ (.B(\i_spi.clock_count[1] ),
    .A(\i_spi.clock_divider[1] ),
    .X(_02872_));
 sg13g2_xor2_1 _08256_ (.B(\i_spi.clock_count[0] ),
    .A(\i_spi.clock_divider[0] ),
    .X(_02873_));
 sg13g2_nor2_2 _08257_ (.A(_02872_),
    .B(_02873_),
    .Y(_02874_));
 sg13g2_o21ai_1 _08258_ (.B1(_02874_),
    .Y(_02875_),
    .A1(_01245_),
    .A2(_02871_));
 sg13g2_a21o_1 _08259_ (.A2(_02875_),
    .A1(net283),
    .B1(net215),
    .X(_02876_));
 sg13g2_nor3_1 _08260_ (.A(_01574_),
    .B(_02869_),
    .C(_02876_),
    .Y(_02877_));
 sg13g2_a21oi_1 _08261_ (.A1(\i_spi.data[0] ),
    .A2(_02869_),
    .Y(_02878_),
    .B1(_02877_));
 sg13g2_nand2_1 _08262_ (.Y(_02879_),
    .A(net283),
    .B(net4));
 sg13g2_nor2_1 _08263_ (.A(_02876_),
    .B(_02879_),
    .Y(_02880_));
 sg13g2_a21oi_1 _08264_ (.A1(\i_spi.data[0] ),
    .A2(_02876_),
    .Y(_02881_),
    .B1(_02880_));
 sg13g2_o21ai_1 _08265_ (.B1(_02881_),
    .Y(_00256_),
    .A1(_02867_),
    .A2(_02878_));
 sg13g2_buf_1 _08266_ (.A(net283),
    .X(_02882_));
 sg13g2_nand2_1 _08267_ (.Y(_02883_),
    .A(net243),
    .B(\i_spi.data[0] ));
 sg13g2_o21ai_1 _08268_ (.B1(_02883_),
    .Y(_02884_),
    .A1(net244),
    .A2(_01601_));
 sg13g2_nand2_1 _08269_ (.Y(_02885_),
    .A(_02207_),
    .B(_02869_));
 sg13g2_nand2_1 _08270_ (.Y(_02886_),
    .A(_01245_),
    .B(_02874_));
 sg13g2_a21oi_1 _08271_ (.A1(net283),
    .A2(_02886_),
    .Y(_02887_),
    .B1(_02861_));
 sg13g2_nand2_1 _08272_ (.Y(_02888_),
    .A(_02885_),
    .B(_02887_));
 sg13g2_buf_2 _08273_ (.A(_02888_),
    .X(_02889_));
 sg13g2_mux2_1 _08274_ (.A0(_02884_),
    .A1(\i_spi.data[1] ),
    .S(_02889_),
    .X(_00257_));
 sg13g2_nand2_1 _08275_ (.Y(_02890_),
    .A(net243),
    .B(\i_spi.data[1] ));
 sg13g2_o21ai_1 _08276_ (.B1(_02890_),
    .Y(_02891_),
    .A1(net244),
    .A2(_01604_));
 sg13g2_mux2_1 _08277_ (.A0(_02891_),
    .A1(\i_spi.data[2] ),
    .S(_02889_),
    .X(_00258_));
 sg13g2_nand2_1 _08278_ (.Y(_02892_),
    .A(net243),
    .B(\i_spi.data[2] ));
 sg13g2_o21ai_1 _08279_ (.B1(_02892_),
    .Y(_02893_),
    .A1(net244),
    .A2(_01607_));
 sg13g2_mux2_1 _08280_ (.A0(_02893_),
    .A1(\i_spi.data[3] ),
    .S(_02889_),
    .X(_00259_));
 sg13g2_nand2_1 _08281_ (.Y(_02894_),
    .A(net243),
    .B(\i_spi.data[3] ));
 sg13g2_o21ai_1 _08282_ (.B1(_02894_),
    .Y(_02895_),
    .A1(net244),
    .A2(_01610_));
 sg13g2_mux2_1 _08283_ (.A0(_02895_),
    .A1(\i_spi.data[4] ),
    .S(_02889_),
    .X(_00260_));
 sg13g2_nand2_1 _08284_ (.Y(_02896_),
    .A(net243),
    .B(\i_spi.data[4] ));
 sg13g2_o21ai_1 _08285_ (.B1(_02896_),
    .Y(_02897_),
    .A1(net244),
    .A2(_01613_));
 sg13g2_mux2_1 _08286_ (.A0(_02897_),
    .A1(\i_spi.data[5] ),
    .S(_02889_),
    .X(_00261_));
 sg13g2_nand2_1 _08287_ (.Y(_02898_),
    .A(net243),
    .B(\i_spi.data[5] ));
 sg13g2_o21ai_1 _08288_ (.B1(_02898_),
    .Y(_02899_),
    .A1(net243),
    .A2(_01617_));
 sg13g2_mux2_1 _08289_ (.A0(_02899_),
    .A1(\i_spi.data[6] ),
    .S(_02889_),
    .X(_00262_));
 sg13g2_nand2_1 _08290_ (.Y(_02900_),
    .A(net283),
    .B(\i_spi.data[6] ));
 sg13g2_o21ai_1 _08291_ (.B1(_02900_),
    .Y(_02901_),
    .A1(net243),
    .A2(_01619_));
 sg13g2_mux2_1 _08292_ (.A0(_02901_),
    .A1(\i_spi.data[7] ),
    .S(_02889_),
    .X(_00263_));
 sg13g2_nand4_1 _08293_ (.B(net261),
    .C(net208),
    .A(_02207_),
    .Y(_02902_),
    .D(net131));
 sg13g2_mux2_1 _08294_ (.A0(\data_to_write[8] ),
    .A1(\i_spi.end_txn_reg ),
    .S(_02902_),
    .X(_00264_));
 sg13g2_mux2_1 _08295_ (.A0(\data_to_write[9] ),
    .A1(\i_spi.spi_dc ),
    .S(_02902_),
    .X(_00267_));
 sg13g2_nand2b_1 _08296_ (.Y(_02903_),
    .B(_01553_),
    .A_N(_01286_));
 sg13g2_buf_1 _08297_ (.A(_02903_),
    .X(_02904_));
 sg13g2_or2_1 _08298_ (.X(_02905_),
    .B(_01289_),
    .A(_01279_));
 sg13g2_and2_1 _08299_ (.A(net172),
    .B(_02905_),
    .X(_02906_));
 sg13g2_buf_1 _08300_ (.A(_02906_),
    .X(_02907_));
 sg13g2_nor2b_1 _08301_ (.A(_01419_),
    .B_N(_02907_),
    .Y(_02908_));
 sg13g2_buf_2 _08302_ (.A(_02908_),
    .X(_02909_));
 sg13g2_nand2_1 _08303_ (.Y(_02910_),
    .A(_02904_),
    .B(_02909_));
 sg13g2_buf_1 _08304_ (.A(_02910_),
    .X(_02911_));
 sg13g2_nor2_1 _08305_ (.A(_01642_),
    .B(net56),
    .Y(_02912_));
 sg13g2_buf_1 _08306_ (.A(_02912_),
    .X(_02913_));
 sg13g2_buf_1 _08307_ (.A(_02913_),
    .X(_02914_));
 sg13g2_buf_1 _08308_ (.A(net43),
    .X(_02915_));
 sg13g2_buf_1 _08309_ (.A(net43),
    .X(_02916_));
 sg13g2_nor2b_1 _08310_ (.A(_01357_),
    .B_N(_01360_),
    .Y(_02917_));
 sg13g2_buf_2 _08311_ (.A(_02917_),
    .X(_02918_));
 sg13g2_nor2_1 _08312_ (.A(_01457_),
    .B(_02918_),
    .Y(_02919_));
 sg13g2_buf_1 _08313_ (.A(_02919_),
    .X(_02920_));
 sg13g2_inv_1 _08314_ (.Y(_02921_),
    .A(_01454_));
 sg13g2_nor2_1 _08315_ (.A(_01345_),
    .B(_01351_),
    .Y(_02922_));
 sg13g2_inv_1 _08316_ (.Y(_02923_),
    .A(_01332_));
 sg13g2_and2_1 _08317_ (.A(_02923_),
    .B(net123),
    .X(_02924_));
 sg13g2_buf_1 _08318_ (.A(_02924_),
    .X(_02925_));
 sg13g2_and2_1 _08319_ (.A(_02922_),
    .B(_02925_),
    .X(_02926_));
 sg13g2_buf_1 _08320_ (.A(_01328_),
    .X(_02927_));
 sg13g2_o21ai_1 _08321_ (.B1(_02927_),
    .Y(_02928_),
    .A1(_01353_),
    .A2(_02926_));
 sg13g2_nand3_1 _08322_ (.B(_02921_),
    .C(_02928_),
    .A(_02920_),
    .Y(_02929_));
 sg13g2_buf_1 _08323_ (.A(_02929_),
    .X(_02930_));
 sg13g2_buf_1 _08324_ (.A(_01465_),
    .X(_02931_));
 sg13g2_buf_1 _08325_ (.A(net117),
    .X(_02932_));
 sg13g2_nor2_2 _08326_ (.A(_01453_),
    .B(_01352_),
    .Y(_02933_));
 sg13g2_nor2b_1 _08327_ (.A(_01347_),
    .B_N(_01349_),
    .Y(_02934_));
 sg13g2_buf_1 _08328_ (.A(_02934_),
    .X(_02935_));
 sg13g2_nand3_1 _08329_ (.B(net123),
    .C(net129),
    .A(_01451_),
    .Y(_02936_));
 sg13g2_buf_1 _08330_ (.A(_02936_),
    .X(_02937_));
 sg13g2_mux2_1 _08331_ (.A0(_00143_),
    .A1(_00144_),
    .S(net152),
    .X(_02938_));
 sg13g2_mux2_1 _08332_ (.A0(_01470_),
    .A1(_02938_),
    .S(_01334_),
    .X(_02939_));
 sg13g2_buf_1 _08333_ (.A(_02939_),
    .X(_02940_));
 sg13g2_nor3_1 _08334_ (.A(net136),
    .B(_02937_),
    .C(_02940_),
    .Y(_02941_));
 sg13g2_nor2_1 _08335_ (.A(_02933_),
    .B(_02941_),
    .Y(_02942_));
 sg13g2_nor2b_1 _08336_ (.A(_01485_),
    .B_N(_01487_),
    .Y(_02943_));
 sg13g2_buf_2 _08337_ (.A(_02943_),
    .X(_02944_));
 sg13g2_buf_1 _08338_ (.A(_02944_),
    .X(_02945_));
 sg13g2_nand2_1 _08339_ (.Y(_02946_),
    .A(net97),
    .B(_02942_));
 sg13g2_o21ai_1 _08340_ (.B1(_02946_),
    .Y(_02947_),
    .A1(net108),
    .A2(_02942_));
 sg13g2_mux4_1 _08341_ (.S0(net159),
    .A0(_00153_),
    .A1(_00152_),
    .A2(_00150_),
    .A3(_00151_),
    .S1(net152),
    .X(_02948_));
 sg13g2_buf_2 _08342_ (.A(_02948_),
    .X(_02949_));
 sg13g2_nor2_1 _08343_ (.A(_01473_),
    .B(_02949_),
    .Y(_02950_));
 sg13g2_nand2_2 _08344_ (.Y(_02951_),
    .A(_01328_),
    .B(_02925_));
 sg13g2_nor2_1 _08345_ (.A(_02944_),
    .B(_02951_),
    .Y(_02952_));
 sg13g2_a21o_1 _08346_ (.A2(_01352_),
    .A1(net97),
    .B1(_02952_),
    .X(_02953_));
 sg13g2_buf_1 _08347_ (.A(_01464_),
    .X(_02954_));
 sg13g2_nor2_1 _08348_ (.A(_01457_),
    .B(_01362_),
    .Y(_02955_));
 sg13g2_buf_1 _08349_ (.A(_02955_),
    .X(_02956_));
 sg13g2_nand2_1 _08350_ (.Y(_02957_),
    .A(_02954_),
    .B(net96));
 sg13g2_a21oi_1 _08351_ (.A1(_02950_),
    .A2(_02953_),
    .Y(_02958_),
    .B1(_02957_));
 sg13g2_buf_1 _08352_ (.A(net107),
    .X(_02959_));
 sg13g2_nor2_1 _08353_ (.A(_01458_),
    .B(net95),
    .Y(_02960_));
 sg13g2_o21ai_1 _08354_ (.B1(_01466_),
    .Y(_02961_),
    .A1(_02958_),
    .A2(_02960_));
 sg13g2_o21ai_1 _08355_ (.B1(_02961_),
    .Y(_02962_),
    .A1(_02930_),
    .A2(_02947_));
 sg13g2_nand2_1 _08356_ (.Y(_02963_),
    .A(net39),
    .B(_02962_));
 sg13g2_o21ai_1 _08357_ (.B1(_02963_),
    .Y(_00272_),
    .A1(_02390_),
    .A2(net40));
 sg13g2_buf_1 _08358_ (.A(net43),
    .X(_02964_));
 sg13g2_nor2b_1 _08359_ (.A(_01318_),
    .B_N(_01320_),
    .Y(_02965_));
 sg13g2_buf_1 _08360_ (.A(_02965_),
    .X(_02966_));
 sg13g2_buf_1 _08361_ (.A(_02966_),
    .X(_02967_));
 sg13g2_buf_1 _08362_ (.A(_01316_),
    .X(_02968_));
 sg13g2_a221oi_1 _08363_ (.B2(_02968_),
    .C1(_02930_),
    .B1(_02942_),
    .A1(net116),
    .Y(_02969_),
    .A2(_02933_));
 sg13g2_nand2_1 _08364_ (.Y(_02970_),
    .A(net95),
    .B(net99));
 sg13g2_nor2_1 _08365_ (.A(_01458_),
    .B(_02970_),
    .Y(_02971_));
 sg13g2_a21oi_1 _08366_ (.A1(net129),
    .A2(net97),
    .Y(_02972_),
    .B1(_02952_));
 sg13g2_nor2_1 _08367_ (.A(_01473_),
    .B(_02972_),
    .Y(_02973_));
 sg13g2_nand3_1 _08368_ (.B(_01466_),
    .C(net96),
    .A(_02954_),
    .Y(_02974_));
 sg13g2_nor3_1 _08369_ (.A(_02949_),
    .B(_02973_),
    .C(_02974_),
    .Y(_02975_));
 sg13g2_nor3_1 _08370_ (.A(_02969_),
    .B(_02971_),
    .C(_02975_),
    .Y(_02976_));
 sg13g2_buf_1 _08371_ (.A(_02913_),
    .X(_02977_));
 sg13g2_nor2_1 _08372_ (.A(_00745_),
    .B(net42),
    .Y(_02978_));
 sg13g2_a21oi_1 _08373_ (.A1(_02964_),
    .A2(_02976_),
    .Y(_00273_),
    .B1(_02978_));
 sg13g2_nor2b_1 _08374_ (.A(_01460_),
    .B_N(_01462_),
    .Y(_02979_));
 sg13g2_buf_1 _08375_ (.A(_02979_),
    .X(_02980_));
 sg13g2_nor2_1 _08376_ (.A(_02980_),
    .B(_02965_),
    .Y(_02981_));
 sg13g2_buf_1 _08377_ (.A(_02981_),
    .X(_02982_));
 sg13g2_and2_1 _08378_ (.A(_02944_),
    .B(_02950_),
    .X(_02983_));
 sg13g2_buf_1 _08379_ (.A(_02983_),
    .X(_02984_));
 sg13g2_nand2_1 _08380_ (.Y(_02985_),
    .A(_02922_),
    .B(_02984_));
 sg13g2_nand2_1 _08381_ (.Y(_02986_),
    .A(net124),
    .B(_02918_));
 sg13g2_nor2_1 _08382_ (.A(_01467_),
    .B(_02986_),
    .Y(_02987_));
 sg13g2_buf_1 _08383_ (.A(_01322_),
    .X(_02988_));
 sg13g2_nand2_1 _08384_ (.Y(_02989_),
    .A(_02988_),
    .B(_02942_));
 sg13g2_buf_1 _08385_ (.A(net152),
    .X(_02990_));
 sg13g2_mux4_1 _08386_ (.S0(net159),
    .A0(_00151_),
    .A1(_00153_),
    .A2(_00152_),
    .A3(_00150_),
    .S1(net127),
    .X(_02991_));
 sg13g2_inv_1 _08387_ (.Y(_02992_),
    .A(_02991_));
 sg13g2_a22oi_1 _08388_ (.Y(_02993_),
    .B1(_02941_),
    .B2(_02992_),
    .A2(_02933_),
    .A1(net116));
 sg13g2_a21oi_1 _08389_ (.A1(_02989_),
    .A2(_02993_),
    .Y(_02994_),
    .B1(_02930_));
 sg13g2_a221oi_1 _08390_ (.B2(_02987_),
    .C1(_02994_),
    .B1(_02985_),
    .A1(_02956_),
    .Y(_02995_),
    .A2(net94));
 sg13g2_nor2_1 _08391_ (.A(net250),
    .B(_02977_),
    .Y(_02996_));
 sg13g2_a21oi_1 _08392_ (.A1(net38),
    .A2(_02995_),
    .Y(_00274_),
    .B1(_02996_));
 sg13g2_a21oi_1 _08393_ (.A1(_02922_),
    .A2(_02945_),
    .Y(_02997_),
    .B1(_02949_));
 sg13g2_nor3_1 _08394_ (.A(_01473_),
    .B(_02974_),
    .C(_02997_),
    .Y(_02998_));
 sg13g2_mux2_1 _08395_ (.A0(_00123_),
    .A1(_00124_),
    .S(_01481_),
    .X(_02999_));
 sg13g2_buf_1 _08396_ (.A(_01334_),
    .X(_03000_));
 sg13g2_mux2_1 _08397_ (.A0(_01317_),
    .A1(_02999_),
    .S(net183),
    .X(_03001_));
 sg13g2_inv_1 _08398_ (.Y(_03002_),
    .A(_03001_));
 sg13g2_o21ai_1 _08399_ (.B1(net136),
    .Y(_03003_),
    .A1(_02932_),
    .A2(net97));
 sg13g2_a21oi_1 _08400_ (.A1(_03002_),
    .A2(_03003_),
    .Y(_03004_),
    .B1(_02941_));
 sg13g2_nor3_1 _08401_ (.A(_02930_),
    .B(_02933_),
    .C(_03004_),
    .Y(_03005_));
 sg13g2_nor3_1 _08402_ (.A(_02971_),
    .B(_02998_),
    .C(_03005_),
    .Y(_03006_));
 sg13g2_nor2_1 _08403_ (.A(net313),
    .B(net42),
    .Y(_03007_));
 sg13g2_a21oi_1 _08404_ (.A1(net38),
    .A2(_03006_),
    .Y(_00275_),
    .B1(_03007_));
 sg13g2_nor2_1 _08405_ (.A(_01642_),
    .B(_01655_),
    .Y(_03008_));
 sg13g2_buf_2 _08406_ (.A(_03008_),
    .X(_03009_));
 sg13g2_buf_1 _08407_ (.A(_03009_),
    .X(_03010_));
 sg13g2_nand4_1 _08408_ (.B(net306),
    .C(_01186_),
    .A(net302),
    .Y(_03011_),
    .D(_01190_));
 sg13g2_buf_1 _08409_ (.A(_03011_),
    .X(_03012_));
 sg13g2_buf_1 _08410_ (.A(_03012_),
    .X(_03013_));
 sg13g2_buf_1 _08411_ (.A(_01276_),
    .X(_03014_));
 sg13g2_and2_1 _08412_ (.A(\i_tinyqv.cpu.i_core.mepc[0] ),
    .B(net148),
    .X(_03015_));
 sg13g2_a21oi_1 _08413_ (.A1(_01765_),
    .A2(net149),
    .Y(_03016_),
    .B1(_03015_));
 sg13g2_nor2_1 _08414_ (.A(\addr[0] ),
    .B(_03009_),
    .Y(_03017_));
 sg13g2_a21oi_1 _08415_ (.A1(net93),
    .A2(_03016_),
    .Y(_00279_),
    .B1(_03017_));
 sg13g2_buf_1 _08416_ (.A(_02108_),
    .X(_03018_));
 sg13g2_mux2_1 _08417_ (.A0(_03018_),
    .A1(\i_tinyqv.cpu.i_core.mepc[10] ),
    .S(net148),
    .X(_03019_));
 sg13g2_mux2_1 _08418_ (.A0(\addr[10] ),
    .A1(_03019_),
    .S(net93),
    .X(_00280_));
 sg13g2_inv_1 _08419_ (.Y(_03020_),
    .A(net291));
 sg13g2_buf_1 _08420_ (.A(_01276_),
    .X(_03021_));
 sg13g2_nand2_1 _08421_ (.Y(_03022_),
    .A(\i_tinyqv.cpu.i_core.mepc[11] ),
    .B(_01276_));
 sg13g2_o21ai_1 _08422_ (.B1(_03022_),
    .Y(_03023_),
    .A1(_03020_),
    .A2(net147));
 sg13g2_mux2_1 _08423_ (.A0(\addr[11] ),
    .A1(_03023_),
    .S(net93),
    .X(_00281_));
 sg13g2_mux2_1 _08424_ (.A0(\i_tinyqv.cpu.i_core.mepc[12] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(net149),
    .X(_03024_));
 sg13g2_mux2_1 _08425_ (.A0(\addr[12] ),
    .A1(_03024_),
    .S(net93),
    .X(_00282_));
 sg13g2_mux2_1 _08426_ (.A0(\i_tinyqv.cpu.i_core.mepc[13] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(net149),
    .X(_03025_));
 sg13g2_mux2_1 _08427_ (.A0(\addr[13] ),
    .A1(_03025_),
    .S(net93),
    .X(_00283_));
 sg13g2_mux2_1 _08428_ (.A0(\i_tinyqv.cpu.i_core.mepc[14] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .S(_03013_),
    .X(_03026_));
 sg13g2_mux2_1 _08429_ (.A0(\addr[14] ),
    .A1(_03026_),
    .S(net93),
    .X(_00284_));
 sg13g2_mux2_1 _08430_ (.A0(\i_tinyqv.cpu.i_core.mepc[15] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .S(_03013_),
    .X(_03027_));
 sg13g2_mux2_1 _08431_ (.A0(\addr[15] ),
    .A1(_03027_),
    .S(net93),
    .X(_00285_));
 sg13g2_mux2_1 _08432_ (.A0(\i_tinyqv.cpu.i_core.mepc[16] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .S(_03012_),
    .X(_03028_));
 sg13g2_mux2_1 _08433_ (.A0(\addr[16] ),
    .A1(_03028_),
    .S(_03010_),
    .X(_00286_));
 sg13g2_mux2_1 _08434_ (.A0(\i_tinyqv.cpu.i_core.mepc[17] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .S(_03012_),
    .X(_03029_));
 sg13g2_mux2_1 _08435_ (.A0(\addr[17] ),
    .A1(_03029_),
    .S(net93),
    .X(_00287_));
 sg13g2_mux2_1 _08436_ (.A0(\i_tinyqv.cpu.i_core.mepc[18] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S(_03012_),
    .X(_03030_));
 sg13g2_buf_1 _08437_ (.A(_03009_),
    .X(_03031_));
 sg13g2_mux2_1 _08438_ (.A0(\addr[18] ),
    .A1(_03030_),
    .S(net92),
    .X(_00288_));
 sg13g2_mux2_1 _08439_ (.A0(\i_tinyqv.cpu.i_core.mepc[19] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .S(net149),
    .X(_03032_));
 sg13g2_mux2_1 _08440_ (.A0(\addr[19] ),
    .A1(_03032_),
    .S(net92),
    .X(_00289_));
 sg13g2_nand2_1 _08441_ (.Y(_03033_),
    .A(\i_tinyqv.cpu.i_core.mepc[1] ),
    .B(_01276_));
 sg13g2_o21ai_1 _08442_ (.B1(_03033_),
    .Y(_03034_),
    .A1(_01809_),
    .A2(_01276_));
 sg13g2_mux2_1 _08443_ (.A0(\addr[1] ),
    .A1(_03034_),
    .S(_03031_),
    .X(_00290_));
 sg13g2_mux2_1 _08444_ (.A0(\i_tinyqv.cpu.i_core.mepc[20] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .S(net149),
    .X(_03035_));
 sg13g2_mux2_1 _08445_ (.A0(\addr[20] ),
    .A1(_03035_),
    .S(net92),
    .X(_00291_));
 sg13g2_mux2_1 _08446_ (.A0(\i_tinyqv.cpu.i_core.mepc[21] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .S(net149),
    .X(_03036_));
 sg13g2_mux2_1 _08447_ (.A0(\addr[21] ),
    .A1(_03036_),
    .S(_03031_),
    .X(_00292_));
 sg13g2_mux2_1 _08448_ (.A0(\i_tinyqv.cpu.i_core.mepc[22] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .S(net149),
    .X(_03037_));
 sg13g2_mux2_1 _08449_ (.A0(\addr[22] ),
    .A1(_03037_),
    .S(net92),
    .X(_00293_));
 sg13g2_mux2_1 _08450_ (.A0(\i_tinyqv.cpu.i_core.mepc[23] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .S(net149),
    .X(_03038_));
 sg13g2_mux2_1 _08451_ (.A0(\addr[23] ),
    .A1(_03038_),
    .S(net92),
    .X(_00294_));
 sg13g2_nand2_1 _08452_ (.Y(_03039_),
    .A(\i_tinyqv.cpu.i_core.mepc[2] ),
    .B(net147));
 sg13g2_o21ai_1 _08453_ (.B1(_03039_),
    .Y(_03040_),
    .A1(_01868_),
    .A2(net147));
 sg13g2_mux2_1 _08454_ (.A0(_01578_),
    .A1(_03040_),
    .S(net92),
    .X(_00299_));
 sg13g2_nand2_1 _08455_ (.Y(_03041_),
    .A(\i_tinyqv.cpu.i_core.mepc[3] ),
    .B(net147));
 sg13g2_o21ai_1 _08456_ (.B1(_03041_),
    .Y(_03042_),
    .A1(_01905_),
    .A2(net148));
 sg13g2_mux2_1 _08457_ (.A0(_01579_),
    .A1(_03042_),
    .S(net92),
    .X(_00300_));
 sg13g2_nand2_1 _08458_ (.Y(_03043_),
    .A(\i_tinyqv.cpu.i_core.mepc[4] ),
    .B(net147));
 sg13g2_o21ai_1 _08459_ (.B1(_03043_),
    .Y(_03044_),
    .A1(_01932_),
    .A2(net147));
 sg13g2_nand2_1 _08460_ (.Y(_03045_),
    .A(_03009_),
    .B(_03044_));
 sg13g2_o21ai_1 _08461_ (.B1(_03045_),
    .Y(_00301_),
    .A1(_02179_),
    .A2(_03010_));
 sg13g2_nand2_1 _08462_ (.Y(_03046_),
    .A(\i_tinyqv.cpu.i_core.mepc[5] ),
    .B(net147));
 sg13g2_o21ai_1 _08463_ (.B1(_03046_),
    .Y(_03047_),
    .A1(_01981_),
    .A2(_03014_));
 sg13g2_mux2_1 _08464_ (.A0(_01576_),
    .A1(_03047_),
    .S(net92),
    .X(_00302_));
 sg13g2_mux2_1 _08465_ (.A0(_01983_),
    .A1(\i_tinyqv.cpu.i_core.mepc[6] ),
    .S(net148),
    .X(_03048_));
 sg13g2_mux2_1 _08466_ (.A0(\addr[6] ),
    .A1(_03048_),
    .S(_03009_),
    .X(_00303_));
 sg13g2_mux2_1 _08467_ (.A0(_02024_),
    .A1(\i_tinyqv.cpu.i_core.mepc[7] ),
    .S(_03021_),
    .X(_03049_));
 sg13g2_mux2_1 _08468_ (.A0(\addr[7] ),
    .A1(_03049_),
    .S(_03009_),
    .X(_00304_));
 sg13g2_mux2_1 _08469_ (.A0(_02045_),
    .A1(\i_tinyqv.cpu.i_core.mepc[8] ),
    .S(net147),
    .X(_03050_));
 sg13g2_mux2_1 _08470_ (.A0(\addr[8] ),
    .A1(_03050_),
    .S(_03009_),
    .X(_00305_));
 sg13g2_mux2_1 _08471_ (.A0(net292),
    .A1(\i_tinyqv.cpu.i_core.mepc[9] ),
    .S(_03021_),
    .X(_03051_));
 sg13g2_mux2_1 _08472_ (.A0(\addr[9] ),
    .A1(_03051_),
    .S(_03009_),
    .X(_00306_));
 sg13g2_nor2_2 _08473_ (.A(_01039_),
    .B(_02254_),
    .Y(_03052_));
 sg13g2_nand4_1 _08474_ (.B(net202),
    .C(_01055_),
    .A(net264),
    .Y(_03053_),
    .D(_01198_));
 sg13g2_buf_2 _08475_ (.A(_03053_),
    .X(_03054_));
 sg13g2_mux2_1 _08476_ (.A0(_03052_),
    .A1(_01573_),
    .S(_03054_),
    .X(_00307_));
 sg13g2_nor2_2 _08477_ (.A(_00916_),
    .B(_02254_),
    .Y(_03055_));
 sg13g2_nand2_1 _08478_ (.Y(_03056_),
    .A(net264),
    .B(_01198_));
 sg13g2_nor2_2 _08479_ (.A(_00805_),
    .B(_03056_),
    .Y(_03057_));
 sg13g2_mux2_1 _08480_ (.A0(\data_to_write[10] ),
    .A1(_03055_),
    .S(_03057_),
    .X(_00308_));
 sg13g2_nand2b_1 _08481_ (.Y(_03058_),
    .B(_02703_),
    .A_N(_00954_));
 sg13g2_inv_1 _08482_ (.Y(_03059_),
    .A(_03058_));
 sg13g2_mux2_1 _08483_ (.A0(\data_to_write[11] ),
    .A1(_03059_),
    .S(_03057_),
    .X(_00309_));
 sg13g2_nand2b_1 _08484_ (.Y(_03060_),
    .B(net201),
    .A_N(net264));
 sg13g2_nand2_1 _08485_ (.Y(_03061_),
    .A(_01055_),
    .B(_03060_));
 sg13g2_nand2_1 _08486_ (.Y(_03062_),
    .A(_03052_),
    .B(_03061_));
 sg13g2_nand2_1 _08487_ (.Y(_03063_),
    .A(net163),
    .B(net264));
 sg13g2_nor2_1 _08488_ (.A(net188),
    .B(_03063_),
    .Y(_03064_));
 sg13g2_nor3_1 _08489_ (.A(net186),
    .B(net163),
    .C(_03060_),
    .Y(_03065_));
 sg13g2_buf_1 _08490_ (.A(_00216_),
    .X(_03066_));
 sg13g2_nor2_1 _08491_ (.A(net282),
    .B(_01649_),
    .Y(_03067_));
 sg13g2_o21ai_1 _08492_ (.B1(_03067_),
    .Y(_03068_),
    .A1(_03064_),
    .A2(_03065_));
 sg13g2_buf_1 _08493_ (.A(_03068_),
    .X(_03069_));
 sg13g2_or2_1 _08494_ (.X(_03070_),
    .B(_03056_),
    .A(_00961_));
 sg13g2_buf_1 _08495_ (.A(_03070_),
    .X(_03071_));
 sg13g2_nand2_1 _08496_ (.Y(_03072_),
    .A(\data_to_write[12] ),
    .B(_03071_));
 sg13g2_o21ai_1 _08497_ (.B1(_03072_),
    .Y(_00310_),
    .A1(_03062_),
    .A2(_03069_));
 sg13g2_nor2_2 _08498_ (.A(_01087_),
    .B(_02254_),
    .Y(_03073_));
 sg13g2_nand2_1 _08499_ (.Y(_03074_),
    .A(_03061_),
    .B(_03073_));
 sg13g2_nand2_1 _08500_ (.Y(_03075_),
    .A(\data_to_write[13] ),
    .B(_03071_));
 sg13g2_o21ai_1 _08501_ (.B1(_03075_),
    .Y(_00311_),
    .A1(_03069_),
    .A2(_03074_));
 sg13g2_nand2_1 _08502_ (.Y(_03076_),
    .A(_03055_),
    .B(_03061_));
 sg13g2_nand2_1 _08503_ (.Y(_03077_),
    .A(\data_to_write[14] ),
    .B(_03071_));
 sg13g2_o21ai_1 _08504_ (.B1(_03077_),
    .Y(_00312_),
    .A1(_03069_),
    .A2(_03076_));
 sg13g2_nand2_1 _08505_ (.Y(_03078_),
    .A(_03059_),
    .B(_03061_));
 sg13g2_nand2_1 _08506_ (.Y(_03079_),
    .A(\data_to_write[15] ),
    .B(_03071_));
 sg13g2_o21ai_1 _08507_ (.B1(_03079_),
    .Y(_00313_),
    .A1(_03069_),
    .A2(_03078_));
 sg13g2_inv_1 _08508_ (.Y(_03080_),
    .A(_03062_));
 sg13g2_nand2b_2 _08509_ (.Y(_03081_),
    .B(_01198_),
    .A_N(net264));
 sg13g2_nor2_2 _08510_ (.A(_02358_),
    .B(_03081_),
    .Y(_03082_));
 sg13g2_mux2_1 _08511_ (.A0(\data_to_write[16] ),
    .A1(_03080_),
    .S(_03082_),
    .X(_00314_));
 sg13g2_inv_1 _08512_ (.Y(_03083_),
    .A(_03074_));
 sg13g2_mux2_1 _08513_ (.A0(\data_to_write[17] ),
    .A1(_03083_),
    .S(_03082_),
    .X(_00315_));
 sg13g2_inv_1 _08514_ (.Y(_03084_),
    .A(_03076_));
 sg13g2_mux2_1 _08515_ (.A0(\data_to_write[18] ),
    .A1(_03084_),
    .S(_03082_),
    .X(_00316_));
 sg13g2_inv_1 _08516_ (.Y(_03085_),
    .A(_03078_));
 sg13g2_mux2_1 _08517_ (.A0(\data_to_write[19] ),
    .A1(_03085_),
    .S(_03082_),
    .X(_00317_));
 sg13g2_mux2_1 _08518_ (.A0(_03073_),
    .A1(_01600_),
    .S(_03054_),
    .X(_00318_));
 sg13g2_nor2_1 _08519_ (.A(_01163_),
    .B(_01649_),
    .Y(_03086_));
 sg13g2_nand2b_1 _08520_ (.Y(_03087_),
    .B(_03052_),
    .A_N(net282));
 sg13g2_nand3_1 _08521_ (.B(_03086_),
    .C(_03087_),
    .A(net163),
    .Y(_03088_));
 sg13g2_o21ai_1 _08522_ (.B1(_03088_),
    .Y(_03089_),
    .A1(net163),
    .A2(\data_to_write[20] ));
 sg13g2_inv_1 _08523_ (.Y(_03090_),
    .A(_00961_));
 sg13g2_nor3_2 _08524_ (.A(net282),
    .B(_03090_),
    .C(_03081_),
    .Y(_03091_));
 sg13g2_a21oi_1 _08525_ (.A1(_03052_),
    .A2(_03091_),
    .Y(_03092_),
    .B1(\data_to_write[20] ));
 sg13g2_a21oi_1 _08526_ (.A1(net188),
    .A2(_03089_),
    .Y(_00319_),
    .B1(_03092_));
 sg13g2_nand2b_1 _08527_ (.Y(_03093_),
    .B(_03073_),
    .A_N(net282));
 sg13g2_nand3_1 _08528_ (.B(_03086_),
    .C(_03093_),
    .A(_02603_),
    .Y(_03094_));
 sg13g2_o21ai_1 _08529_ (.B1(_03094_),
    .Y(_03095_),
    .A1(net163),
    .A2(\data_to_write[21] ));
 sg13g2_a21oi_1 _08530_ (.A1(_03073_),
    .A2(_03091_),
    .Y(_03096_),
    .B1(\data_to_write[21] ));
 sg13g2_a21oi_1 _08531_ (.A1(net188),
    .A2(_03095_),
    .Y(_00320_),
    .B1(_03096_));
 sg13g2_nand2b_1 _08532_ (.Y(_03097_),
    .B(_03055_),
    .A_N(net282));
 sg13g2_nand3_1 _08533_ (.B(_03086_),
    .C(_03097_),
    .A(net163),
    .Y(_03098_));
 sg13g2_o21ai_1 _08534_ (.B1(_03098_),
    .Y(_03099_),
    .A1(net163),
    .A2(\data_to_write[22] ));
 sg13g2_a21oi_1 _08535_ (.A1(_03055_),
    .A2(_03091_),
    .Y(_03100_),
    .B1(\data_to_write[22] ));
 sg13g2_a21oi_1 _08536_ (.A1(net188),
    .A2(_03099_),
    .Y(_00321_),
    .B1(_03100_));
 sg13g2_o21ai_1 _08537_ (.B1(_03086_),
    .Y(_03101_),
    .A1(net282),
    .A2(_03058_));
 sg13g2_or2_1 _08538_ (.X(_03102_),
    .B(\data_to_write[23] ),
    .A(net163));
 sg13g2_o21ai_1 _08539_ (.B1(_03102_),
    .Y(_03103_),
    .A1(net207),
    .A2(_03101_));
 sg13g2_a21oi_1 _08540_ (.A1(_03059_),
    .A2(_03091_),
    .Y(_03104_),
    .B1(\data_to_write[23] ));
 sg13g2_a21oi_1 _08541_ (.A1(_02178_),
    .A2(_03103_),
    .Y(_00322_),
    .B1(_03104_));
 sg13g2_nor2_2 _08542_ (.A(_00805_),
    .B(_03081_),
    .Y(_03105_));
 sg13g2_mux2_1 _08543_ (.A0(\data_to_write[24] ),
    .A1(_03052_),
    .S(_03105_),
    .X(_00323_));
 sg13g2_mux2_1 _08544_ (.A0(\data_to_write[25] ),
    .A1(_03073_),
    .S(_03105_),
    .X(_00324_));
 sg13g2_mux2_1 _08545_ (.A0(\data_to_write[26] ),
    .A1(_03055_),
    .S(_03105_),
    .X(_00325_));
 sg13g2_mux2_1 _08546_ (.A0(\data_to_write[27] ),
    .A1(_03059_),
    .S(_03105_),
    .X(_00326_));
 sg13g2_and3_1 _08547_ (.X(_03106_),
    .A(_01163_),
    .B(net201),
    .C(_01055_));
 sg13g2_o21ai_1 _08548_ (.B1(_03067_),
    .Y(_03107_),
    .A1(net160),
    .A2(_03106_));
 sg13g2_buf_1 _08549_ (.A(_03107_),
    .X(_03108_));
 sg13g2_nand2_1 _08550_ (.Y(_03109_),
    .A(_01166_),
    .B(_01198_));
 sg13g2_nand2_1 _08551_ (.Y(_03110_),
    .A(\data_to_write[28] ),
    .B(_03109_));
 sg13g2_o21ai_1 _08552_ (.B1(_03110_),
    .Y(_00327_),
    .A1(_03062_),
    .A2(_03108_));
 sg13g2_nand2_1 _08553_ (.Y(_03111_),
    .A(\data_to_write[29] ),
    .B(_03109_));
 sg13g2_o21ai_1 _08554_ (.B1(_03111_),
    .Y(_00328_),
    .A1(_03074_),
    .A2(_03108_));
 sg13g2_mux2_1 _08555_ (.A0(_03055_),
    .A1(_01603_),
    .S(_03054_),
    .X(_00329_));
 sg13g2_nand2_1 _08556_ (.Y(_03112_),
    .A(\data_to_write[30] ),
    .B(_03109_));
 sg13g2_o21ai_1 _08557_ (.B1(_03112_),
    .Y(_00330_),
    .A1(_03076_),
    .A2(_03108_));
 sg13g2_nand2_1 _08558_ (.Y(_03113_),
    .A(\data_to_write[31] ),
    .B(_03109_));
 sg13g2_o21ai_1 _08559_ (.B1(_03113_),
    .Y(_00331_),
    .A1(_03078_),
    .A2(_03108_));
 sg13g2_nand2_1 _08560_ (.Y(_03114_),
    .A(_01606_),
    .B(_03054_));
 sg13g2_o21ai_1 _08561_ (.B1(_03114_),
    .Y(_00332_),
    .A1(_03054_),
    .A2(_03058_));
 sg13g2_nor2_1 _08562_ (.A(_00893_),
    .B(_01145_),
    .Y(_03115_));
 sg13g2_or3_1 _08563_ (.A(_03066_),
    .B(_03056_),
    .C(_03115_),
    .X(_03116_));
 sg13g2_buf_1 _08564_ (.A(_03116_),
    .X(_03117_));
 sg13g2_nand2_1 _08565_ (.Y(_03118_),
    .A(_01198_),
    .B(_02364_));
 sg13g2_nand2_1 _08566_ (.Y(_03119_),
    .A(_01609_),
    .B(_03118_));
 sg13g2_o21ai_1 _08567_ (.B1(_03119_),
    .Y(_00333_),
    .A1(_03062_),
    .A2(_03117_));
 sg13g2_nand2_1 _08568_ (.Y(_03120_),
    .A(_01612_),
    .B(_03118_));
 sg13g2_o21ai_1 _08569_ (.B1(_03120_),
    .Y(_00334_),
    .A1(_03074_),
    .A2(_03117_));
 sg13g2_nand2_1 _08570_ (.Y(_03121_),
    .A(_01616_),
    .B(_03118_));
 sg13g2_o21ai_1 _08571_ (.B1(_03121_),
    .Y(_00335_),
    .A1(_03076_),
    .A2(_03117_));
 sg13g2_nand2_1 _08572_ (.Y(_03122_),
    .A(\data_to_write[7] ),
    .B(_03118_));
 sg13g2_o21ai_1 _08573_ (.B1(_03122_),
    .Y(_00336_),
    .A1(_03078_),
    .A2(_03117_));
 sg13g2_mux2_1 _08574_ (.A0(\data_to_write[8] ),
    .A1(_03052_),
    .S(_03057_),
    .X(_00337_));
 sg13g2_mux2_1 _08575_ (.A0(\data_to_write[9] ),
    .A1(_03073_),
    .S(_03057_),
    .X(_00338_));
 sg13g2_or2_1 _08576_ (.X(_03123_),
    .B(_01194_),
    .A(net173));
 sg13g2_buf_1 _08577_ (.A(_03123_),
    .X(_03124_));
 sg13g2_nand2_1 _08578_ (.Y(_03125_),
    .A(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .B(net173));
 sg13g2_o21ai_1 _08579_ (.B1(_03125_),
    .Y(_00357_),
    .A1(_02728_),
    .A2(_03124_));
 sg13g2_inv_1 _08580_ (.Y(_03126_),
    .A(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ));
 sg13g2_nor2_1 _08581_ (.A(_01642_),
    .B(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .Y(_03127_));
 sg13g2_o21ai_1 _08582_ (.B1(_03127_),
    .Y(_03128_),
    .A1(_02728_),
    .A2(_03124_));
 sg13g2_buf_1 _08583_ (.A(_03128_),
    .X(_03129_));
 sg13g2_nor4_2 _08584_ (.A(_02232_),
    .B(_02193_),
    .C(_02247_),
    .Y(_03130_),
    .D(net105));
 sg13g2_nand2_1 _08585_ (.Y(_03131_),
    .A(\i_tinyqv.cpu.i_core.interrupt_req[0] ),
    .B(_03130_));
 sg13g2_o21ai_1 _08586_ (.B1(_03131_),
    .Y(_00358_),
    .A1(_03126_),
    .A2(_03130_));
 sg13g2_inv_1 _08587_ (.Y(_03132_),
    .A(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ));
 sg13g2_nand2_1 _08588_ (.Y(_03133_),
    .A(\i_tinyqv.cpu.i_core.interrupt_req[1] ),
    .B(_03130_));
 sg13g2_o21ai_1 _08589_ (.B1(_03133_),
    .Y(_00359_),
    .A1(_03132_),
    .A2(_03130_));
 sg13g2_inv_1 _08590_ (.Y(_03134_),
    .A(\i_tinyqv.cpu.i_core.load_done ));
 sg13g2_nand3_1 _08591_ (.B(\i_tinyqv.cpu.data_ready_core ),
    .C(net157),
    .A(_01647_),
    .Y(_03135_));
 sg13g2_o21ai_1 _08592_ (.B1(_03135_),
    .Y(_00360_),
    .A1(_03134_),
    .A2(net157));
 sg13g2_and2_1 _08593_ (.A(\i_tinyqv.cpu.i_core.load_top_bit ),
    .B(_01060_),
    .X(_03136_));
 sg13g2_nor4_1 _08594_ (.A(_02250_),
    .B(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .C(_01535_),
    .D(_02251_),
    .Y(_03137_));
 sg13g2_a21oi_1 _08595_ (.A1(net188),
    .A2(_01263_),
    .Y(_03138_),
    .B1(_03063_));
 sg13g2_nand2_1 _08596_ (.Y(_03139_),
    .A(_03137_),
    .B(_03138_));
 sg13g2_mux2_1 _08597_ (.A0(_02813_),
    .A1(_03136_),
    .S(_03139_),
    .X(_00361_));
 sg13g2_nand2_1 _08598_ (.Y(_03140_),
    .A(net218),
    .B(\i_tinyqv.cpu.is_alu_imm ));
 sg13g2_buf_2 _08599_ (.A(_03140_),
    .X(_03141_));
 sg13g2_and3_1 _08600_ (.X(_03142_),
    .A(net218),
    .B(\i_tinyqv.cpu.is_alu_imm ),
    .C(_01049_));
 sg13g2_a21oi_1 _08601_ (.A1(_01039_),
    .A2(_03141_),
    .Y(_03143_),
    .B1(_03142_));
 sg13g2_nand2_1 _08602_ (.Y(_03144_),
    .A(net157),
    .B(_01648_));
 sg13g2_buf_2 _08603_ (.A(_03144_),
    .X(_03145_));
 sg13g2_mux2_1 _08604_ (.A0(_03143_),
    .A1(net249),
    .S(_03145_),
    .X(_00397_));
 sg13g2_nand2_1 _08605_ (.Y(_03146_),
    .A(_01087_),
    .B(_03141_));
 sg13g2_o21ai_1 _08606_ (.B1(_03146_),
    .Y(_03147_),
    .A1(_01096_),
    .A2(_03141_));
 sg13g2_nand2_1 _08607_ (.Y(_03148_),
    .A(_02437_),
    .B(_03145_));
 sg13g2_o21ai_1 _08608_ (.B1(_03148_),
    .Y(_00398_),
    .A1(_03145_),
    .A2(_03147_));
 sg13g2_nand2_1 _08609_ (.Y(_03149_),
    .A(_00916_),
    .B(_03141_));
 sg13g2_o21ai_1 _08610_ (.B1(_03149_),
    .Y(_03150_),
    .A1(_00924_),
    .A2(_03141_));
 sg13g2_nand2_1 _08611_ (.Y(_03151_),
    .A(_02416_),
    .B(_03145_));
 sg13g2_o21ai_1 _08612_ (.B1(_03151_),
    .Y(_00399_),
    .A1(_03145_),
    .A2(_03150_));
 sg13g2_nor2_1 _08613_ (.A(_00975_),
    .B(_03141_),
    .Y(_03152_));
 sg13g2_a21oi_1 _08614_ (.A1(_00954_),
    .A2(_03141_),
    .Y(_03153_),
    .B1(_03152_));
 sg13g2_mux2_1 _08615_ (.A0(_03153_),
    .A1(_02438_),
    .S(_03145_),
    .X(_00400_));
 sg13g2_nor4_1 _08616_ (.A(_01646_),
    .B(_01647_),
    .C(net282),
    .D(_02363_),
    .Y(_03154_));
 sg13g2_mux2_1 _08617_ (.A0(_02466_),
    .A1(_03143_),
    .S(_03154_),
    .X(_00401_));
 sg13g2_nand3_1 _08618_ (.B(net129),
    .C(_02925_),
    .A(_01328_),
    .Y(_03155_));
 sg13g2_nand2_1 _08619_ (.Y(_03156_),
    .A(_02920_),
    .B(_03155_));
 sg13g2_buf_2 _08620_ (.A(_03156_),
    .X(_03157_));
 sg13g2_inv_1 _08621_ (.Y(_03158_),
    .A(_01491_));
 sg13g2_nor3_2 _08622_ (.A(_01453_),
    .B(net136),
    .C(_01351_),
    .Y(_03159_));
 sg13g2_nor2_1 _08623_ (.A(_01453_),
    .B(net136),
    .Y(_03160_));
 sg13g2_buf_2 _08624_ (.A(_03160_),
    .X(_03161_));
 sg13g2_mux2_1 _08625_ (.A0(_00107_),
    .A1(_00108_),
    .S(net152),
    .X(_03162_));
 sg13g2_mux2_1 _08626_ (.A0(_01335_),
    .A1(_03162_),
    .S(_01334_),
    .X(_03163_));
 sg13g2_buf_1 _08627_ (.A(_03163_),
    .X(_03164_));
 sg13g2_nor3_1 _08628_ (.A(_01355_),
    .B(_03161_),
    .C(_03164_),
    .Y(_03165_));
 sg13g2_a21oi_1 _08629_ (.A1(_03158_),
    .A2(_03159_),
    .Y(_03166_),
    .B1(_03165_));
 sg13g2_nor2_1 _08630_ (.A(_03157_),
    .B(_03166_),
    .Y(_03167_));
 sg13g2_nor2_2 _08631_ (.A(net124),
    .B(_02918_),
    .Y(_03168_));
 sg13g2_nor2_2 _08632_ (.A(_01464_),
    .B(_01322_),
    .Y(_03169_));
 sg13g2_nor2_1 _08633_ (.A(_01362_),
    .B(net94),
    .Y(_03170_));
 sg13g2_a22oi_1 _08634_ (.Y(_03171_),
    .B1(_03170_),
    .B2(net124),
    .A2(_03169_),
    .A1(_03168_));
 sg13g2_or2_1 _08635_ (.X(_03172_),
    .B(_03171_),
    .A(net117));
 sg13g2_buf_1 _08636_ (.A(_03172_),
    .X(_03173_));
 sg13g2_nand2b_1 _08637_ (.Y(_03174_),
    .B(net130),
    .A_N(_03173_));
 sg13g2_nand3_1 _08638_ (.B(_02950_),
    .C(_02987_),
    .A(_01489_),
    .Y(_03175_));
 sg13g2_buf_1 _08639_ (.A(_03175_),
    .X(_03176_));
 sg13g2_and4_1 _08640_ (.A(_01480_),
    .B(net122),
    .C(_01491_),
    .D(_02949_),
    .X(_03177_));
 sg13g2_buf_1 _08641_ (.A(_03177_),
    .X(_03178_));
 sg13g2_nand2_2 _08642_ (.Y(_03179_),
    .A(_01457_),
    .B(_02918_));
 sg13g2_nor3_1 _08643_ (.A(_02935_),
    .B(_01467_),
    .C(_03179_),
    .Y(_03180_));
 sg13g2_a22oi_1 _08644_ (.Y(_03181_),
    .B1(_03180_),
    .B2(_01473_),
    .A2(_03178_),
    .A1(_01468_));
 sg13g2_nand3_1 _08645_ (.B(_03176_),
    .C(_03181_),
    .A(_03174_),
    .Y(_03182_));
 sg13g2_buf_1 _08646_ (.A(_02913_),
    .X(_03183_));
 sg13g2_o21ai_1 _08647_ (.B1(net41),
    .Y(_03184_),
    .A1(_03167_),
    .A2(_03182_));
 sg13g2_o21ai_1 _08648_ (.B1(_03184_),
    .Y(_00437_),
    .A1(_02325_),
    .A2(_02915_));
 sg13g2_nand2_1 _08649_ (.Y(_03185_),
    .A(net107),
    .B(_01322_));
 sg13g2_buf_2 _08650_ (.A(_03185_),
    .X(_03186_));
 sg13g2_nand3_1 _08651_ (.B(_02950_),
    .C(_02951_),
    .A(_01464_),
    .Y(_03187_));
 sg13g2_o21ai_1 _08652_ (.B1(net106),
    .Y(_03188_),
    .A1(_01332_),
    .A2(_03187_));
 sg13g2_nand2_1 _08653_ (.Y(_03189_),
    .A(_03186_),
    .B(_03188_));
 sg13g2_a22oi_1 _08654_ (.Y(_03190_),
    .B1(_03189_),
    .B2(net96),
    .A2(_02960_),
    .A1(_01466_));
 sg13g2_buf_1 _08655_ (.A(_02980_),
    .X(_03191_));
 sg13g2_nand2_2 _08656_ (.Y(_03192_),
    .A(_02931_),
    .B(_01322_));
 sg13g2_nor3_2 _08657_ (.A(net104),
    .B(_03179_),
    .C(_03192_),
    .Y(_03193_));
 sg13g2_nand2_1 _08658_ (.Y(_03194_),
    .A(_02980_),
    .B(net99));
 sg13g2_nor2_2 _08659_ (.A(_01316_),
    .B(net128),
    .Y(_03195_));
 sg13g2_nand3_1 _08660_ (.B(net96),
    .C(_03195_),
    .A(_02980_),
    .Y(_03196_));
 sg13g2_buf_1 _08661_ (.A(_03196_),
    .X(_03197_));
 sg13g2_nor4_2 _08662_ (.A(_01474_),
    .B(_01479_),
    .C(net122),
    .Y(_03198_),
    .D(_03158_));
 sg13g2_nand2b_1 _08663_ (.Y(_03199_),
    .B(_03198_),
    .A_N(_03197_));
 sg13g2_o21ai_1 _08664_ (.B1(_03199_),
    .Y(_03200_),
    .A1(_01458_),
    .A2(_03194_));
 sg13g2_buf_1 _08665_ (.A(_03200_),
    .X(_03201_));
 sg13g2_nor2_1 _08666_ (.A(_03193_),
    .B(_03201_),
    .Y(_03202_));
 sg13g2_a21oi_1 _08667_ (.A1(_03190_),
    .A2(_03202_),
    .Y(_03203_),
    .B1(net97));
 sg13g2_buf_1 _08668_ (.A(_01362_),
    .X(_03204_));
 sg13g2_buf_1 _08669_ (.A(net114),
    .X(_03205_));
 sg13g2_nand2_1 _08670_ (.Y(_03206_),
    .A(_02931_),
    .B(net128));
 sg13g2_nor3_1 _08671_ (.A(net103),
    .B(net122),
    .C(_03206_),
    .Y(_03207_));
 sg13g2_buf_1 _08672_ (.A(_02918_),
    .X(_03208_));
 sg13g2_buf_1 _08673_ (.A(net113),
    .X(_03209_));
 sg13g2_nor2_2 _08674_ (.A(_01351_),
    .B(_02951_),
    .Y(_03210_));
 sg13g2_nor3_1 _08675_ (.A(net102),
    .B(_03001_),
    .C(_03210_),
    .Y(_03211_));
 sg13g2_buf_1 _08676_ (.A(net124),
    .X(_03212_));
 sg13g2_buf_1 _08677_ (.A(net101),
    .X(_03213_));
 sg13g2_buf_1 _08678_ (.A(net91),
    .X(_03214_));
 sg13g2_o21ai_1 _08679_ (.B1(_03214_),
    .Y(_03215_),
    .A1(_03207_),
    .A2(_03211_));
 sg13g2_nor2b_1 _08680_ (.A(_03203_),
    .B_N(_03215_),
    .Y(_03216_));
 sg13g2_nor2_1 _08681_ (.A(net285),
    .B(net42),
    .Y(_03217_));
 sg13g2_a21oi_1 _08682_ (.A1(net38),
    .A2(_03216_),
    .Y(_00438_),
    .B1(_03217_));
 sg13g2_mux2_1 _08683_ (.A0(_00127_),
    .A1(_00128_),
    .S(net152),
    .X(_03218_));
 sg13g2_mux2_1 _08684_ (.A0(_01459_),
    .A1(_03218_),
    .S(net183),
    .X(_03219_));
 sg13g2_inv_1 _08685_ (.Y(_03220_),
    .A(_03219_));
 sg13g2_nand2_1 _08686_ (.Y(_03221_),
    .A(net129),
    .B(_03220_));
 sg13g2_o21ai_1 _08687_ (.B1(_03221_),
    .Y(_03222_),
    .A1(net129),
    .A2(_01491_));
 sg13g2_nand2_1 _08688_ (.Y(_03223_),
    .A(_01355_),
    .B(_03164_));
 sg13g2_o21ai_1 _08689_ (.B1(_03223_),
    .Y(_03224_),
    .A1(_01355_),
    .A2(_03220_));
 sg13g2_nor2_1 _08690_ (.A(_03161_),
    .B(_03224_),
    .Y(_03225_));
 sg13g2_a21oi_1 _08691_ (.A1(_03161_),
    .A2(_03222_),
    .Y(_03226_),
    .B1(_03225_));
 sg13g2_a21oi_1 _08692_ (.A1(_01310_),
    .A2(net128),
    .Y(_03227_),
    .B1(net94));
 sg13g2_nor2_1 _08693_ (.A(_01457_),
    .B(net117),
    .Y(_03228_));
 sg13g2_o21ai_1 _08694_ (.B1(_03228_),
    .Y(_03229_),
    .A1(_01322_),
    .A2(_03187_));
 sg13g2_o21ai_1 _08695_ (.B1(_03229_),
    .Y(_03230_),
    .A1(_01316_),
    .A2(_03227_));
 sg13g2_a22oi_1 _08696_ (.Y(_03231_),
    .B1(_03230_),
    .B2(_02918_),
    .A2(_03169_),
    .A1(_03168_));
 sg13g2_nand2_1 _08697_ (.Y(_03232_),
    .A(_03199_),
    .B(_03231_));
 sg13g2_nor2_1 _08698_ (.A(_02923_),
    .B(_02974_),
    .Y(_03233_));
 sg13g2_o21ai_1 _08699_ (.B1(_01489_),
    .Y(_03234_),
    .A1(_03232_),
    .A2(_03233_));
 sg13g2_buf_1 _08700_ (.A(_03234_),
    .X(_03235_));
 sg13g2_o21ai_1 _08701_ (.B1(_03235_),
    .Y(_03236_),
    .A1(_03157_),
    .A2(_03226_));
 sg13g2_buf_1 _08702_ (.A(_02914_),
    .X(_03237_));
 sg13g2_mux2_1 _08703_ (.A0(net310),
    .A1(_03236_),
    .S(net37),
    .X(_00439_));
 sg13g2_nor2_2 _08704_ (.A(_03197_),
    .B(_03198_),
    .Y(_03238_));
 sg13g2_nand2_1 _08705_ (.Y(_03239_),
    .A(net130),
    .B(_03238_));
 sg13g2_nor2_1 _08706_ (.A(_01355_),
    .B(_03210_),
    .Y(_03240_));
 sg13g2_buf_1 _08707_ (.A(_03240_),
    .X(_03241_));
 sg13g2_buf_1 _08708_ (.A(_01395_),
    .X(_03242_));
 sg13g2_a21oi_1 _08709_ (.A1(_03219_),
    .A2(net87),
    .Y(_03243_),
    .B1(_03242_));
 sg13g2_buf_2 _08710_ (.A(_03243_),
    .X(_03244_));
 sg13g2_o21ai_1 _08711_ (.B1(_03244_),
    .Y(_03245_),
    .A1(_01489_),
    .A2(_03241_));
 sg13g2_nand4_1 _08712_ (.B(_03235_),
    .C(_03239_),
    .A(net43),
    .Y(_03246_),
    .D(_03245_));
 sg13g2_o21ai_1 _08713_ (.B1(_03246_),
    .Y(_03247_),
    .A1(_01043_),
    .A2(net41));
 sg13g2_inv_1 _08714_ (.Y(_00440_),
    .A(_03247_));
 sg13g2_nand2_1 _08715_ (.Y(_03248_),
    .A(_01332_),
    .B(_03238_));
 sg13g2_o21ai_1 _08716_ (.B1(_03244_),
    .Y(_03249_),
    .A1(net108),
    .A2(net87));
 sg13g2_nand4_1 _08717_ (.B(_03235_),
    .C(_03248_),
    .A(net43),
    .Y(_03250_),
    .D(_03249_));
 sg13g2_o21ai_1 _08718_ (.B1(_03250_),
    .Y(_03251_),
    .A1(_01088_),
    .A2(net41));
 sg13g2_inv_1 _08719_ (.Y(_00441_),
    .A(_03251_));
 sg13g2_nand2_1 _08720_ (.Y(_03252_),
    .A(net123),
    .B(_03238_));
 sg13g2_o21ai_1 _08721_ (.B1(_03244_),
    .Y(_03253_),
    .A1(net115),
    .A2(net87));
 sg13g2_nand4_1 _08722_ (.B(_03235_),
    .C(_03252_),
    .A(net43),
    .Y(_03254_),
    .D(_03253_));
 sg13g2_o21ai_1 _08723_ (.B1(_03254_),
    .Y(_03255_),
    .A1(_00917_),
    .A2(net41));
 sg13g2_inv_1 _08724_ (.Y(_00442_),
    .A(_03255_));
 sg13g2_nand2_1 _08725_ (.Y(_03256_),
    .A(_01345_),
    .B(_03238_));
 sg13g2_o21ai_1 _08726_ (.B1(_03244_),
    .Y(_03257_),
    .A1(net95),
    .A2(net87));
 sg13g2_nand4_1 _08727_ (.B(_03235_),
    .C(_03256_),
    .A(net43),
    .Y(_03258_),
    .D(_03257_));
 sg13g2_o21ai_1 _08728_ (.B1(_03258_),
    .Y(_03259_),
    .A1(_00959_),
    .A2(net41));
 sg13g2_inv_1 _08729_ (.Y(_00443_),
    .A(_03259_));
 sg13g2_inv_1 _08730_ (.Y(_03260_),
    .A(_03238_));
 sg13g2_mux2_1 _08731_ (.A0(\i_tinyqv.cpu.instr_data[0][0] ),
    .A1(\i_tinyqv.cpu.instr_data[2][0] ),
    .S(net152),
    .X(_03261_));
 sg13g2_mux2_1 _08732_ (.A0(_01305_),
    .A1(_03261_),
    .S(net183),
    .X(_03262_));
 sg13g2_o21ai_1 _08733_ (.B1(_03244_),
    .Y(_03263_),
    .A1(net87),
    .A2(_03262_));
 sg13g2_o21ai_1 _08734_ (.B1(_03263_),
    .Y(_03264_),
    .A1(net129),
    .A2(_03260_));
 sg13g2_a21oi_1 _08735_ (.A1(_01489_),
    .A2(_03232_),
    .Y(_03265_),
    .B1(_03264_));
 sg13g2_buf_1 _08736_ (.A(net43),
    .X(_03266_));
 sg13g2_nor2_1 _08737_ (.A(_01045_),
    .B(net36),
    .Y(_03267_));
 sg13g2_a21oi_1 _08738_ (.A1(net38),
    .A2(_03265_),
    .Y(_00444_),
    .B1(_03267_));
 sg13g2_a21oi_2 _08739_ (.B1(_02944_),
    .Y(_03268_),
    .A2(_03231_),
    .A1(_03197_));
 sg13g2_mux4_1 _08740_ (.S0(net127),
    .A0(\i_tinyqv.cpu.instr_data[0][1] ),
    .A1(\i_tinyqv.cpu.instr_data[2][1] ),
    .A2(\i_tinyqv.cpu.instr_data[3][1] ),
    .A3(\i_tinyqv.cpu.instr_data[1][1] ),
    .S1(_01397_),
    .X(_03269_));
 sg13g2_o21ai_1 _08741_ (.B1(_03244_),
    .Y(_03270_),
    .A1(net87),
    .A2(_03269_));
 sg13g2_nor2b_1 _08742_ (.A(_03268_),
    .B_N(_03270_),
    .Y(_03271_));
 sg13g2_nor2_1 _08743_ (.A(_01092_),
    .B(net36),
    .Y(_03272_));
 sg13g2_a21oi_1 _08744_ (.A1(net38),
    .A2(_03271_),
    .Y(_00445_),
    .B1(_03272_));
 sg13g2_mux2_1 _08745_ (.A0(\i_tinyqv.cpu.instr_data[0][2] ),
    .A1(\i_tinyqv.cpu.instr_data[2][2] ),
    .S(net152),
    .X(_03273_));
 sg13g2_mux2_1 _08746_ (.A0(_01325_),
    .A1(_03273_),
    .S(net183),
    .X(_03274_));
 sg13g2_o21ai_1 _08747_ (.B1(_03244_),
    .Y(_03275_),
    .A1(net87),
    .A2(_03274_));
 sg13g2_nor2b_1 _08748_ (.A(_03268_),
    .B_N(_03275_),
    .Y(_03276_));
 sg13g2_nor2_1 _08749_ (.A(_00921_),
    .B(net36),
    .Y(_03277_));
 sg13g2_a21oi_1 _08750_ (.A1(net38),
    .A2(_03276_),
    .Y(_00446_),
    .B1(_03277_));
 sg13g2_mux2_1 _08751_ (.A0(\i_tinyqv.cpu.instr_data[0][3] ),
    .A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .S(net127),
    .X(_03278_));
 sg13g2_mux2_1 _08752_ (.A0(_01329_),
    .A1(_03278_),
    .S(net183),
    .X(_03279_));
 sg13g2_o21ai_1 _08753_ (.B1(_03244_),
    .Y(_03280_),
    .A1(net87),
    .A2(_03279_));
 sg13g2_nor2b_1 _08754_ (.A(_03268_),
    .B_N(_03280_),
    .Y(_03281_));
 sg13g2_nor2_1 _08755_ (.A(_00965_),
    .B(net36),
    .Y(_03282_));
 sg13g2_a21oi_1 _08756_ (.A1(net38),
    .A2(_03281_),
    .Y(_00447_),
    .B1(_03282_));
 sg13g2_nor2_1 _08757_ (.A(net106),
    .B(net107),
    .Y(_03283_));
 sg13g2_inv_1 _08758_ (.Y(_03284_),
    .A(_03283_));
 sg13g2_o21ai_1 _08759_ (.B1(net96),
    .Y(_03285_),
    .A1(net99),
    .A2(_02982_));
 sg13g2_a22oi_1 _08760_ (.Y(_03286_),
    .B1(_03285_),
    .B2(_03173_),
    .A2(_03176_),
    .A1(_02923_));
 sg13g2_nor3_1 _08761_ (.A(net136),
    .B(_01467_),
    .C(_03179_),
    .Y(_03287_));
 sg13g2_nor2_1 _08762_ (.A(_03286_),
    .B(_03287_),
    .Y(_03288_));
 sg13g2_o21ai_1 _08763_ (.B1(_03288_),
    .Y(_03289_),
    .A1(net89),
    .A2(_03284_));
 sg13g2_mux2_1 _08764_ (.A0(_00111_),
    .A1(_00112_),
    .S(net127),
    .X(_03290_));
 sg13g2_mux2_1 _08765_ (.A0(_01340_),
    .A1(_03290_),
    .S(net183),
    .X(_03291_));
 sg13g2_nor2b_1 _08766_ (.A(_03161_),
    .B_N(_03291_),
    .Y(_03292_));
 sg13g2_a21oi_1 _08767_ (.A1(_01483_),
    .A2(_03161_),
    .Y(_03293_),
    .B1(_03292_));
 sg13g2_nor2_2 _08768_ (.A(_01395_),
    .B(_03210_),
    .Y(_03294_));
 sg13g2_a21oi_1 _08769_ (.A1(_02970_),
    .A2(_03288_),
    .Y(_03295_),
    .B1(_03214_));
 sg13g2_a221oi_1 _08770_ (.B2(_03294_),
    .C1(_03295_),
    .B1(_03293_),
    .A1(net102),
    .Y(_03296_),
    .A2(_03289_));
 sg13g2_nor2_1 _08771_ (.A(_01090_),
    .B(net36),
    .Y(_03297_));
 sg13g2_a21oi_1 _08772_ (.A1(_02964_),
    .A2(_03296_),
    .Y(_00448_),
    .B1(_03297_));
 sg13g2_nand2_1 _08773_ (.Y(_03298_),
    .A(_02920_),
    .B(_03210_));
 sg13g2_buf_1 _08774_ (.A(_03298_),
    .X(_03299_));
 sg13g2_a21oi_1 _08775_ (.A1(_03294_),
    .A2(_03220_),
    .Y(_03300_),
    .B1(_03268_));
 sg13g2_buf_1 _08776_ (.A(_03300_),
    .X(_03301_));
 sg13g2_o21ai_1 _08777_ (.B1(net84),
    .Y(_03302_),
    .A1(_03164_),
    .A2(net86));
 sg13g2_mux2_1 _08778_ (.A0(_01046_),
    .A1(_03302_),
    .S(net37),
    .X(_00449_));
 sg13g2_o21ai_1 _08779_ (.B1(net84),
    .Y(_03303_),
    .A1(_03291_),
    .A2(net86));
 sg13g2_mux2_1 _08780_ (.A0(_01093_),
    .A1(_03303_),
    .S(net37),
    .X(_00450_));
 sg13g2_inv_2 _08781_ (.Y(_03304_),
    .A(\i_tinyqv.cpu.imm[22] ));
 sg13g2_mux2_1 _08782_ (.A0(_00115_),
    .A1(_00116_),
    .S(net127),
    .X(_03305_));
 sg13g2_mux2_1 _08783_ (.A0(_01346_),
    .A1(_03305_),
    .S(net183),
    .X(_03306_));
 sg13g2_o21ai_1 _08784_ (.B1(net84),
    .Y(_03307_),
    .A1(net86),
    .A2(_03306_));
 sg13g2_nand2_1 _08785_ (.Y(_03308_),
    .A(_02977_),
    .B(_03307_));
 sg13g2_o21ai_1 _08786_ (.B1(_03308_),
    .Y(_00451_),
    .A1(_03304_),
    .A2(net40));
 sg13g2_mux4_1 _08787_ (.S0(net159),
    .A0(_00131_),
    .A1(_00133_),
    .A2(_00132_),
    .A3(_00130_),
    .S1(net127),
    .X(_03309_));
 sg13g2_o21ai_1 _08788_ (.B1(_03301_),
    .Y(_03310_),
    .A1(_03299_),
    .A2(_03309_));
 sg13g2_mux2_1 _08789_ (.A0(\i_tinyqv.cpu.imm[23] ),
    .A1(_03310_),
    .S(net37),
    .X(_00452_));
 sg13g2_mux4_1 _08790_ (.S0(net159),
    .A0(_00135_),
    .A1(_00137_),
    .A2(_00136_),
    .A3(_00134_),
    .S1(_02990_),
    .X(_03311_));
 sg13g2_o21ai_1 _08791_ (.B1(net84),
    .Y(_03312_),
    .A1(net86),
    .A2(_03311_));
 sg13g2_mux2_1 _08792_ (.A0(\i_tinyqv.cpu.imm[24] ),
    .A1(_03312_),
    .S(net39),
    .X(_00453_));
 sg13g2_mux2_1 _08793_ (.A0(_00139_),
    .A1(_00140_),
    .S(_02990_),
    .X(_03313_));
 sg13g2_mux2_1 _08794_ (.A0(_01475_),
    .A1(_03313_),
    .S(net183),
    .X(_03314_));
 sg13g2_nor2_1 _08795_ (.A(net90),
    .B(_03314_),
    .Y(_03315_));
 sg13g2_inv_1 _08796_ (.Y(_03316_),
    .A(_03300_));
 sg13g2_a21oi_1 _08797_ (.A1(_03210_),
    .A2(_03315_),
    .Y(_03317_),
    .B1(_03316_));
 sg13g2_nor2_1 _08798_ (.A(\i_tinyqv.cpu.imm[25] ),
    .B(net36),
    .Y(_03318_));
 sg13g2_a21oi_1 _08799_ (.A1(net38),
    .A2(_03317_),
    .Y(_00454_),
    .B1(_03318_));
 sg13g2_o21ai_1 _08800_ (.B1(net84),
    .Y(_03319_),
    .A1(_02940_),
    .A2(net86));
 sg13g2_mux2_1 _08801_ (.A0(\i_tinyqv.cpu.imm[26] ),
    .A1(_03319_),
    .S(net39),
    .X(_00455_));
 sg13g2_o21ai_1 _08802_ (.B1(net84),
    .Y(_03320_),
    .A1(_02991_),
    .A2(net86));
 sg13g2_mux2_1 _08803_ (.A0(\i_tinyqv.cpu.imm[27] ),
    .A1(_03320_),
    .S(net39),
    .X(_00456_));
 sg13g2_mux2_1 _08804_ (.A0(_00147_),
    .A1(_00148_),
    .S(net127),
    .X(_03321_));
 sg13g2_mux2_1 _08805_ (.A0(_01484_),
    .A1(_03321_),
    .S(_03000_),
    .X(_03322_));
 sg13g2_o21ai_1 _08806_ (.B1(net84),
    .Y(_03323_),
    .A1(net86),
    .A2(_03322_));
 sg13g2_mux2_1 _08807_ (.A0(\i_tinyqv.cpu.imm[28] ),
    .A1(_03323_),
    .S(net39),
    .X(_00457_));
 sg13g2_mux2_1 _08808_ (.A0(_00119_),
    .A1(_00120_),
    .S(net127),
    .X(_03324_));
 sg13g2_mux2_1 _08809_ (.A0(_01311_),
    .A1(_03324_),
    .S(_03000_),
    .X(_03325_));
 sg13g2_o21ai_1 _08810_ (.B1(net84),
    .Y(_03326_),
    .A1(net86),
    .A2(_03325_));
 sg13g2_mux2_1 _08811_ (.A0(\i_tinyqv.cpu.imm[29] ),
    .A1(_03326_),
    .S(net39),
    .X(_00458_));
 sg13g2_a22oi_1 _08812_ (.Y(_03327_),
    .B1(_03294_),
    .B2(_03161_),
    .A2(net94),
    .A1(_03168_));
 sg13g2_o21ai_1 _08813_ (.B1(net96),
    .Y(_03328_),
    .A1(net95),
    .A2(_03192_));
 sg13g2_buf_1 _08814_ (.A(_01457_),
    .X(_03329_));
 sg13g2_nor2_1 _08815_ (.A(net113),
    .B(net107),
    .Y(_03330_));
 sg13g2_nand3_1 _08816_ (.B(_03206_),
    .C(_03330_),
    .A(net100),
    .Y(_03331_));
 sg13g2_nor2b_1 _08817_ (.A(net123),
    .B_N(_03176_),
    .Y(_03332_));
 sg13g2_a21oi_1 _08818_ (.A1(_03328_),
    .A2(_03331_),
    .Y(_03333_),
    .B1(_03332_));
 sg13g2_o21ai_1 _08819_ (.B1(net106),
    .Y(_03334_),
    .A1(net104),
    .A2(net115));
 sg13g2_nor3_1 _08820_ (.A(net129),
    .B(_03179_),
    .C(_03334_),
    .Y(_03335_));
 sg13g2_or2_1 _08821_ (.X(_03336_),
    .B(_03161_),
    .A(_03157_));
 sg13g2_buf_1 _08822_ (.A(_03336_),
    .X(_03337_));
 sg13g2_nor2_1 _08823_ (.A(_03306_),
    .B(_03337_),
    .Y(_03338_));
 sg13g2_nor3_1 _08824_ (.A(_03333_),
    .B(_03335_),
    .C(_03338_),
    .Y(_03339_));
 sg13g2_o21ai_1 _08825_ (.B1(_03339_),
    .Y(_03340_),
    .A1(_01478_),
    .A2(_03327_));
 sg13g2_nand2_1 _08826_ (.Y(_03341_),
    .A(net42),
    .B(_03340_));
 sg13g2_o21ai_1 _08827_ (.B1(_03341_),
    .Y(_00459_),
    .A1(_02317_),
    .A2(net40));
 sg13g2_o21ai_1 _08828_ (.B1(_03301_),
    .Y(_03342_),
    .A1(_03001_),
    .A2(_03299_));
 sg13g2_mux2_1 _08829_ (.A0(\i_tinyqv.cpu.imm[30] ),
    .A1(_03342_),
    .S(_02916_),
    .X(_00460_));
 sg13g2_buf_1 _08830_ (.A(_02920_),
    .X(_03343_));
 sg13g2_a21oi_1 _08831_ (.A1(_03343_),
    .A2(_03220_),
    .Y(_03344_),
    .B1(_03268_));
 sg13g2_nor2_1 _08832_ (.A(\i_tinyqv.cpu.imm[31] ),
    .B(net36),
    .Y(_03345_));
 sg13g2_a21oi_1 _08833_ (.A1(net40),
    .A2(_03344_),
    .Y(_00461_),
    .B1(_03345_));
 sg13g2_nand2_1 _08834_ (.Y(_03346_),
    .A(net106),
    .B(_02980_));
 sg13g2_a21oi_1 _08835_ (.A1(net115),
    .A2(_03346_),
    .Y(_03347_),
    .B1(net114));
 sg13g2_a22oi_1 _08836_ (.Y(_03348_),
    .B1(_03206_),
    .B2(net114),
    .A2(_01466_),
    .A1(_01345_));
 sg13g2_nor3_1 _08837_ (.A(net91),
    .B(net95),
    .C(_03348_),
    .Y(_03349_));
 sg13g2_a21oi_1 _08838_ (.A1(net89),
    .A2(_03347_),
    .Y(_03350_),
    .B1(_03349_));
 sg13g2_a21oi_1 _08839_ (.A1(net136),
    .A2(_03176_),
    .Y(_03351_),
    .B1(_03350_));
 sg13g2_nor2_1 _08840_ (.A(_01362_),
    .B(net117),
    .Y(_03352_));
 sg13g2_nor2_1 _08841_ (.A(_02918_),
    .B(_02980_),
    .Y(_03353_));
 sg13g2_nor2_1 _08842_ (.A(_03352_),
    .B(_03353_),
    .Y(_03354_));
 sg13g2_o21ai_1 _08843_ (.B1(_02957_),
    .Y(_03355_),
    .A1(net101),
    .A2(_03354_));
 sg13g2_a22oi_1 _08844_ (.Y(_03356_),
    .B1(_03355_),
    .B2(net115),
    .A2(_03161_),
    .A1(_03294_));
 sg13g2_nand2b_1 _08845_ (.Y(_03357_),
    .B(_01474_),
    .A_N(_03356_));
 sg13g2_o21ai_1 _08846_ (.B1(_03357_),
    .Y(_03358_),
    .A1(_03309_),
    .A2(_03337_));
 sg13g2_o21ai_1 _08847_ (.B1(_03183_),
    .Y(_03359_),
    .A1(_03351_),
    .A2(_03358_));
 sg13g2_o21ai_1 _08848_ (.B1(_03359_),
    .Y(_00462_),
    .A1(_02338_),
    .A2(_02915_));
 sg13g2_nor2_1 _08849_ (.A(net117),
    .B(net107),
    .Y(_03360_));
 sg13g2_a22oi_1 _08850_ (.Y(_03361_),
    .B1(_03195_),
    .B2(net107),
    .A2(_03360_),
    .A1(net128));
 sg13g2_nor2_1 _08851_ (.A(net101),
    .B(_03361_),
    .Y(_03362_));
 sg13g2_a21oi_1 _08852_ (.A1(net101),
    .A2(net99),
    .Y(_03363_),
    .B1(_03362_));
 sg13g2_nor2_1 _08853_ (.A(net114),
    .B(_03363_),
    .Y(_03364_));
 sg13g2_inv_1 _08854_ (.Y(_03365_),
    .A(_03364_));
 sg13g2_a21oi_1 _08855_ (.A1(_03356_),
    .A2(_03365_),
    .Y(_03366_),
    .B1(_02949_));
 sg13g2_nor2_1 _08856_ (.A(_03311_),
    .B(_03337_),
    .Y(_03367_));
 sg13g2_a21oi_1 _08857_ (.A1(net115),
    .A2(_02960_),
    .Y(_03368_),
    .B1(_03201_));
 sg13g2_a22oi_1 _08858_ (.Y(_03369_),
    .B1(_03368_),
    .B2(_03173_),
    .A2(_03176_),
    .A1(net129));
 sg13g2_nor3_1 _08859_ (.A(_03366_),
    .B(_03367_),
    .C(_03369_),
    .Y(_03370_));
 sg13g2_nor2_1 _08860_ (.A(_01041_),
    .B(net36),
    .Y(_03371_));
 sg13g2_a21oi_1 _08861_ (.A1(net40),
    .A2(_03370_),
    .Y(_00463_),
    .B1(_03371_));
 sg13g2_o21ai_1 _08862_ (.B1(net108),
    .Y(_03372_),
    .A1(net102),
    .A2(net116));
 sg13g2_nand2_1 _08863_ (.Y(_03373_),
    .A(net113),
    .B(_03186_));
 sg13g2_nor2_1 _08864_ (.A(_03212_),
    .B(_03191_),
    .Y(_03374_));
 sg13g2_a221oi_1 _08865_ (.B2(net116),
    .C1(net97),
    .B1(_03374_),
    .A1(_03213_),
    .Y(_03375_),
    .A2(_03373_));
 sg13g2_nand2_1 _08866_ (.Y(_03376_),
    .A(_03372_),
    .B(_03375_));
 sg13g2_a22oi_1 _08867_ (.Y(_03377_),
    .B1(_03315_),
    .B2(_03155_),
    .A2(_03193_),
    .A1(_01474_));
 sg13g2_a21oi_1 _08868_ (.A1(_03206_),
    .A2(_03186_),
    .Y(_03378_),
    .B1(_02986_));
 sg13g2_o21ai_1 _08869_ (.B1(net130),
    .Y(_03379_),
    .A1(_03201_),
    .A2(_03378_));
 sg13g2_nand4_1 _08870_ (.B(_03376_),
    .C(_03377_),
    .A(_02914_),
    .Y(_03380_),
    .D(_03379_));
 sg13g2_o21ai_1 _08871_ (.B1(_03380_),
    .Y(_03381_),
    .A1(_01091_),
    .A2(_03183_));
 sg13g2_inv_1 _08872_ (.Y(_00464_),
    .A(_03381_));
 sg13g2_nor2_1 _08873_ (.A(net97),
    .B(_03173_),
    .Y(_03382_));
 sg13g2_nand3_1 _08874_ (.B(net115),
    .C(_02960_),
    .A(net130),
    .Y(_03383_));
 sg13g2_o21ai_1 _08875_ (.B1(_03383_),
    .Y(_03384_),
    .A1(_02940_),
    .A2(_03157_));
 sg13g2_a21oi_1 _08876_ (.A1(_03168_),
    .A2(net94),
    .Y(_03385_),
    .B1(_03364_));
 sg13g2_nor2_1 _08877_ (.A(_01491_),
    .B(_03385_),
    .Y(_03386_));
 sg13g2_a21o_1 _08878_ (.A2(_03198_),
    .A1(net108),
    .B1(net95),
    .X(_03387_));
 sg13g2_nand3_1 _08879_ (.B(net96),
    .C(_03387_),
    .A(net115),
    .Y(_03388_));
 sg13g2_nor2_1 _08880_ (.A(net117),
    .B(net128),
    .Y(_03389_));
 sg13g2_a22oi_1 _08881_ (.Y(_03390_),
    .B1(_03389_),
    .B2(net113),
    .A2(_03330_),
    .A1(net99));
 sg13g2_nand2b_1 _08882_ (.Y(_03391_),
    .B(net100),
    .A_N(_03390_));
 sg13g2_a21oi_1 _08883_ (.A1(_03388_),
    .A2(_03391_),
    .Y(_03392_),
    .B1(net136));
 sg13g2_nor4_1 _08884_ (.A(_03382_),
    .B(_03384_),
    .C(_03386_),
    .D(_03392_),
    .Y(_03393_));
 sg13g2_nor2_1 _08885_ (.A(_00920_),
    .B(_03266_),
    .Y(_03394_));
 sg13g2_a21oi_1 _08886_ (.A1(net40),
    .A2(_03393_),
    .Y(_00465_),
    .B1(_03394_));
 sg13g2_inv_1 _08887_ (.Y(_03395_),
    .A(_00956_));
 sg13g2_nor2_1 _08888_ (.A(_03186_),
    .B(_03352_),
    .Y(_03396_));
 sg13g2_a21oi_1 _08889_ (.A1(_03169_),
    .A2(_03352_),
    .Y(_03397_),
    .B1(_03396_));
 sg13g2_nor3_1 _08890_ (.A(net101),
    .B(net122),
    .C(_03397_),
    .Y(_03398_));
 sg13g2_a21oi_1 _08891_ (.A1(_01351_),
    .A2(_03378_),
    .Y(_03399_),
    .B1(_03398_));
 sg13g2_o21ai_1 _08892_ (.B1(_03399_),
    .Y(_03400_),
    .A1(_02991_),
    .A2(_03157_));
 sg13g2_nor2_1 _08893_ (.A(_03382_),
    .B(_03400_),
    .Y(_03401_));
 sg13g2_o21ai_1 _08894_ (.B1(_03401_),
    .Y(_03402_),
    .A1(_02923_),
    .A2(_03368_));
 sg13g2_nand2_1 _08895_ (.Y(_03403_),
    .A(net42),
    .B(_03402_));
 sg13g2_o21ai_1 _08896_ (.B1(_03403_),
    .Y(_00466_),
    .A1(_03395_),
    .A2(_03237_));
 sg13g2_nor2_1 _08897_ (.A(_03157_),
    .B(_03322_),
    .Y(_03404_));
 sg13g2_a221oi_1 _08898_ (.B2(_01479_),
    .C1(_03404_),
    .B1(_03364_),
    .A1(net123),
    .Y(_03405_),
    .A2(_03201_));
 sg13g2_o21ai_1 _08899_ (.B1(_03405_),
    .Y(_03406_),
    .A1(net97),
    .A2(_03190_));
 sg13g2_mux2_1 _08900_ (.A0(net306),
    .A1(_03406_),
    .S(net39),
    .X(_00467_));
 sg13g2_nor2_1 _08901_ (.A(net91),
    .B(_03346_),
    .Y(_03407_));
 sg13g2_a21oi_1 _08902_ (.A1(net91),
    .A2(net108),
    .Y(_03408_),
    .B1(_03407_));
 sg13g2_nand2_1 _08903_ (.Y(_03409_),
    .A(net116),
    .B(_01474_));
 sg13g2_nor3_1 _08904_ (.A(_03205_),
    .B(_03408_),
    .C(_03409_),
    .Y(_03410_));
 sg13g2_nor2_1 _08905_ (.A(_03157_),
    .B(_03325_),
    .Y(_03411_));
 sg13g2_nor3_1 _08906_ (.A(_03203_),
    .B(_03410_),
    .C(_03411_),
    .Y(_03412_));
 sg13g2_nor2_1 _08907_ (.A(net302),
    .B(_03266_),
    .Y(_03413_));
 sg13g2_a21oi_1 _08908_ (.A1(net40),
    .A2(_03412_),
    .Y(_00468_),
    .B1(_03413_));
 sg13g2_inv_1 _08909_ (.Y(_03414_),
    .A(_01282_));
 sg13g2_nand2_2 _08910_ (.Y(_03415_),
    .A(_01165_),
    .B(_01279_));
 sg13g2_nand2b_1 _08911_ (.Y(_03416_),
    .B(_03415_),
    .A_N(_01529_));
 sg13g2_buf_2 _08912_ (.A(_03416_),
    .X(_03417_));
 sg13g2_nor4_2 _08913_ (.A(_01431_),
    .B(_03414_),
    .C(_01433_),
    .Y(_03418_),
    .D(_03417_));
 sg13g2_nor2b_1 _08914_ (.A(net298),
    .B_N(_03418_),
    .Y(_03419_));
 sg13g2_nand2b_1 _08915_ (.Y(_03420_),
    .B(_03419_),
    .A_N(_01396_));
 sg13g2_buf_2 _08916_ (.A(_03420_),
    .X(_03421_));
 sg13g2_buf_1 _08917_ (.A(_03421_),
    .X(_03422_));
 sg13g2_o21ai_1 _08918_ (.B1(_03421_),
    .Y(_03423_),
    .A1(\i_tinyqv.cpu.instr_data[0][0] ),
    .A2(net260));
 sg13g2_o21ai_1 _08919_ (.B1(_03423_),
    .Y(_00469_),
    .A1(_02234_),
    .A2(net51));
 sg13g2_buf_2 _08920_ (.A(_00209_),
    .X(_03424_));
 sg13g2_buf_1 _08921_ (.A(_03421_),
    .X(_03425_));
 sg13g2_nand2_1 _08922_ (.Y(_03426_),
    .A(\i_tinyqv.cpu.instr_data[0][10] ),
    .B(net50));
 sg13g2_o21ai_1 _08923_ (.B1(_03426_),
    .Y(_00470_),
    .A1(_03424_),
    .A2(net51));
 sg13g2_buf_2 _08924_ (.A(_00210_),
    .X(_03427_));
 sg13g2_nand2_1 _08925_ (.Y(_03428_),
    .A(\i_tinyqv.cpu.instr_data[0][11] ),
    .B(net50));
 sg13g2_o21ai_1 _08926_ (.B1(_03428_),
    .Y(_00471_),
    .A1(_03427_),
    .A2(net51));
 sg13g2_buf_2 _08927_ (.A(_00204_),
    .X(_03429_));
 sg13g2_nand2_1 _08928_ (.Y(_03430_),
    .A(\i_tinyqv.cpu.instr_data[0][12] ),
    .B(net50));
 sg13g2_o21ai_1 _08929_ (.B1(_03430_),
    .Y(_00472_),
    .A1(_03429_),
    .A2(net51));
 sg13g2_buf_2 _08930_ (.A(_00205_),
    .X(_03431_));
 sg13g2_nand2_1 _08931_ (.Y(_03432_),
    .A(\i_tinyqv.cpu.instr_data[0][13] ),
    .B(_03425_));
 sg13g2_o21ai_1 _08932_ (.B1(_03432_),
    .Y(_00473_),
    .A1(_03431_),
    .A2(net51));
 sg13g2_buf_2 _08933_ (.A(_00211_),
    .X(_03433_));
 sg13g2_nand2_1 _08934_ (.Y(_03434_),
    .A(\i_tinyqv.cpu.instr_data[0][14] ),
    .B(_03421_));
 sg13g2_o21ai_1 _08935_ (.B1(_03434_),
    .Y(_00474_),
    .A1(_03433_),
    .A2(_03422_));
 sg13g2_buf_2 _08936_ (.A(_00206_),
    .X(_03435_));
 sg13g2_nand2_1 _08937_ (.Y(_03436_),
    .A(\i_tinyqv.cpu.instr_data[0][15] ),
    .B(_03421_));
 sg13g2_o21ai_1 _08938_ (.B1(_03436_),
    .Y(_00475_),
    .A1(_03435_),
    .A2(net51));
 sg13g2_o21ai_1 _08939_ (.B1(_03421_),
    .Y(_03437_),
    .A1(net260),
    .A2(\i_tinyqv.cpu.instr_data[0][1] ));
 sg13g2_o21ai_1 _08940_ (.B1(_03437_),
    .Y(_00476_),
    .A1(_02590_),
    .A2(_03422_));
 sg13g2_mux2_1 _08941_ (.A0(_02681_),
    .A1(\i_tinyqv.cpu.instr_data[0][2] ),
    .S(net50),
    .X(_00477_));
 sg13g2_mux2_1 _08942_ (.A0(_02791_),
    .A1(\i_tinyqv.cpu.instr_data[0][3] ),
    .S(net50),
    .X(_00478_));
 sg13g2_mux2_1 _08943_ (.A0(_02235_),
    .A1(\i_tinyqv.cpu.instr_data[0][4] ),
    .S(_03425_),
    .X(_00479_));
 sg13g2_mux2_1 _08944_ (.A0(_02591_),
    .A1(\i_tinyqv.cpu.instr_data[0][5] ),
    .S(net50),
    .X(_00480_));
 sg13g2_mux2_1 _08945_ (.A0(_02682_),
    .A1(\i_tinyqv.cpu.instr_data[0][6] ),
    .S(net50),
    .X(_00481_));
 sg13g2_mux2_1 _08946_ (.A0(_02781_),
    .A1(\i_tinyqv.cpu.instr_data[0][7] ),
    .S(net50),
    .X(_00482_));
 sg13g2_buf_2 _08947_ (.A(_00207_),
    .X(_03438_));
 sg13g2_nand2_1 _08948_ (.Y(_03439_),
    .A(\i_tinyqv.cpu.instr_data[0][8] ),
    .B(_03421_));
 sg13g2_o21ai_1 _08949_ (.B1(_03439_),
    .Y(_00483_),
    .A1(_03438_),
    .A2(net51));
 sg13g2_buf_2 _08950_ (.A(_00208_),
    .X(_03440_));
 sg13g2_nand2_1 _08951_ (.Y(_03441_),
    .A(\i_tinyqv.cpu.instr_data[0][9] ),
    .B(_03421_));
 sg13g2_o21ai_1 _08952_ (.B1(_03441_),
    .Y(_00484_),
    .A1(_03440_),
    .A2(net51));
 sg13g2_nand2_1 _08953_ (.Y(_03442_),
    .A(_01396_),
    .B(_03419_));
 sg13g2_buf_2 _08954_ (.A(_03442_),
    .X(_03443_));
 sg13g2_buf_1 _08955_ (.A(_03443_),
    .X(_03444_));
 sg13g2_o21ai_1 _08956_ (.B1(_03443_),
    .Y(_03445_),
    .A1(\i_tinyqv.cpu.instr_data[1][0] ),
    .A2(net260));
 sg13g2_o21ai_1 _08957_ (.B1(_03445_),
    .Y(_00485_),
    .A1(_02234_),
    .A2(_03444_));
 sg13g2_buf_1 _08958_ (.A(_03443_),
    .X(_03446_));
 sg13g2_nand2_1 _08959_ (.Y(_03447_),
    .A(\i_tinyqv.cpu.instr_data[1][10] ),
    .B(net48));
 sg13g2_o21ai_1 _08960_ (.B1(_03447_),
    .Y(_00486_),
    .A1(_03424_),
    .A2(net49));
 sg13g2_nand2_1 _08961_ (.Y(_03448_),
    .A(\i_tinyqv.cpu.instr_data[1][11] ),
    .B(net48));
 sg13g2_o21ai_1 _08962_ (.B1(_03448_),
    .Y(_00487_),
    .A1(_03427_),
    .A2(net49));
 sg13g2_nand2_1 _08963_ (.Y(_03449_),
    .A(\i_tinyqv.cpu.instr_data[1][12] ),
    .B(net48));
 sg13g2_o21ai_1 _08964_ (.B1(_03449_),
    .Y(_00488_),
    .A1(_03429_),
    .A2(net49));
 sg13g2_nand2_1 _08965_ (.Y(_03450_),
    .A(\i_tinyqv.cpu.instr_data[1][13] ),
    .B(_03446_));
 sg13g2_o21ai_1 _08966_ (.B1(_03450_),
    .Y(_00489_),
    .A1(_03431_),
    .A2(net49));
 sg13g2_nand2_1 _08967_ (.Y(_03451_),
    .A(\i_tinyqv.cpu.instr_data[1][14] ),
    .B(_03443_));
 sg13g2_o21ai_1 _08968_ (.B1(_03451_),
    .Y(_00490_),
    .A1(_03433_),
    .A2(net49));
 sg13g2_nand2_1 _08969_ (.Y(_03452_),
    .A(\i_tinyqv.cpu.instr_data[1][15] ),
    .B(_03443_));
 sg13g2_o21ai_1 _08970_ (.B1(_03452_),
    .Y(_00491_),
    .A1(_03435_),
    .A2(net49));
 sg13g2_o21ai_1 _08971_ (.B1(_03443_),
    .Y(_03453_),
    .A1(net260),
    .A2(\i_tinyqv.cpu.instr_data[1][1] ));
 sg13g2_o21ai_1 _08972_ (.B1(_03453_),
    .Y(_00492_),
    .A1(_02590_),
    .A2(_03444_));
 sg13g2_mux2_1 _08973_ (.A0(_02681_),
    .A1(\i_tinyqv.cpu.instr_data[1][2] ),
    .S(net48),
    .X(_00493_));
 sg13g2_mux2_1 _08974_ (.A0(_02791_),
    .A1(\i_tinyqv.cpu.instr_data[1][3] ),
    .S(net48),
    .X(_00494_));
 sg13g2_mux2_1 _08975_ (.A0(_02235_),
    .A1(\i_tinyqv.cpu.instr_data[1][4] ),
    .S(_03446_),
    .X(_00495_));
 sg13g2_mux2_1 _08976_ (.A0(_02591_),
    .A1(\i_tinyqv.cpu.instr_data[1][5] ),
    .S(net48),
    .X(_00496_));
 sg13g2_mux2_1 _08977_ (.A0(_02682_),
    .A1(\i_tinyqv.cpu.instr_data[1][6] ),
    .S(net48),
    .X(_00497_));
 sg13g2_mux2_1 _08978_ (.A0(_02781_),
    .A1(\i_tinyqv.cpu.instr_data[1][7] ),
    .S(net48),
    .X(_00498_));
 sg13g2_nand2_1 _08979_ (.Y(_03454_),
    .A(\i_tinyqv.cpu.instr_data[1][8] ),
    .B(_03443_));
 sg13g2_o21ai_1 _08980_ (.B1(_03454_),
    .Y(_00499_),
    .A1(_03438_),
    .A2(net49));
 sg13g2_nand2_1 _08981_ (.Y(_03455_),
    .A(\i_tinyqv.cpu.instr_data[1][9] ),
    .B(_03443_));
 sg13g2_o21ai_1 _08982_ (.B1(_03455_),
    .Y(_00500_),
    .A1(_03440_),
    .A2(net49));
 sg13g2_nand3b_1 _08983_ (.B(_03418_),
    .C(net298),
    .Y(_03456_),
    .A_N(_01396_));
 sg13g2_buf_2 _08984_ (.A(_03456_),
    .X(_03457_));
 sg13g2_buf_1 _08985_ (.A(_03457_),
    .X(_03458_));
 sg13g2_o21ai_1 _08986_ (.B1(_03457_),
    .Y(_03459_),
    .A1(\i_tinyqv.cpu.instr_data[2][0] ),
    .A2(net260));
 sg13g2_o21ai_1 _08987_ (.B1(_03459_),
    .Y(_00501_),
    .A1(_02234_),
    .A2(net55));
 sg13g2_buf_1 _08988_ (.A(_03457_),
    .X(_03460_));
 sg13g2_nand2_1 _08989_ (.Y(_03461_),
    .A(\i_tinyqv.cpu.instr_data[2][10] ),
    .B(net54));
 sg13g2_o21ai_1 _08990_ (.B1(_03461_),
    .Y(_00502_),
    .A1(_03424_),
    .A2(net55));
 sg13g2_nand2_1 _08991_ (.Y(_03462_),
    .A(\i_tinyqv.cpu.instr_data[2][11] ),
    .B(net54));
 sg13g2_o21ai_1 _08992_ (.B1(_03462_),
    .Y(_00503_),
    .A1(_03427_),
    .A2(net55));
 sg13g2_nand2_1 _08993_ (.Y(_03463_),
    .A(\i_tinyqv.cpu.instr_data[2][12] ),
    .B(net54));
 sg13g2_o21ai_1 _08994_ (.B1(_03463_),
    .Y(_00504_),
    .A1(_03429_),
    .A2(net55));
 sg13g2_nand2_1 _08995_ (.Y(_03464_),
    .A(\i_tinyqv.cpu.instr_data[2][13] ),
    .B(_03460_));
 sg13g2_o21ai_1 _08996_ (.B1(_03464_),
    .Y(_00505_),
    .A1(_03431_),
    .A2(net55));
 sg13g2_nand2_1 _08997_ (.Y(_03465_),
    .A(\i_tinyqv.cpu.instr_data[2][14] ),
    .B(_03457_));
 sg13g2_o21ai_1 _08998_ (.B1(_03465_),
    .Y(_00506_),
    .A1(_03433_),
    .A2(_03458_));
 sg13g2_nand2_1 _08999_ (.Y(_03466_),
    .A(\i_tinyqv.cpu.instr_data[2][15] ),
    .B(_03457_));
 sg13g2_o21ai_1 _09000_ (.B1(_03466_),
    .Y(_00507_),
    .A1(_03435_),
    .A2(net55));
 sg13g2_o21ai_1 _09001_ (.B1(_03457_),
    .Y(_03467_),
    .A1(net260),
    .A2(\i_tinyqv.cpu.instr_data[2][1] ));
 sg13g2_o21ai_1 _09002_ (.B1(_03467_),
    .Y(_00508_),
    .A1(_02590_),
    .A2(_03458_));
 sg13g2_mux2_1 _09003_ (.A0(_02681_),
    .A1(\i_tinyqv.cpu.instr_data[2][2] ),
    .S(net54),
    .X(_00509_));
 sg13g2_mux2_1 _09004_ (.A0(_02791_),
    .A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .S(net54),
    .X(_00510_));
 sg13g2_mux2_1 _09005_ (.A0(_02235_),
    .A1(\i_tinyqv.cpu.instr_data[2][4] ),
    .S(_03460_),
    .X(_00511_));
 sg13g2_mux2_1 _09006_ (.A0(_02591_),
    .A1(\i_tinyqv.cpu.instr_data[2][5] ),
    .S(net54),
    .X(_00512_));
 sg13g2_mux2_1 _09007_ (.A0(_02682_),
    .A1(\i_tinyqv.cpu.instr_data[2][6] ),
    .S(net54),
    .X(_00513_));
 sg13g2_mux2_1 _09008_ (.A0(_02781_),
    .A1(\i_tinyqv.cpu.instr_data[2][7] ),
    .S(net54),
    .X(_00514_));
 sg13g2_nand2_1 _09009_ (.Y(_03468_),
    .A(\i_tinyqv.cpu.instr_data[2][8] ),
    .B(_03457_));
 sg13g2_o21ai_1 _09010_ (.B1(_03468_),
    .Y(_00515_),
    .A1(_03438_),
    .A2(net55));
 sg13g2_nand2_1 _09011_ (.Y(_03469_),
    .A(\i_tinyqv.cpu.instr_data[2][9] ),
    .B(_03457_));
 sg13g2_o21ai_1 _09012_ (.B1(_03469_),
    .Y(_00516_),
    .A1(_03440_),
    .A2(net55));
 sg13g2_buf_1 _09013_ (.A(_01282_),
    .X(_03470_));
 sg13g2_buf_1 _09014_ (.A(_01529_),
    .X(_03471_));
 sg13g2_nor2_1 _09015_ (.A(net81),
    .B(net83),
    .Y(_03472_));
 sg13g2_buf_1 _09016_ (.A(_03472_),
    .X(_03473_));
 sg13g2_nand4_1 _09017_ (.B(_01396_),
    .C(_01439_),
    .A(net298),
    .Y(_03474_),
    .D(_03473_));
 sg13g2_buf_1 _09018_ (.A(_03474_),
    .X(_03475_));
 sg13g2_nand2_1 _09019_ (.Y(_03476_),
    .A(\i_tinyqv.cpu.instr_data[3][0] ),
    .B(_03475_));
 sg13g2_or2_1 _09020_ (.X(_03477_),
    .B(_03475_),
    .A(_02234_));
 sg13g2_nand3_1 _09021_ (.B(_03476_),
    .C(_03477_),
    .A(net241),
    .Y(_00517_));
 sg13g2_nand3_1 _09022_ (.B(_01396_),
    .C(_03418_),
    .A(net298),
    .Y(_03478_));
 sg13g2_buf_1 _09023_ (.A(_03478_),
    .X(_03479_));
 sg13g2_buf_1 _09024_ (.A(_03479_),
    .X(_03480_));
 sg13g2_buf_1 _09025_ (.A(_03479_),
    .X(_03481_));
 sg13g2_nand2_1 _09026_ (.Y(_03482_),
    .A(\i_tinyqv.cpu.instr_data[3][10] ),
    .B(net52));
 sg13g2_o21ai_1 _09027_ (.B1(_03482_),
    .Y(_00518_),
    .A1(_03424_),
    .A2(net53));
 sg13g2_nand2_1 _09028_ (.Y(_03483_),
    .A(\i_tinyqv.cpu.instr_data[3][11] ),
    .B(net52));
 sg13g2_o21ai_1 _09029_ (.B1(_03483_),
    .Y(_00519_),
    .A1(_03427_),
    .A2(net53));
 sg13g2_nand2_1 _09030_ (.Y(_03484_),
    .A(\i_tinyqv.cpu.instr_data[3][12] ),
    .B(net52));
 sg13g2_o21ai_1 _09031_ (.B1(_03484_),
    .Y(_00520_),
    .A1(_03429_),
    .A2(_03480_));
 sg13g2_nand2_1 _09032_ (.Y(_03485_),
    .A(\i_tinyqv.cpu.instr_data[3][13] ),
    .B(net52));
 sg13g2_o21ai_1 _09033_ (.B1(_03485_),
    .Y(_00521_),
    .A1(_03431_),
    .A2(net53));
 sg13g2_nand2_1 _09034_ (.Y(_03486_),
    .A(\i_tinyqv.cpu.instr_data[3][14] ),
    .B(_03481_));
 sg13g2_o21ai_1 _09035_ (.B1(_03486_),
    .Y(_00522_),
    .A1(_03433_),
    .A2(net53));
 sg13g2_nand2_1 _09036_ (.Y(_03487_),
    .A(\i_tinyqv.cpu.instr_data[3][15] ),
    .B(net52));
 sg13g2_o21ai_1 _09037_ (.B1(_03487_),
    .Y(_00523_),
    .A1(_03435_),
    .A2(_03480_));
 sg13g2_or2_1 _09038_ (.X(_03488_),
    .B(_03475_),
    .A(_02590_));
 sg13g2_nand2_1 _09039_ (.Y(_03489_),
    .A(\i_tinyqv.cpu.instr_data[3][1] ),
    .B(_03475_));
 sg13g2_nand3_1 _09040_ (.B(_03488_),
    .C(_03489_),
    .A(net241),
    .Y(_00524_));
 sg13g2_mux2_1 _09041_ (.A0(_02681_),
    .A1(\i_tinyqv.cpu.instr_data[3][2] ),
    .S(net53),
    .X(_00525_));
 sg13g2_mux2_1 _09042_ (.A0(_02791_),
    .A1(\i_tinyqv.cpu.instr_data[3][3] ),
    .S(net53),
    .X(_00526_));
 sg13g2_mux2_1 _09043_ (.A0(_02235_),
    .A1(\i_tinyqv.cpu.instr_data[3][4] ),
    .S(_03481_),
    .X(_00527_));
 sg13g2_mux2_1 _09044_ (.A0(_02591_),
    .A1(\i_tinyqv.cpu.instr_data[3][5] ),
    .S(net52),
    .X(_00528_));
 sg13g2_mux2_1 _09045_ (.A0(_02682_),
    .A1(\i_tinyqv.cpu.instr_data[3][6] ),
    .S(net52),
    .X(_00529_));
 sg13g2_mux2_1 _09046_ (.A0(_02781_),
    .A1(\i_tinyqv.cpu.instr_data[3][7] ),
    .S(net52),
    .X(_00530_));
 sg13g2_nand2_1 _09047_ (.Y(_03490_),
    .A(\i_tinyqv.cpu.instr_data[3][8] ),
    .B(_03479_));
 sg13g2_o21ai_1 _09048_ (.B1(_03490_),
    .Y(_00531_),
    .A1(_03438_),
    .A2(net53));
 sg13g2_nand2_1 _09049_ (.Y(_03491_),
    .A(\i_tinyqv.cpu.instr_data[3][9] ),
    .B(_03479_));
 sg13g2_o21ai_1 _09050_ (.B1(_03491_),
    .Y(_00532_),
    .A1(_03440_),
    .A2(net53));
 sg13g2_nand2_1 _09051_ (.Y(_03492_),
    .A(_03208_),
    .B(net95));
 sg13g2_nand2_1 _09052_ (.Y(_03493_),
    .A(_01454_),
    .B(net108));
 sg13g2_nand3_1 _09053_ (.B(_01489_),
    .C(_03493_),
    .A(net103),
    .Y(_03494_));
 sg13g2_o21ai_1 _09054_ (.B1(_03494_),
    .Y(_03495_),
    .A1(_03492_),
    .A2(_03192_));
 sg13g2_nand2_1 _09055_ (.Y(_03496_),
    .A(_03329_),
    .B(_03284_));
 sg13g2_o21ai_1 _09056_ (.B1(net104),
    .Y(_03497_),
    .A1(_03212_),
    .A2(net108));
 sg13g2_a22oi_1 _09057_ (.Y(_03498_),
    .B1(_03497_),
    .B2(_02988_),
    .A2(_03496_),
    .A1(net103));
 sg13g2_a22oi_1 _09058_ (.Y(_03499_),
    .B1(_03498_),
    .B2(_01474_),
    .A2(_03495_),
    .A1(net89));
 sg13g2_nor2_1 _09059_ (.A(_01263_),
    .B(net41),
    .Y(_03500_));
 sg13g2_a21oi_1 _09060_ (.A1(net40),
    .A2(_03499_),
    .Y(_00573_),
    .B1(_03500_));
 sg13g2_nor2_1 _09061_ (.A(_02967_),
    .B(_03496_),
    .Y(_03501_));
 sg13g2_nor3_1 _09062_ (.A(_03209_),
    .B(net106),
    .C(_03374_),
    .Y(_03502_));
 sg13g2_o21ai_1 _09063_ (.B1(net41),
    .Y(_03503_),
    .A1(_03501_),
    .A2(_03502_));
 sg13g2_o21ai_1 _09064_ (.B1(_03503_),
    .Y(_00574_),
    .A1(_02702_),
    .A2(_03237_));
 sg13g2_nand2_1 _09065_ (.Y(_03504_),
    .A(_02966_),
    .B(_02944_));
 sg13g2_nor2_1 _09066_ (.A(_01455_),
    .B(_02944_),
    .Y(_03505_));
 sg13g2_a21oi_1 _09067_ (.A1(_03159_),
    .A2(_03504_),
    .Y(_03506_),
    .B1(_03505_));
 sg13g2_o21ai_1 _09068_ (.B1(net88),
    .Y(_03507_),
    .A1(_02968_),
    .A2(_03506_));
 sg13g2_nand2_1 _09069_ (.Y(_03508_),
    .A(_01351_),
    .B(_01474_));
 sg13g2_nand3_1 _09070_ (.B(_03498_),
    .C(_03508_),
    .A(_02949_),
    .Y(_03509_));
 sg13g2_o21ai_1 _09071_ (.B1(_03509_),
    .Y(_03510_),
    .A1(_02967_),
    .A2(_03507_));
 sg13g2_mux2_1 _09072_ (.A0(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .A1(_03510_),
    .S(_02916_),
    .X(_00575_));
 sg13g2_buf_1 _09073_ (.A(\i_tinyqv.cpu.mem_op_increment_reg ),
    .X(_03511_));
 sg13g2_nand4_1 _09074_ (.B(_02945_),
    .C(_03159_),
    .A(net88),
    .Y(_03512_),
    .D(_03195_));
 sg13g2_mux2_1 _09075_ (.A0(_03511_),
    .A1(_03512_),
    .S(net39),
    .X(_00576_));
 sg13g2_nor2b_1 _09076_ (.A(_01286_),
    .B_N(_01553_),
    .Y(_03513_));
 sg13g2_buf_2 _09077_ (.A(_03513_),
    .X(_03514_));
 sg13g2_buf_1 _09078_ (.A(_03514_),
    .X(_03515_));
 sg13g2_a221oi_1 _09079_ (.B2(net104),
    .C1(net94),
    .B1(net99),
    .A1(_01469_),
    .Y(_03516_),
    .A2(_01489_));
 sg13g2_a21oi_1 _09080_ (.A1(_03186_),
    .A2(_03179_),
    .Y(_03517_),
    .B1(net130));
 sg13g2_a21oi_1 _09081_ (.A1(net103),
    .A2(_03516_),
    .Y(_03518_),
    .B1(_03517_));
 sg13g2_o21ai_1 _09082_ (.B1(_03213_),
    .Y(_03519_),
    .A1(net103),
    .A2(_03516_));
 sg13g2_o21ai_1 _09083_ (.B1(net128),
    .Y(_03520_),
    .A1(_01455_),
    .A2(net117));
 sg13g2_nand2_1 _09084_ (.Y(_03521_),
    .A(net107),
    .B(_03520_));
 sg13g2_o21ai_1 _09085_ (.B1(net114),
    .Y(_03522_),
    .A1(net124),
    .A2(net107));
 sg13g2_nand2_1 _09086_ (.Y(_03523_),
    .A(net124),
    .B(_03186_));
 sg13g2_a22oi_1 _09087_ (.Y(_03524_),
    .B1(_03523_),
    .B2(net113),
    .A2(_03522_),
    .A1(net99));
 sg13g2_o21ai_1 _09088_ (.B1(_03524_),
    .Y(_03525_),
    .A1(net101),
    .A2(_03521_));
 sg13g2_nor2_1 _09089_ (.A(_01491_),
    .B(_03525_),
    .Y(_03526_));
 sg13g2_a21oi_1 _09090_ (.A1(_03518_),
    .A2(_03519_),
    .Y(_03527_),
    .B1(_03526_));
 sg13g2_nand2_1 _09091_ (.Y(_03528_),
    .A(_00213_),
    .B(_03514_));
 sg13g2_o21ai_1 _09092_ (.B1(_03528_),
    .Y(_03529_),
    .A1(net80),
    .A2(_03527_));
 sg13g2_nor2_1 _09093_ (.A(_03514_),
    .B(_02909_),
    .Y(_03530_));
 sg13g2_nor2_1 _09094_ (.A(_01643_),
    .B(_03530_),
    .Y(_03531_));
 sg13g2_buf_1 _09095_ (.A(_03531_),
    .X(_03532_));
 sg13g2_buf_1 _09096_ (.A(_03532_),
    .X(_03533_));
 sg13g2_mux2_1 _09097_ (.A0(_02521_),
    .A1(_03529_),
    .S(net45),
    .X(_00580_));
 sg13g2_buf_1 _09098_ (.A(_02904_),
    .X(_03534_));
 sg13g2_o21ai_1 _09099_ (.B1(_03532_),
    .Y(_03535_),
    .A1(_02521_),
    .A2(net79));
 sg13g2_nand2_1 _09100_ (.Y(_03536_),
    .A(_02522_),
    .B(_03514_));
 sg13g2_nor2_1 _09101_ (.A(net114),
    .B(_03186_),
    .Y(_03537_));
 sg13g2_o21ai_1 _09102_ (.B1(_03329_),
    .Y(_03538_),
    .A1(_03208_),
    .A2(net94));
 sg13g2_nand2b_1 _09103_ (.Y(_03539_),
    .B(_03538_),
    .A_N(_03537_));
 sg13g2_nand2_1 _09104_ (.Y(_03540_),
    .A(_01332_),
    .B(_03539_));
 sg13g2_o21ai_1 _09105_ (.B1(_03540_),
    .Y(_03541_),
    .A1(net122),
    .A2(_03525_));
 sg13g2_nand2_1 _09106_ (.Y(_03542_),
    .A(net79),
    .B(_03541_));
 sg13g2_and2_1 _09107_ (.A(_03536_),
    .B(_03542_),
    .X(_03543_));
 sg13g2_a22oi_1 _09108_ (.Y(_00581_),
    .B1(_03543_),
    .B2(net45),
    .A2(_03535_),
    .A1(_02838_));
 sg13g2_nand2_1 _09109_ (.Y(_03544_),
    .A(_03532_),
    .B(_03536_));
 sg13g2_nand2_1 _09110_ (.Y(_03545_),
    .A(net123),
    .B(_03539_));
 sg13g2_o21ai_1 _09111_ (.B1(_03545_),
    .Y(_03546_),
    .A1(_01478_),
    .A2(_03525_));
 sg13g2_nand4_1 _09112_ (.B(_02521_),
    .C(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .A(_02520_),
    .Y(_03547_),
    .D(_03514_));
 sg13g2_o21ai_1 _09113_ (.B1(_03547_),
    .Y(_03548_),
    .A1(net80),
    .A2(_03546_));
 sg13g2_a22oi_1 _09114_ (.Y(_00582_),
    .B1(_03548_),
    .B2(net45),
    .A2(_03544_),
    .A1(_02523_));
 sg13g2_nor2_1 _09115_ (.A(net113),
    .B(_03521_),
    .Y(_03549_));
 sg13g2_a21oi_1 _09116_ (.A1(net102),
    .A2(net104),
    .Y(_03550_),
    .B1(_03549_));
 sg13g2_a22oi_1 _09117_ (.Y(_03551_),
    .B1(_03492_),
    .B2(_01473_),
    .A2(net99),
    .A1(net102));
 sg13g2_o21ai_1 _09118_ (.B1(_03551_),
    .Y(_03552_),
    .A1(net91),
    .A2(_03550_));
 sg13g2_nand3_1 _09119_ (.B(_03538_),
    .C(_03552_),
    .A(net79),
    .Y(_03553_));
 sg13g2_o21ai_1 _09120_ (.B1(_03553_),
    .Y(_03554_),
    .A1(_02525_),
    .A2(_03547_));
 sg13g2_o21ai_1 _09121_ (.B1(net80),
    .Y(_03555_),
    .A1(_02523_),
    .A2(_02522_));
 sg13g2_a21oi_1 _09122_ (.A1(_03532_),
    .A2(_03555_),
    .Y(_03556_),
    .B1(_02524_));
 sg13g2_a21oi_1 _09123_ (.A1(net45),
    .A2(_03554_),
    .Y(_00583_),
    .B1(_03556_));
 sg13g2_and3_1 _09124_ (.X(_03557_),
    .A(_01455_),
    .B(net106),
    .C(_02944_));
 sg13g2_o21ai_1 _09125_ (.B1(_03346_),
    .Y(_03558_),
    .A1(net104),
    .A2(_03557_));
 sg13g2_a22oi_1 _09126_ (.Y(_03559_),
    .B1(_03558_),
    .B2(_03168_),
    .A2(_03360_),
    .A1(net96));
 sg13g2_inv_1 _09127_ (.Y(_03560_),
    .A(_03559_));
 sg13g2_o21ai_1 _09128_ (.B1(net117),
    .Y(_03561_),
    .A1(net100),
    .A2(net128));
 sg13g2_a22oi_1 _09129_ (.Y(_03562_),
    .B1(_03561_),
    .B2(net95),
    .A2(_03389_),
    .A1(net100));
 sg13g2_inv_1 _09130_ (.Y(_03563_),
    .A(_03562_));
 sg13g2_a22oi_1 _09131_ (.Y(_03564_),
    .B1(_03563_),
    .B2(net102),
    .A2(_03560_),
    .A1(net116));
 sg13g2_a21o_1 _09132_ (.A2(_03169_),
    .A1(_03205_),
    .B1(_03537_),
    .X(_03565_));
 sg13g2_nor2_1 _09133_ (.A(net101),
    .B(net106),
    .Y(_03566_));
 sg13g2_a22oi_1 _09134_ (.Y(_03567_),
    .B1(_03565_),
    .B2(_03566_),
    .A2(_03353_),
    .A1(net89));
 sg13g2_o21ai_1 _09135_ (.B1(_03567_),
    .Y(_03568_),
    .A1(_01491_),
    .A2(_03564_));
 sg13g2_nand2_1 _09136_ (.Y(_03569_),
    .A(net42),
    .B(_03568_));
 sg13g2_o21ai_1 _09137_ (.B1(_03569_),
    .Y(_00584_),
    .A1(_01721_),
    .A2(net37));
 sg13g2_nor2_1 _09138_ (.A(net113),
    .B(_03389_),
    .Y(_03570_));
 sg13g2_a22oi_1 _09139_ (.Y(_03571_),
    .B1(_03570_),
    .B2(_03194_),
    .A2(_03361_),
    .A1(net102));
 sg13g2_nand3_1 _09140_ (.B(net104),
    .C(_03195_),
    .A(net113),
    .Y(_03572_));
 sg13g2_nand2_1 _09141_ (.Y(_03573_),
    .A(net114),
    .B(_03262_));
 sg13g2_a21oi_1 _09142_ (.A1(_03572_),
    .A2(_03573_),
    .Y(_03574_),
    .B1(net100));
 sg13g2_a21oi_1 _09143_ (.A1(net100),
    .A2(_03571_),
    .Y(_03575_),
    .B1(_03574_));
 sg13g2_o21ai_1 _09144_ (.B1(_03575_),
    .Y(_03576_),
    .A1(net122),
    .A2(_03564_));
 sg13g2_nand2_1 _09145_ (.Y(_03577_),
    .A(net42),
    .B(_03576_));
 sg13g2_o21ai_1 _09146_ (.B1(_03577_),
    .Y(_00585_),
    .A1(_00840_),
    .A2(net37));
 sg13g2_nor2_1 _09147_ (.A(_01478_),
    .B(_03564_),
    .Y(_03578_));
 sg13g2_nor2_1 _09148_ (.A(net91),
    .B(_03192_),
    .Y(_03579_));
 sg13g2_a21oi_1 _09149_ (.A1(net89),
    .A2(_03269_),
    .Y(_03580_),
    .B1(_03579_));
 sg13g2_nor2_1 _09150_ (.A(net102),
    .B(_03580_),
    .Y(_03581_));
 sg13g2_o21ai_1 _09151_ (.B1(net41),
    .Y(_03582_),
    .A1(_03578_),
    .A2(_03581_));
 sg13g2_o21ai_1 _09152_ (.B1(_03582_),
    .Y(_00586_),
    .A1(_00794_),
    .A2(net37));
 sg13g2_o21ai_1 _09153_ (.B1(net104),
    .Y(_03583_),
    .A1(net91),
    .A2(net116));
 sg13g2_a21o_1 _09154_ (.A2(_03274_),
    .A1(net114),
    .B1(_03537_),
    .X(_03584_));
 sg13g2_a22oi_1 _09155_ (.Y(_03585_),
    .B1(_03584_),
    .B2(net89),
    .A2(_03583_),
    .A1(_03352_));
 sg13g2_o21ai_1 _09156_ (.B1(_03585_),
    .Y(_03586_),
    .A1(_03409_),
    .A2(_03559_));
 sg13g2_nand2_1 _09157_ (.Y(_03587_),
    .A(net42),
    .B(_03586_));
 sg13g2_o21ai_1 _09158_ (.B1(_03587_),
    .Y(_00587_),
    .A1(_00799_),
    .A2(net37));
 sg13g2_o21ai_1 _09159_ (.B1(_03532_),
    .Y(_03588_),
    .A1(_03511_),
    .A2(net79));
 sg13g2_nor2_1 _09160_ (.A(_03204_),
    .B(_03191_),
    .Y(_03589_));
 sg13g2_a21oi_1 _09161_ (.A1(_03589_),
    .A2(_03195_),
    .Y(_03590_),
    .B1(net130));
 sg13g2_inv_1 _09162_ (.Y(_03591_),
    .A(_03164_));
 sg13g2_a22oi_1 _09163_ (.Y(_03592_),
    .B1(_03170_),
    .B2(_02927_),
    .A2(_03591_),
    .A1(_03343_));
 sg13g2_o21ai_1 _09164_ (.B1(_03592_),
    .Y(_03593_),
    .A1(net89),
    .A2(_03590_));
 sg13g2_nand3_1 _09165_ (.B(_03511_),
    .C(_03514_),
    .A(net221),
    .Y(_03594_));
 sg13g2_o21ai_1 _09166_ (.B1(_03594_),
    .Y(_03595_),
    .A1(net80),
    .A2(_03593_));
 sg13g2_a22oi_1 _09167_ (.Y(_00588_),
    .B1(_03595_),
    .B2(net45),
    .A2(_03588_),
    .A1(_00910_));
 sg13g2_o21ai_1 _09168_ (.B1(net100),
    .Y(_03596_),
    .A1(_03204_),
    .A2(net106));
 sg13g2_nand2_1 _09169_ (.Y(_03597_),
    .A(_03373_),
    .B(_03596_));
 sg13g2_nand2_1 _09170_ (.Y(_03598_),
    .A(_01332_),
    .B(_03597_));
 sg13g2_o21ai_1 _09171_ (.B1(_03598_),
    .Y(_03599_),
    .A1(net90),
    .A2(_03291_));
 sg13g2_or2_1 _09172_ (.X(_03600_),
    .B(_03594_),
    .A(_00902_));
 sg13g2_o21ai_1 _09173_ (.B1(_03600_),
    .Y(_03601_),
    .A1(net80),
    .A2(_03599_));
 sg13g2_a21oi_1 _09174_ (.A1(net221),
    .A2(_03511_),
    .Y(_03602_),
    .B1(net79));
 sg13g2_nand2b_1 _09175_ (.Y(_03603_),
    .B(net45),
    .A_N(_03602_));
 sg13g2_a22oi_1 _09176_ (.Y(_00589_),
    .B1(_03603_),
    .B2(_00902_),
    .A2(_03601_),
    .A1(net45));
 sg13g2_nand2_1 _09177_ (.Y(_03604_),
    .A(_01339_),
    .B(_03597_));
 sg13g2_o21ai_1 _09178_ (.B1(_03604_),
    .Y(_03605_),
    .A1(net90),
    .A2(_03306_));
 sg13g2_nand3_1 _09179_ (.B(net221),
    .C(_03511_),
    .A(_00882_),
    .Y(_03606_));
 sg13g2_nor2_1 _09180_ (.A(_00875_),
    .B(_03606_),
    .Y(_03607_));
 sg13g2_nand2_1 _09181_ (.Y(_03608_),
    .A(net80),
    .B(_03607_));
 sg13g2_o21ai_1 _09182_ (.B1(_03608_),
    .Y(_03609_),
    .A1(net80),
    .A2(_03605_));
 sg13g2_nand2_1 _09183_ (.Y(_03610_),
    .A(_03515_),
    .B(_03606_));
 sg13g2_a21oi_1 _09184_ (.A1(_03532_),
    .A2(_03610_),
    .Y(_03611_),
    .B1(net224));
 sg13g2_a21oi_1 _09185_ (.A1(net45),
    .A2(_03609_),
    .Y(_00590_),
    .B1(_03611_));
 sg13g2_a21o_1 _09186_ (.A2(_03309_),
    .A1(net103),
    .B1(_03537_),
    .X(_03612_));
 sg13g2_nand2_1 _09187_ (.Y(_03613_),
    .A(_01450_),
    .B(_03374_));
 sg13g2_a21oi_1 _09188_ (.A1(_03209_),
    .A2(_03192_),
    .Y(_03614_),
    .B1(_03613_));
 sg13g2_a21oi_1 _09189_ (.A1(net89),
    .A2(_03612_),
    .Y(_03615_),
    .B1(_03614_));
 sg13g2_nand3_1 _09190_ (.B(_03514_),
    .C(_03607_),
    .A(net222),
    .Y(_03616_));
 sg13g2_o21ai_1 _09191_ (.B1(_03616_),
    .Y(_03617_),
    .A1(net80),
    .A2(_03615_));
 sg13g2_o21ai_1 _09192_ (.B1(_03533_),
    .Y(_03618_),
    .A1(net79),
    .A2(_03607_));
 sg13g2_a22oi_1 _09193_ (.Y(_00591_),
    .B1(_03618_),
    .B2(_00889_),
    .A2(_03617_),
    .A1(_03533_));
 sg13g2_nand2_1 _09194_ (.Y(_03619_),
    .A(_00154_),
    .B(_01520_));
 sg13g2_a21oi_1 _09195_ (.A1(_01501_),
    .A2(_01509_),
    .Y(_03620_),
    .B1(_03619_));
 sg13g2_buf_2 _09196_ (.A(_03620_),
    .X(_03621_));
 sg13g2_and4_1 _09197_ (.A(_01431_),
    .B(_01500_),
    .C(_01509_),
    .D(_01522_),
    .X(_03622_));
 sg13g2_buf_2 _09198_ (.A(_03622_),
    .X(_03623_));
 sg13g2_nor2_1 _09199_ (.A(_01423_),
    .B(_03623_),
    .Y(_03624_));
 sg13g2_buf_1 _09200_ (.A(_03624_),
    .X(_03625_));
 sg13g2_buf_1 _09201_ (.A(net71),
    .X(_03626_));
 sg13g2_nand3_1 _09202_ (.B(_03621_),
    .C(net62),
    .A(\addr[0] ),
    .Y(_03627_));
 sg13g2_a21o_1 _09203_ (.A2(_01509_),
    .A1(_01501_),
    .B1(_03619_),
    .X(_03628_));
 sg13g2_buf_2 _09204_ (.A(_03628_),
    .X(_03629_));
 sg13g2_buf_1 _09205_ (.A(_03629_),
    .X(_03630_));
 sg13g2_buf_2 _09206_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .X(_03631_));
 sg13g2_buf_1 _09207_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .X(_03632_));
 sg13g2_inv_1 _09208_ (.Y(_03633_),
    .A(net281));
 sg13g2_nor2_1 _09209_ (.A(_03633_),
    .B(_01517_),
    .Y(_03634_));
 sg13g2_buf_1 _09210_ (.A(_03634_),
    .X(_03635_));
 sg13g2_nand3_1 _09211_ (.B(_03631_),
    .C(net200),
    .A(_01518_),
    .Y(_03636_));
 sg13g2_buf_1 _09212_ (.A(_03636_),
    .X(_03637_));
 sg13g2_buf_1 _09213_ (.A(_03637_),
    .X(_03638_));
 sg13g2_nand3_1 _09214_ (.B(net70),
    .C(net156),
    .A(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .Y(_03639_));
 sg13g2_nand2_1 _09215_ (.Y(_00597_),
    .A(_03627_),
    .B(_03639_));
 sg13g2_buf_1 _09216_ (.A(_03629_),
    .X(_03640_));
 sg13g2_buf_1 _09217_ (.A(net71),
    .X(_03641_));
 sg13g2_buf_1 _09218_ (.A(\i_tinyqv.cpu.was_early_branch ),
    .X(_03642_));
 sg13g2_buf_1 _09219_ (.A(net280),
    .X(_03643_));
 sg13g2_xnor2_1 _09220_ (.Y(_03644_),
    .A(net257),
    .B(net285));
 sg13g2_a21o_1 _09221_ (.A2(_01090_),
    .A1(net309),
    .B1(net311),
    .X(_03645_));
 sg13g2_and3_1 _09222_ (.X(_03646_),
    .A(net309),
    .B(net311),
    .C(_01090_));
 sg13g2_a21oi_2 _09223_ (.B1(_03646_),
    .Y(_03647_),
    .A2(_03645_),
    .A1(_00758_));
 sg13g2_a22oi_1 _09224_ (.Y(_03648_),
    .B1(net303),
    .B2(_01041_),
    .A2(_00955_),
    .A1(net312));
 sg13g2_nor2_1 _09225_ (.A(net312),
    .B(_00955_),
    .Y(_03649_));
 sg13g2_nand2_1 _09226_ (.Y(_03650_),
    .A(net303),
    .B(_01041_));
 sg13g2_nor2_1 _09227_ (.A(net303),
    .B(_01041_),
    .Y(_03651_));
 sg13g2_a221oi_1 _09228_ (.B2(_03650_),
    .C1(_03651_),
    .B1(_03649_),
    .A1(_03647_),
    .Y(_03652_),
    .A2(_03648_));
 sg13g2_buf_2 _09229_ (.A(_03652_),
    .X(_03653_));
 sg13g2_inv_1 _09230_ (.Y(_03654_),
    .A(_00988_));
 sg13g2_inv_1 _09231_ (.Y(_03655_),
    .A(_01091_));
 sg13g2_nor2_1 _09232_ (.A(_00759_),
    .B(_00920_),
    .Y(_03656_));
 sg13g2_a21oi_1 _09233_ (.A1(_03654_),
    .A2(_03655_),
    .Y(_03657_),
    .B1(_03656_));
 sg13g2_a21o_1 _09234_ (.A2(_01091_),
    .A1(_00988_),
    .B1(_00920_),
    .X(_03658_));
 sg13g2_and3_1 _09235_ (.X(_03659_),
    .A(_00920_),
    .B(_00988_),
    .C(_01091_));
 sg13g2_a221oi_1 _09236_ (.B2(_00759_),
    .C1(_03659_),
    .B1(_03658_),
    .A1(_03653_),
    .Y(_03660_),
    .A2(_03657_));
 sg13g2_buf_2 _09237_ (.A(_03660_),
    .X(_03661_));
 sg13g2_or2_1 _09238_ (.X(_03662_),
    .B(net306),
    .A(net304));
 sg13g2_or2_1 _09239_ (.X(_03663_),
    .B(_00956_),
    .A(_00858_));
 sg13g2_and2_1 _09240_ (.A(net304),
    .B(net306),
    .X(_03664_));
 sg13g2_a21oi_2 _09241_ (.B1(_03664_),
    .Y(_03665_),
    .A2(_03663_),
    .A1(_03662_));
 sg13g2_nor2_1 _09242_ (.A(net287),
    .B(net302),
    .Y(_03666_));
 sg13g2_or2_1 _09243_ (.X(_03667_),
    .B(_03666_),
    .A(_03665_));
 sg13g2_and2_1 _09244_ (.A(net287),
    .B(net302),
    .X(_03668_));
 sg13g2_a21oi_2 _09245_ (.B1(_03664_),
    .Y(_03669_),
    .A2(_00956_),
    .A1(_00858_));
 sg13g2_nor3_1 _09246_ (.A(_03665_),
    .B(_03669_),
    .C(_03666_),
    .Y(_03670_));
 sg13g2_nor2_1 _09247_ (.A(_03668_),
    .B(_03670_),
    .Y(_03671_));
 sg13g2_o21ai_1 _09248_ (.B1(_03671_),
    .Y(_03672_),
    .A1(_03661_),
    .A2(_03667_));
 sg13g2_xnor2_1 _09249_ (.Y(_03673_),
    .A(_03644_),
    .B(_03672_));
 sg13g2_buf_1 _09250_ (.A(net280),
    .X(_03674_));
 sg13g2_nand2_2 _09251_ (.Y(_03675_),
    .A(net312),
    .B(_01399_));
 sg13g2_or2_1 _09252_ (.X(_03676_),
    .B(_03675_),
    .A(_02270_));
 sg13g2_buf_1 _09253_ (.A(_03676_),
    .X(_03677_));
 sg13g2_nor3_1 _09254_ (.A(_02707_),
    .B(_02267_),
    .C(_03677_),
    .Y(_03678_));
 sg13g2_xnor2_1 _09255_ (.Y(_03679_),
    .A(net257),
    .B(_03678_));
 sg13g2_nor2_1 _09256_ (.A(_03674_),
    .B(_03679_),
    .Y(_03680_));
 sg13g2_a21oi_1 _09257_ (.A1(net240),
    .A2(_03673_),
    .Y(_03681_),
    .B1(_03680_));
 sg13g2_nor2_1 _09258_ (.A(net61),
    .B(_03681_),
    .Y(_03682_));
 sg13g2_a21oi_1 _09259_ (.A1(\addr[10] ),
    .A2(net62),
    .Y(_03683_),
    .B1(_03682_));
 sg13g2_buf_1 _09260_ (.A(_01518_),
    .X(_03684_));
 sg13g2_and3_1 _09261_ (.X(_03685_),
    .A(net238),
    .B(_03631_),
    .C(net200));
 sg13g2_buf_2 _09262_ (.A(_03685_),
    .X(_03686_));
 sg13g2_nor2_1 _09263_ (.A(_03621_),
    .B(_03686_),
    .Y(_03687_));
 sg13g2_a22oi_1 _09264_ (.Y(_03688_),
    .B1(_03687_),
    .B2(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .A2(_03686_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[6] ));
 sg13g2_o21ai_1 _09265_ (.B1(_03688_),
    .Y(_00598_),
    .A1(net69),
    .A2(_03683_));
 sg13g2_nand2_1 _09266_ (.Y(_03689_),
    .A(net257),
    .B(net302));
 sg13g2_nand2_1 _09267_ (.Y(_03690_),
    .A(_00768_),
    .B(net287));
 sg13g2_a221oi_1 _09268_ (.B2(_03690_),
    .C1(_03665_),
    .B1(_03689_),
    .A1(_03661_),
    .Y(_03691_),
    .A2(_03669_));
 sg13g2_nand2_1 _09269_ (.Y(_03692_),
    .A(net285),
    .B(net302));
 sg13g2_nand2_1 _09270_ (.Y(_03693_),
    .A(net285),
    .B(net287));
 sg13g2_a221oi_1 _09271_ (.B2(_03693_),
    .C1(_03665_),
    .B1(_03692_),
    .A1(_03661_),
    .Y(_03694_),
    .A2(_03669_));
 sg13g2_nand2_1 _09272_ (.Y(_03695_),
    .A(net257),
    .B(net285));
 sg13g2_o21ai_1 _09273_ (.B1(_03668_),
    .Y(_03696_),
    .A1(net257),
    .A2(net285));
 sg13g2_nand2_1 _09274_ (.Y(_03697_),
    .A(_03695_),
    .B(_03696_));
 sg13g2_or3_1 _09275_ (.A(_03691_),
    .B(_03694_),
    .C(_03697_),
    .X(_03698_));
 sg13g2_buf_1 _09276_ (.A(_03698_),
    .X(_03699_));
 sg13g2_xnor2_1 _09277_ (.Y(_03700_),
    .A(net288),
    .B(net310));
 sg13g2_xnor2_1 _09278_ (.Y(_03701_),
    .A(_03699_),
    .B(_03700_));
 sg13g2_nor2_1 _09279_ (.A(_02284_),
    .B(_03675_),
    .Y(_03702_));
 sg13g2_and2_1 _09280_ (.A(_02618_),
    .B(_03702_),
    .X(_03703_));
 sg13g2_buf_1 _09281_ (.A(_03703_),
    .X(_03704_));
 sg13g2_xnor2_1 _09282_ (.Y(_03705_),
    .A(net288),
    .B(_03704_));
 sg13g2_nor2_1 _09283_ (.A(net239),
    .B(_03705_),
    .Y(_03706_));
 sg13g2_a21oi_1 _09284_ (.A1(net240),
    .A2(_03701_),
    .Y(_03707_),
    .B1(_03706_));
 sg13g2_nor2_1 _09285_ (.A(net61),
    .B(_03707_),
    .Y(_03708_));
 sg13g2_a21oi_1 _09286_ (.A1(\addr[11] ),
    .A2(net62),
    .Y(_03709_),
    .B1(_03708_));
 sg13g2_a22oi_1 _09287_ (.Y(_03710_),
    .B1(_03687_),
    .B2(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .A2(_03686_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[7] ));
 sg13g2_o21ai_1 _09288_ (.B1(_03710_),
    .Y(_00599_),
    .A1(net69),
    .A2(_03709_));
 sg13g2_buf_1 _09289_ (.A(net280),
    .X(_03711_));
 sg13g2_nor2_1 _09290_ (.A(_02267_),
    .B(_03677_),
    .Y(_03712_));
 sg13g2_nand2b_1 _09291_ (.Y(_03713_),
    .B(_03712_),
    .A_N(_02279_));
 sg13g2_xnor2_1 _09292_ (.Y(_03714_),
    .A(_02265_),
    .B(_03713_));
 sg13g2_buf_1 _09293_ (.A(_03642_),
    .X(_03715_));
 sg13g2_xnor2_1 _09294_ (.Y(_03716_),
    .A(net289),
    .B(_01043_));
 sg13g2_a21o_1 _09295_ (.A2(_03699_),
    .A1(net310),
    .B1(_02274_),
    .X(_03717_));
 sg13g2_o21ai_1 _09296_ (.B1(_03717_),
    .Y(_03718_),
    .A1(net310),
    .A2(_03699_));
 sg13g2_xnor2_1 _09297_ (.Y(_03719_),
    .A(_03716_),
    .B(_03718_));
 sg13g2_nand2_1 _09298_ (.Y(_03720_),
    .A(_03715_),
    .B(_03719_));
 sg13g2_o21ai_1 _09299_ (.B1(_03720_),
    .Y(_03721_),
    .A1(_03711_),
    .A2(_03714_));
 sg13g2_nor2_1 _09300_ (.A(net61),
    .B(_03721_),
    .Y(_03722_));
 sg13g2_a21oi_1 _09301_ (.A1(\addr[12] ),
    .A2(net62),
    .Y(_03723_),
    .B1(_03722_));
 sg13g2_buf_1 _09302_ (.A(_03629_),
    .X(_03724_));
 sg13g2_mux2_1 _09303_ (.A0(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .S(net156),
    .X(_03725_));
 sg13g2_nand2_1 _09304_ (.Y(_03726_),
    .A(net68),
    .B(_03725_));
 sg13g2_o21ai_1 _09305_ (.B1(_03726_),
    .Y(_00600_),
    .A1(net69),
    .A2(_03723_));
 sg13g2_nand2b_1 _09306_ (.Y(_03727_),
    .B(_03704_),
    .A_N(_02616_));
 sg13g2_xnor2_1 _09307_ (.Y(_03728_),
    .A(_02308_),
    .B(_03727_));
 sg13g2_a21o_1 _09308_ (.A2(_01043_),
    .A1(net289),
    .B1(net310),
    .X(_03729_));
 sg13g2_nor4_2 _09309_ (.A(_03691_),
    .B(_03694_),
    .C(_03697_),
    .Y(_03730_),
    .D(_03729_));
 sg13g2_nor2_2 _09310_ (.A(net289),
    .B(_01043_),
    .Y(_03731_));
 sg13g2_nor2_1 _09311_ (.A(net257),
    .B(_02318_),
    .Y(_03732_));
 sg13g2_nor2b_1 _09312_ (.A(_03732_),
    .B_N(_00969_),
    .Y(_03733_));
 sg13g2_a21oi_1 _09313_ (.A1(net289),
    .A2(_01043_),
    .Y(_03734_),
    .B1(_02274_));
 sg13g2_nand3_1 _09314_ (.B(_02275_),
    .C(_02318_),
    .A(_00969_),
    .Y(_03735_));
 sg13g2_nand2_1 _09315_ (.Y(_03736_),
    .A(_03734_),
    .B(_03735_));
 sg13g2_a21oi_2 _09316_ (.B1(_03736_),
    .Y(_03737_),
    .A2(_03733_),
    .A1(_03672_));
 sg13g2_nor3_2 _09317_ (.A(_03730_),
    .B(_03731_),
    .C(_03737_),
    .Y(_03738_));
 sg13g2_xor2_1 _09318_ (.B(_01088_),
    .A(net252),
    .X(_03739_));
 sg13g2_xnor2_1 _09319_ (.Y(_03740_),
    .A(_03738_),
    .B(_03739_));
 sg13g2_nand2_1 _09320_ (.Y(_03741_),
    .A(net236),
    .B(_03740_));
 sg13g2_o21ai_1 _09321_ (.B1(_03741_),
    .Y(_03742_),
    .A1(net237),
    .A2(_03728_));
 sg13g2_nor2_1 _09322_ (.A(net61),
    .B(_03742_),
    .Y(_03743_));
 sg13g2_a21oi_1 _09323_ (.A1(\addr[13] ),
    .A2(net62),
    .Y(_03744_),
    .B1(_03743_));
 sg13g2_mux2_1 _09324_ (.A0(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .S(_03638_),
    .X(_03745_));
 sg13g2_nand2_1 _09325_ (.Y(_03746_),
    .A(net68),
    .B(_03745_));
 sg13g2_o21ai_1 _09326_ (.B1(_03746_),
    .Y(_00601_),
    .A1(net69),
    .A2(_03744_));
 sg13g2_and2_1 _09327_ (.A(_02294_),
    .B(_03712_),
    .X(_03747_));
 sg13g2_buf_1 _09328_ (.A(_03747_),
    .X(_03748_));
 sg13g2_xnor2_1 _09329_ (.Y(_03749_),
    .A(_02292_),
    .B(_03748_));
 sg13g2_xnor2_1 _09330_ (.Y(_03750_),
    .A(_02292_),
    .B(_00917_));
 sg13g2_a21o_1 _09331_ (.A2(_03738_),
    .A1(net252),
    .B1(_01088_),
    .X(_03751_));
 sg13g2_o21ai_1 _09332_ (.B1(_03751_),
    .Y(_03752_),
    .A1(net252),
    .A2(_03738_));
 sg13g2_xnor2_1 _09333_ (.Y(_03753_),
    .A(_03750_),
    .B(_03752_));
 sg13g2_mux2_1 _09334_ (.A0(_03749_),
    .A1(_03753_),
    .S(_03715_),
    .X(_03754_));
 sg13g2_nor2_1 _09335_ (.A(net61),
    .B(_03754_),
    .Y(_03755_));
 sg13g2_a21oi_1 _09336_ (.A1(\addr[14] ),
    .A2(net62),
    .Y(_03756_),
    .B1(_03755_));
 sg13g2_mux2_1 _09337_ (.A0(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .S(_03638_),
    .X(_03757_));
 sg13g2_nand2_1 _09338_ (.Y(_03758_),
    .A(net68),
    .B(_03757_));
 sg13g2_o21ai_1 _09339_ (.B1(_03758_),
    .Y(_00602_),
    .A1(net69),
    .A2(_03756_));
 sg13g2_and2_1 _09340_ (.A(_02310_),
    .B(_03704_),
    .X(_03759_));
 sg13g2_buf_1 _09341_ (.A(_03759_),
    .X(_03760_));
 sg13g2_nand2_1 _09342_ (.Y(_03761_),
    .A(_00769_),
    .B(_01088_));
 sg13g2_nor4_1 _09343_ (.A(_03730_),
    .B(_03731_),
    .C(_03737_),
    .D(_03761_),
    .Y(_03762_));
 sg13g2_nand2_1 _09344_ (.Y(_03763_),
    .A(_00769_),
    .B(net252));
 sg13g2_nor4_1 _09345_ (.A(_03730_),
    .B(_03731_),
    .C(_03737_),
    .D(_03763_),
    .Y(_03764_));
 sg13g2_nand2_1 _09346_ (.Y(_03765_),
    .A(_00917_),
    .B(_01088_));
 sg13g2_nor4_1 _09347_ (.A(_03730_),
    .B(_03731_),
    .C(_03737_),
    .D(_03765_),
    .Y(_03766_));
 sg13g2_nand2_1 _09348_ (.Y(_03767_),
    .A(_00917_),
    .B(net252));
 sg13g2_nor4_1 _09349_ (.A(_03730_),
    .B(_03731_),
    .C(_03737_),
    .D(_03767_),
    .Y(_03768_));
 sg13g2_nor4_2 _09350_ (.A(_03762_),
    .B(_03764_),
    .C(_03766_),
    .Y(_03769_),
    .D(_03768_));
 sg13g2_nand2_1 _09351_ (.Y(_03770_),
    .A(net254),
    .B(_00917_));
 sg13g2_and2_1 _09352_ (.A(_02308_),
    .B(_01088_),
    .X(_03771_));
 sg13g2_o21ai_1 _09353_ (.B1(_03771_),
    .Y(_03772_),
    .A1(net254),
    .A2(_00917_));
 sg13g2_and2_1 _09354_ (.A(_03770_),
    .B(_03772_),
    .X(_03773_));
 sg13g2_buf_1 _09355_ (.A(_03773_),
    .X(_03774_));
 sg13g2_nand2_1 _09356_ (.Y(_03775_),
    .A(_03769_),
    .B(_03774_));
 sg13g2_xor2_1 _09357_ (.B(_03775_),
    .A(_00959_),
    .X(_03776_));
 sg13g2_mux2_1 _09358_ (.A0(_03760_),
    .A1(_03776_),
    .S(net280),
    .X(_03777_));
 sg13g2_xnor2_1 _09359_ (.Y(_03778_),
    .A(_02306_),
    .B(_03777_));
 sg13g2_nor2_1 _09360_ (.A(_03641_),
    .B(_03778_),
    .Y(_03779_));
 sg13g2_a21oi_1 _09361_ (.A1(\addr[15] ),
    .A2(_03626_),
    .Y(_03780_),
    .B1(_03779_));
 sg13g2_buf_1 _09362_ (.A(_03637_),
    .X(_03781_));
 sg13g2_mux2_1 _09363_ (.A0(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .S(net155),
    .X(_03782_));
 sg13g2_nand2_1 _09364_ (.Y(_03783_),
    .A(net68),
    .B(_03782_));
 sg13g2_o21ai_1 _09365_ (.B1(_03783_),
    .Y(_00603_),
    .A1(net69),
    .A2(_03780_));
 sg13g2_nor2_1 _09366_ (.A(_00959_),
    .B(_03775_),
    .Y(_03784_));
 sg13g2_a21oi_1 _09367_ (.A1(_00959_),
    .A2(_03775_),
    .Y(_03785_),
    .B1(net253));
 sg13g2_nor2_1 _09368_ (.A(_03784_),
    .B(_03785_),
    .Y(_03786_));
 sg13g2_xnor2_1 _09369_ (.Y(_03787_),
    .A(net305),
    .B(_01045_));
 sg13g2_xnor2_1 _09370_ (.Y(_03788_),
    .A(_03786_),
    .B(_03787_));
 sg13g2_nand3_1 _09371_ (.B(net254),
    .C(_03748_),
    .A(net253),
    .Y(_03789_));
 sg13g2_xor2_1 _09372_ (.B(_03789_),
    .A(_01137_),
    .X(_03790_));
 sg13g2_nor2_1 _09373_ (.A(_03674_),
    .B(_03790_),
    .Y(_03791_));
 sg13g2_a21oi_1 _09374_ (.A1(net240),
    .A2(_03788_),
    .Y(_03792_),
    .B1(_03791_));
 sg13g2_nor2_1 _09375_ (.A(_03641_),
    .B(_03792_),
    .Y(_03793_));
 sg13g2_a21oi_1 _09376_ (.A1(\addr[16] ),
    .A2(net62),
    .Y(_03794_),
    .B1(_03793_));
 sg13g2_mux2_1 _09377_ (.A0(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .S(net155),
    .X(_03795_));
 sg13g2_nand2_1 _09378_ (.Y(_03796_),
    .A(_03724_),
    .B(_03795_));
 sg13g2_o21ai_1 _09379_ (.B1(_03796_),
    .Y(_00604_),
    .A1(_03640_),
    .A2(_03794_));
 sg13g2_nand2_1 _09380_ (.Y(_03797_),
    .A(_02299_),
    .B(_03760_));
 sg13g2_xnor2_1 _09381_ (.Y(_03798_),
    .A(_00989_),
    .B(_03797_));
 sg13g2_xnor2_1 _09382_ (.Y(_03799_),
    .A(net308),
    .B(_01092_));
 sg13g2_nand2_1 _09383_ (.Y(_03800_),
    .A(_00959_),
    .B(net305));
 sg13g2_a22oi_1 _09384_ (.Y(_03801_),
    .B1(_03800_),
    .B2(_02635_),
    .A2(_03774_),
    .A1(_03769_));
 sg13g2_nand2_1 _09385_ (.Y(_03802_),
    .A(_00959_),
    .B(_01045_));
 sg13g2_nand2_1 _09386_ (.Y(_03803_),
    .A(net253),
    .B(_01045_));
 sg13g2_a22oi_1 _09387_ (.Y(_03804_),
    .B1(_03802_),
    .B2(_03803_),
    .A2(_03774_),
    .A1(_03769_));
 sg13g2_nand2_1 _09388_ (.Y(_03805_),
    .A(net305),
    .B(_01045_));
 sg13g2_and2_1 _09389_ (.A(net253),
    .B(_00959_),
    .X(_03806_));
 sg13g2_o21ai_1 _09390_ (.B1(_03806_),
    .Y(_03807_),
    .A1(net305),
    .A2(_01045_));
 sg13g2_nand2_1 _09391_ (.Y(_03808_),
    .A(_03805_),
    .B(_03807_));
 sg13g2_nor3_2 _09392_ (.A(_03801_),
    .B(_03804_),
    .C(_03808_),
    .Y(_03809_));
 sg13g2_xnor2_1 _09393_ (.Y(_03810_),
    .A(_03799_),
    .B(_03809_));
 sg13g2_nand2_1 _09394_ (.Y(_03811_),
    .A(net236),
    .B(_03810_));
 sg13g2_o21ai_1 _09395_ (.B1(_03811_),
    .Y(_03812_),
    .A1(_03711_),
    .A2(_03798_));
 sg13g2_nor2_1 _09396_ (.A(net61),
    .B(_03812_),
    .Y(_03813_));
 sg13g2_a21oi_1 _09397_ (.A1(\addr[17] ),
    .A2(_03626_),
    .Y(_03814_),
    .B1(_03813_));
 sg13g2_mux2_1 _09398_ (.A0(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .S(net155),
    .X(_03815_));
 sg13g2_nand2_1 _09399_ (.Y(_03816_),
    .A(net68),
    .B(_03815_));
 sg13g2_o21ai_1 _09400_ (.B1(_03816_),
    .Y(_00605_),
    .A1(_03640_),
    .A2(_03814_));
 sg13g2_buf_1 _09401_ (.A(net71),
    .X(_03817_));
 sg13g2_buf_1 _09402_ (.A(net71),
    .X(_03818_));
 sg13g2_nand4_1 _09403_ (.B(_00989_),
    .C(_02299_),
    .A(net254),
    .Y(_03819_),
    .D(_03748_));
 sg13g2_xnor2_1 _09404_ (.Y(_03820_),
    .A(_02297_),
    .B(_03819_));
 sg13g2_nand2_1 _09405_ (.Y(_03821_),
    .A(net308),
    .B(_01092_));
 sg13g2_nor2_1 _09406_ (.A(net308),
    .B(_01092_),
    .Y(_03822_));
 sg13g2_a21oi_2 _09407_ (.B1(_03822_),
    .Y(_03823_),
    .A2(_03821_),
    .A1(_03809_));
 sg13g2_xor2_1 _09408_ (.B(_00921_),
    .A(net286),
    .X(_03824_));
 sg13g2_xnor2_1 _09409_ (.Y(_03825_),
    .A(_03823_),
    .B(_03824_));
 sg13g2_nand2_1 _09410_ (.Y(_03826_),
    .A(net236),
    .B(_03825_));
 sg13g2_o21ai_1 _09411_ (.B1(_03826_),
    .Y(_03827_),
    .A1(net237),
    .A2(_03820_));
 sg13g2_nor2_1 _09412_ (.A(net59),
    .B(_03827_),
    .Y(_03828_));
 sg13g2_a21oi_1 _09413_ (.A1(\addr[18] ),
    .A2(_03817_),
    .Y(_03829_),
    .B1(_03828_));
 sg13g2_mux2_1 _09414_ (.A0(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .S(_03781_),
    .X(_03830_));
 sg13g2_nand2_1 _09415_ (.Y(_03831_),
    .A(_03724_),
    .B(_03830_));
 sg13g2_o21ai_1 _09416_ (.B1(_03831_),
    .Y(_00606_),
    .A1(net69),
    .A2(_03829_));
 sg13g2_buf_1 _09417_ (.A(_03629_),
    .X(_03832_));
 sg13g2_xor2_1 _09418_ (.B(_00965_),
    .A(_00859_),
    .X(_03833_));
 sg13g2_a21o_1 _09419_ (.A2(_03823_),
    .A1(net286),
    .B1(_00921_),
    .X(_03834_));
 sg13g2_o21ai_1 _09420_ (.B1(_03834_),
    .Y(_03835_),
    .A1(net286),
    .A2(_03823_));
 sg13g2_xnor2_1 _09421_ (.Y(_03836_),
    .A(_03833_),
    .B(_03835_));
 sg13g2_nand2_1 _09422_ (.Y(_03837_),
    .A(_02301_),
    .B(_03760_));
 sg13g2_xor2_1 _09423_ (.B(_03837_),
    .A(_00859_),
    .X(_03838_));
 sg13g2_nor2_1 _09424_ (.A(net239),
    .B(_03838_),
    .Y(_03839_));
 sg13g2_a21oi_1 _09425_ (.A1(net240),
    .A2(_03836_),
    .Y(_03840_),
    .B1(_03839_));
 sg13g2_nor2_1 _09426_ (.A(net59),
    .B(_03840_),
    .Y(_03841_));
 sg13g2_a21oi_1 _09427_ (.A1(\addr[19] ),
    .A2(net60),
    .Y(_03842_),
    .B1(_03841_));
 sg13g2_mux2_1 _09428_ (.A0(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .S(_03781_),
    .X(_03843_));
 sg13g2_nand2_1 _09429_ (.Y(_03844_),
    .A(net68),
    .B(_03843_));
 sg13g2_o21ai_1 _09430_ (.B1(_03844_),
    .Y(_00607_),
    .A1(net67),
    .A2(_03842_));
 sg13g2_xnor2_1 _09431_ (.Y(_03845_),
    .A(net309),
    .B(_01090_));
 sg13g2_nand2_1 _09432_ (.Y(_03846_),
    .A(net236),
    .B(_03845_));
 sg13g2_o21ai_1 _09433_ (.B1(_03846_),
    .Y(_03847_),
    .A1(_01396_),
    .A2(net237));
 sg13g2_nor2_1 _09434_ (.A(net59),
    .B(_03847_),
    .Y(_03848_));
 sg13g2_a21oi_1 _09435_ (.A1(\addr[1] ),
    .A2(net60),
    .Y(_03849_),
    .B1(_03848_));
 sg13g2_nand3_1 _09436_ (.B(net70),
    .C(net156),
    .A(\i_tinyqv.mem.q_ctrl.addr[1] ),
    .Y(_03850_));
 sg13g2_o21ai_1 _09437_ (.B1(_03850_),
    .Y(_00608_),
    .A1(net67),
    .A2(_03849_));
 sg13g2_and2_1 _09438_ (.A(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .B(_03686_),
    .X(_03851_));
 sg13g2_a21oi_1 _09439_ (.A1(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .A2(net156),
    .Y(_03852_),
    .B1(_03851_));
 sg13g2_a21oi_1 _09440_ (.A1(\addr[20] ),
    .A2(net62),
    .Y(_03853_),
    .B1(net70));
 sg13g2_nand2b_1 _09441_ (.Y(_03854_),
    .B(_00097_),
    .A_N(_03623_));
 sg13g2_buf_1 _09442_ (.A(_03854_),
    .X(_03855_));
 sg13g2_nand2_1 _09443_ (.Y(_03856_),
    .A(_00859_),
    .B(_00965_));
 sg13g2_and2_1 _09444_ (.A(_03821_),
    .B(_03856_),
    .X(_03857_));
 sg13g2_nand2b_1 _09445_ (.Y(_03858_),
    .B(_03857_),
    .A_N(_00921_));
 sg13g2_nor4_1 _09446_ (.A(_03801_),
    .B(_03804_),
    .C(_03808_),
    .D(_03858_),
    .Y(_03859_));
 sg13g2_nand2b_1 _09447_ (.Y(_03860_),
    .B(_03857_),
    .A_N(net286));
 sg13g2_nor4_1 _09448_ (.A(_03801_),
    .B(_03804_),
    .C(_03808_),
    .D(_03860_),
    .Y(_03861_));
 sg13g2_nor2_1 _09449_ (.A(net286),
    .B(_00921_),
    .Y(_03862_));
 sg13g2_nand2_1 _09450_ (.Y(_03863_),
    .A(_03822_),
    .B(_03856_));
 sg13g2_a21oi_1 _09451_ (.A1(net286),
    .A2(_00921_),
    .Y(_03864_),
    .B1(_03863_));
 sg13g2_a21o_1 _09452_ (.A2(_03862_),
    .A1(_03856_),
    .B1(_03864_),
    .X(_03865_));
 sg13g2_nor2_1 _09453_ (.A(_00859_),
    .B(_00965_),
    .Y(_03866_));
 sg13g2_nor4_2 _09454_ (.A(_03859_),
    .B(_03861_),
    .C(_03865_),
    .Y(_03867_),
    .D(_03866_));
 sg13g2_xnor2_1 _09455_ (.Y(_03868_),
    .A(_01046_),
    .B(_03867_));
 sg13g2_nor2b_1 _09456_ (.A(_03868_),
    .B_N(net280),
    .Y(_03869_));
 sg13g2_nor3_1 _09457_ (.A(net280),
    .B(_02303_),
    .C(_03675_),
    .Y(_03870_));
 sg13g2_nor2_1 _09458_ (.A(_03869_),
    .B(_03870_),
    .Y(_03871_));
 sg13g2_xnor2_1 _09459_ (.Y(_03872_),
    .A(_01138_),
    .B(_03871_));
 sg13g2_nand2_1 _09460_ (.Y(_03873_),
    .A(_03855_),
    .B(_03872_));
 sg13g2_a22oi_1 _09461_ (.Y(_00609_),
    .B1(_03853_),
    .B2(_03873_),
    .A2(_03852_),
    .A1(net69));
 sg13g2_xor2_1 _09462_ (.B(_01093_),
    .A(net307),
    .X(_03874_));
 sg13g2_a21oi_1 _09463_ (.A1(_01138_),
    .A2(_03867_),
    .Y(_03875_),
    .B1(_01046_));
 sg13g2_nor2_1 _09464_ (.A(_01138_),
    .B(_03867_),
    .Y(_03876_));
 sg13g2_nor2_1 _09465_ (.A(_03875_),
    .B(_03876_),
    .Y(_03877_));
 sg13g2_xnor2_1 _09466_ (.Y(_03878_),
    .A(_03874_),
    .B(_03877_));
 sg13g2_or2_1 _09467_ (.X(_03879_),
    .B(_03675_),
    .A(_02284_));
 sg13g2_nor2_1 _09468_ (.A(_02632_),
    .B(_03879_),
    .Y(_03880_));
 sg13g2_xor2_1 _09469_ (.B(_03880_),
    .A(net307),
    .X(_03881_));
 sg13g2_o21ai_1 _09470_ (.B1(_03855_),
    .Y(_03882_),
    .A1(net236),
    .A2(_03881_));
 sg13g2_a21oi_1 _09471_ (.A1(net240),
    .A2(_03878_),
    .Y(_03883_),
    .B1(_03882_));
 sg13g2_a21oi_1 _09472_ (.A1(\addr[21] ),
    .A2(_03817_),
    .Y(_03884_),
    .B1(_03883_));
 sg13g2_mux2_1 _09473_ (.A0(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .S(_03686_),
    .X(_03885_));
 sg13g2_nand2_1 _09474_ (.Y(_03886_),
    .A(net68),
    .B(_03885_));
 sg13g2_o21ai_1 _09475_ (.B1(_03886_),
    .Y(_00610_),
    .A1(net67),
    .A2(_03884_));
 sg13g2_and2_1 _09476_ (.A(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .B(_03686_),
    .X(_03887_));
 sg13g2_a21oi_1 _09477_ (.A1(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .A2(net156),
    .Y(_03888_),
    .B1(_03887_));
 sg13g2_and2_1 _09478_ (.A(net307),
    .B(_01093_),
    .X(_03889_));
 sg13g2_or2_1 _09479_ (.X(_03890_),
    .B(_01093_),
    .A(net307));
 sg13g2_o21ai_1 _09480_ (.B1(_03890_),
    .Y(_03891_),
    .A1(_03877_),
    .A2(_03889_));
 sg13g2_buf_2 _09481_ (.A(_03891_),
    .X(_03892_));
 sg13g2_xnor2_1 _09482_ (.Y(_03893_),
    .A(_03304_),
    .B(_03892_));
 sg13g2_nand3_1 _09483_ (.B(_02296_),
    .C(_02631_),
    .A(net307),
    .Y(_03894_));
 sg13g2_nor2_1 _09484_ (.A(_03894_),
    .B(_03677_),
    .Y(_03895_));
 sg13g2_nor2_1 _09485_ (.A(net280),
    .B(_03895_),
    .Y(_03896_));
 sg13g2_a21oi_1 _09486_ (.A1(net280),
    .A2(_03893_),
    .Y(_03897_),
    .B1(_03896_));
 sg13g2_xnor2_1 _09487_ (.Y(_03898_),
    .A(_00760_),
    .B(_03897_));
 sg13g2_o21ai_1 _09488_ (.B1(_03621_),
    .Y(_03899_),
    .A1(\addr[22] ),
    .A2(_03855_));
 sg13g2_a21o_1 _09489_ (.A2(_03898_),
    .A1(_03855_),
    .B1(_03899_),
    .X(_03900_));
 sg13g2_o21ai_1 _09490_ (.B1(_03900_),
    .Y(_00611_),
    .A1(_03621_),
    .A2(_03888_));
 sg13g2_and2_1 _09491_ (.A(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .B(_03686_),
    .X(_03901_));
 sg13g2_a21oi_1 _09492_ (.A1(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .A2(net156),
    .Y(_03902_),
    .B1(_03901_));
 sg13g2_buf_1 _09493_ (.A(_00159_),
    .X(_03903_));
 sg13g2_nor2b_1 _09494_ (.A(_02759_),
    .B_N(_03760_),
    .Y(_03904_));
 sg13g2_xnor2_1 _09495_ (.Y(_03905_),
    .A(_00160_),
    .B(_03904_));
 sg13g2_nor3_1 _09496_ (.A(net237),
    .B(_03625_),
    .C(_03905_),
    .Y(_03906_));
 sg13g2_a21oi_1 _09497_ (.A1(_03903_),
    .A2(net71),
    .Y(_03907_),
    .B1(_03906_));
 sg13g2_xnor2_1 _09498_ (.Y(_03908_),
    .A(\i_tinyqv.cpu.instr_data_start[23] ),
    .B(\i_tinyqv.cpu.imm[23] ));
 sg13g2_a21oi_1 _09499_ (.A1(_03304_),
    .A2(_03892_),
    .Y(_03909_),
    .B1(_02719_));
 sg13g2_nor2_1 _09500_ (.A(_03304_),
    .B(_03892_),
    .Y(_03910_));
 sg13g2_nor2_1 _09501_ (.A(_03909_),
    .B(_03910_),
    .Y(_03911_));
 sg13g2_xnor2_1 _09502_ (.Y(_03912_),
    .A(_03908_),
    .B(_03911_));
 sg13g2_nand3_1 _09503_ (.B(_03855_),
    .C(_03912_),
    .A(_03643_),
    .Y(_03913_));
 sg13g2_nand3_1 _09504_ (.B(_03907_),
    .C(_03913_),
    .A(_03621_),
    .Y(_03914_));
 sg13g2_o21ai_1 _09505_ (.B1(_03914_),
    .Y(_00612_),
    .A1(_03621_),
    .A2(_03902_));
 sg13g2_nand2_1 _09506_ (.Y(_03915_),
    .A(net309),
    .B(_01090_));
 sg13g2_xor2_1 _09507_ (.B(_00919_),
    .A(_00758_),
    .X(_03916_));
 sg13g2_xnor2_1 _09508_ (.Y(_03917_),
    .A(_03915_),
    .B(_03916_));
 sg13g2_nor2b_1 _09509_ (.A(net239),
    .B_N(_01406_),
    .Y(_03918_));
 sg13g2_a21oi_1 _09510_ (.A1(_03643_),
    .A2(_03917_),
    .Y(_03919_),
    .B1(_03918_));
 sg13g2_nor2_1 _09511_ (.A(net59),
    .B(_03919_),
    .Y(_03920_));
 sg13g2_a21oi_1 _09512_ (.A1(_01578_),
    .A2(net60),
    .Y(_03921_),
    .B1(_03920_));
 sg13g2_nand3_1 _09513_ (.B(net70),
    .C(net156),
    .A(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .Y(_03922_));
 sg13g2_o21ai_1 _09514_ (.B1(_03922_),
    .Y(_00613_),
    .A1(net67),
    .A2(_03921_));
 sg13g2_xor2_1 _09515_ (.B(_01399_),
    .A(_00857_),
    .X(_03923_));
 sg13g2_xnor2_1 _09516_ (.Y(_03924_),
    .A(net312),
    .B(_00955_));
 sg13g2_xnor2_1 _09517_ (.Y(_03925_),
    .A(_03647_),
    .B(_03924_));
 sg13g2_nand2_1 _09518_ (.Y(_03926_),
    .A(net236),
    .B(_03925_));
 sg13g2_o21ai_1 _09519_ (.B1(_03926_),
    .Y(_03927_),
    .A1(net237),
    .A2(_03923_));
 sg13g2_nor2_1 _09520_ (.A(net59),
    .B(_03927_),
    .Y(_03928_));
 sg13g2_a21oi_1 _09521_ (.A1(net295),
    .A2(net60),
    .Y(_03929_),
    .B1(_03928_));
 sg13g2_nand3_1 _09522_ (.B(_03630_),
    .C(net156),
    .A(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .Y(_03930_));
 sg13g2_o21ai_1 _09523_ (.B1(_03930_),
    .Y(_00614_),
    .A1(net67),
    .A2(_03929_));
 sg13g2_xnor2_1 _09524_ (.Y(_03931_),
    .A(_01146_),
    .B(_03675_));
 sg13g2_nor2_1 _09525_ (.A(_02338_),
    .B(_03647_),
    .Y(_03932_));
 sg13g2_nand2_1 _09526_ (.Y(_03933_),
    .A(_02338_),
    .B(_03647_));
 sg13g2_o21ai_1 _09527_ (.B1(_03933_),
    .Y(_03934_),
    .A1(net312),
    .A2(_03932_));
 sg13g2_xnor2_1 _09528_ (.Y(_03935_),
    .A(net303),
    .B(_01041_));
 sg13g2_xnor2_1 _09529_ (.Y(_03936_),
    .A(_03934_),
    .B(_03935_));
 sg13g2_nand2_1 _09530_ (.Y(_03937_),
    .A(net239),
    .B(_03936_));
 sg13g2_o21ai_1 _09531_ (.B1(_03937_),
    .Y(_03938_),
    .A1(net237),
    .A2(_03931_));
 sg13g2_nor2_1 _09532_ (.A(net59),
    .B(_03938_),
    .Y(_03939_));
 sg13g2_a21oi_1 _09533_ (.A1(_01575_),
    .A2(net60),
    .Y(_03940_),
    .B1(_03939_));
 sg13g2_mux2_1 _09534_ (.A0(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[4] ),
    .S(net155),
    .X(_03941_));
 sg13g2_nand2_1 _09535_ (.Y(_03942_),
    .A(net70),
    .B(_03941_));
 sg13g2_o21ai_1 _09536_ (.B1(_03942_),
    .Y(_00615_),
    .A1(net67),
    .A2(_03940_));
 sg13g2_xnor2_1 _09537_ (.Y(_03943_),
    .A(_03654_),
    .B(_03702_));
 sg13g2_xor2_1 _09538_ (.B(_01091_),
    .A(net256),
    .X(_03944_));
 sg13g2_xnor2_1 _09539_ (.Y(_03945_),
    .A(_03653_),
    .B(_03944_));
 sg13g2_nand2_1 _09540_ (.Y(_03946_),
    .A(net239),
    .B(_03945_));
 sg13g2_o21ai_1 _09541_ (.B1(_03946_),
    .Y(_03947_),
    .A1(net237),
    .A2(_03943_));
 sg13g2_nor2_1 _09542_ (.A(net59),
    .B(_03947_),
    .Y(_03948_));
 sg13g2_a21oi_1 _09543_ (.A1(_01576_),
    .A2(net60),
    .Y(_03949_),
    .B1(_03948_));
 sg13g2_mux2_1 _09544_ (.A0(\i_tinyqv.mem.q_ctrl.addr[1] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .S(net155),
    .X(_03950_));
 sg13g2_nand2_1 _09545_ (.Y(_03951_),
    .A(net70),
    .B(_03950_));
 sg13g2_o21ai_1 _09546_ (.B1(_03951_),
    .Y(_00616_),
    .A1(net67),
    .A2(_03949_));
 sg13g2_a21o_1 _09547_ (.A2(_03653_),
    .A1(net256),
    .B1(_01091_),
    .X(_03952_));
 sg13g2_o21ai_1 _09548_ (.B1(_03952_),
    .Y(_03953_),
    .A1(_02290_),
    .A2(_03653_));
 sg13g2_xor2_1 _09549_ (.B(_00920_),
    .A(net258),
    .X(_03954_));
 sg13g2_xnor2_1 _09550_ (.Y(_03955_),
    .A(_03953_),
    .B(_03954_));
 sg13g2_xor2_1 _09551_ (.B(_03677_),
    .A(_02266_),
    .X(_03956_));
 sg13g2_nor2_1 _09552_ (.A(net239),
    .B(_03956_),
    .Y(_03957_));
 sg13g2_a21oi_1 _09553_ (.A1(net240),
    .A2(_03955_),
    .Y(_03958_),
    .B1(_03957_));
 sg13g2_nor2_1 _09554_ (.A(net59),
    .B(_03958_),
    .Y(_03959_));
 sg13g2_a21oi_1 _09555_ (.A1(\addr[6] ),
    .A2(net60),
    .Y(_03960_),
    .B1(_03959_));
 sg13g2_mux2_1 _09556_ (.A0(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[6] ),
    .S(net155),
    .X(_03961_));
 sg13g2_nand2_1 _09557_ (.Y(_03962_),
    .A(net70),
    .B(_03961_));
 sg13g2_o21ai_1 _09558_ (.B1(_03962_),
    .Y(_00617_),
    .A1(net67),
    .A2(_03960_));
 sg13g2_nand3_1 _09559_ (.B(_02290_),
    .C(_03702_),
    .A(_02266_),
    .Y(_03963_));
 sg13g2_xnor2_1 _09560_ (.Y(_03964_),
    .A(_02291_),
    .B(_03963_));
 sg13g2_xnor2_1 _09561_ (.Y(_03965_),
    .A(net255),
    .B(_00956_));
 sg13g2_xnor2_1 _09562_ (.Y(_03966_),
    .A(_03661_),
    .B(_03965_));
 sg13g2_nand2_1 _09563_ (.Y(_03967_),
    .A(net239),
    .B(_03966_));
 sg13g2_o21ai_1 _09564_ (.B1(_03967_),
    .Y(_03968_),
    .A1(net236),
    .A2(_03964_));
 sg13g2_nor2_1 _09565_ (.A(_03818_),
    .B(_03968_),
    .Y(_03969_));
 sg13g2_a21oi_1 _09566_ (.A1(\addr[7] ),
    .A2(net60),
    .Y(_03970_),
    .B1(_03969_));
 sg13g2_mux2_1 _09567_ (.A0(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[7] ),
    .S(net155),
    .X(_03971_));
 sg13g2_nand2_1 _09568_ (.Y(_03972_),
    .A(net70),
    .B(_03971_));
 sg13g2_o21ai_1 _09569_ (.B1(_03972_),
    .Y(_00618_),
    .A1(_03832_),
    .A2(_03970_));
 sg13g2_nand2_1 _09570_ (.Y(_03973_),
    .A(_03395_),
    .B(_03661_));
 sg13g2_nor2_1 _09571_ (.A(_03395_),
    .B(_03661_),
    .Y(_03974_));
 sg13g2_a21oi_1 _09572_ (.A1(net255),
    .A2(_03973_),
    .Y(_03975_),
    .B1(_03974_));
 sg13g2_xor2_1 _09573_ (.B(_01042_),
    .A(net304),
    .X(_03976_));
 sg13g2_xnor2_1 _09574_ (.Y(_03977_),
    .A(_03975_),
    .B(_03976_));
 sg13g2_xnor2_1 _09575_ (.Y(_03978_),
    .A(_01142_),
    .B(_03712_));
 sg13g2_nor2_1 _09576_ (.A(_03642_),
    .B(_03978_),
    .Y(_03979_));
 sg13g2_a21oi_1 _09577_ (.A1(net237),
    .A2(_03977_),
    .Y(_03980_),
    .B1(_03979_));
 sg13g2_nor2_1 _09578_ (.A(_03818_),
    .B(_03980_),
    .Y(_03981_));
 sg13g2_a21oi_1 _09579_ (.A1(\addr[8] ),
    .A2(net61),
    .Y(_03982_),
    .B1(_03981_));
 sg13g2_a22oi_1 _09580_ (.Y(_03983_),
    .B1(_03687_),
    .B2(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .A2(_03686_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[4] ));
 sg13g2_o21ai_1 _09581_ (.B1(_03983_),
    .Y(_00619_),
    .A1(_03832_),
    .A2(_03982_));
 sg13g2_nor2_1 _09582_ (.A(_02622_),
    .B(_03879_),
    .Y(_03984_));
 sg13g2_xor2_1 _09583_ (.B(_03984_),
    .A(net287),
    .X(_03985_));
 sg13g2_a21oi_1 _09584_ (.A1(_03661_),
    .A2(_03669_),
    .Y(_03986_),
    .B1(_03665_));
 sg13g2_xor2_1 _09585_ (.B(_01191_),
    .A(net287),
    .X(_03987_));
 sg13g2_xnor2_1 _09586_ (.Y(_03988_),
    .A(_03986_),
    .B(_03987_));
 sg13g2_nand2_1 _09587_ (.Y(_03989_),
    .A(net239),
    .B(_03988_));
 sg13g2_o21ai_1 _09588_ (.B1(_03989_),
    .Y(_03990_),
    .A1(net236),
    .A2(_03985_));
 sg13g2_nor2_1 _09589_ (.A(_03625_),
    .B(_03990_),
    .Y(_03991_));
 sg13g2_a21oi_1 _09590_ (.A1(\addr[9] ),
    .A2(net61),
    .Y(_03992_),
    .B1(_03991_));
 sg13g2_mux2_1 _09591_ (.A0(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .S(net155),
    .X(_03993_));
 sg13g2_nand2_1 _09592_ (.Y(_03994_),
    .A(_03630_),
    .B(_03993_));
 sg13g2_o21ai_1 _09593_ (.B1(_03994_),
    .Y(_00620_),
    .A1(net68),
    .A2(_03992_));
 sg13g2_buf_1 _09594_ (.A(\i_tinyqv.mem.q_ctrl.is_writing ),
    .X(_03995_));
 sg13g2_inv_1 _09595_ (.Y(_03996_),
    .A(_03995_));
 sg13g2_buf_2 _09596_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .X(_03997_));
 sg13g2_buf_1 _09597_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ),
    .X(_03998_));
 sg13g2_buf_1 _09598_ (.A(net281),
    .X(_03999_));
 sg13g2_buf_2 _09599_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .X(_04000_));
 sg13g2_nor2b_1 _09600_ (.A(net235),
    .B_N(_04000_),
    .Y(_04001_));
 sg13g2_buf_1 _09601_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .X(_04002_));
 sg13g2_nand2_1 _09602_ (.Y(_04003_),
    .A(_01517_),
    .B(net279));
 sg13g2_nor4_1 _09603_ (.A(_03997_),
    .B(_03998_),
    .C(_04001_),
    .D(_04003_),
    .Y(_04004_));
 sg13g2_nand2_1 _09604_ (.Y(_04005_),
    .A(net279),
    .B(net200));
 sg13g2_buf_2 _09605_ (.A(_04005_),
    .X(_04006_));
 sg13g2_buf_2 _09606_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .X(_04007_));
 sg13g2_buf_1 _09607_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .X(_04008_));
 sg13g2_nor3_2 _09608_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .B(_04007_),
    .C(_04008_),
    .Y(_04009_));
 sg13g2_nor2_2 _09609_ (.A(net281),
    .B(_04003_),
    .Y(_04010_));
 sg13g2_o21ai_1 _09610_ (.B1(_03631_),
    .Y(_04011_),
    .A1(_04009_),
    .A2(_04010_));
 sg13g2_a21oi_1 _09611_ (.A1(_04006_),
    .A2(_04011_),
    .Y(_04012_),
    .B1(_03996_));
 sg13g2_a21oi_1 _09612_ (.A1(_03996_),
    .A2(_04004_),
    .Y(_04013_),
    .B1(_04012_));
 sg13g2_buf_1 _09613_ (.A(_04013_),
    .X(_04014_));
 sg13g2_buf_1 _09614_ (.A(_04014_),
    .X(_04015_));
 sg13g2_buf_1 _09615_ (.A(_03995_),
    .X(_04016_));
 sg13g2_xnor2_1 _09616_ (.Y(_04017_),
    .A(_01424_),
    .B(_01240_));
 sg13g2_buf_4 _09617_ (.X(_04018_),
    .A(_04017_));
 sg13g2_buf_1 _09618_ (.A(_01230_),
    .X(_04019_));
 sg13g2_nand2_1 _09619_ (.Y(_04020_),
    .A(_01424_),
    .B(_01240_));
 sg13g2_xor2_1 _09620_ (.B(_04020_),
    .A(net233),
    .X(_04021_));
 sg13g2_buf_4 _09621_ (.X(_04022_),
    .A(_04021_));
 sg13g2_mux4_1 _09622_ (.S0(_04018_),
    .A0(\data_to_write[24] ),
    .A1(\data_to_write[16] ),
    .A2(\data_to_write[8] ),
    .A3(_01573_),
    .S1(_04022_),
    .X(_04023_));
 sg13g2_nor2_1 _09623_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .B(_04007_),
    .Y(_04024_));
 sg13g2_nand2b_1 _09624_ (.Y(_04025_),
    .B(_04024_),
    .A_N(_04008_));
 sg13g2_buf_2 _09625_ (.A(_04025_),
    .X(_04026_));
 sg13g2_nand2_2 _09626_ (.Y(_04027_),
    .A(_04006_),
    .B(_04026_));
 sg13g2_mux2_1 _09627_ (.A0(net8),
    .A1(_04023_),
    .S(_04027_),
    .X(_04028_));
 sg13g2_nor3_1 _09628_ (.A(_03997_),
    .B(_04000_),
    .C(_03998_),
    .Y(_04029_));
 sg13g2_and2_1 _09629_ (.A(_04010_),
    .B(_04029_),
    .X(_04030_));
 sg13g2_buf_2 _09630_ (.A(_04030_),
    .X(_04031_));
 sg13g2_nor2b_1 _09631_ (.A(net8),
    .B_N(_04031_),
    .Y(_04032_));
 sg13g2_nor2_1 _09632_ (.A(_03997_),
    .B(_03998_),
    .Y(_04033_));
 sg13g2_and2_1 _09633_ (.A(_01517_),
    .B(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .X(_04034_));
 sg13g2_buf_2 _09634_ (.A(_04034_),
    .X(_04035_));
 sg13g2_nand4_1 _09635_ (.B(_04000_),
    .C(_04033_),
    .A(_03632_),
    .Y(_04036_),
    .D(_04035_));
 sg13g2_buf_1 _09636_ (.A(_04036_),
    .X(_04037_));
 sg13g2_mux2_1 _09637_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .S(_04037_),
    .X(_04038_));
 sg13g2_nor2_1 _09638_ (.A(_04031_),
    .B(_04038_),
    .Y(_04039_));
 sg13g2_nor3_1 _09639_ (.A(net234),
    .B(_04032_),
    .C(_04039_),
    .Y(_04040_));
 sg13g2_a21oi_1 _09640_ (.A1(net234),
    .A2(_04028_),
    .Y(_04041_),
    .B1(_04040_));
 sg13g2_nand2_1 _09641_ (.Y(_04042_),
    .A(_02226_),
    .B(net112));
 sg13g2_o21ai_1 _09642_ (.B1(_04042_),
    .Y(_00621_),
    .A1(_04015_),
    .A2(_04041_));
 sg13g2_mux4_1 _09643_ (.S0(_04018_),
    .A0(\data_to_write[25] ),
    .A1(\data_to_write[17] ),
    .A2(\data_to_write[9] ),
    .A3(_01600_),
    .S1(_04022_),
    .X(_04043_));
 sg13g2_mux2_1 _09644_ (.A0(net9),
    .A1(_04043_),
    .S(_04027_),
    .X(_04044_));
 sg13g2_nor2b_1 _09645_ (.A(net9),
    .B_N(_04031_),
    .Y(_04045_));
 sg13g2_mux2_1 _09646_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .S(_04037_),
    .X(_04046_));
 sg13g2_nor2_1 _09647_ (.A(_04031_),
    .B(_04046_),
    .Y(_04047_));
 sg13g2_nor3_1 _09648_ (.A(net234),
    .B(_04045_),
    .C(_04047_),
    .Y(_04048_));
 sg13g2_a21oi_1 _09649_ (.A1(net234),
    .A2(_04044_),
    .Y(_04049_),
    .B1(_04048_));
 sg13g2_nand2_1 _09650_ (.Y(_04050_),
    .A(_02582_),
    .B(net112));
 sg13g2_o21ai_1 _09651_ (.B1(_04050_),
    .Y(_00622_),
    .A1(_04015_),
    .A2(_04049_));
 sg13g2_mux4_1 _09652_ (.S0(_04018_),
    .A0(\data_to_write[26] ),
    .A1(\data_to_write[18] ),
    .A2(\data_to_write[10] ),
    .A3(_01603_),
    .S1(_04022_),
    .X(_04051_));
 sg13g2_mux2_1 _09653_ (.A0(net10),
    .A1(_04051_),
    .S(_04027_),
    .X(_04052_));
 sg13g2_nor2b_1 _09654_ (.A(net10),
    .B_N(_04031_),
    .Y(_04053_));
 sg13g2_mux2_1 _09655_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .S(_04037_),
    .X(_04054_));
 sg13g2_nor2_1 _09656_ (.A(_04031_),
    .B(_04054_),
    .Y(_04055_));
 sg13g2_nor3_1 _09657_ (.A(_04016_),
    .B(_04053_),
    .C(_04055_),
    .Y(_04056_));
 sg13g2_a21oi_1 _09658_ (.A1(net234),
    .A2(_04052_),
    .Y(_04057_),
    .B1(_04056_));
 sg13g2_nand2_1 _09659_ (.Y(_04058_),
    .A(_02675_),
    .B(_04014_));
 sg13g2_o21ai_1 _09660_ (.B1(_04058_),
    .Y(_00623_),
    .A1(net112),
    .A2(_04057_));
 sg13g2_mux4_1 _09661_ (.S0(_04018_),
    .A0(\data_to_write[27] ),
    .A1(\data_to_write[19] ),
    .A2(\data_to_write[11] ),
    .A3(_01606_),
    .S1(_04022_),
    .X(_04059_));
 sg13g2_mux2_1 _09662_ (.A0(net11),
    .A1(_04059_),
    .S(_04027_),
    .X(_04060_));
 sg13g2_nor2b_1 _09663_ (.A(net11),
    .B_N(_04031_),
    .Y(_04061_));
 sg13g2_mux2_1 _09664_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .S(_04037_),
    .X(_04062_));
 sg13g2_nor2_1 _09665_ (.A(_04031_),
    .B(_04062_),
    .Y(_04063_));
 sg13g2_nor3_1 _09666_ (.A(_04016_),
    .B(_04061_),
    .C(_04063_),
    .Y(_04064_));
 sg13g2_a21oi_1 _09667_ (.A1(net234),
    .A2(_04060_),
    .Y(_04065_),
    .B1(_04064_));
 sg13g2_nand2_1 _09668_ (.Y(_04066_),
    .A(_02790_),
    .B(_04014_));
 sg13g2_o21ai_1 _09669_ (.B1(_04066_),
    .Y(_00624_),
    .A1(net112),
    .A2(_04065_));
 sg13g2_mux4_1 _09670_ (.S0(_04018_),
    .A0(\data_to_write[28] ),
    .A1(\data_to_write[20] ),
    .A2(\data_to_write[12] ),
    .A3(_01609_),
    .S1(_04022_),
    .X(_04067_));
 sg13g2_a21oi_1 _09671_ (.A1(_04006_),
    .A2(_04026_),
    .Y(_04068_),
    .B1(_03996_));
 sg13g2_buf_2 _09672_ (.A(_04068_),
    .X(_04069_));
 sg13g2_nor2b_1 _09673_ (.A(_04069_),
    .B_N(_02226_),
    .Y(_04070_));
 sg13g2_a21oi_1 _09674_ (.A1(_04067_),
    .A2(_04069_),
    .Y(_04071_),
    .B1(_04070_));
 sg13g2_nand2_1 _09675_ (.Y(_04072_),
    .A(\i_tinyqv.cpu.instr_data_in[12] ),
    .B(_04014_));
 sg13g2_o21ai_1 _09676_ (.B1(_04072_),
    .Y(_00625_),
    .A1(net112),
    .A2(_04071_));
 sg13g2_mux4_1 _09677_ (.S0(_04018_),
    .A0(\data_to_write[29] ),
    .A1(\data_to_write[21] ),
    .A2(\data_to_write[13] ),
    .A3(_01612_),
    .S1(_04022_),
    .X(_04073_));
 sg13g2_nor2b_1 _09678_ (.A(_04069_),
    .B_N(_02582_),
    .Y(_04074_));
 sg13g2_a21oi_1 _09679_ (.A1(_04069_),
    .A2(_04073_),
    .Y(_04075_),
    .B1(_04074_));
 sg13g2_nand2_1 _09680_ (.Y(_04076_),
    .A(\i_tinyqv.cpu.instr_data_in[13] ),
    .B(_04014_));
 sg13g2_o21ai_1 _09681_ (.B1(_04076_),
    .Y(_00626_),
    .A1(net112),
    .A2(_04075_));
 sg13g2_mux4_1 _09682_ (.S0(_04018_),
    .A0(\data_to_write[30] ),
    .A1(\data_to_write[22] ),
    .A2(\data_to_write[14] ),
    .A3(_01616_),
    .S1(_04022_),
    .X(_04077_));
 sg13g2_nor2b_1 _09683_ (.A(_04069_),
    .B_N(_02675_),
    .Y(_04078_));
 sg13g2_a21oi_1 _09684_ (.A1(_04069_),
    .A2(_04077_),
    .Y(_04079_),
    .B1(_04078_));
 sg13g2_nand2_1 _09685_ (.Y(_04080_),
    .A(_02676_),
    .B(_04014_));
 sg13g2_o21ai_1 _09686_ (.B1(_04080_),
    .Y(_00627_),
    .A1(net112),
    .A2(_04079_));
 sg13g2_mux4_1 _09687_ (.S0(_04018_),
    .A0(\data_to_write[31] ),
    .A1(\data_to_write[23] ),
    .A2(\data_to_write[15] ),
    .A3(\data_to_write[7] ),
    .S1(_04022_),
    .X(_04081_));
 sg13g2_nor2b_1 _09688_ (.A(_04069_),
    .B_N(_02790_),
    .Y(_04082_));
 sg13g2_a21oi_1 _09689_ (.A1(_04069_),
    .A2(_04081_),
    .Y(_04083_),
    .B1(_04082_));
 sg13g2_nand2_1 _09690_ (.Y(_04084_),
    .A(_02780_),
    .B(_04014_));
 sg13g2_o21ai_1 _09691_ (.B1(_04084_),
    .Y(_00628_),
    .A1(net112),
    .A2(_04083_));
 sg13g2_buf_1 _09692_ (.A(_01517_),
    .X(_04085_));
 sg13g2_nor2_1 _09693_ (.A(net281),
    .B(_01519_),
    .Y(_04086_));
 sg13g2_nand2b_1 _09694_ (.Y(_04087_),
    .B(_04086_),
    .A_N(net232));
 sg13g2_buf_1 _09695_ (.A(_04087_),
    .X(_04088_));
 sg13g2_o21ai_1 _09696_ (.B1(_01514_),
    .Y(_04089_),
    .A1(_01501_),
    .A2(_01502_));
 sg13g2_and2_1 _09697_ (.A(_04089_),
    .B(_01526_),
    .X(_04090_));
 sg13g2_buf_1 _09698_ (.A(_04090_),
    .X(_04091_));
 sg13g2_nand2b_1 _09699_ (.Y(_04092_),
    .B(_03995_),
    .A_N(_03631_));
 sg13g2_or2_1 _09700_ (.X(_04093_),
    .B(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .A(_02861_));
 sg13g2_a21oi_1 _09701_ (.A1(_04091_),
    .A2(_04092_),
    .Y(_04094_),
    .B1(_04093_));
 sg13g2_buf_2 _09702_ (.A(_04094_),
    .X(_04095_));
 sg13g2_nand2_1 _09703_ (.Y(_04096_),
    .A(_04088_),
    .B(_04095_));
 sg13g2_buf_2 _09704_ (.A(_04096_),
    .X(_04097_));
 sg13g2_o21ai_1 _09705_ (.B1(_04035_),
    .Y(_04098_),
    .A1(_03632_),
    .A2(_00162_));
 sg13g2_nor4_1 _09706_ (.A(_03997_),
    .B(_04000_),
    .C(_03998_),
    .D(_04098_),
    .Y(_04099_));
 sg13g2_a21o_1 _09707_ (.A2(_04098_),
    .A1(_03631_),
    .B1(_04099_),
    .X(_04100_));
 sg13g2_buf_1 _09708_ (.A(_04100_),
    .X(_04101_));
 sg13g2_buf_1 _09709_ (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ),
    .X(_04102_));
 sg13g2_nand3_1 _09710_ (.B(_04102_),
    .C(_04035_),
    .A(net281),
    .Y(_04103_));
 sg13g2_buf_1 _09711_ (.A(_04103_),
    .X(_04104_));
 sg13g2_nand2_1 _09712_ (.Y(_04105_),
    .A(_04026_),
    .B(_04104_));
 sg13g2_nand3_1 _09713_ (.B(_04101_),
    .C(_04105_),
    .A(net279),
    .Y(_04106_));
 sg13g2_nor2_2 _09714_ (.A(\i_tinyqv.mem.data_stall ),
    .B(_01446_),
    .Y(_04107_));
 sg13g2_nand2_1 _09715_ (.Y(_04108_),
    .A(_04085_),
    .B(_04107_));
 sg13g2_nand2b_1 _09716_ (.Y(_04109_),
    .B(_04108_),
    .A_N(_04106_));
 sg13g2_nor2_1 _09717_ (.A(_00165_),
    .B(_04029_),
    .Y(_04110_));
 sg13g2_nand2_1 _09718_ (.Y(_04111_),
    .A(_04109_),
    .B(_04110_));
 sg13g2_a21oi_2 _09719_ (.B1(_04099_),
    .Y(_04112_),
    .A2(_04098_),
    .A1(_03631_));
 sg13g2_nor3_1 _09720_ (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .B(_04026_),
    .C(_04112_),
    .Y(_04113_));
 sg13g2_buf_1 _09721_ (.A(net279),
    .X(_04114_));
 sg13g2_nor2b_1 _09722_ (.A(net232),
    .B_N(_04114_),
    .Y(_04115_));
 sg13g2_o21ai_1 _09723_ (.B1(_04115_),
    .Y(_04116_),
    .A1(_03999_),
    .A2(_04113_));
 sg13g2_nor2_1 _09724_ (.A(_04000_),
    .B(_03998_),
    .Y(_04117_));
 sg13g2_nand2_1 _09725_ (.Y(_04118_),
    .A(_04117_),
    .B(_04107_));
 sg13g2_a21oi_1 _09726_ (.A1(_03996_),
    .A2(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .Y(_04119_),
    .B1(_04118_));
 sg13g2_a21oi_1 _09727_ (.A1(_04110_),
    .A2(_04118_),
    .Y(_04120_),
    .B1(_04119_));
 sg13g2_and2_1 _09728_ (.A(net279),
    .B(net200),
    .X(_04121_));
 sg13g2_buf_1 _09729_ (.A(_04121_),
    .X(_04122_));
 sg13g2_a22oi_1 _09730_ (.Y(_04123_),
    .B1(_04120_),
    .B2(_04122_),
    .A2(_04116_),
    .A1(_04111_));
 sg13g2_nand2_1 _09731_ (.Y(_04124_),
    .A(_03997_),
    .B(_04097_));
 sg13g2_o21ai_1 _09732_ (.B1(_04124_),
    .Y(_00643_),
    .A1(_04097_),
    .A2(_04123_));
 sg13g2_nor2_1 _09733_ (.A(net200),
    .B(_04109_),
    .Y(_04125_));
 sg13g2_nor3_1 _09734_ (.A(_03995_),
    .B(_04006_),
    .C(_04118_),
    .Y(_04126_));
 sg13g2_nor2_1 _09735_ (.A(_03997_),
    .B(_04000_),
    .Y(_04127_));
 sg13g2_nand2_1 _09736_ (.Y(_04128_),
    .A(_03998_),
    .B(_04127_));
 sg13g2_nand2_1 _09737_ (.Y(_04129_),
    .A(_03997_),
    .B(_04000_));
 sg13g2_a21oi_1 _09738_ (.A1(_04128_),
    .A2(_04129_),
    .Y(_04130_),
    .B1(_04125_));
 sg13g2_a221oi_1 _09739_ (.B2(_04102_),
    .C1(_04130_),
    .B1(_04126_),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .Y(_04131_),
    .A2(_04125_));
 sg13g2_nand2_1 _09740_ (.Y(_04132_),
    .A(_04000_),
    .B(_04097_));
 sg13g2_o21ai_1 _09741_ (.B1(_04132_),
    .Y(_00644_),
    .A1(_04097_),
    .A2(_04131_));
 sg13g2_nand2_1 _09742_ (.Y(_04133_),
    .A(_04102_),
    .B(_04125_));
 sg13g2_nor2_1 _09743_ (.A(_04125_),
    .B(_04127_),
    .Y(_04134_));
 sg13g2_o21ai_1 _09744_ (.B1(_03998_),
    .Y(_04135_),
    .A1(_04097_),
    .A2(_04134_));
 sg13g2_o21ai_1 _09745_ (.B1(_04135_),
    .Y(_00645_),
    .A1(_04097_),
    .A2(_04133_));
 sg13g2_inv_1 _09746_ (.Y(_04136_),
    .A(_00162_));
 sg13g2_inv_1 _09747_ (.Y(_04137_),
    .A(_00165_));
 sg13g2_nor4_1 _09748_ (.A(_04136_),
    .B(_04137_),
    .C(_04006_),
    .D(_04117_),
    .Y(_04138_));
 sg13g2_buf_4 _09749_ (.X(_04139_),
    .A(_04138_));
 sg13g2_mux2_1 _09750_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .A1(net8),
    .S(_04139_),
    .X(_00649_));
 sg13g2_mux2_1 _09751_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .A1(net9),
    .S(_04139_),
    .X(_00650_));
 sg13g2_mux2_1 _09752_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .A1(net10),
    .S(_04139_),
    .X(_00651_));
 sg13g2_mux2_1 _09753_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .A1(net11),
    .S(_04139_),
    .X(_00652_));
 sg13g2_mux2_1 _09754_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .S(_04139_),
    .X(_00653_));
 sg13g2_mux2_1 _09755_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .S(_04139_),
    .X(_00654_));
 sg13g2_mux2_1 _09756_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .S(_04139_),
    .X(_00655_));
 sg13g2_mux2_1 _09757_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .S(_04139_),
    .X(_00656_));
 sg13g2_buf_1 _09758_ (.A(_01424_),
    .X(_04140_));
 sg13g2_nor2_1 _09759_ (.A(net233),
    .B(net230),
    .Y(_04141_));
 sg13g2_nand2_1 _09760_ (.Y(_04142_),
    .A(net297),
    .B(_04141_));
 sg13g2_buf_4 _09761_ (.X(_04143_),
    .A(_04142_));
 sg13g2_mux2_1 _09762_ (.A0(_02226_),
    .A1(\i_tinyqv.cpu.instr_data_in[0] ),
    .S(_04143_),
    .X(_00660_));
 sg13g2_nor2b_1 _09763_ (.A(net230),
    .B_N(net233),
    .Y(_04144_));
 sg13g2_buf_1 _09764_ (.A(_01231_),
    .X(_04145_));
 sg13g2_nor2b_1 _09765_ (.A(_04145_),
    .B_N(net297),
    .Y(_04146_));
 sg13g2_o21ai_1 _09766_ (.B1(_04146_),
    .Y(_04147_),
    .A1(_01426_),
    .A2(_04144_));
 sg13g2_buf_2 _09767_ (.A(_04147_),
    .X(_04148_));
 sg13g2_nand2_1 _09768_ (.Y(_04149_),
    .A(\i_tinyqv.mem.qspi_data_buf[10] ),
    .B(_01512_));
 sg13g2_o21ai_1 _09769_ (.B1(_04149_),
    .Y(_00661_),
    .A1(_03424_),
    .A2(_04148_));
 sg13g2_nand2_1 _09770_ (.Y(_04150_),
    .A(\i_tinyqv.mem.qspi_data_buf[11] ),
    .B(net190));
 sg13g2_o21ai_1 _09771_ (.B1(_04150_),
    .Y(_00662_),
    .A1(_03427_),
    .A2(_04148_));
 sg13g2_nand2_1 _09772_ (.Y(_04151_),
    .A(\i_tinyqv.mem.qspi_data_buf[12] ),
    .B(net190));
 sg13g2_o21ai_1 _09773_ (.B1(_04151_),
    .Y(_00663_),
    .A1(_03429_),
    .A2(_04148_));
 sg13g2_nand2_1 _09774_ (.Y(_04152_),
    .A(\i_tinyqv.mem.qspi_data_buf[13] ),
    .B(net190));
 sg13g2_o21ai_1 _09775_ (.B1(_04152_),
    .Y(_00664_),
    .A1(_03431_),
    .A2(_04148_));
 sg13g2_nand2_1 _09776_ (.Y(_04153_),
    .A(\i_tinyqv.mem.qspi_data_buf[14] ),
    .B(net190));
 sg13g2_o21ai_1 _09777_ (.B1(_04153_),
    .Y(_00665_),
    .A1(_03433_),
    .A2(_04148_));
 sg13g2_nand2_1 _09778_ (.Y(_04154_),
    .A(\i_tinyqv.mem.qspi_data_buf[15] ),
    .B(net190));
 sg13g2_o21ai_1 _09779_ (.B1(_04154_),
    .Y(_00666_),
    .A1(_03435_),
    .A2(_04148_));
 sg13g2_nand3b_1 _09780_ (.B(net233),
    .C(net297),
    .Y(_04155_),
    .A_N(net230));
 sg13g2_buf_2 _09781_ (.A(_04155_),
    .X(_04156_));
 sg13g2_buf_1 _09782_ (.A(_04156_),
    .X(_04157_));
 sg13g2_nand2_1 _09783_ (.Y(_04158_),
    .A(\i_tinyqv.mem.data_from_read[16] ),
    .B(net182));
 sg13g2_o21ai_1 _09784_ (.B1(_04158_),
    .Y(_00667_),
    .A1(_03438_),
    .A2(net182));
 sg13g2_nand2_1 _09785_ (.Y(_04159_),
    .A(\i_tinyqv.mem.data_from_read[17] ),
    .B(_04157_));
 sg13g2_o21ai_1 _09786_ (.B1(_04159_),
    .Y(_00668_),
    .A1(_03440_),
    .A2(_04157_));
 sg13g2_nand2_1 _09787_ (.Y(_04160_),
    .A(\i_tinyqv.mem.data_from_read[18] ),
    .B(_04156_));
 sg13g2_o21ai_1 _09788_ (.B1(_04160_),
    .Y(_00669_),
    .A1(_03424_),
    .A2(net182));
 sg13g2_nand2_1 _09789_ (.Y(_04161_),
    .A(\i_tinyqv.mem.data_from_read[19] ),
    .B(_04156_));
 sg13g2_o21ai_1 _09790_ (.B1(_04161_),
    .Y(_00670_),
    .A1(_03427_),
    .A2(net182));
 sg13g2_mux2_1 _09791_ (.A0(_02582_),
    .A1(\i_tinyqv.cpu.instr_data_in[1] ),
    .S(_04143_),
    .X(_00671_));
 sg13g2_nand2_1 _09792_ (.Y(_04162_),
    .A(\i_tinyqv.mem.data_from_read[20] ),
    .B(_04156_));
 sg13g2_o21ai_1 _09793_ (.B1(_04162_),
    .Y(_00672_),
    .A1(_03429_),
    .A2(net182));
 sg13g2_nand2_1 _09794_ (.Y(_04163_),
    .A(\i_tinyqv.mem.data_from_read[21] ),
    .B(_04156_));
 sg13g2_o21ai_1 _09795_ (.B1(_04163_),
    .Y(_00673_),
    .A1(_03431_),
    .A2(net182));
 sg13g2_nand2_1 _09796_ (.Y(_04164_),
    .A(\i_tinyqv.mem.data_from_read[22] ),
    .B(_04156_));
 sg13g2_o21ai_1 _09797_ (.B1(_04164_),
    .Y(_00674_),
    .A1(_03433_),
    .A2(net182));
 sg13g2_nand2_1 _09798_ (.Y(_04165_),
    .A(\i_tinyqv.mem.data_from_read[23] ),
    .B(_04156_));
 sg13g2_o21ai_1 _09799_ (.B1(_04165_),
    .Y(_00675_),
    .A1(_03435_),
    .A2(net182));
 sg13g2_nand3_1 _09800_ (.B(net233),
    .C(net230),
    .A(net297),
    .Y(_04166_));
 sg13g2_buf_1 _09801_ (.A(_04166_),
    .X(_04167_));
 sg13g2_buf_1 _09802_ (.A(_04167_),
    .X(_04168_));
 sg13g2_nor3_1 _09803_ (.A(net229),
    .B(_03438_),
    .C(net181),
    .Y(_04169_));
 sg13g2_a21o_1 _09804_ (.A2(net181),
    .A1(\i_tinyqv.mem.qspi_data_buf[24] ),
    .B1(_04169_),
    .X(_00676_));
 sg13g2_nor3_1 _09805_ (.A(net229),
    .B(_03440_),
    .C(net181),
    .Y(_04170_));
 sg13g2_a21o_1 _09806_ (.A2(net181),
    .A1(\i_tinyqv.mem.qspi_data_buf[25] ),
    .B1(_04170_),
    .X(_00677_));
 sg13g2_nor3_1 _09807_ (.A(net229),
    .B(_03424_),
    .C(_04167_),
    .Y(_04171_));
 sg13g2_a21o_1 _09808_ (.A2(net181),
    .A1(\i_tinyqv.mem.qspi_data_buf[26] ),
    .B1(_04171_),
    .X(_00678_));
 sg13g2_nor3_1 _09809_ (.A(net229),
    .B(_03427_),
    .C(_04167_),
    .Y(_04172_));
 sg13g2_a21o_1 _09810_ (.A2(net181),
    .A1(\i_tinyqv.mem.qspi_data_buf[27] ),
    .B1(_04172_),
    .X(_00679_));
 sg13g2_nor3_1 _09811_ (.A(net229),
    .B(_03429_),
    .C(_04167_),
    .Y(_04173_));
 sg13g2_a21o_1 _09812_ (.A2(net181),
    .A1(\i_tinyqv.mem.qspi_data_buf[28] ),
    .B1(_04173_),
    .X(_00680_));
 sg13g2_nor3_1 _09813_ (.A(net229),
    .B(_03431_),
    .C(_04167_),
    .Y(_04174_));
 sg13g2_a21o_1 _09814_ (.A2(_04168_),
    .A1(\i_tinyqv.mem.qspi_data_buf[29] ),
    .B1(_04174_),
    .X(_00681_));
 sg13g2_mux2_1 _09815_ (.A0(_02675_),
    .A1(_02681_),
    .S(_04143_),
    .X(_00682_));
 sg13g2_nor3_1 _09816_ (.A(net229),
    .B(_03433_),
    .C(_04167_),
    .Y(_04175_));
 sg13g2_a21o_1 _09817_ (.A2(_04168_),
    .A1(\i_tinyqv.mem.qspi_data_buf[30] ),
    .B1(_04175_),
    .X(_00683_));
 sg13g2_nor3_1 _09818_ (.A(net229),
    .B(_03435_),
    .C(_04167_),
    .Y(_04176_));
 sg13g2_a21o_1 _09819_ (.A2(net181),
    .A1(\i_tinyqv.mem.qspi_data_buf[31] ),
    .B1(_04176_),
    .X(_00684_));
 sg13g2_mux2_1 _09820_ (.A0(_02790_),
    .A1(_02791_),
    .S(_04143_),
    .X(_00685_));
 sg13g2_mux2_1 _09821_ (.A0(\i_tinyqv.cpu.instr_data_in[12] ),
    .A1(_02235_),
    .S(_04143_),
    .X(_00686_));
 sg13g2_mux2_1 _09822_ (.A0(\i_tinyqv.cpu.instr_data_in[13] ),
    .A1(_02591_),
    .S(_04143_),
    .X(_00687_));
 sg13g2_mux2_1 _09823_ (.A0(_02676_),
    .A1(_02682_),
    .S(_04143_),
    .X(_00688_));
 sg13g2_mux2_1 _09824_ (.A0(_02780_),
    .A1(_02781_),
    .S(_04143_),
    .X(_00689_));
 sg13g2_nand2_1 _09825_ (.Y(_04177_),
    .A(\i_tinyqv.mem.qspi_data_buf[8] ),
    .B(net190));
 sg13g2_o21ai_1 _09826_ (.B1(_04177_),
    .Y(_00690_),
    .A1(_03438_),
    .A2(_04148_));
 sg13g2_nand2_1 _09827_ (.Y(_04178_),
    .A(\i_tinyqv.mem.qspi_data_buf[9] ),
    .B(net190));
 sg13g2_o21ai_1 _09828_ (.B1(_04178_),
    .Y(_00691_),
    .A1(_03440_),
    .A2(_04148_));
 sg13g2_buf_1 _09829_ (.A(\i_uart_rx.cycle_counter[5] ),
    .X(_04179_));
 sg13g2_buf_1 _09830_ (.A(\i_uart_rx.cycle_counter[1] ),
    .X(_04180_));
 sg13g2_buf_1 _09831_ (.A(\i_uart_rx.cycle_counter[0] ),
    .X(_04181_));
 sg13g2_and3_1 _09832_ (.X(_04182_),
    .A(_04180_),
    .B(_04181_),
    .C(\i_uart_rx.cycle_counter[3] ));
 sg13g2_buf_1 _09833_ (.A(_04182_),
    .X(_04183_));
 sg13g2_buf_1 _09834_ (.A(\i_uart_rx.cycle_counter[7] ),
    .X(_04184_));
 sg13g2_buf_1 _09835_ (.A(\i_uart_rx.cycle_counter[6] ),
    .X(_04185_));
 sg13g2_nor3_1 _09836_ (.A(_04184_),
    .B(_04185_),
    .C(\i_uart_rx.cycle_counter[10] ),
    .Y(_04186_));
 sg13g2_buf_2 _09837_ (.A(\i_uart_rx.cycle_counter[2] ),
    .X(_04187_));
 sg13g2_buf_1 _09838_ (.A(\i_uart_rx.cycle_counter[4] ),
    .X(_04188_));
 sg13g2_inv_1 _09839_ (.Y(_04189_),
    .A(\i_uart_rx.cycle_counter[9] ));
 sg13g2_nor4_1 _09840_ (.A(_04187_),
    .B(_04188_),
    .C(_04189_),
    .D(\i_uart_rx.cycle_counter[8] ),
    .Y(_04190_));
 sg13g2_and4_1 _09841_ (.A(_04179_),
    .B(_04183_),
    .C(_04186_),
    .D(_04190_),
    .X(_04191_));
 sg13g2_buf_1 _09842_ (.A(_04191_),
    .X(_04192_));
 sg13g2_buf_1 _09843_ (.A(\i_uart_rx.fsm_state[3] ),
    .X(_04193_));
 sg13g2_nor2_1 _09844_ (.A(_01377_),
    .B(net299),
    .Y(_04194_));
 sg13g2_xnor2_1 _09845_ (.Y(_04195_),
    .A(net278),
    .B(_04194_));
 sg13g2_nand2_1 _09846_ (.Y(_04196_),
    .A(_04192_),
    .B(_04195_));
 sg13g2_buf_4 _09847_ (.X(_04197_),
    .A(_04196_));
 sg13g2_mux2_1 _09848_ (.A0(\i_uart_rx.recieved_data[1] ),
    .A1(\i_uart_rx.recieved_data[0] ),
    .S(_04197_),
    .X(_00710_));
 sg13g2_mux2_1 _09849_ (.A0(\i_uart_rx.recieved_data[2] ),
    .A1(\i_uart_rx.recieved_data[1] ),
    .S(_04197_),
    .X(_00711_));
 sg13g2_mux2_1 _09850_ (.A0(\i_uart_rx.recieved_data[3] ),
    .A1(\i_uart_rx.recieved_data[2] ),
    .S(_04197_),
    .X(_00712_));
 sg13g2_mux2_1 _09851_ (.A0(\i_uart_rx.recieved_data[4] ),
    .A1(\i_uart_rx.recieved_data[3] ),
    .S(_04197_),
    .X(_00713_));
 sg13g2_mux2_1 _09852_ (.A0(\i_uart_rx.recieved_data[5] ),
    .A1(\i_uart_rx.recieved_data[4] ),
    .S(_04197_),
    .X(_00714_));
 sg13g2_mux2_1 _09853_ (.A0(\i_uart_rx.recieved_data[6] ),
    .A1(\i_uart_rx.recieved_data[5] ),
    .S(_04197_),
    .X(_00715_));
 sg13g2_mux2_1 _09854_ (.A0(\i_uart_rx.recieved_data[7] ),
    .A1(\i_uart_rx.recieved_data[6] ),
    .S(_04197_),
    .X(_00716_));
 sg13g2_mux2_1 _09855_ (.A0(\i_uart_rx.bit_sample ),
    .A1(\i_uart_rx.recieved_data[7] ),
    .S(_04197_),
    .X(_00717_));
 sg13g2_nand2_1 _09856_ (.Y(_04198_),
    .A(_02232_),
    .B(_02264_));
 sg13g2_buf_1 _09857_ (.A(_04198_),
    .X(_04199_));
 sg13g2_buf_1 _09858_ (.A(_04199_),
    .X(_04200_));
 sg13g2_mux2_1 _09859_ (.A0(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[4] ),
    .S(net146),
    .X(_00366_));
 sg13g2_mux2_1 _09860_ (.A0(\i_tinyqv.cpu.i_core.mepc[10] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[14] ),
    .S(net146),
    .X(_00367_));
 sg13g2_mux2_1 _09861_ (.A0(\i_tinyqv.cpu.i_core.mepc[11] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[15] ),
    .S(net146),
    .X(_00368_));
 sg13g2_mux2_1 _09862_ (.A0(\i_tinyqv.cpu.i_core.mepc[12] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[16] ),
    .S(net146),
    .X(_00369_));
 sg13g2_mux2_1 _09863_ (.A0(\i_tinyqv.cpu.i_core.mepc[13] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[17] ),
    .S(net146),
    .X(_00370_));
 sg13g2_mux2_1 _09864_ (.A0(\i_tinyqv.cpu.i_core.mepc[14] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[18] ),
    .S(_04200_),
    .X(_00371_));
 sg13g2_mux2_1 _09865_ (.A0(\i_tinyqv.cpu.i_core.mepc[15] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[19] ),
    .S(net146),
    .X(_00372_));
 sg13g2_mux2_1 _09866_ (.A0(\i_tinyqv.cpu.i_core.mepc[16] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[20] ),
    .S(_04200_),
    .X(_00373_));
 sg13g2_mux2_1 _09867_ (.A0(\i_tinyqv.cpu.i_core.mepc[17] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[21] ),
    .S(net146),
    .X(_00374_));
 sg13g2_mux2_1 _09868_ (.A0(\i_tinyqv.cpu.i_core.mepc[18] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[22] ),
    .S(net146),
    .X(_00375_));
 sg13g2_buf_1 _09869_ (.A(_04199_),
    .X(_04201_));
 sg13g2_mux2_1 _09870_ (.A0(\i_tinyqv.cpu.i_core.mepc[19] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[23] ),
    .S(net145),
    .X(_00376_));
 sg13g2_mux2_1 _09871_ (.A0(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[5] ),
    .S(net145),
    .X(_00377_));
 sg13g2_and2_1 _09872_ (.A(_01185_),
    .B(_01194_),
    .X(_04202_));
 sg13g2_buf_1 _09873_ (.A(_04202_),
    .X(_04203_));
 sg13g2_nand2_1 _09874_ (.Y(_04204_),
    .A(net218),
    .B(\i_tinyqv.cpu.is_system ));
 sg13g2_nor2_2 _09875_ (.A(_01179_),
    .B(_04204_),
    .Y(_04205_));
 sg13g2_nor2b_1 _09876_ (.A(_02355_),
    .B_N(_04205_),
    .Y(_04206_));
 sg13g2_buf_1 _09877_ (.A(_04206_),
    .X(_04207_));
 sg13g2_mux2_1 _09878_ (.A0(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A1(net133),
    .S(_04207_),
    .X(_04208_));
 sg13g2_nor2_1 _09879_ (.A(_01148_),
    .B(_04203_),
    .Y(_04209_));
 sg13g2_a21oi_1 _09880_ (.A1(_04203_),
    .A2(_04208_),
    .Y(_04210_),
    .B1(_04209_));
 sg13g2_nand2_1 _09881_ (.Y(_04211_),
    .A(_01282_),
    .B(_04199_));
 sg13g2_nand2_1 _09882_ (.Y(_04212_),
    .A(\i_tinyqv.cpu.i_core.mepc[20] ),
    .B(_02354_));
 sg13g2_o21ai_1 _09883_ (.B1(_04212_),
    .Y(_00378_),
    .A1(_04210_),
    .A2(_04211_));
 sg13g2_mux2_1 _09884_ (.A0(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A1(net151),
    .S(_04207_),
    .X(_04213_));
 sg13g2_nand2_1 _09885_ (.Y(_04214_),
    .A(_00994_),
    .B(net137));
 sg13g2_o21ai_1 _09886_ (.B1(_04214_),
    .Y(_04215_),
    .A1(net137),
    .A2(_04213_));
 sg13g2_nand2_1 _09887_ (.Y(_04216_),
    .A(\i_tinyqv.cpu.i_core.mepc[21] ),
    .B(_02354_));
 sg13g2_o21ai_1 _09888_ (.B1(_04216_),
    .Y(_00379_),
    .A1(_04211_),
    .A2(_04215_));
 sg13g2_mux2_1 _09889_ (.A0(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A1(_01696_),
    .S(_04207_),
    .X(_04217_));
 sg13g2_nand2_1 _09890_ (.Y(_04218_),
    .A(_00773_),
    .B(net137));
 sg13g2_o21ai_1 _09891_ (.B1(_04218_),
    .Y(_04219_),
    .A1(net137),
    .A2(_04217_));
 sg13g2_nand2_1 _09892_ (.Y(_04220_),
    .A(\i_tinyqv.cpu.i_core.mepc[22] ),
    .B(_02354_));
 sg13g2_o21ai_1 _09893_ (.B1(_04220_),
    .Y(_00380_),
    .A1(_04211_),
    .A2(_04219_));
 sg13g2_inv_1 _09894_ (.Y(_04221_),
    .A(net154));
 sg13g2_mux2_1 _09895_ (.A0(\i_tinyqv.cpu.i_core.mepc[3] ),
    .A1(_04221_),
    .S(_04207_),
    .X(_04222_));
 sg13g2_nand2_1 _09896_ (.Y(_04223_),
    .A(_00863_),
    .B(_01221_));
 sg13g2_o21ai_1 _09897_ (.B1(_04223_),
    .Y(_04224_),
    .A1(_01221_),
    .A2(_04222_));
 sg13g2_nand2_1 _09898_ (.Y(_04225_),
    .A(\i_tinyqv.cpu.i_core.mepc[23] ),
    .B(_02354_));
 sg13g2_o21ai_1 _09899_ (.B1(_04225_),
    .Y(_00381_),
    .A1(_04211_),
    .A2(_04224_));
 sg13g2_mux2_1 _09900_ (.A0(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[6] ),
    .S(net145),
    .X(_00382_));
 sg13g2_mux2_1 _09901_ (.A0(\i_tinyqv.cpu.i_core.mepc[3] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[7] ),
    .S(net145),
    .X(_00383_));
 sg13g2_mux2_1 _09902_ (.A0(\i_tinyqv.cpu.i_core.mepc[4] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[8] ),
    .S(net145),
    .X(_00384_));
 sg13g2_mux2_1 _09903_ (.A0(\i_tinyqv.cpu.i_core.mepc[5] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[9] ),
    .S(net145),
    .X(_00385_));
 sg13g2_mux2_1 _09904_ (.A0(\i_tinyqv.cpu.i_core.mepc[6] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[10] ),
    .S(net145),
    .X(_00386_));
 sg13g2_mux2_1 _09905_ (.A0(\i_tinyqv.cpu.i_core.mepc[7] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[11] ),
    .S(net145),
    .X(_00387_));
 sg13g2_mux2_1 _09906_ (.A0(\i_tinyqv.cpu.i_core.mepc[8] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[12] ),
    .S(_04201_),
    .X(_00388_));
 sg13g2_mux2_1 _09907_ (.A0(\i_tinyqv.cpu.i_core.mepc[9] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[13] ),
    .S(_04201_),
    .X(_00389_));
 sg13g2_a21oi_1 _09908_ (.A1(_01179_),
    .A2(net184),
    .Y(_04226_),
    .B1(_02379_));
 sg13g2_buf_1 _09909_ (.A(_04226_),
    .X(_04227_));
 sg13g2_buf_1 _09910_ (.A(_04227_),
    .X(_04228_));
 sg13g2_mux2_1 _09911_ (.A0(_01765_),
    .A1(net259),
    .S(net144),
    .X(_00405_));
 sg13g2_mux2_1 _09912_ (.A0(net242),
    .A1(_01983_),
    .S(_04228_),
    .X(_00406_));
 sg13g2_buf_1 _09913_ (.A(_04227_),
    .X(_04229_));
 sg13g2_nand2_1 _09914_ (.Y(_04230_),
    .A(net293),
    .B(_04229_));
 sg13g2_o21ai_1 _09915_ (.B1(_04230_),
    .Y(_00407_),
    .A1(_03020_),
    .A2(_04228_));
 sg13g2_buf_1 _09916_ (.A(_04227_),
    .X(_04231_));
 sg13g2_mux2_1 _09917_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .A1(_02045_),
    .S(net142),
    .X(_00408_));
 sg13g2_mux2_1 _09918_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .A1(_02085_),
    .S(net142),
    .X(_00409_));
 sg13g2_mux2_1 _09919_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .A1(_03018_),
    .S(net142),
    .X(_00410_));
 sg13g2_mux2_1 _09920_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A1(_02162_),
    .S(net142),
    .X(_00411_));
 sg13g2_mux2_1 _09921_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(_04231_),
    .X(_00412_));
 sg13g2_mux2_1 _09922_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(_04231_),
    .X(_00413_));
 sg13g2_mux2_1 _09923_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .S(net142),
    .X(_00414_));
 sg13g2_mux2_1 _09924_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .S(net142),
    .X(_00415_));
 sg13g2_nand2_1 _09925_ (.Y(_04232_),
    .A(_01662_),
    .B(net143));
 sg13g2_o21ai_1 _09926_ (.B1(_04232_),
    .Y(_00416_),
    .A1(_01809_),
    .A2(net144));
 sg13g2_mux2_1 _09927_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .S(net142),
    .X(_00417_));
 sg13g2_mux2_1 _09928_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .S(net142),
    .X(_00418_));
 sg13g2_buf_1 _09929_ (.A(_04227_),
    .X(_04233_));
 sg13g2_mux2_1 _09930_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S(net141),
    .X(_00419_));
 sg13g2_mux2_1 _09931_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .S(net141),
    .X(_00420_));
 sg13g2_mux2_1 _09932_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .S(net141),
    .X(_00421_));
 sg13g2_mux2_1 _09933_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .S(net141),
    .X(_00422_));
 sg13g2_mux2_1 _09934_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .S(_04233_),
    .X(_00423_));
 sg13g2_mux2_1 _09935_ (.A0(_02445_),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .S(_04233_),
    .X(_00424_));
 sg13g2_nand2_1 _09936_ (.Y(_04234_),
    .A(_01167_),
    .B(_01179_));
 sg13g2_buf_2 _09937_ (.A(_04234_),
    .X(_04235_));
 sg13g2_and2_1 _09938_ (.A(_02386_),
    .B(_01648_),
    .X(_04236_));
 sg13g2_buf_2 _09939_ (.A(_04236_),
    .X(_04237_));
 sg13g2_nor2_1 _09940_ (.A(_01039_),
    .B(_04237_),
    .Y(_04238_));
 sg13g2_a21oi_1 _09941_ (.A1(_02404_),
    .A2(_04237_),
    .Y(_04239_),
    .B1(_04238_));
 sg13g2_nor2_1 _09942_ (.A(_04235_),
    .B(_04239_),
    .Y(_04240_));
 sg13g2_a21oi_1 _09943_ (.A1(_01709_),
    .A2(_04235_),
    .Y(_04241_),
    .B1(_04240_));
 sg13g2_nand2b_1 _09944_ (.Y(_04242_),
    .B(_04203_),
    .A_N(_04227_));
 sg13g2_nand2_1 _09945_ (.Y(_04243_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .B(net143));
 sg13g2_o21ai_1 _09946_ (.B1(_04243_),
    .Y(_00425_),
    .A1(_04241_),
    .A2(_04242_));
 sg13g2_nor2_1 _09947_ (.A(_01087_),
    .B(_04237_),
    .Y(_04244_));
 sg13g2_a21oi_1 _09948_ (.A1(_02543_),
    .A2(_04237_),
    .Y(_04245_),
    .B1(_04244_));
 sg13g2_nor2_1 _09949_ (.A(_04235_),
    .B(_04245_),
    .Y(_04246_));
 sg13g2_a21oi_1 _09950_ (.A1(net151),
    .A2(_04235_),
    .Y(_04247_),
    .B1(_04246_));
 sg13g2_nand2_1 _09951_ (.Y(_04248_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .B(net143));
 sg13g2_o21ai_1 _09952_ (.B1(_04248_),
    .Y(_00426_),
    .A1(_04242_),
    .A2(_04247_));
 sg13g2_nand2_1 _09953_ (.Y(_04249_),
    .A(_01664_),
    .B(net143));
 sg13g2_o21ai_1 _09954_ (.B1(_04249_),
    .Y(_00427_),
    .A1(_01868_),
    .A2(net144));
 sg13g2_nor2_1 _09955_ (.A(net173),
    .B(_01194_),
    .Y(_04250_));
 sg13g2_nor2_1 _09956_ (.A(_00916_),
    .B(_04237_),
    .Y(_04251_));
 sg13g2_a21oi_1 _09957_ (.A1(_02668_),
    .A2(_04237_),
    .Y(_04252_),
    .B1(_04251_));
 sg13g2_nand2_1 _09958_ (.Y(_04253_),
    .A(_01696_),
    .B(_04235_));
 sg13g2_o21ai_1 _09959_ (.B1(_04253_),
    .Y(_04254_),
    .A1(_04235_),
    .A2(_04252_));
 sg13g2_a22oi_1 _09960_ (.Y(_04255_),
    .B1(_04254_),
    .B2(_04203_),
    .A2(_04250_),
    .A1(_02728_));
 sg13g2_nand2_1 _09961_ (.Y(_04256_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .B(net143));
 sg13g2_o21ai_1 _09962_ (.B1(_04256_),
    .Y(_00428_),
    .A1(net144),
    .A2(_04255_));
 sg13g2_nor2b_1 _09963_ (.A(_04237_),
    .B_N(_00954_),
    .Y(_04257_));
 sg13g2_a21oi_1 _09964_ (.A1(_02822_),
    .A2(_04237_),
    .Y(_04258_),
    .B1(_04257_));
 sg13g2_nor2_1 _09965_ (.A(_04235_),
    .B(_04258_),
    .Y(_04259_));
 sg13g2_a21oi_1 _09966_ (.A1(net154),
    .A2(_04235_),
    .Y(_04260_),
    .B1(_04259_));
 sg13g2_nor2_2 _09967_ (.A(_01185_),
    .B(net173),
    .Y(_04261_));
 sg13g2_a21oi_1 _09968_ (.A1(_04203_),
    .A2(_04260_),
    .Y(_04262_),
    .B1(_04261_));
 sg13g2_nand2_1 _09969_ (.Y(_04263_),
    .A(_02445_),
    .B(net143));
 sg13g2_o21ai_1 _09970_ (.B1(_04263_),
    .Y(_00429_),
    .A1(net144),
    .A2(_04262_));
 sg13g2_nand2_1 _09971_ (.Y(_04264_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net143));
 sg13g2_o21ai_1 _09972_ (.B1(_04264_),
    .Y(_00430_),
    .A1(_01905_),
    .A2(net144));
 sg13g2_nand2_1 _09973_ (.Y(_04265_),
    .A(_01765_),
    .B(_04229_));
 sg13g2_o21ai_1 _09974_ (.B1(_04265_),
    .Y(_00431_),
    .A1(_01932_),
    .A2(net144));
 sg13g2_nand2_1 _09975_ (.Y(_04266_),
    .A(_01808_),
    .B(net143));
 sg13g2_o21ai_1 _09976_ (.B1(_04266_),
    .Y(_00432_),
    .A1(_01981_),
    .A2(net144));
 sg13g2_mux2_1 _09977_ (.A0(net294),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .S(net141),
    .X(_00433_));
 sg13g2_mux2_1 _09978_ (.A0(net293),
    .A1(_01872_),
    .S(net141),
    .X(_00434_));
 sg13g2_mux2_1 _09979_ (.A0(_02045_),
    .A1(_01910_),
    .S(net141),
    .X(_00435_));
 sg13g2_mux2_1 _09980_ (.A0(net292),
    .A1(_01934_),
    .S(net141),
    .X(_00436_));
 sg13g2_mux2_1 _09981_ (.A0(net8),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .S(net217),
    .X(_00631_));
 sg13g2_mux2_1 _09982_ (.A0(net9),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .S(net217),
    .X(_00632_));
 sg13g2_mux2_1 _09983_ (.A0(net10),
    .A1(_04102_),
    .S(net217),
    .X(_00633_));
 sg13g2_a21oi_1 _09984_ (.A1(\i_tinyqv.cpu.i_core.interrupt_req[1] ),
    .A2(_03132_),
    .Y(_04267_),
    .B1(_01370_));
 sg13g2_o21ai_1 _09985_ (.B1(_02193_),
    .Y(_04268_),
    .A1(_01537_),
    .A2(_02349_));
 sg13g2_nand2_1 _09986_ (.Y(_04269_),
    .A(_00968_),
    .B(_04268_));
 sg13g2_nand2_1 _09987_ (.Y(_04270_),
    .A(_00745_),
    .B(_02390_));
 sg13g2_a21oi_1 _09988_ (.A1(_01179_),
    .A2(_04270_),
    .Y(_04271_),
    .B1(_04204_));
 sg13g2_a21oi_1 _09989_ (.A1(net151),
    .A2(_04271_),
    .Y(_04272_),
    .B1(_02358_));
 sg13g2_or2_1 _09990_ (.X(_04273_),
    .B(_04272_),
    .A(_04269_));
 sg13g2_nor2_1 _09991_ (.A(_01699_),
    .B(_04205_),
    .Y(_04274_));
 sg13g2_o21ai_1 _09992_ (.B1(_01370_),
    .Y(_04275_),
    .A1(_04269_),
    .A2(_04274_));
 sg13g2_a221oi_1 _09993_ (.B2(_04275_),
    .C1(net105),
    .B1(_04273_),
    .A1(_02358_),
    .Y(_00222_),
    .A2(_04267_));
 sg13g2_a21oi_1 _09994_ (.A1(net133),
    .A2(_04271_),
    .Y(_04276_),
    .B1(_02358_));
 sg13g2_or2_1 _09995_ (.X(_04277_),
    .B(_04276_),
    .A(_04269_));
 sg13g2_nor2_1 _09996_ (.A(_01709_),
    .B(_04205_),
    .Y(_04278_));
 sg13g2_o21ai_1 _09997_ (.B1(\i_tinyqv.cpu.i_core.mip[16] ),
    .Y(_04279_),
    .A1(_04269_),
    .A2(_04278_));
 sg13g2_a21oi_1 _09998_ (.A1(\i_tinyqv.cpu.i_core.interrupt_req[0] ),
    .A2(_03126_),
    .Y(_04280_),
    .B1(\i_tinyqv.cpu.i_core.mip[16] ));
 sg13g2_a221oi_1 _09999_ (.B2(_02358_),
    .C1(net105),
    .B1(_04280_),
    .A1(_04277_),
    .Y(_00223_),
    .A2(_04279_));
 sg13g2_nor2_1 _10000_ (.A(_04221_),
    .B(_04205_),
    .Y(_04281_));
 sg13g2_nand2b_1 _10001_ (.Y(_04282_),
    .B(_02369_),
    .A_N(_01537_));
 sg13g2_buf_1 _10002_ (.A(_04282_),
    .X(_04283_));
 sg13g2_o21ai_1 _10003_ (.B1(_01390_),
    .Y(_04284_),
    .A1(_04281_),
    .A2(_04283_));
 sg13g2_a21o_1 _10004_ (.A2(_04270_),
    .A1(_01179_),
    .B1(_04204_),
    .X(_04285_));
 sg13g2_nor2_1 _10005_ (.A(_04285_),
    .B(_04283_),
    .Y(_04286_));
 sg13g2_nand2_1 _10006_ (.Y(_04287_),
    .A(_04221_),
    .B(_04286_));
 sg13g2_a21oi_1 _10007_ (.A1(_04284_),
    .A2(_04287_),
    .Y(_00224_),
    .B1(net105));
 sg13g2_nor2_1 _10008_ (.A(_01696_),
    .B(_04205_),
    .Y(_04288_));
 sg13g2_o21ai_1 _10009_ (.B1(_01374_),
    .Y(_04289_),
    .A1(_04283_),
    .A2(_04288_));
 sg13g2_nand2_1 _10010_ (.Y(_04290_),
    .A(_01696_),
    .B(_04286_));
 sg13g2_a21oi_1 _10011_ (.A1(_04289_),
    .A2(_04290_),
    .Y(_00225_),
    .B1(net105));
 sg13g2_o21ai_1 _10012_ (.B1(\i_tinyqv.cpu.i_core.mie[17] ),
    .Y(_04291_),
    .A1(_04274_),
    .A2(_04283_));
 sg13g2_nand2_1 _10013_ (.Y(_04292_),
    .A(_01699_),
    .B(_04286_));
 sg13g2_a21oi_1 _10014_ (.A1(_04291_),
    .A2(_04292_),
    .Y(_00226_),
    .B1(_03129_));
 sg13g2_o21ai_1 _10015_ (.B1(\i_tinyqv.cpu.i_core.mie[16] ),
    .Y(_04293_),
    .A1(_04278_),
    .A2(_04283_));
 sg13g2_nand2_1 _10016_ (.Y(_04294_),
    .A(net133),
    .B(_04286_));
 sg13g2_a21oi_1 _10017_ (.A1(_04293_),
    .A2(_04294_),
    .Y(_00227_),
    .B1(net105));
 sg13g2_and3_1 _10018_ (.X(_04295_),
    .A(\i_debug_uart_tx.cycle_counter[1] ),
    .B(\i_debug_uart_tx.cycle_counter[0] ),
    .C(\i_debug_uart_tx.cycle_counter[2] ));
 sg13g2_buf_1 _10019_ (.A(_04295_),
    .X(_04296_));
 sg13g2_and3_1 _10020_ (.X(_04297_),
    .A(\i_debug_uart_tx.cycle_counter[3] ),
    .B(_00166_),
    .C(_04296_));
 sg13g2_buf_1 _10021_ (.A(_04297_),
    .X(_04298_));
 sg13g2_buf_1 _10022_ (.A(_04298_),
    .X(_04299_));
 sg13g2_nor3_1 _10023_ (.A(net290),
    .B(_02199_),
    .C(_02196_),
    .Y(_04300_));
 sg13g2_nor2b_1 _10024_ (.A(_02198_),
    .B_N(_04300_),
    .Y(_04301_));
 sg13g2_and2_1 _10025_ (.A(\i_debug_uart_tx.cycle_counter[0] ),
    .B(_04301_),
    .X(_04302_));
 sg13g2_a21oi_1 _10026_ (.A1(_00217_),
    .A2(net206),
    .Y(_04303_),
    .B1(_04302_));
 sg13g2_nor3_1 _10027_ (.A(net215),
    .B(_04299_),
    .C(_04303_),
    .Y(_00229_));
 sg13g2_nand2_1 _10028_ (.Y(_04304_),
    .A(\i_debug_uart_tx.cycle_counter[0] ),
    .B(net206));
 sg13g2_xor2_1 _10029_ (.B(_04304_),
    .A(\i_debug_uart_tx.cycle_counter[1] ),
    .X(_04305_));
 sg13g2_nor3_1 _10030_ (.A(net215),
    .B(_04299_),
    .C(_04305_),
    .Y(_00230_));
 sg13g2_nand3_1 _10031_ (.B(\i_debug_uart_tx.cycle_counter[0] ),
    .C(net206),
    .A(\i_debug_uart_tx.cycle_counter[1] ),
    .Y(_04306_));
 sg13g2_xor2_1 _10032_ (.B(_04306_),
    .A(\i_debug_uart_tx.cycle_counter[2] ),
    .X(_04307_));
 sg13g2_nor3_1 _10033_ (.A(net215),
    .B(net180),
    .C(_04307_),
    .Y(_00231_));
 sg13g2_o21ai_1 _10034_ (.B1(_04296_),
    .Y(_04308_),
    .A1(_00166_),
    .A2(net206));
 sg13g2_nand2_1 _10035_ (.Y(_04309_),
    .A(\i_debug_uart_tx.cycle_counter[3] ),
    .B(_04308_));
 sg13g2_nand3b_1 _10036_ (.B(net206),
    .C(_04296_),
    .Y(_04310_),
    .A_N(\i_debug_uart_tx.cycle_counter[3] ));
 sg13g2_a21oi_1 _10037_ (.A1(_04309_),
    .A2(_04310_),
    .Y(_00232_),
    .B1(_02862_));
 sg13g2_nor2_1 _10038_ (.A(_00166_),
    .B(net206),
    .Y(_04311_));
 sg13g2_nor2_1 _10039_ (.A(\i_debug_uart_tx.cycle_counter[4] ),
    .B(net206),
    .Y(_04312_));
 sg13g2_a221oi_1 _10040_ (.B2(\i_debug_uart_tx.cycle_counter[3] ),
    .C1(_04312_),
    .B1(_04296_),
    .A1(_00166_),
    .Y(_04313_),
    .A2(_02202_));
 sg13g2_a21oi_1 _10041_ (.A1(\i_debug_uart_tx.cycle_counter[4] ),
    .A2(_04311_),
    .Y(_04314_),
    .B1(_04313_));
 sg13g2_nor2_1 _10042_ (.A(net215),
    .B(_04314_),
    .Y(_00233_));
 sg13g2_nand2_1 _10043_ (.Y(_04315_),
    .A(_01170_),
    .B(net85));
 sg13g2_a21oi_1 _10044_ (.A1(\i_tinyqv.cpu.load_started ),
    .A2(_01565_),
    .Y(_04316_),
    .B1(_04315_));
 sg13g2_nand2_1 _10045_ (.Y(_04317_),
    .A(_01263_),
    .B(_01652_));
 sg13g2_nand2_1 _10046_ (.Y(_04318_),
    .A(_01233_),
    .B(net134));
 sg13g2_nand3_1 _10047_ (.B(_04317_),
    .C(_04318_),
    .A(_04316_),
    .Y(_00339_));
 sg13g2_nand2_1 _10048_ (.Y(_04319_),
    .A(\i_tinyqv.cpu.data_read_n[1] ),
    .B(net134));
 sg13g2_nand2_1 _10049_ (.Y(_04320_),
    .A(_02250_),
    .B(_01652_));
 sg13g2_nand3_1 _10050_ (.B(_04319_),
    .C(_04320_),
    .A(_04316_),
    .Y(_00340_));
 sg13g2_nor2_1 _10051_ (.A(\i_tinyqv.cpu.data_ready_latch ),
    .B(_01565_),
    .Y(_04321_));
 sg13g2_nor3_1 _10052_ (.A(_01643_),
    .B(_01166_),
    .C(_04321_),
    .Y(_00342_));
 sg13g2_a21oi_2 _10053_ (.B1(net173),
    .Y(_04322_),
    .A2(_01194_),
    .A1(_01185_));
 sg13g2_nor3_1 _10054_ (.A(net154),
    .B(_04285_),
    .C(_04322_),
    .Y(_04323_));
 sg13g2_nand2b_1 _10055_ (.Y(_04324_),
    .B(_02344_),
    .A_N(_01537_));
 sg13g2_a21oi_1 _10056_ (.A1(_00745_),
    .A2(net154),
    .Y(_04325_),
    .B1(_04324_));
 sg13g2_o21ai_1 _10057_ (.B1(_02381_),
    .Y(_04326_),
    .A1(net137),
    .A2(_04325_));
 sg13g2_mux2_1 _10058_ (.A0(_04323_),
    .A1(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .S(_04326_),
    .X(_04327_));
 sg13g2_nor2_2 _10059_ (.A(_04250_),
    .B(_04261_),
    .Y(_04328_));
 sg13g2_a21oi_1 _10060_ (.A1(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .A2(_04328_),
    .Y(_04329_),
    .B1(_04323_));
 sg13g2_nand2_1 _10061_ (.Y(_04330_),
    .A(net148),
    .B(_04329_));
 sg13g2_o21ai_1 _10062_ (.B1(_04330_),
    .Y(_04331_),
    .A1(net148),
    .A2(_04327_));
 sg13g2_nand2b_1 _10063_ (.Y(_00390_),
    .B(_04331_),
    .A_N(net105));
 sg13g2_nor2_1 _10064_ (.A(net148),
    .B(_02363_),
    .Y(_04332_));
 sg13g2_a21oi_1 _10065_ (.A1(_04325_),
    .A2(_04332_),
    .Y(_04333_),
    .B1(_04322_));
 sg13g2_nand2_1 _10066_ (.Y(_04334_),
    .A(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .B(_04333_));
 sg13g2_nand3_1 _10067_ (.B(_02381_),
    .C(net137),
    .A(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .Y(_04335_));
 sg13g2_nand2b_1 _10068_ (.Y(_04336_),
    .B(_04335_),
    .A_N(_04323_));
 sg13g2_nand2b_1 _10069_ (.Y(_04337_),
    .B(_04336_),
    .A_N(_04333_));
 sg13g2_a21oi_1 _10070_ (.A1(_04334_),
    .A2(_04337_),
    .Y(_00391_),
    .B1(net105));
 sg13g2_o21ai_1 _10071_ (.B1(_04328_),
    .Y(_04338_),
    .A1(_02728_),
    .A2(net148));
 sg13g2_nand2b_1 _10072_ (.Y(_00392_),
    .B(_04338_),
    .A_N(_03129_));
 sg13g2_nor2_1 _10073_ (.A(_02168_),
    .B(_02165_),
    .Y(_04339_));
 sg13g2_nor2_1 _10074_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .B(_04339_),
    .Y(_04340_));
 sg13g2_a21oi_1 _10075_ (.A1(_02168_),
    .A2(_02165_),
    .Y(_04341_),
    .B1(_04340_));
 sg13g2_nand2_1 _10076_ (.Y(_04342_),
    .A(net292),
    .B(net109));
 sg13g2_nand2b_1 _10077_ (.Y(_04343_),
    .B(net132),
    .A_N(_02108_));
 sg13g2_inv_1 _10078_ (.Y(_04344_),
    .A(net119));
 sg13g2_nand2_1 _10079_ (.Y(_04345_),
    .A(_02108_),
    .B(net291));
 sg13g2_or4_1 _10080_ (.A(_04344_),
    .B(_02046_),
    .C(net132),
    .D(_04345_),
    .X(_04346_));
 sg13g2_a21oi_1 _10081_ (.A1(_04343_),
    .A2(_04346_),
    .Y(_04347_),
    .B1(net292));
 sg13g2_o21ai_1 _10082_ (.B1(net291),
    .Y(_04348_),
    .A1(_02046_),
    .A2(_02083_));
 sg13g2_nor2b_1 _10083_ (.A(net242),
    .B_N(_04348_),
    .Y(_04349_));
 sg13g2_a21o_1 _10084_ (.A2(_02106_),
    .A1(net119),
    .B1(net291),
    .X(_04350_));
 sg13g2_o21ai_1 _10085_ (.B1(_04350_),
    .Y(_04351_),
    .A1(net119),
    .A2(_02083_));
 sg13g2_nand3b_1 _10086_ (.B(net119),
    .C(net118),
    .Y(_04352_),
    .A_N(_02108_));
 sg13g2_o21ai_1 _10087_ (.B1(_04352_),
    .Y(_04353_),
    .A1(net118),
    .A2(_04345_));
 sg13g2_a22oi_1 _10088_ (.Y(_04354_),
    .B1(_04353_),
    .B2(net292),
    .A2(_04344_),
    .A1(net242));
 sg13g2_nor2_1 _10089_ (.A(_01736_),
    .B(_04354_),
    .Y(_04355_));
 sg13g2_nor4_2 _10090_ (.A(_04347_),
    .B(_04349_),
    .C(_04351_),
    .Y(_04356_),
    .D(_04355_));
 sg13g2_xor2_1 _10091_ (.B(_04356_),
    .A(_04342_),
    .X(_04357_));
 sg13g2_xnor2_1 _10092_ (.Y(_04358_),
    .A(_04341_),
    .B(_04357_));
 sg13g2_buf_2 _10093_ (.A(_04358_),
    .X(_04359_));
 sg13g2_inv_1 _10094_ (.Y(_04360_),
    .A(_02159_));
 sg13g2_nand2_1 _10095_ (.Y(_04361_),
    .A(_02155_),
    .B(_04360_));
 sg13g2_nor2_1 _10096_ (.A(_02155_),
    .B(_04360_),
    .Y(_04362_));
 sg13g2_nand2_1 _10097_ (.Y(_04363_),
    .A(_02172_),
    .B(_04362_));
 sg13g2_o21ai_1 _10098_ (.B1(_04363_),
    .Y(_04364_),
    .A1(_02174_),
    .A2(_04361_));
 sg13g2_a21oi_1 _10099_ (.A1(_02159_),
    .A2(_02174_),
    .Y(_04365_),
    .B1(_02172_));
 sg13g2_nand2_1 _10100_ (.Y(_04366_),
    .A(_02159_),
    .B(_02172_));
 sg13g2_o21ai_1 _10101_ (.B1(_04366_),
    .Y(_04367_),
    .A1(_02155_),
    .A2(_04365_));
 sg13g2_nand2_1 _10102_ (.Y(_04368_),
    .A(_02155_),
    .B(_04365_));
 sg13g2_o21ai_1 _10103_ (.B1(_04368_),
    .Y(_04369_),
    .A1(_02159_),
    .A2(_02174_));
 sg13g2_mux2_1 _10104_ (.A0(_04367_),
    .A1(_04369_),
    .S(_02150_),
    .X(_04370_));
 sg13g2_nor2_1 _10105_ (.A(_04364_),
    .B(_04370_),
    .Y(_04371_));
 sg13g2_xor2_1 _10106_ (.B(_04371_),
    .A(_04359_),
    .X(_00393_));
 sg13g2_o21ai_1 _10107_ (.B1(_02174_),
    .Y(_04372_),
    .A1(_04359_),
    .A2(_04362_));
 sg13g2_nand3_1 _10108_ (.B(_04359_),
    .C(_04361_),
    .A(_02174_),
    .Y(_04373_));
 sg13g2_o21ai_1 _10109_ (.B1(_04373_),
    .Y(_04374_),
    .A1(_02150_),
    .A2(_04372_));
 sg13g2_buf_1 _10110_ (.A(_04374_),
    .X(_04375_));
 sg13g2_o21ai_1 _10111_ (.B1(_04361_),
    .Y(_04376_),
    .A1(_02172_),
    .A2(_04359_));
 sg13g2_nor2_1 _10112_ (.A(_02172_),
    .B(_04359_),
    .Y(_04377_));
 sg13g2_nor2_1 _10113_ (.A(_02155_),
    .B(_04377_),
    .Y(_04378_));
 sg13g2_a22oi_1 _10114_ (.Y(_04379_),
    .B1(_04378_),
    .B2(_02159_),
    .A2(_04359_),
    .A1(_02172_));
 sg13g2_o21ai_1 _10115_ (.B1(_04379_),
    .Y(_04380_),
    .A1(_02150_),
    .A2(_04376_));
 sg13g2_buf_2 _10116_ (.A(_04380_),
    .X(_04381_));
 sg13g2_nor2_1 _10117_ (.A(_04375_),
    .B(_04381_),
    .Y(_04382_));
 sg13g2_nand2b_1 _10118_ (.Y(_04383_),
    .B(_04341_),
    .A_N(_04357_));
 sg13g2_buf_1 _10119_ (.A(_04383_),
    .X(_04384_));
 sg13g2_nor2_1 _10120_ (.A(net132),
    .B(net109),
    .Y(_04385_));
 sg13g2_nand4_1 _10121_ (.B(_02081_),
    .C(_01814_),
    .A(net291),
    .Y(_04386_),
    .D(net109));
 sg13g2_nand2b_1 _10122_ (.Y(_04387_),
    .B(_04386_),
    .A_N(_04385_));
 sg13g2_a22oi_1 _10123_ (.Y(_04388_),
    .B1(net109),
    .B2(net242),
    .A2(net119),
    .A1(net291));
 sg13g2_a21o_1 _10124_ (.A2(_04387_),
    .A1(net242),
    .B1(_04388_),
    .X(_04389_));
 sg13g2_buf_1 _10125_ (.A(_04389_),
    .X(_04390_));
 sg13g2_nand2b_1 _10126_ (.Y(_04391_),
    .B(_04356_),
    .A_N(_04342_));
 sg13g2_a21oi_1 _10127_ (.A1(net120),
    .A2(net132),
    .Y(_04392_),
    .B1(_03020_));
 sg13g2_a21oi_1 _10128_ (.A1(_03020_),
    .A2(net132),
    .Y(_04393_),
    .B1(_04392_));
 sg13g2_nor3_1 _10129_ (.A(net242),
    .B(_03020_),
    .C(_01682_),
    .Y(_04394_));
 sg13g2_a21oi_1 _10130_ (.A1(net242),
    .A2(_04393_),
    .Y(_04395_),
    .B1(_04394_));
 sg13g2_nor2_1 _10131_ (.A(_02161_),
    .B(_04395_),
    .Y(_04396_));
 sg13g2_nor3_1 _10132_ (.A(net119),
    .B(_01682_),
    .C(_04345_),
    .Y(_04397_));
 sg13g2_nor2_1 _10133_ (.A(_04396_),
    .B(_04397_),
    .Y(_04398_));
 sg13g2_nand2_1 _10134_ (.Y(_04399_),
    .A(_04391_),
    .B(_04398_));
 sg13g2_nand2b_1 _10135_ (.Y(_04400_),
    .B(_04399_),
    .A_N(_04390_));
 sg13g2_inv_1 _10136_ (.Y(_04401_),
    .A(_04399_));
 sg13g2_nand2_1 _10137_ (.Y(_04402_),
    .A(_04390_),
    .B(_04401_));
 sg13g2_nand2_1 _10138_ (.Y(_04403_),
    .A(_04400_),
    .B(_04402_));
 sg13g2_xor2_1 _10139_ (.B(_04403_),
    .A(_04384_),
    .X(_04404_));
 sg13g2_xnor2_1 _10140_ (.Y(_00394_),
    .A(_04382_),
    .B(_04404_));
 sg13g2_nand2_1 _10141_ (.Y(_04405_),
    .A(net242),
    .B(_02081_));
 sg13g2_mux2_1 _10142_ (.A0(_04385_),
    .A1(net109),
    .S(_04405_),
    .X(_04406_));
 sg13g2_nand2_1 _10143_ (.Y(_04407_),
    .A(net291),
    .B(_04406_));
 sg13g2_or3_1 _10144_ (.A(_04375_),
    .B(_04381_),
    .C(_04402_),
    .X(_04408_));
 sg13g2_nor3_1 _10145_ (.A(_04384_),
    .B(_04390_),
    .C(_04401_),
    .Y(_04409_));
 sg13g2_o21ai_1 _10146_ (.B1(_04409_),
    .Y(_04410_),
    .A1(_04375_),
    .A2(_04381_));
 sg13g2_nand3_1 _10147_ (.B(_04390_),
    .C(_04401_),
    .A(_04384_),
    .Y(_04411_));
 sg13g2_nand2_1 _10148_ (.Y(_04412_),
    .A(_04384_),
    .B(_04400_));
 sg13g2_or3_1 _10149_ (.A(_04375_),
    .B(_04381_),
    .C(_04412_),
    .X(_04413_));
 sg13g2_nand4_1 _10150_ (.B(_04410_),
    .C(_04411_),
    .A(_04408_),
    .Y(_04414_),
    .D(_04413_));
 sg13g2_xor2_1 _10151_ (.B(_04414_),
    .A(_04407_),
    .X(_00395_));
 sg13g2_nor4_1 _10152_ (.A(_01174_),
    .B(_01686_),
    .C(_00856_),
    .D(_04345_),
    .Y(_04415_));
 sg13g2_o21ai_1 _10153_ (.B1(_04399_),
    .Y(_04416_),
    .A1(_04375_),
    .A2(_04381_));
 sg13g2_nor2_1 _10154_ (.A(_04407_),
    .B(_04416_),
    .Y(_04417_));
 sg13g2_nor2b_1 _10155_ (.A(_04399_),
    .B_N(_04384_),
    .Y(_04418_));
 sg13g2_a21o_1 _10156_ (.A2(_04407_),
    .A1(_04384_),
    .B1(_04390_),
    .X(_04419_));
 sg13g2_a221oi_1 _10157_ (.B2(_04416_),
    .C1(_04419_),
    .B1(_04407_),
    .A1(_04382_),
    .Y(_04420_),
    .A2(_04418_));
 sg13g2_or3_1 _10158_ (.A(_04415_),
    .B(_04417_),
    .C(_04420_),
    .X(_00396_));
 sg13g2_nor3_1 _10159_ (.A(net260),
    .B(_01438_),
    .C(_03417_),
    .Y(_00560_));
 sg13g2_a21oi_1 _10160_ (.A1(_01428_),
    .A2(_04088_),
    .Y(_04421_),
    .B1(_03623_));
 sg13g2_nor3_1 _10161_ (.A(net215),
    .B(_04091_),
    .C(_04421_),
    .Y(_00594_));
 sg13g2_inv_1 _10162_ (.Y(_04422_),
    .A(_04095_));
 sg13g2_nand3_1 _10163_ (.B(_04009_),
    .C(_04010_),
    .A(net234),
    .Y(_04423_));
 sg13g2_nor3_1 _10164_ (.A(net47),
    .B(_04101_),
    .C(_04423_),
    .Y(_00630_));
 sg13g2_buf_1 _10165_ (.A(net232),
    .X(_04424_));
 sg13g2_nand2_1 _10166_ (.Y(_04425_),
    .A(net232),
    .B(_04112_));
 sg13g2_nor2_1 _10167_ (.A(_04026_),
    .B(_04112_),
    .Y(_04426_));
 sg13g2_a21o_1 _10168_ (.A2(_04425_),
    .A1(_04002_),
    .B1(_04426_),
    .X(_04427_));
 sg13g2_nand2b_1 _10169_ (.Y(_04428_),
    .B(_01518_),
    .A_N(net232));
 sg13g2_inv_1 _10170_ (.Y(_04429_),
    .A(\addr[24] ));
 sg13g2_nor3_2 _10171_ (.A(_01423_),
    .B(_04429_),
    .C(_03623_),
    .Y(_04430_));
 sg13g2_nand2b_1 _10172_ (.Y(_04431_),
    .B(_03903_),
    .A_N(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ));
 sg13g2_o21ai_1 _10173_ (.B1(_04431_),
    .Y(_04432_),
    .A1(_03903_),
    .A2(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ));
 sg13g2_a21oi_2 _10174_ (.B1(_03629_),
    .Y(_04433_),
    .A2(_04432_),
    .A1(_04430_));
 sg13g2_a221oi_1 _10175_ (.B2(_04426_),
    .C1(_04433_),
    .B1(_04428_),
    .A1(_03999_),
    .Y(_04434_),
    .A2(_04427_));
 sg13g2_buf_1 _10176_ (.A(_04434_),
    .X(_04435_));
 sg13g2_nand2_1 _10177_ (.Y(_04436_),
    .A(net214),
    .B(_04435_));
 sg13g2_a21oi_1 _10178_ (.A1(_04122_),
    .A2(_04118_),
    .Y(_04437_),
    .B1(_04435_));
 sg13g2_nand2_1 _10179_ (.Y(_04438_),
    .A(\addr[24] ),
    .B(net71));
 sg13g2_nand2_1 _10180_ (.Y(_04439_),
    .A(_01520_),
    .B(_04438_));
 sg13g2_a21oi_1 _10181_ (.A1(net238),
    .A2(net200),
    .Y(_04440_),
    .B1(_00163_));
 sg13g2_nand2b_1 _10182_ (.Y(_04441_),
    .B(net281),
    .A_N(net232));
 sg13g2_nand2b_1 _10183_ (.Y(_04442_),
    .B(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .A_N(_03995_));
 sg13g2_nor3_1 _10184_ (.A(_01519_),
    .B(_04441_),
    .C(_04442_),
    .Y(_04443_));
 sg13g2_nor3_1 _10185_ (.A(_04035_),
    .B(_04440_),
    .C(_04443_),
    .Y(_04444_));
 sg13g2_a21oi_1 _10186_ (.A1(_04035_),
    .A2(_04107_),
    .Y(_04445_),
    .B1(_04444_));
 sg13g2_nand4_1 _10187_ (.B(_04006_),
    .C(_04105_),
    .A(_04088_),
    .Y(_04446_),
    .D(_04445_));
 sg13g2_nand3_1 _10188_ (.B(_04439_),
    .C(_04446_),
    .A(_04437_),
    .Y(_04447_));
 sg13g2_a21oi_1 _10189_ (.A1(_04436_),
    .A2(_04447_),
    .Y(_00634_),
    .B1(net47));
 sg13g2_nor2_1 _10190_ (.A(net235),
    .B(_04437_),
    .Y(_04448_));
 sg13g2_o21ai_1 _10191_ (.B1(net214),
    .Y(_04449_),
    .A1(_03633_),
    .A2(net231));
 sg13g2_a21oi_1 _10192_ (.A1(net231),
    .A2(_04107_),
    .Y(_04450_),
    .B1(_04449_));
 sg13g2_or2_1 _10193_ (.X(_04451_),
    .B(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .A(_03995_));
 sg13g2_or2_1 _10194_ (.X(_04452_),
    .B(_04441_),
    .A(net279));
 sg13g2_buf_1 _10195_ (.A(_04452_),
    .X(_04453_));
 sg13g2_a21oi_1 _10196_ (.A1(net238),
    .A2(_04451_),
    .Y(_04454_),
    .B1(_04453_));
 sg13g2_o21ai_1 _10197_ (.B1(_04105_),
    .Y(_04455_),
    .A1(_04450_),
    .A2(_04454_));
 sg13g2_or2_1 _10198_ (.X(_04456_),
    .B(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .A(_04102_));
 sg13g2_nand3_1 _10199_ (.B(_04122_),
    .C(_04456_),
    .A(_00162_),
    .Y(_04457_));
 sg13g2_and4_1 _10200_ (.A(_04437_),
    .B(_04439_),
    .C(_04455_),
    .D(_04457_),
    .X(_04458_));
 sg13g2_nor3_1 _10201_ (.A(net47),
    .B(_04448_),
    .C(_04458_),
    .Y(_00635_));
 sg13g2_nor2b_1 _10202_ (.A(net231),
    .B_N(_04435_),
    .Y(_04459_));
 sg13g2_nand2b_1 _10203_ (.Y(_04460_),
    .B(_04009_),
    .A_N(net279));
 sg13g2_nor3_1 _10204_ (.A(net214),
    .B(_04451_),
    .C(_04460_),
    .Y(_04461_));
 sg13g2_a21oi_1 _10205_ (.A1(_04424_),
    .A2(_04460_),
    .Y(_04462_),
    .B1(net235));
 sg13g2_o21ai_1 _10206_ (.B1(net238),
    .Y(_04463_),
    .A1(_04461_),
    .A2(_04462_));
 sg13g2_nor2_1 _10207_ (.A(net279),
    .B(_04026_),
    .Y(_04464_));
 sg13g2_nand4_1 _10208_ (.B(net214),
    .C(_01519_),
    .A(net235),
    .Y(_04465_),
    .D(_04464_));
 sg13g2_a21oi_1 _10209_ (.A1(_04463_),
    .A2(_04465_),
    .Y(_04466_),
    .B1(_04435_));
 sg13g2_nor3_1 _10210_ (.A(net47),
    .B(_04459_),
    .C(_04466_),
    .Y(_00636_));
 sg13g2_a21o_1 _10211_ (.A2(_04432_),
    .A1(_04430_),
    .B1(_03629_),
    .X(_04467_));
 sg13g2_buf_2 _10212_ (.A(_04467_),
    .X(_04468_));
 sg13g2_a21oi_1 _10213_ (.A1(_01233_),
    .A2(\i_tinyqv.cpu.data_read_n[1] ),
    .Y(_04469_),
    .B1(_01227_));
 sg13g2_and2_1 _10214_ (.A(_01522_),
    .B(_04469_),
    .X(_04470_));
 sg13g2_nor4_1 _10215_ (.A(_03623_),
    .B(_04438_),
    .C(_04468_),
    .D(_04470_),
    .Y(_04471_));
 sg13g2_a21oi_1 _10216_ (.A1(net234),
    .A2(_04468_),
    .Y(_04472_),
    .B1(_04471_));
 sg13g2_nor2_1 _10217_ (.A(_04422_),
    .B(_04472_),
    .Y(_00637_));
 sg13g2_nand2_1 _10218_ (.Y(_04473_),
    .A(_04088_),
    .B(_04006_));
 sg13g2_nand2_1 _10219_ (.Y(_04474_),
    .A(_04101_),
    .B(_04460_));
 sg13g2_a22oi_1 _10220_ (.Y(_04475_),
    .B1(_04474_),
    .B2(_03633_),
    .A2(_04464_),
    .A1(_04085_));
 sg13g2_nor2_1 _10221_ (.A(_03633_),
    .B(_04002_),
    .Y(_04476_));
 sg13g2_o21ai_1 _10222_ (.B1(_04112_),
    .Y(_04477_),
    .A1(net232),
    .A2(_04476_));
 sg13g2_o21ai_1 _10223_ (.B1(_04477_),
    .Y(_04478_),
    .A1(net238),
    .A2(_04475_));
 sg13g2_a21o_1 _10224_ (.A2(_04473_),
    .A1(_04468_),
    .B1(_04478_),
    .X(_04479_));
 sg13g2_buf_2 _10225_ (.A(_04479_),
    .X(_04480_));
 sg13g2_nand3_1 _10226_ (.B(_04088_),
    .C(_04104_),
    .A(_04007_),
    .Y(_04481_));
 sg13g2_nor2_1 _10227_ (.A(_04480_),
    .B(_04481_),
    .Y(_04482_));
 sg13g2_nor2b_1 _10228_ (.A(_04007_),
    .B_N(_04480_),
    .Y(_04483_));
 sg13g2_nor3_1 _10229_ (.A(net47),
    .B(_04482_),
    .C(_04483_),
    .Y(_00640_));
 sg13g2_nand2b_1 _10230_ (.Y(_04484_),
    .B(_04481_),
    .A_N(_04480_));
 sg13g2_nor2_1 _10231_ (.A(_03633_),
    .B(_01519_),
    .Y(_04485_));
 sg13g2_nand2b_1 _10232_ (.Y(_04486_),
    .B(net214),
    .A_N(net231));
 sg13g2_o21ai_1 _10233_ (.B1(_04486_),
    .Y(_04487_),
    .A1(net214),
    .A2(_04442_));
 sg13g2_a21oi_1 _10234_ (.A1(_04485_),
    .A2(_04487_),
    .Y(_04488_),
    .B1(_04008_));
 sg13g2_nand3_1 _10235_ (.B(_04024_),
    .C(_04104_),
    .A(_04088_),
    .Y(_04489_));
 sg13g2_nor3_1 _10236_ (.A(_04480_),
    .B(_04488_),
    .C(_04489_),
    .Y(_04490_));
 sg13g2_a21oi_1 _10237_ (.A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .A2(_04484_),
    .Y(_04491_),
    .B1(_04490_));
 sg13g2_nor2_1 _10238_ (.A(net47),
    .B(_04491_),
    .Y(_00641_));
 sg13g2_nand2_1 _10239_ (.Y(_04492_),
    .A(_04008_),
    .B(_04480_));
 sg13g2_nor2b_1 _10240_ (.A(_04024_),
    .B_N(_04008_),
    .Y(_04493_));
 sg13g2_a22oi_1 _10241_ (.Y(_04494_),
    .B1(_04493_),
    .B2(_04104_),
    .A2(_04464_),
    .A1(_04086_));
 sg13g2_o21ai_1 _10242_ (.B1(_04439_),
    .Y(_04495_),
    .A1(_01520_),
    .A2(_04494_));
 sg13g2_nand2b_1 _10243_ (.Y(_04496_),
    .B(_04495_),
    .A_N(_04480_));
 sg13g2_a21oi_1 _10244_ (.A1(_04492_),
    .A2(_04496_),
    .Y(_00642_),
    .B1(net47));
 sg13g2_nand3_1 _10245_ (.B(_01520_),
    .C(_04468_),
    .A(_03631_),
    .Y(_04497_));
 sg13g2_o21ai_1 _10246_ (.B1(_04497_),
    .Y(_04498_),
    .A1(_03631_),
    .A2(_04473_));
 sg13g2_and2_1 _10247_ (.A(_04095_),
    .B(_04498_),
    .X(_00646_));
 sg13g2_a22oi_1 _10248_ (.Y(_04499_),
    .B1(_04441_),
    .B2(_01518_),
    .A2(_00163_),
    .A1(net281));
 sg13g2_nor4_1 _10249_ (.A(_04136_),
    .B(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .C(_03637_),
    .D(_04035_),
    .Y(_04500_));
 sg13g2_a21o_1 _10250_ (.A2(_04499_),
    .A1(_04101_),
    .B1(_04500_),
    .X(_04501_));
 sg13g2_nand2_1 _10251_ (.Y(_04502_),
    .A(_04105_),
    .B(_04501_));
 sg13g2_o21ai_1 _10252_ (.B1(_04502_),
    .Y(_04503_),
    .A1(_04101_),
    .A2(_04473_));
 sg13g2_nor2b_1 _10253_ (.A(net281),
    .B_N(net232),
    .Y(_04504_));
 sg13g2_a21oi_1 _10254_ (.A1(_04136_),
    .A2(_03635_),
    .Y(_04505_),
    .B1(_04504_));
 sg13g2_nor2_1 _10255_ (.A(_04035_),
    .B(_04026_),
    .Y(_04506_));
 sg13g2_o21ai_1 _10256_ (.B1(_04506_),
    .Y(_04507_),
    .A1(_01519_),
    .A2(_04505_));
 sg13g2_a22oi_1 _10257_ (.Y(_04508_),
    .B1(_04507_),
    .B2(_04101_),
    .A2(_04115_),
    .A1(net235));
 sg13g2_or2_1 _10258_ (.X(_04509_),
    .B(net231),
    .A(net214));
 sg13g2_nor2_1 _10259_ (.A(net235),
    .B(_04509_),
    .Y(_04510_));
 sg13g2_nor2_1 _10260_ (.A(_04508_),
    .B(_04510_),
    .Y(_04511_));
 sg13g2_nor3_1 _10261_ (.A(_01520_),
    .B(_04503_),
    .C(_04511_),
    .Y(_04512_));
 sg13g2_nor2_1 _10262_ (.A(_04503_),
    .B(_04511_),
    .Y(_04513_));
 sg13g2_a21oi_1 _10263_ (.A1(_04433_),
    .A2(_04513_),
    .Y(_04514_),
    .B1(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ));
 sg13g2_nor3_1 _10264_ (.A(net47),
    .B(_04512_),
    .C(_04514_),
    .Y(_00647_));
 sg13g2_nor2_1 _10265_ (.A(_03629_),
    .B(_04430_),
    .Y(_04515_));
 sg13g2_nor2_1 _10266_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .B(_04433_),
    .Y(_04516_));
 sg13g2_o21ai_1 _10267_ (.B1(_04095_),
    .Y(_00648_),
    .A1(_04515_),
    .A2(_04516_));
 sg13g2_nand3_1 _10268_ (.B(_04430_),
    .C(_04433_),
    .A(_03903_),
    .Y(_04517_));
 sg13g2_o21ai_1 _10269_ (.B1(_04517_),
    .Y(_04518_),
    .A1(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .A2(_04433_));
 sg13g2_nand2_1 _10270_ (.Y(_00657_),
    .A(_04095_),
    .B(_04518_));
 sg13g2_nor2_1 _10271_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .B(_04433_),
    .Y(_04519_));
 sg13g2_nor3_1 _10272_ (.A(_03903_),
    .B(_04438_),
    .C(_04468_),
    .Y(_04520_));
 sg13g2_o21ai_1 _10273_ (.B1(_04095_),
    .Y(_00658_),
    .A1(_04519_),
    .A2(_04520_));
 sg13g2_nand2_1 _10274_ (.Y(_04521_),
    .A(net210),
    .B(_04141_));
 sg13g2_nand3b_1 _10275_ (.B(net230),
    .C(net233),
    .Y(_04522_),
    .A_N(net210));
 sg13g2_o21ai_1 _10276_ (.B1(_04522_),
    .Y(_04523_),
    .A1(_01235_),
    .A2(_04521_));
 sg13g2_o21ai_1 _10277_ (.B1(net210),
    .Y(_04524_),
    .A1(_01227_),
    .A2(_01235_));
 sg13g2_nand2_1 _10278_ (.Y(_04525_),
    .A(net71),
    .B(_04524_));
 sg13g2_a22oi_1 _10279_ (.Y(_04526_),
    .B1(_04525_),
    .B2(_01426_),
    .A2(_04523_),
    .A1(net71));
 sg13g2_nor2b_1 _10280_ (.A(_01523_),
    .B_N(_04145_),
    .Y(_04527_));
 sg13g2_a22oi_1 _10281_ (.Y(_04528_),
    .B1(_04526_),
    .B2(_04527_),
    .A2(_01523_),
    .A1(net230));
 sg13g2_nor3_1 _10282_ (.A(net215),
    .B(_03621_),
    .C(_04528_),
    .Y(_00692_));
 sg13g2_o21ai_1 _10283_ (.B1(net230),
    .Y(_04529_),
    .A1(net297),
    .A2(_01240_));
 sg13g2_nor2_1 _10284_ (.A(net233),
    .B(_04529_),
    .Y(_04530_));
 sg13g2_and2_1 _10285_ (.A(net233),
    .B(_04529_),
    .X(_04531_));
 sg13g2_a21oi_1 _10286_ (.A1(_04526_),
    .A2(_04530_),
    .Y(_04532_),
    .B1(_04531_));
 sg13g2_nor3_1 _10287_ (.A(net215),
    .B(_03621_),
    .C(_04532_),
    .Y(_00693_));
 sg13g2_inv_1 _10288_ (.Y(_04533_),
    .A(_00220_));
 sg13g2_inv_1 _10289_ (.Y(_04534_),
    .A(_01377_));
 sg13g2_nor2_1 _10290_ (.A(net300),
    .B(net278),
    .Y(_04535_));
 sg13g2_nand2_1 _10291_ (.Y(_04536_),
    .A(_04534_),
    .B(_04535_));
 sg13g2_nand3_1 _10292_ (.B(net300),
    .C(net278),
    .A(_01377_),
    .Y(_04537_));
 sg13g2_a21oi_1 _10293_ (.A1(_04536_),
    .A2(_04537_),
    .Y(_04538_),
    .B1(_01376_));
 sg13g2_or3_1 _10294_ (.A(_02861_),
    .B(_04192_),
    .C(_04538_),
    .X(_04539_));
 sg13g2_buf_1 _10295_ (.A(_04539_),
    .X(_04540_));
 sg13g2_buf_1 _10296_ (.A(_04540_),
    .X(_04541_));
 sg13g2_nor2_1 _10297_ (.A(_04533_),
    .B(net140),
    .Y(_00695_));
 sg13g2_and4_1 _10298_ (.A(_04187_),
    .B(_04179_),
    .C(_04188_),
    .D(_04183_),
    .X(_04542_));
 sg13g2_and2_1 _10299_ (.A(_04185_),
    .B(_04542_),
    .X(_04543_));
 sg13g2_buf_1 _10300_ (.A(_04543_),
    .X(_04544_));
 sg13g2_nand3_1 _10301_ (.B(\i_uart_rx.cycle_counter[8] ),
    .C(_04544_),
    .A(_04184_),
    .Y(_04545_));
 sg13g2_nor2_1 _10302_ (.A(_04189_),
    .B(_04545_),
    .Y(_04546_));
 sg13g2_xnor2_1 _10303_ (.Y(_04547_),
    .A(\i_uart_rx.cycle_counter[10] ),
    .B(_04546_));
 sg13g2_nor2_1 _10304_ (.A(net140),
    .B(_04547_),
    .Y(_00696_));
 sg13g2_xnor2_1 _10305_ (.Y(_04548_),
    .A(_04180_),
    .B(_04181_));
 sg13g2_nor2_1 _10306_ (.A(net140),
    .B(_04548_),
    .Y(_00697_));
 sg13g2_nand2_1 _10307_ (.Y(_04549_),
    .A(_04180_),
    .B(_04181_));
 sg13g2_xor2_1 _10308_ (.B(_04549_),
    .A(_04187_),
    .X(_04550_));
 sg13g2_nor2_1 _10309_ (.A(_04541_),
    .B(_04550_),
    .Y(_00698_));
 sg13g2_nand3_1 _10310_ (.B(_04181_),
    .C(_04187_),
    .A(_04180_),
    .Y(_04551_));
 sg13g2_xor2_1 _10311_ (.B(_04551_),
    .A(\i_uart_rx.cycle_counter[3] ),
    .X(_04552_));
 sg13g2_nor2_1 _10312_ (.A(net140),
    .B(_04552_),
    .Y(_00699_));
 sg13g2_nand2_1 _10313_ (.Y(_04553_),
    .A(_04187_),
    .B(_04183_));
 sg13g2_xor2_1 _10314_ (.B(_04553_),
    .A(_04188_),
    .X(_04554_));
 sg13g2_nor2_1 _10315_ (.A(net140),
    .B(_04554_),
    .Y(_00700_));
 sg13g2_nand3_1 _10316_ (.B(_04188_),
    .C(_04183_),
    .A(_04187_),
    .Y(_04555_));
 sg13g2_xor2_1 _10317_ (.B(_04555_),
    .A(_04179_),
    .X(_04556_));
 sg13g2_nor2_1 _10318_ (.A(net140),
    .B(_04556_),
    .Y(_00701_));
 sg13g2_xnor2_1 _10319_ (.Y(_04557_),
    .A(_04185_),
    .B(_04542_));
 sg13g2_nor2_1 _10320_ (.A(_04541_),
    .B(_04557_),
    .Y(_00702_));
 sg13g2_xnor2_1 _10321_ (.Y(_04558_),
    .A(_04184_),
    .B(_04544_));
 sg13g2_nor2_1 _10322_ (.A(net140),
    .B(_04558_),
    .Y(_00703_));
 sg13g2_inv_1 _10323_ (.Y(_04559_),
    .A(\i_uart_rx.cycle_counter[8] ));
 sg13g2_nand2_1 _10324_ (.Y(_04560_),
    .A(_04184_),
    .B(_04544_));
 sg13g2_xnor2_1 _10325_ (.Y(_04561_),
    .A(_04559_),
    .B(_04560_));
 sg13g2_nor2_1 _10326_ (.A(net140),
    .B(_04561_),
    .Y(_00704_));
 sg13g2_xnor2_1 _10327_ (.Y(_04562_),
    .A(_04189_),
    .B(_04545_));
 sg13g2_nor2_1 _10328_ (.A(_04540_),
    .B(_04562_),
    .Y(_00705_));
 sg13g2_inv_1 _10329_ (.Y(_04563_),
    .A(\i_uart_tx.cycle_counter[4] ));
 sg13g2_buf_1 _10330_ (.A(\i_uart_tx.cycle_counter[5] ),
    .X(_04564_));
 sg13g2_buf_1 _10331_ (.A(\i_uart_tx.cycle_counter[2] ),
    .X(_04565_));
 sg13g2_buf_1 _10332_ (.A(\i_uart_tx.cycle_counter[8] ),
    .X(_04566_));
 sg13g2_inv_1 _10333_ (.Y(_04567_),
    .A(\i_uart_tx.cycle_counter[9] ));
 sg13g2_or4_1 _10334_ (.A(\i_uart_tx.cycle_counter[7] ),
    .B(\i_uart_tx.cycle_counter[6] ),
    .C(_04566_),
    .D(_04567_),
    .X(_04568_));
 sg13g2_nand2_1 _10335_ (.Y(_04569_),
    .A(\i_uart_tx.cycle_counter[1] ),
    .B(\i_uart_tx.cycle_counter[0] ));
 sg13g2_nor4_1 _10336_ (.A(_04565_),
    .B(\i_uart_tx.cycle_counter[10] ),
    .C(_04568_),
    .D(_04569_),
    .Y(_04570_));
 sg13g2_and4_1 _10337_ (.A(\i_uart_tx.cycle_counter[3] ),
    .B(_04563_),
    .C(_04564_),
    .D(_04570_),
    .X(_04571_));
 sg13g2_buf_1 _10338_ (.A(_04571_),
    .X(_04572_));
 sg13g2_or2_1 _10339_ (.X(_04573_),
    .B(_04572_),
    .A(_02861_));
 sg13g2_buf_1 _10340_ (.A(_04573_),
    .X(_04574_));
 sg13g2_buf_1 _10341_ (.A(_04574_),
    .X(_04575_));
 sg13g2_nor2b_1 _10342_ (.A(net209),
    .B_N(_00219_),
    .Y(_04576_));
 sg13g2_a21oi_1 _10343_ (.A1(\i_uart_tx.cycle_counter[0] ),
    .A2(net209),
    .Y(_04577_),
    .B1(_04576_));
 sg13g2_nor2_1 _10344_ (.A(net139),
    .B(_04577_),
    .Y(_00721_));
 sg13g2_inv_1 _10345_ (.Y(_04578_),
    .A(\i_uart_tx.cycle_counter[7] ));
 sg13g2_nor2_1 _10346_ (.A(net209),
    .B(_04569_),
    .Y(_04579_));
 sg13g2_nand3_1 _10347_ (.B(\i_uart_tx.cycle_counter[3] ),
    .C(_04579_),
    .A(_04565_),
    .Y(_04580_));
 sg13g2_nor2_1 _10348_ (.A(_04563_),
    .B(_04580_),
    .Y(_04581_));
 sg13g2_nand3_1 _10349_ (.B(\i_uart_tx.cycle_counter[6] ),
    .C(_04581_),
    .A(_04564_),
    .Y(_04582_));
 sg13g2_nor2_1 _10350_ (.A(_04578_),
    .B(_04582_),
    .Y(_04583_));
 sg13g2_nand3_1 _10351_ (.B(\i_uart_tx.cycle_counter[9] ),
    .C(_04583_),
    .A(_04566_),
    .Y(_04584_));
 sg13g2_xor2_1 _10352_ (.B(_04584_),
    .A(\i_uart_tx.cycle_counter[10] ),
    .X(_04585_));
 sg13g2_nor2_1 _10353_ (.A(net139),
    .B(_04585_),
    .Y(_00722_));
 sg13g2_nor2b_1 _10354_ (.A(_01389_),
    .B_N(\i_uart_tx.cycle_counter[0] ),
    .Y(_04586_));
 sg13g2_xnor2_1 _10355_ (.Y(_04587_),
    .A(\i_uart_tx.cycle_counter[1] ),
    .B(_04586_));
 sg13g2_nor2_1 _10356_ (.A(net139),
    .B(_04587_),
    .Y(_00723_));
 sg13g2_xnor2_1 _10357_ (.Y(_04588_),
    .A(_04565_),
    .B(_04579_));
 sg13g2_nor2_1 _10358_ (.A(net139),
    .B(_04588_),
    .Y(_00724_));
 sg13g2_nand2_1 _10359_ (.Y(_04589_),
    .A(_04565_),
    .B(_04579_));
 sg13g2_xor2_1 _10360_ (.B(_04589_),
    .A(\i_uart_tx.cycle_counter[3] ),
    .X(_04590_));
 sg13g2_nor2_1 _10361_ (.A(net139),
    .B(_04590_),
    .Y(_00725_));
 sg13g2_xnor2_1 _10362_ (.Y(_04591_),
    .A(_04563_),
    .B(_04580_));
 sg13g2_nor2_1 _10363_ (.A(net139),
    .B(_04591_),
    .Y(_00726_));
 sg13g2_xnor2_1 _10364_ (.Y(_04592_),
    .A(_04564_),
    .B(_04581_));
 sg13g2_nor2_1 _10365_ (.A(net139),
    .B(_04592_),
    .Y(_00727_));
 sg13g2_nand2_1 _10366_ (.Y(_04593_),
    .A(_04564_),
    .B(_04581_));
 sg13g2_xor2_1 _10367_ (.B(_04593_),
    .A(\i_uart_tx.cycle_counter[6] ),
    .X(_04594_));
 sg13g2_nor2_1 _10368_ (.A(net139),
    .B(_04594_),
    .Y(_00728_));
 sg13g2_xnor2_1 _10369_ (.Y(_04595_),
    .A(_04578_),
    .B(_04582_));
 sg13g2_nor2_1 _10370_ (.A(_04575_),
    .B(_04595_),
    .Y(_00729_));
 sg13g2_xnor2_1 _10371_ (.Y(_04596_),
    .A(_04566_),
    .B(_04583_));
 sg13g2_nor2_1 _10372_ (.A(_04575_),
    .B(_04596_),
    .Y(_00730_));
 sg13g2_nand2_1 _10373_ (.Y(_04597_),
    .A(_04566_),
    .B(_04583_));
 sg13g2_xnor2_1 _10374_ (.Y(_04598_),
    .A(_04567_),
    .B(_04597_));
 sg13g2_nor2_1 _10375_ (.A(_04574_),
    .B(_04598_),
    .Y(_00731_));
 sg13g2_inv_1 _10376_ (.Y(_04599_),
    .A(_01597_));
 sg13g2_buf_1 _10377_ (.A(_04599_),
    .X(_04600_));
 sg13g2_buf_1 _10378_ (.A(_04600_),
    .X(_04601_));
 sg13g2_nor2b_1 _10379_ (.A(_01578_),
    .B_N(net295),
    .Y(_04602_));
 sg13g2_nand4_1 _10380_ (.B(_02180_),
    .C(_04301_),
    .A(_01567_),
    .Y(_04603_),
    .D(_04602_));
 sg13g2_buf_1 _10381_ (.A(_04603_),
    .X(_04604_));
 sg13g2_buf_1 _10382_ (.A(net138),
    .X(_04605_));
 sg13g2_nor2_1 _10383_ (.A(_01573_),
    .B(net126),
    .Y(_04606_));
 sg13g2_o21ai_1 _10384_ (.B1(_02199_),
    .Y(_04607_),
    .A1(net290),
    .A2(_02196_));
 sg13g2_nand3b_1 _10385_ (.B(_04298_),
    .C(_04607_),
    .Y(_04608_),
    .A_N(_04300_));
 sg13g2_buf_2 _10386_ (.A(_04608_),
    .X(_04609_));
 sg13g2_mux2_1 _10387_ (.A0(\i_debug_uart_tx.data_to_send[1] ),
    .A1(\i_debug_uart_tx.data_to_send[0] ),
    .S(_04609_),
    .X(_04610_));
 sg13g2_nor2b_1 _10388_ (.A(_04610_),
    .B_N(_04605_),
    .Y(_04611_));
 sg13g2_nor3_1 _10389_ (.A(net178),
    .B(_04606_),
    .C(_04611_),
    .Y(_00234_));
 sg13g2_nor2_1 _10390_ (.A(_01600_),
    .B(net126),
    .Y(_04612_));
 sg13g2_mux2_1 _10391_ (.A0(\i_debug_uart_tx.data_to_send[2] ),
    .A1(\i_debug_uart_tx.data_to_send[1] ),
    .S(_04609_),
    .X(_04613_));
 sg13g2_nor2b_1 _10392_ (.A(_04613_),
    .B_N(net126),
    .Y(_04614_));
 sg13g2_nor3_1 _10393_ (.A(_04601_),
    .B(_04612_),
    .C(_04614_),
    .Y(_00235_));
 sg13g2_nor2_1 _10394_ (.A(_01603_),
    .B(net126),
    .Y(_04615_));
 sg13g2_mux2_1 _10395_ (.A0(\i_debug_uart_tx.data_to_send[3] ),
    .A1(\i_debug_uart_tx.data_to_send[2] ),
    .S(_04609_),
    .X(_04616_));
 sg13g2_nor2b_1 _10396_ (.A(_04616_),
    .B_N(net138),
    .Y(_04617_));
 sg13g2_nor3_1 _10397_ (.A(net178),
    .B(_04615_),
    .C(_04617_),
    .Y(_00236_));
 sg13g2_nor2_1 _10398_ (.A(_01606_),
    .B(_04605_),
    .Y(_04618_));
 sg13g2_mux2_1 _10399_ (.A0(\i_debug_uart_tx.data_to_send[4] ),
    .A1(\i_debug_uart_tx.data_to_send[3] ),
    .S(_04609_),
    .X(_04619_));
 sg13g2_nor2b_1 _10400_ (.A(_04619_),
    .B_N(net138),
    .Y(_04620_));
 sg13g2_nor3_1 _10401_ (.A(net178),
    .B(_04618_),
    .C(_04620_),
    .Y(_00237_));
 sg13g2_nor2_1 _10402_ (.A(_01609_),
    .B(net126),
    .Y(_04621_));
 sg13g2_mux2_1 _10403_ (.A0(\i_debug_uart_tx.data_to_send[5] ),
    .A1(\i_debug_uart_tx.data_to_send[4] ),
    .S(_04609_),
    .X(_04622_));
 sg13g2_nor2b_1 _10404_ (.A(_04622_),
    .B_N(net138),
    .Y(_04623_));
 sg13g2_nor3_1 _10405_ (.A(net178),
    .B(_04621_),
    .C(_04623_),
    .Y(_00238_));
 sg13g2_nor2_1 _10406_ (.A(_01612_),
    .B(net126),
    .Y(_04624_));
 sg13g2_mux2_1 _10407_ (.A0(\i_debug_uart_tx.data_to_send[6] ),
    .A1(\i_debug_uart_tx.data_to_send[5] ),
    .S(_04609_),
    .X(_04625_));
 sg13g2_nor2b_1 _10408_ (.A(_04625_),
    .B_N(net138),
    .Y(_04626_));
 sg13g2_nor3_1 _10409_ (.A(net178),
    .B(_04624_),
    .C(_04626_),
    .Y(_00239_));
 sg13g2_nor2_1 _10410_ (.A(_01616_),
    .B(net126),
    .Y(_04627_));
 sg13g2_mux2_1 _10411_ (.A0(\i_debug_uart_tx.data_to_send[7] ),
    .A1(\i_debug_uart_tx.data_to_send[6] ),
    .S(_04609_),
    .X(_04628_));
 sg13g2_nor2b_1 _10412_ (.A(_04628_),
    .B_N(net138),
    .Y(_04629_));
 sg13g2_nor3_1 _10413_ (.A(_04600_),
    .B(_04627_),
    .C(_04629_),
    .Y(_00240_));
 sg13g2_or2_1 _10414_ (.X(_04630_),
    .B(net138),
    .A(_00201_));
 sg13g2_nand3_1 _10415_ (.B(net126),
    .C(_04609_),
    .A(\i_debug_uart_tx.data_to_send[7] ),
    .Y(_04631_));
 sg13g2_buf_1 _10416_ (.A(_04600_),
    .X(_04632_));
 sg13g2_a21oi_1 _10417_ (.A1(_04630_),
    .A2(_04631_),
    .Y(_00241_),
    .B1(net177));
 sg13g2_buf_1 _10418_ (.A(_04600_),
    .X(_04633_));
 sg13g2_nand2b_1 _10419_ (.Y(_04634_),
    .B(net180),
    .A_N(_04300_));
 sg13g2_inv_1 _10420_ (.Y(_04635_),
    .A(_02199_));
 sg13g2_nor2_1 _10421_ (.A(_04635_),
    .B(_02196_),
    .Y(_04636_));
 sg13g2_nand2b_1 _10422_ (.Y(_04637_),
    .B(net180),
    .A_N(_04636_));
 sg13g2_a22oi_1 _10423_ (.Y(_04638_),
    .B1(_04637_),
    .B2(net290),
    .A2(_04634_),
    .A1(net138));
 sg13g2_nand3_1 _10424_ (.B(net180),
    .C(_04604_),
    .A(_02198_),
    .Y(_04639_));
 sg13g2_o21ai_1 _10425_ (.B1(_04639_),
    .Y(_04640_),
    .A1(_02198_),
    .A2(_04638_));
 sg13g2_nor2_1 _10426_ (.A(net176),
    .B(_04640_),
    .Y(_00242_));
 sg13g2_o21ai_1 _10427_ (.B1(net180),
    .Y(_04641_),
    .A1(_02198_),
    .A2(_04636_));
 sg13g2_nor2_1 _10428_ (.A(net290),
    .B(_04639_),
    .Y(_04642_));
 sg13g2_a21oi_1 _10429_ (.A1(net290),
    .A2(_04641_),
    .Y(_04643_),
    .B1(_04642_));
 sg13g2_nor2_1 _10430_ (.A(net176),
    .B(_04643_),
    .Y(_00243_));
 sg13g2_nand3_1 _10431_ (.B(net290),
    .C(net180),
    .A(_02198_),
    .Y(_04644_));
 sg13g2_xor2_1 _10432_ (.B(_04644_),
    .A(_02196_),
    .X(_04645_));
 sg13g2_nor2_1 _10433_ (.A(net176),
    .B(_04645_),
    .Y(_00244_));
 sg13g2_nand2b_1 _10434_ (.Y(_04646_),
    .B(_02196_),
    .A_N(_02198_));
 sg13g2_nand3_1 _10435_ (.B(net180),
    .C(_04646_),
    .A(net290),
    .Y(_04647_));
 sg13g2_nand4_1 _10436_ (.B(_04635_),
    .C(_02196_),
    .A(_02195_),
    .Y(_04648_),
    .D(net180));
 sg13g2_nand2b_1 _10437_ (.Y(_04649_),
    .B(_04648_),
    .A_N(_04636_));
 sg13g2_a22oi_1 _10438_ (.Y(_04650_),
    .B1(_04649_),
    .B2(_02198_),
    .A2(_04647_),
    .A1(_02199_));
 sg13g2_nor2_1 _10439_ (.A(net176),
    .B(_04650_),
    .Y(_00245_));
 sg13g2_a21oi_1 _10440_ (.A1(_02199_),
    .A2(\i_debug_uart_tx.data_to_send[0] ),
    .Y(_04651_),
    .B1(_02200_));
 sg13g2_nor3_1 _10441_ (.A(_02199_),
    .B(\i_debug_uart_tx.data_to_send[0] ),
    .C(_02197_),
    .Y(_04652_));
 sg13g2_a21oi_1 _10442_ (.A1(_02197_),
    .A2(_04651_),
    .Y(_04653_),
    .B1(_04652_));
 sg13g2_buf_1 _10443_ (.A(net261),
    .X(_04654_));
 sg13g2_nand2b_1 _10444_ (.Y(_00246_),
    .B(net213),
    .A_N(_04653_));
 sg13g2_nor3_1 _10445_ (.A(\i_spi.bits_remaining[0] ),
    .B(\i_spi.bits_remaining[1] ),
    .C(\i_spi.bits_remaining[2] ),
    .Y(_04655_));
 sg13g2_nor2b_1 _10446_ (.A(_02870_),
    .B_N(_04655_),
    .Y(_04656_));
 sg13g2_nor2b_1 _10447_ (.A(_04656_),
    .B_N(_02874_),
    .Y(_04657_));
 sg13g2_nand2_1 _10448_ (.Y(_04658_),
    .A(_01245_),
    .B(_04657_));
 sg13g2_nand2_1 _10449_ (.Y(_04659_),
    .A(net283),
    .B(_04658_));
 sg13g2_and2_1 _10450_ (.A(_02885_),
    .B(_04659_),
    .X(_04660_));
 sg13g2_buf_1 _10451_ (.A(_04660_),
    .X(_04661_));
 sg13g2_nand2b_1 _10452_ (.Y(_04662_),
    .B(\i_spi.bits_remaining[0] ),
    .A_N(_04661_));
 sg13g2_nand2b_1 _10453_ (.Y(_04663_),
    .B(_04661_),
    .A_N(\i_spi.bits_remaining[0] ));
 sg13g2_a21oi_1 _10454_ (.A1(_02207_),
    .A2(_02869_),
    .Y(_04664_),
    .B1(net283));
 sg13g2_nand2b_1 _10455_ (.Y(_04665_),
    .B(_01614_),
    .A_N(_04664_));
 sg13g2_a21oi_1 _10456_ (.A1(_04662_),
    .A2(_04663_),
    .Y(_00247_),
    .B1(_04665_));
 sg13g2_xor2_1 _10457_ (.B(_04663_),
    .A(\i_spi.bits_remaining[1] ),
    .X(_04666_));
 sg13g2_nor2_1 _10458_ (.A(_04665_),
    .B(_04666_),
    .Y(_00248_));
 sg13g2_nor2_1 _10459_ (.A(\i_spi.bits_remaining[1] ),
    .B(_04663_),
    .Y(_04667_));
 sg13g2_xnor2_1 _10460_ (.Y(_04668_),
    .A(\i_spi.bits_remaining[2] ),
    .B(_04667_));
 sg13g2_nor2_1 _10461_ (.A(_04665_),
    .B(_04668_),
    .Y(_00249_));
 sg13g2_nand3_1 _10462_ (.B(_04655_),
    .C(_04659_),
    .A(_02870_),
    .Y(_04669_));
 sg13g2_or2_1 _10463_ (.X(_04670_),
    .B(_04655_),
    .A(_02870_));
 sg13g2_a21oi_1 _10464_ (.A1(_04669_),
    .A2(_04670_),
    .Y(_04671_),
    .B1(_02207_));
 sg13g2_nor2_1 _10465_ (.A(_02870_),
    .B(_04661_),
    .Y(_04672_));
 sg13g2_nor3_1 _10466_ (.A(_04600_),
    .B(_04671_),
    .C(_04672_),
    .Y(_00250_));
 sg13g2_a21oi_1 _10467_ (.A1(net208),
    .A2(_02186_),
    .Y(_04673_),
    .B1(net244));
 sg13g2_nand4_1 _10468_ (.B(_01246_),
    .C(_02874_),
    .A(_02866_),
    .Y(_04674_),
    .D(_04656_));
 sg13g2_inv_1 _10469_ (.Y(_04675_),
    .A(_04674_));
 sg13g2_nor3_1 _10470_ (.A(_04600_),
    .B(_04673_),
    .C(_04675_),
    .Y(_00251_));
 sg13g2_o21ai_1 _10471_ (.B1(_02866_),
    .Y(_04676_),
    .A1(_02872_),
    .A2(_02873_));
 sg13g2_inv_1 _10472_ (.Y(_04677_),
    .A(\i_spi.clock_count[0] ));
 sg13g2_mux2_1 _10473_ (.A0(_02867_),
    .A1(_04676_),
    .S(_04677_),
    .X(_04678_));
 sg13g2_nor2_1 _10474_ (.A(net176),
    .B(_04678_),
    .Y(_00252_));
 sg13g2_o21ai_1 _10475_ (.B1(_02882_),
    .Y(_04679_),
    .A1(\i_spi.clock_count[0] ),
    .A2(_02874_));
 sg13g2_nor3_1 _10476_ (.A(_04677_),
    .B(\i_spi.clock_count[1] ),
    .C(_04676_),
    .Y(_04680_));
 sg13g2_a21oi_1 _10477_ (.A1(\i_spi.clock_count[1] ),
    .A2(_04679_),
    .Y(_04681_),
    .B1(_04680_));
 sg13g2_nor2_1 _10478_ (.A(net176),
    .B(_04681_),
    .Y(_00253_));
 sg13g2_and3_1 _10479_ (.X(_04682_),
    .A(net208),
    .B(_02183_),
    .C(_02190_));
 sg13g2_buf_1 _10480_ (.A(_04682_),
    .X(_04683_));
 sg13g2_nand2b_1 _10481_ (.Y(_04684_),
    .B(\i_spi.clock_divider[0] ),
    .A_N(_04683_));
 sg13g2_nand2_1 _10482_ (.Y(_04685_),
    .A(_01573_),
    .B(_04683_));
 sg13g2_nand3_1 _10483_ (.B(_04684_),
    .C(_04685_),
    .A(net213),
    .Y(_00254_));
 sg13g2_nand2_1 _10484_ (.Y(_04686_),
    .A(_01600_),
    .B(_04683_));
 sg13g2_nand2b_1 _10485_ (.Y(_04687_),
    .B(\i_spi.clock_divider[1] ),
    .A_N(_04683_));
 sg13g2_a21oi_1 _10486_ (.A1(_04686_),
    .A2(_04687_),
    .Y(_00255_),
    .B1(net177));
 sg13g2_nand2_1 _10487_ (.Y(_04688_),
    .A(_01603_),
    .B(_04683_));
 sg13g2_nand2b_1 _10488_ (.Y(_04689_),
    .B(\i_spi.read_latency ),
    .A_N(_04683_));
 sg13g2_a21oi_1 _10489_ (.A1(_04688_),
    .A2(_04689_),
    .Y(_00265_),
    .B1(net177));
 sg13g2_nand2_1 _10490_ (.Y(_04690_),
    .A(_01246_),
    .B(_04657_));
 sg13g2_o21ai_1 _10491_ (.B1(_04690_),
    .Y(_04691_),
    .A1(_01246_),
    .A2(_02874_));
 sg13g2_nor2_1 _10492_ (.A(_02882_),
    .B(_01246_),
    .Y(_04692_));
 sg13g2_a22oi_1 _10493_ (.Y(_04693_),
    .B1(_04692_),
    .B2(_02869_),
    .A2(_04691_),
    .A1(net244));
 sg13g2_nor2_1 _10494_ (.A(net176),
    .B(_04693_),
    .Y(_00266_));
 sg13g2_nor2_1 _10495_ (.A(net244),
    .B(_02869_),
    .Y(_04694_));
 sg13g2_nand2_1 _10496_ (.Y(_04695_),
    .A(\i_spi.spi_select ),
    .B(_04674_));
 sg13g2_a21oi_1 _10497_ (.A1(\i_spi.end_txn_reg ),
    .A2(_04675_),
    .Y(_04696_),
    .B1(_04600_));
 sg13g2_o21ai_1 _10498_ (.B1(_04696_),
    .Y(_00268_),
    .A1(_04694_),
    .A2(_04695_));
 sg13g2_buf_1 _10499_ (.A(_03414_),
    .X(_04697_));
 sg13g2_buf_1 _10500_ (.A(net212),
    .X(_04698_));
 sg13g2_nor2_1 _10501_ (.A(_00212_),
    .B(net79),
    .Y(_04699_));
 sg13g2_nor2_1 _10502_ (.A(_01458_),
    .B(_03194_),
    .Y(_04700_));
 sg13g2_a22oi_1 _10503_ (.Y(_04701_),
    .B1(_04700_),
    .B2(_03158_),
    .A2(_03193_),
    .A1(net130));
 sg13g2_nand2_1 _10504_ (.Y(_04702_),
    .A(net90),
    .B(_04701_));
 sg13g2_and3_1 _10505_ (.X(_04703_),
    .A(_02909_),
    .B(_03507_),
    .C(_04702_));
 sg13g2_nor2b_1 _10506_ (.A(_02909_),
    .B_N(_01283_),
    .Y(_04704_));
 sg13g2_nor3_1 _10507_ (.A(_03515_),
    .B(_04703_),
    .C(_04704_),
    .Y(_04705_));
 sg13g2_nor3_1 _10508_ (.A(net199),
    .B(_04699_),
    .C(_04705_),
    .Y(_00269_));
 sg13g2_o21ai_1 _10509_ (.B1(_03195_),
    .Y(_04706_),
    .A1(_03159_),
    .A2(_03505_));
 sg13g2_inv_1 _10510_ (.Y(_04707_),
    .A(net122));
 sg13g2_a221oi_1 _10511_ (.B2(_04707_),
    .C1(_02920_),
    .B1(_04700_),
    .A1(_01332_),
    .Y(_04708_),
    .A2(_03193_));
 sg13g2_a21oi_1 _10512_ (.A1(_02920_),
    .A2(_04706_),
    .Y(_04709_),
    .B1(_04708_));
 sg13g2_nor3_1 _10513_ (.A(_01553_),
    .B(_03530_),
    .C(_04709_),
    .Y(_04710_));
 sg13g2_xor2_1 _10514_ (.B(_01284_),
    .A(_01283_),
    .X(_04711_));
 sg13g2_and2_1 _10515_ (.A(_01553_),
    .B(_04711_),
    .X(_04712_));
 sg13g2_nor2_1 _10516_ (.A(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .B(_04709_),
    .Y(_04713_));
 sg13g2_nor2_1 _10517_ (.A(_03530_),
    .B(_04713_),
    .Y(_04714_));
 sg13g2_o21ai_1 _10518_ (.B1(net241),
    .Y(_04715_),
    .A1(_01284_),
    .A2(_04714_));
 sg13g2_nor3_1 _10519_ (.A(_04710_),
    .B(_04712_),
    .C(_04715_),
    .Y(_00270_));
 sg13g2_buf_1 _10520_ (.A(net212),
    .X(_04716_));
 sg13g2_and2_1 _10521_ (.A(_02904_),
    .B(_02909_),
    .X(_04717_));
 sg13g2_buf_2 _10522_ (.A(_04717_),
    .X(_04718_));
 sg13g2_a22oi_1 _10523_ (.Y(_04719_),
    .B1(_04700_),
    .B2(_01479_),
    .A2(_03193_),
    .A1(_01339_));
 sg13g2_inv_1 _10524_ (.Y(_04720_),
    .A(_04719_));
 sg13g2_o21ai_1 _10525_ (.B1(_01553_),
    .Y(_04721_),
    .A1(_01283_),
    .A2(_01284_));
 sg13g2_o21ai_1 _10526_ (.B1(_04721_),
    .Y(_04722_),
    .A1(_01553_),
    .A2(_02909_));
 sg13g2_a22oi_1 _10527_ (.Y(_04723_),
    .B1(_04722_),
    .B2(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .A2(_04720_),
    .A1(_04718_));
 sg13g2_nor2_1 _10528_ (.A(net198),
    .B(_04723_),
    .Y(_00271_));
 sg13g2_and2_1 _10529_ (.A(_03470_),
    .B(net282),
    .X(_00276_));
 sg13g2_nor2_1 _10530_ (.A(net198),
    .B(_03115_),
    .Y(_00277_));
 sg13g2_xnor2_1 _10531_ (.Y(_04724_),
    .A(net202),
    .B(_00961_));
 sg13g2_nor2_1 _10532_ (.A(net198),
    .B(_04724_),
    .Y(_00278_));
 sg13g2_nor2_2 _10533_ (.A(_03014_),
    .B(net134),
    .Y(_04725_));
 sg13g2_a22oi_1 _10534_ (.Y(_04726_),
    .B1(_04725_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A2(net134),
    .A1(\addr[24] ));
 sg13g2_nor2_1 _10535_ (.A(net198),
    .B(_04726_),
    .Y(_00295_));
 sg13g2_a22oi_1 _10536_ (.Y(_04727_),
    .B1(_04725_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .A2(net134),
    .A1(\addr[25] ));
 sg13g2_nor2_1 _10537_ (.A(net198),
    .B(_04727_),
    .Y(_00296_));
 sg13g2_a22oi_1 _10538_ (.Y(_04728_),
    .B1(_04725_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A2(_01655_),
    .A1(\addr[26] ));
 sg13g2_nor2_1 _10539_ (.A(_04716_),
    .B(_04728_),
    .Y(_00297_));
 sg13g2_a22oi_1 _10540_ (.Y(_04729_),
    .B1(_04725_),
    .B2(_02445_),
    .A2(net134),
    .A1(\addr[27] ));
 sg13g2_nor2_1 _10541_ (.A(_04716_),
    .B(_04729_),
    .Y(_00298_));
 sg13g2_nor2_1 _10542_ (.A(net168),
    .B(_04321_),
    .Y(_04730_));
 sg13g2_a21oi_1 _10543_ (.A1(\i_tinyqv.cpu.data_ready_core ),
    .A2(net168),
    .Y(_04731_),
    .B1(_04730_));
 sg13g2_nor2_1 _10544_ (.A(net198),
    .B(_04731_),
    .Y(_00341_));
 sg13g2_nand2_1 _10545_ (.Y(_04732_),
    .A(_01196_),
    .B(_01652_));
 sg13g2_nor2_1 _10546_ (.A(_01263_),
    .B(_04732_),
    .Y(_04733_));
 sg13g2_and2_1 _10547_ (.A(_01196_),
    .B(_01652_),
    .X(_04734_));
 sg13g2_nor3_1 _10548_ (.A(_01232_),
    .B(_01565_),
    .C(_04734_),
    .Y(_04735_));
 sg13g2_o21ai_1 _10549_ (.B1(net241),
    .Y(_00343_),
    .A1(_04733_),
    .A2(_04735_));
 sg13g2_nor2_1 _10550_ (.A(_02250_),
    .B(_04732_),
    .Y(_04736_));
 sg13g2_nor3_1 _10551_ (.A(\i_tinyqv.cpu.data_write_n[1] ),
    .B(_01565_),
    .C(_04734_),
    .Y(_04737_));
 sg13g2_o21ai_1 _10552_ (.B1(net241),
    .Y(_00344_),
    .A1(_04736_),
    .A2(_04737_));
 sg13g2_nand2_1 _10553_ (.Y(_04738_),
    .A(net160),
    .B(_02379_));
 sg13g2_a21oi_1 _10554_ (.A1(_01210_),
    .A2(_01223_),
    .Y(_04739_),
    .B1(_04738_));
 sg13g2_a21oi_1 _10555_ (.A1(_01646_),
    .A2(net168),
    .Y(_04740_),
    .B1(_04739_));
 sg13g2_nor2_1 _10556_ (.A(net198),
    .B(_04740_),
    .Y(_00345_));
 sg13g2_a21oi_1 _10557_ (.A1(_01646_),
    .A2(net160),
    .Y(_04741_),
    .B1(_01647_));
 sg13g2_nor3_1 _10558_ (.A(net199),
    .B(_01369_),
    .C(_04741_),
    .Y(_00346_));
 sg13g2_nor2_1 _10559_ (.A(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .B(net157),
    .Y(_04742_));
 sg13g2_nor2b_1 _10560_ (.A(_04742_),
    .B_N(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .Y(_04743_));
 sg13g2_buf_1 _10561_ (.A(_04743_),
    .X(_04744_));
 sg13g2_nand4_1 _10562_ (.B(_02366_),
    .C(_02644_),
    .A(_02733_),
    .Y(_04745_),
    .D(_04744_));
 sg13g2_nor2_1 _10563_ (.A(net198),
    .B(_04745_),
    .Y(_00347_));
 sg13g2_nor3_1 _10564_ (.A(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .B(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .C(net157),
    .Y(_04746_));
 sg13g2_nor3_1 _10565_ (.A(net199),
    .B(_04744_),
    .C(_04746_),
    .Y(_00348_));
 sg13g2_buf_1 _10566_ (.A(net212),
    .X(_04747_));
 sg13g2_xnor2_1 _10567_ (.Y(_04748_),
    .A(_02644_),
    .B(_04744_));
 sg13g2_nor2_1 _10568_ (.A(net197),
    .B(_04748_),
    .Y(_00349_));
 sg13g2_nand2_1 _10569_ (.Y(_04749_),
    .A(_02644_),
    .B(_04744_));
 sg13g2_xor2_1 _10570_ (.B(_04749_),
    .A(_02733_),
    .X(_04750_));
 sg13g2_nor2_1 _10571_ (.A(_04747_),
    .B(_04750_),
    .Y(_00350_));
 sg13g2_nand3_1 _10572_ (.B(_02644_),
    .C(_04744_),
    .A(_02733_),
    .Y(_04751_));
 sg13g2_xor2_1 _10573_ (.B(_04751_),
    .A(_02366_),
    .X(_04752_));
 sg13g2_nor2_1 _10574_ (.A(_04747_),
    .B(_04752_),
    .Y(_00351_));
 sg13g2_inv_1 _10575_ (.Y(_04753_),
    .A(\i_tinyqv.cpu.i_core.i_instrret.data[2] ));
 sg13g2_and2_1 _10576_ (.A(_00214_),
    .B(net157),
    .X(_04754_));
 sg13g2_a21oi_2 _10577_ (.B1(_04754_),
    .Y(_04755_),
    .A2(net173),
    .A1(_00215_));
 sg13g2_nand3_1 _10578_ (.B(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .C(_04755_),
    .A(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .Y(_04756_));
 sg13g2_nor2_1 _10579_ (.A(_04753_),
    .B(_04756_),
    .Y(_04757_));
 sg13g2_and3_1 _10580_ (.X(_00352_),
    .A(net241),
    .B(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .C(_04757_));
 sg13g2_xnor2_1 _10581_ (.Y(_04758_),
    .A(_02368_),
    .B(_04755_));
 sg13g2_nor2_1 _10582_ (.A(net197),
    .B(_04758_),
    .Y(_00353_));
 sg13g2_nand2_1 _10583_ (.Y(_04759_),
    .A(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .B(_04755_));
 sg13g2_xor2_1 _10584_ (.B(_04759_),
    .A(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .X(_04760_));
 sg13g2_nor2_1 _10585_ (.A(net197),
    .B(_04760_),
    .Y(_00354_));
 sg13g2_xnor2_1 _10586_ (.Y(_04761_),
    .A(_04753_),
    .B(_04756_));
 sg13g2_nor2_1 _10587_ (.A(net197),
    .B(_04761_),
    .Y(_00355_));
 sg13g2_xnor2_1 _10588_ (.Y(_04762_),
    .A(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .B(_04757_));
 sg13g2_nor2_1 _10589_ (.A(net197),
    .B(_04762_),
    .Y(_00356_));
 sg13g2_buf_1 _10590_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .X(_04763_));
 sg13g2_nor4_1 _10591_ (.A(_04763_),
    .B(_00924_),
    .C(_00975_),
    .D(_01096_),
    .Y(_04764_));
 sg13g2_nor2_1 _10592_ (.A(_04328_),
    .B(_04764_),
    .Y(_04765_));
 sg13g2_nand2_1 _10593_ (.Y(_04766_),
    .A(_01374_),
    .B(_01381_));
 sg13g2_nand3_1 _10594_ (.B(_04766_),
    .C(net209),
    .A(_01390_),
    .Y(_04767_));
 sg13g2_nand2_1 _10595_ (.Y(_04768_),
    .A(_01371_),
    .B(_04767_));
 sg13g2_nand3_1 _10596_ (.B(_01372_),
    .C(_04768_),
    .A(_04763_),
    .Y(_04769_));
 sg13g2_o21ai_1 _10597_ (.B1(_03470_),
    .Y(_04770_),
    .A1(\i_tinyqv.cpu.i_core.mcause[0] ),
    .A2(_04322_));
 sg13g2_a21oi_1 _10598_ (.A1(_04765_),
    .A2(_04769_),
    .Y(_00362_),
    .B1(_04770_));
 sg13g2_or2_1 _10599_ (.X(_04771_),
    .B(_01391_),
    .A(_01373_));
 sg13g2_nor2_1 _10600_ (.A(\i_tinyqv.cpu.i_core.mcause[1] ),
    .B(_04261_),
    .Y(_04772_));
 sg13g2_a221oi_1 _10601_ (.B2(_03124_),
    .C1(_04698_),
    .B1(_04772_),
    .A1(_04261_),
    .Y(_00363_),
    .A2(_04771_));
 sg13g2_buf_1 _10602_ (.A(net212),
    .X(_04773_));
 sg13g2_and2_1 _10603_ (.A(_01049_),
    .B(_04322_),
    .X(_04774_));
 sg13g2_a21oi_1 _10604_ (.A1(\i_tinyqv.cpu.i_core.mcause[3] ),
    .A2(_04328_),
    .Y(_04775_),
    .B1(_04774_));
 sg13g2_nor3_1 _10605_ (.A(net196),
    .B(_04765_),
    .C(_04775_),
    .Y(_00364_));
 sg13g2_nand2_1 _10606_ (.Y(_04776_),
    .A(\i_tinyqv.cpu.i_core.mcause[4] ),
    .B(_04328_));
 sg13g2_nand2_1 _10607_ (.Y(_04777_),
    .A(_04763_),
    .B(_04322_));
 sg13g2_buf_1 _10608_ (.A(net212),
    .X(_04778_));
 sg13g2_a21oi_1 _10609_ (.A1(_04776_),
    .A2(_04777_),
    .Y(_00365_),
    .B1(_04778_));
 sg13g2_nor2_1 _10610_ (.A(net168),
    .B(_04745_),
    .Y(_04779_));
 sg13g2_nand2_1 _10611_ (.Y(_04780_),
    .A(_00218_),
    .B(_04779_));
 sg13g2_o21ai_1 _10612_ (.B1(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .Y(_04781_),
    .A1(net168),
    .A2(_04745_));
 sg13g2_a21oi_1 _10613_ (.A1(_04780_),
    .A2(_04781_),
    .Y(_00402_),
    .B1(net195));
 sg13g2_nand2_1 _10614_ (.Y(_04782_),
    .A(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .B(_04779_));
 sg13g2_xor2_1 _10615_ (.B(_04782_),
    .A(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .X(_04783_));
 sg13g2_nor2_1 _10616_ (.A(net197),
    .B(_04783_),
    .Y(_00403_));
 sg13g2_nand3_1 _10617_ (.B(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .C(_04779_),
    .A(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .Y(_04784_));
 sg13g2_xor2_1 _10618_ (.B(_04784_),
    .A(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .X(_04785_));
 sg13g2_nor2_1 _10619_ (.A(net197),
    .B(_04785_),
    .Y(_00404_));
 sg13g2_and2_1 _10620_ (.A(_01286_),
    .B(_01553_),
    .X(_04786_));
 sg13g2_buf_1 _10621_ (.A(_04786_),
    .X(_04787_));
 sg13g2_nor2_1 _10622_ (.A(_04787_),
    .B(_03417_),
    .Y(_04788_));
 sg13g2_buf_1 _10623_ (.A(_04788_),
    .X(_04789_));
 sg13g2_buf_1 _10624_ (.A(_01200_),
    .X(_04790_));
 sg13g2_buf_1 _10625_ (.A(net175),
    .X(_04791_));
 sg13g2_nor2_1 _10626_ (.A(net162),
    .B(_03042_),
    .Y(_04792_));
 sg13g2_a21oi_1 _10627_ (.A1(net162),
    .A2(_03925_),
    .Y(_04793_),
    .B1(_04792_));
 sg13g2_buf_1 _10628_ (.A(net83),
    .X(_04794_));
 sg13g2_buf_1 _10629_ (.A(net83),
    .X(_04795_));
 sg13g2_buf_1 _10630_ (.A(net81),
    .X(_04796_));
 sg13g2_buf_1 _10631_ (.A(net81),
    .X(_04797_));
 sg13g2_nor3_1 _10632_ (.A(net85),
    .B(net74),
    .C(_02750_),
    .Y(_04798_));
 sg13g2_a21oi_1 _10633_ (.A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .A2(net75),
    .Y(_04799_),
    .B1(_04798_));
 sg13g2_nor2_1 _10634_ (.A(net76),
    .B(_04799_),
    .Y(_04800_));
 sg13g2_a221oi_1 _10635_ (.B2(net77),
    .C1(_04800_),
    .B1(_04793_),
    .A1(net312),
    .Y(_04801_),
    .A2(net66));
 sg13g2_nor2_1 _10636_ (.A(net197),
    .B(_04801_),
    .Y(_00533_));
 sg13g2_nand2_1 _10637_ (.Y(_04802_),
    .A(_01554_),
    .B(_03473_));
 sg13g2_buf_1 _10638_ (.A(_04802_),
    .X(_04803_));
 sg13g2_nor2_1 _10639_ (.A(net252),
    .B(net58),
    .Y(_04804_));
 sg13g2_buf_1 _10640_ (.A(_03473_),
    .X(_04805_));
 sg13g2_buf_1 _10641_ (.A(net81),
    .X(_04806_));
 sg13g2_mux2_1 _10642_ (.A0(_02621_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .S(net73),
    .X(_04807_));
 sg13g2_buf_1 _10643_ (.A(_03415_),
    .X(_04808_));
 sg13g2_buf_1 _10644_ (.A(net78),
    .X(_04809_));
 sg13g2_buf_1 _10645_ (.A(_01262_),
    .X(_04810_));
 sg13g2_buf_1 _10646_ (.A(_04810_),
    .X(_04811_));
 sg13g2_nor2_1 _10647_ (.A(net174),
    .B(_03740_),
    .Y(_04812_));
 sg13g2_a21oi_1 _10648_ (.A1(net161),
    .A2(_03025_),
    .Y(_04813_),
    .B1(_04812_));
 sg13g2_nor2_1 _10649_ (.A(net78),
    .B(_04813_),
    .Y(_04814_));
 sg13g2_a221oi_1 _10650_ (.B2(net72),
    .C1(_04814_),
    .B1(_04807_),
    .A1(net82),
    .Y(_04815_),
    .A2(net65));
 sg13g2_nor3_1 _10651_ (.A(net196),
    .B(_04804_),
    .C(_04815_),
    .Y(_00534_));
 sg13g2_nor2_1 _10652_ (.A(net254),
    .B(net58),
    .Y(_04816_));
 sg13g2_mux2_1 _10653_ (.A0(_02711_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .S(net73),
    .X(_04817_));
 sg13g2_nor2_1 _10654_ (.A(net174),
    .B(_03753_),
    .Y(_04818_));
 sg13g2_a21oi_1 _10655_ (.A1(net161),
    .A2(_03026_),
    .Y(_04819_),
    .B1(_04818_));
 sg13g2_nor2_1 _10656_ (.A(net78),
    .B(_04819_),
    .Y(_04820_));
 sg13g2_a221oi_1 _10657_ (.B2(net72),
    .C1(_04820_),
    .B1(_04817_),
    .A1(net82),
    .Y(_04821_),
    .A2(net65));
 sg13g2_nor3_1 _10658_ (.A(_04773_),
    .B(_04816_),
    .C(_04821_),
    .Y(_00535_));
 sg13g2_buf_1 _10659_ (.A(net212),
    .X(_04822_));
 sg13g2_xnor2_1 _10660_ (.Y(_04823_),
    .A(_02306_),
    .B(_03776_));
 sg13g2_nand2_1 _10661_ (.Y(_04824_),
    .A(net175),
    .B(_04823_));
 sg13g2_o21ai_1 _10662_ (.B1(_04824_),
    .Y(_04825_),
    .A1(net175),
    .A2(_03027_));
 sg13g2_inv_1 _10663_ (.Y(_04826_),
    .A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_mux2_1 _10664_ (.A0(_02746_),
    .A1(_04826_),
    .S(net81),
    .X(_04827_));
 sg13g2_mux2_1 _10665_ (.A0(_04825_),
    .A1(_04827_),
    .S(_03415_),
    .X(_04828_));
 sg13g2_nand2_1 _10666_ (.Y(_04829_),
    .A(_04802_),
    .B(_04828_));
 sg13g2_o21ai_1 _10667_ (.B1(_04829_),
    .Y(_04830_),
    .A1(net253),
    .A2(net58));
 sg13g2_nor2_1 _10668_ (.A(net194),
    .B(_04830_),
    .Y(_00536_));
 sg13g2_nand2b_1 _10669_ (.Y(_04831_),
    .B(_04810_),
    .A_N(_03028_));
 sg13g2_o21ai_1 _10670_ (.B1(_04831_),
    .Y(_04832_),
    .A1(net174),
    .A2(_03788_));
 sg13g2_mux2_1 _10671_ (.A0(_02312_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .S(_03471_),
    .X(_04833_));
 sg13g2_nor2_1 _10672_ (.A(net83),
    .B(_04833_),
    .Y(_04834_));
 sg13g2_a221oi_1 _10673_ (.B2(net83),
    .C1(_04834_),
    .B1(_04832_),
    .A1(net82),
    .Y(_04835_),
    .A2(_03473_));
 sg13g2_a21oi_1 _10674_ (.A1(net305),
    .A2(net66),
    .Y(_04836_),
    .B1(_04835_));
 sg13g2_nor2_1 _10675_ (.A(net194),
    .B(_04836_),
    .Y(_00537_));
 sg13g2_nand2b_1 _10676_ (.Y(_04837_),
    .B(net81),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_o21ai_1 _10677_ (.B1(_04837_),
    .Y(_04838_),
    .A1(net74),
    .A2(_02639_));
 sg13g2_nand2_1 _10678_ (.Y(_04839_),
    .A(_01262_),
    .B(_03029_));
 sg13g2_o21ai_1 _10679_ (.B1(_04839_),
    .Y(_04840_),
    .A1(net174),
    .A2(_03810_));
 sg13g2_nor2_1 _10680_ (.A(net78),
    .B(_04840_),
    .Y(_04841_));
 sg13g2_a221oi_1 _10681_ (.B2(net78),
    .C1(_04841_),
    .B1(_04838_),
    .A1(net85),
    .Y(_04842_),
    .A2(_03473_));
 sg13g2_a21oi_1 _10682_ (.A1(net308),
    .A2(net66),
    .Y(_04843_),
    .B1(_04842_));
 sg13g2_nor2_1 _10683_ (.A(net194),
    .B(_04843_),
    .Y(_00538_));
 sg13g2_nand2b_1 _10684_ (.Y(_04844_),
    .B(_03471_),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_o21ai_1 _10685_ (.B1(_04844_),
    .Y(_04845_),
    .A1(net74),
    .A2(_02723_));
 sg13g2_nand2_1 _10686_ (.Y(_04846_),
    .A(_01262_),
    .B(_03030_));
 sg13g2_o21ai_1 _10687_ (.B1(_04846_),
    .Y(_04847_),
    .A1(net174),
    .A2(_03825_));
 sg13g2_nor2_1 _10688_ (.A(_03415_),
    .B(_04847_),
    .Y(_04848_));
 sg13g2_a221oi_1 _10689_ (.B2(net78),
    .C1(_04848_),
    .B1(_04845_),
    .A1(net85),
    .Y(_04849_),
    .A2(_03473_));
 sg13g2_a21oi_1 _10690_ (.A1(net286),
    .A2(net66),
    .Y(_04850_),
    .B1(_04849_));
 sg13g2_nor2_1 _10691_ (.A(net194),
    .B(_04850_),
    .Y(_00539_));
 sg13g2_nor2_1 _10692_ (.A(_00859_),
    .B(_04802_),
    .Y(_04851_));
 sg13g2_mux2_1 _10693_ (.A0(_03032_),
    .A1(_03836_),
    .S(_04791_),
    .X(_04852_));
 sg13g2_nor2_1 _10694_ (.A(net72),
    .B(_04852_),
    .Y(_04853_));
 sg13g2_nand2_1 _10695_ (.Y(_04854_),
    .A(_04787_),
    .B(_02758_));
 sg13g2_mux2_1 _10696_ (.A0(_04854_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .S(_04796_),
    .X(_04855_));
 sg13g2_nor2_1 _10697_ (.A(_04794_),
    .B(_04855_),
    .Y(_04856_));
 sg13g2_nor4_1 _10698_ (.A(net212),
    .B(_04851_),
    .C(_04853_),
    .D(_04856_),
    .Y(_00540_));
 sg13g2_xor2_1 _10699_ (.B(_03868_),
    .A(_01138_),
    .X(_04857_));
 sg13g2_nor2_1 _10700_ (.A(net162),
    .B(_03035_),
    .Y(_04858_));
 sg13g2_a21oi_1 _10701_ (.A1(net162),
    .A2(_04857_),
    .Y(_04859_),
    .B1(_04858_));
 sg13g2_nor2_1 _10702_ (.A(net72),
    .B(_04859_),
    .Y(_04860_));
 sg13g2_a21oi_1 _10703_ (.A1(_04787_),
    .A2(_02305_),
    .Y(_04861_),
    .B1(net75));
 sg13g2_a221oi_1 _10704_ (.B2(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .C1(_04861_),
    .B1(net75),
    .A1(net160),
    .Y(_04862_),
    .A2(_01279_));
 sg13g2_o21ai_1 _10705_ (.B1(net241),
    .Y(_04863_),
    .A1(_01138_),
    .A2(net58));
 sg13g2_nor3_1 _10706_ (.A(_04860_),
    .B(_04862_),
    .C(_04863_),
    .Y(_00541_));
 sg13g2_nand2_1 _10707_ (.Y(_04864_),
    .A(_04787_),
    .B(_02634_));
 sg13g2_nand2b_1 _10708_ (.Y(_04865_),
    .B(net75),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_o21ai_1 _10709_ (.B1(_04865_),
    .Y(_04866_),
    .A1(net75),
    .A2(_04864_));
 sg13g2_nand2b_1 _10710_ (.Y(_04867_),
    .B(net162),
    .A_N(_03878_));
 sg13g2_a21oi_1 _10711_ (.A1(net161),
    .A2(_03036_),
    .Y(_04868_),
    .B1(net72));
 sg13g2_o21ai_1 _10712_ (.B1(_01282_),
    .Y(_04869_),
    .A1(_00990_),
    .A2(_04803_));
 sg13g2_a221oi_1 _10713_ (.B2(_04868_),
    .C1(_04869_),
    .B1(_04867_),
    .A1(net72),
    .Y(_00542_),
    .A2(_04866_));
 sg13g2_nand2b_1 _10714_ (.Y(_04870_),
    .B(_04796_),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_nand3b_1 _10715_ (.B(_02721_),
    .C(_04787_),
    .Y(_04871_),
    .A_N(net75));
 sg13g2_nand3_1 _10716_ (.B(_04870_),
    .C(_04871_),
    .A(net72),
    .Y(_04872_));
 sg13g2_xnor2_1 _10717_ (.Y(_04873_),
    .A(_02719_),
    .B(_03893_));
 sg13g2_nand2_1 _10718_ (.Y(_04874_),
    .A(net161),
    .B(_03037_));
 sg13g2_o21ai_1 _10719_ (.B1(_04874_),
    .Y(_04875_),
    .A1(net161),
    .A2(_04873_));
 sg13g2_nand2_1 _10720_ (.Y(_04876_),
    .A(net77),
    .B(_04875_));
 sg13g2_a221oi_1 _10721_ (.B2(_04876_),
    .C1(_04698_),
    .B1(_04872_),
    .A1(_02719_),
    .Y(_00543_),
    .A2(net66));
 sg13g2_nor2_1 _10722_ (.A(net175),
    .B(_03044_),
    .Y(_04877_));
 sg13g2_a21oi_1 _10723_ (.A1(net162),
    .A2(_03936_),
    .Y(_04878_),
    .B1(_04877_));
 sg13g2_nor4_1 _10724_ (.A(_01554_),
    .B(net81),
    .C(_02286_),
    .D(_02287_),
    .Y(_04879_));
 sg13g2_a21oi_1 _10725_ (.A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .A2(_04806_),
    .Y(_04880_),
    .B1(_04879_));
 sg13g2_nor2_1 _10726_ (.A(net76),
    .B(_04880_),
    .Y(_04881_));
 sg13g2_a221oi_1 _10727_ (.B2(net77),
    .C1(_04881_),
    .B1(_04878_),
    .A1(net303),
    .Y(_04882_),
    .A2(net66));
 sg13g2_nor2_1 _10728_ (.A(net194),
    .B(_04882_),
    .Y(_00544_));
 sg13g2_nand2b_1 _10729_ (.Y(_04883_),
    .B(net75),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_or3_1 _10730_ (.A(net85),
    .B(net73),
    .C(_02761_),
    .X(_04884_));
 sg13g2_a21oi_1 _10731_ (.A1(_04883_),
    .A2(_04884_),
    .Y(_04885_),
    .B1(_04794_));
 sg13g2_nand4_1 _10732_ (.B(_03304_),
    .C(net175),
    .A(_02719_),
    .Y(_04886_),
    .D(_03908_));
 sg13g2_o21ai_1 _10733_ (.B1(_04886_),
    .Y(_04887_),
    .A1(net175),
    .A2(_03038_));
 sg13g2_a21oi_1 _10734_ (.A1(net76),
    .A2(_04887_),
    .Y(_04888_),
    .B1(_04697_));
 sg13g2_o21ai_1 _10735_ (.B1(_04888_),
    .Y(_04889_),
    .A1(\i_tinyqv.cpu.instr_data_start[23] ),
    .A2(_04802_));
 sg13g2_and2_1 _10736_ (.A(_03304_),
    .B(_03892_),
    .X(_04890_));
 sg13g2_o21ai_1 _10737_ (.B1(_03892_),
    .Y(_04891_),
    .A1(_02719_),
    .A2(_03304_));
 sg13g2_mux2_1 _10738_ (.A0(_04890_),
    .A1(_04891_),
    .S(_03908_),
    .X(_04892_));
 sg13g2_and2_1 _10739_ (.A(_03892_),
    .B(_03908_),
    .X(_04893_));
 sg13g2_nor3_1 _10740_ (.A(_00760_),
    .B(_03910_),
    .C(_04893_),
    .Y(_04894_));
 sg13g2_nor4_1 _10741_ (.A(net161),
    .B(net72),
    .C(_04892_),
    .D(_04894_),
    .Y(_04895_));
 sg13g2_nor3_1 _10742_ (.A(_04885_),
    .B(_04889_),
    .C(_04895_),
    .Y(_00545_));
 sg13g2_nor2_1 _10743_ (.A(net175),
    .B(_03047_),
    .Y(_04896_));
 sg13g2_a21oi_1 _10744_ (.A1(net162),
    .A2(_03945_),
    .Y(_04897_),
    .B1(_04896_));
 sg13g2_nor3_1 _10745_ (.A(net85),
    .B(net74),
    .C(_02626_),
    .Y(_04898_));
 sg13g2_a21oi_1 _10746_ (.A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .A2(net73),
    .Y(_04899_),
    .B1(_04898_));
 sg13g2_nor2_1 _10747_ (.A(net76),
    .B(_04899_),
    .Y(_04900_));
 sg13g2_a221oi_1 _10748_ (.B2(net77),
    .C1(_04900_),
    .B1(_04897_),
    .A1(net256),
    .Y(_04901_),
    .A2(_04789_));
 sg13g2_nor2_1 _10749_ (.A(net194),
    .B(_04901_),
    .Y(_00546_));
 sg13g2_mux2_1 _10750_ (.A0(_03048_),
    .A1(_03955_),
    .S(_04791_),
    .X(_04902_));
 sg13g2_nor3_1 _10751_ (.A(_01644_),
    .B(net74),
    .C(_02714_),
    .Y(_04903_));
 sg13g2_a21oi_1 _10752_ (.A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .A2(net73),
    .Y(_04904_),
    .B1(_04903_));
 sg13g2_nor2_1 _10753_ (.A(net76),
    .B(_04904_),
    .Y(_04905_));
 sg13g2_a221oi_1 _10754_ (.B2(net77),
    .C1(_04905_),
    .B1(_04902_),
    .A1(net258),
    .Y(_04906_),
    .A2(_04789_));
 sg13g2_nor2_1 _10755_ (.A(_04822_),
    .B(_04906_),
    .Y(_00547_));
 sg13g2_nor2_1 _10756_ (.A(net255),
    .B(net58),
    .Y(_04907_));
 sg13g2_nand2_1 _10757_ (.Y(_04908_),
    .A(net161),
    .B(_03049_));
 sg13g2_o21ai_1 _10758_ (.B1(_04908_),
    .Y(_04909_),
    .A1(net161),
    .A2(_03966_));
 sg13g2_xor2_1 _10759_ (.B(_02753_),
    .A(net255),
    .X(_04910_));
 sg13g2_nor2_1 _10760_ (.A(net74),
    .B(_04910_),
    .Y(_04911_));
 sg13g2_a21oi_1 _10761_ (.A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .A2(_04806_),
    .Y(_04912_),
    .B1(_04911_));
 sg13g2_nor2_1 _10762_ (.A(net76),
    .B(_04912_),
    .Y(_04913_));
 sg13g2_a221oi_1 _10763_ (.B2(net77),
    .C1(_04913_),
    .B1(_04909_),
    .A1(net82),
    .Y(_04914_),
    .A2(net65));
 sg13g2_nor3_1 _10764_ (.A(net196),
    .B(_04907_),
    .C(_04914_),
    .Y(_00548_));
 sg13g2_nor2_1 _10765_ (.A(net304),
    .B(net58),
    .Y(_04915_));
 sg13g2_mux2_1 _10766_ (.A0(_02282_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .S(net73),
    .X(_04916_));
 sg13g2_nor2_1 _10767_ (.A(net174),
    .B(_03977_),
    .Y(_04917_));
 sg13g2_nor2_1 _10768_ (.A(net175),
    .B(_03050_),
    .Y(_04918_));
 sg13g2_nor3_1 _10769_ (.A(net78),
    .B(_04917_),
    .C(_04918_),
    .Y(_04919_));
 sg13g2_a221oi_1 _10770_ (.B2(_04809_),
    .C1(_04919_),
    .B1(_04916_),
    .A1(net82),
    .Y(_04920_),
    .A2(net65));
 sg13g2_nor3_1 _10771_ (.A(_04773_),
    .B(_04915_),
    .C(_04920_),
    .Y(_00549_));
 sg13g2_nor2_1 _10772_ (.A(net287),
    .B(net58),
    .Y(_04921_));
 sg13g2_mux2_1 _10773_ (.A0(_02624_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .S(net73),
    .X(_04922_));
 sg13g2_nor2_1 _10774_ (.A(net174),
    .B(_03988_),
    .Y(_04923_));
 sg13g2_a21oi_1 _10775_ (.A1(_04811_),
    .A2(_03051_),
    .Y(_04924_),
    .B1(_04923_));
 sg13g2_nor2_1 _10776_ (.A(_04808_),
    .B(_04924_),
    .Y(_04925_));
 sg13g2_a221oi_1 _10777_ (.B2(_04809_),
    .C1(_04925_),
    .B1(_04922_),
    .A1(_01658_),
    .Y(_04926_),
    .A2(_04805_));
 sg13g2_nor3_1 _10778_ (.A(net196),
    .B(_04921_),
    .C(_04926_),
    .Y(_00550_));
 sg13g2_mux2_1 _10779_ (.A0(_03019_),
    .A1(_03673_),
    .S(net162),
    .X(_04927_));
 sg13g2_nor3_1 _10780_ (.A(_01644_),
    .B(_04797_),
    .C(_02709_),
    .Y(_04928_));
 sg13g2_a21oi_1 _10781_ (.A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .A2(net73),
    .Y(_04929_),
    .B1(_04928_));
 sg13g2_nor2_1 _10782_ (.A(_04795_),
    .B(_04929_),
    .Y(_04930_));
 sg13g2_a221oi_1 _10783_ (.B2(net77),
    .C1(_04930_),
    .B1(_04927_),
    .A1(net257),
    .Y(_04931_),
    .A2(_04788_));
 sg13g2_nor2_1 _10784_ (.A(_04822_),
    .B(_04931_),
    .Y(_00551_));
 sg13g2_nand2_1 _10785_ (.Y(_04932_),
    .A(net288),
    .B(net66));
 sg13g2_nand2b_1 _10786_ (.Y(_04933_),
    .B(net81),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_o21ai_1 _10787_ (.B1(_04933_),
    .Y(_04934_),
    .A1(_04797_),
    .A2(_02747_));
 sg13g2_mux2_1 _10788_ (.A0(_03023_),
    .A1(_03701_),
    .S(_04790_),
    .X(_04935_));
 sg13g2_nand2_1 _10789_ (.Y(_04936_),
    .A(net83),
    .B(_04935_));
 sg13g2_o21ai_1 _10790_ (.B1(_04936_),
    .Y(_04937_),
    .A1(_04795_),
    .A2(_04934_));
 sg13g2_nand2_1 _10791_ (.Y(_04938_),
    .A(net58),
    .B(_04937_));
 sg13g2_a21oi_1 _10792_ (.A1(_04932_),
    .A2(_04938_),
    .Y(_00552_),
    .B1(_04778_));
 sg13g2_nor2_1 _10793_ (.A(net289),
    .B(_04803_),
    .Y(_04939_));
 sg13g2_mux2_1 _10794_ (.A0(_02281_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .S(net74),
    .X(_04940_));
 sg13g2_nor2_1 _10795_ (.A(net174),
    .B(_03719_),
    .Y(_04941_));
 sg13g2_a21oi_1 _10796_ (.A1(_04811_),
    .A2(_03024_),
    .Y(_04942_),
    .B1(_04941_));
 sg13g2_nor2_1 _10797_ (.A(_04808_),
    .B(_04942_),
    .Y(_04943_));
 sg13g2_a221oi_1 _10798_ (.B2(net78),
    .C1(_04943_),
    .B1(_04940_),
    .A1(_01658_),
    .Y(_04944_),
    .A2(_04805_));
 sg13g2_nor3_1 _10799_ (.A(net196),
    .B(_04939_),
    .C(_04944_),
    .Y(_00553_));
 sg13g2_nor3_1 _10800_ (.A(net83),
    .B(_01365_),
    .C(_01419_),
    .Y(_04945_));
 sg13g2_nor2_1 _10801_ (.A(_04945_),
    .B(_03417_),
    .Y(_04946_));
 sg13g2_nor3_1 _10802_ (.A(\i_tinyqv.cpu.instr_fetch_started ),
    .B(\i_tinyqv.cpu.instr_fetch_stopped ),
    .C(\i_tinyqv.cpu.instr_fetch_running ),
    .Y(_04947_));
 sg13g2_and2_1 _10803_ (.A(_04946_),
    .B(_04947_),
    .X(_04948_));
 sg13g2_nand2b_1 _10804_ (.Y(_04949_),
    .B(\i_tinyqv.cpu.instr_fetch_stopped ),
    .A_N(\i_tinyqv.cpu.instr_fetch_started ));
 sg13g2_a22oi_1 _10805_ (.Y(_04950_),
    .B1(_04946_),
    .B2(_04949_),
    .A2(net77),
    .A1(net240));
 sg13g2_nor3_1 _10806_ (.A(net196),
    .B(_04948_),
    .C(_04950_),
    .Y(_00554_));
 sg13g2_inv_1 _10807_ (.Y(_04951_),
    .A(_01290_));
 sg13g2_buf_1 _10808_ (.A(net56),
    .X(_04952_));
 sg13g2_o21ai_1 _10809_ (.B1(_01282_),
    .Y(_04953_),
    .A1(net90),
    .A2(net56));
 sg13g2_a21oi_1 _10810_ (.A1(_04951_),
    .A2(_04952_),
    .Y(_00555_),
    .B1(_04953_));
 sg13g2_a21o_1 _10811_ (.A2(_04952_),
    .A1(\i_tinyqv.cpu.instr_len[2] ),
    .B1(_04953_),
    .X(_00556_));
 sg13g2_nor2_1 _10812_ (.A(_01224_),
    .B(_01393_),
    .Y(_04954_));
 sg13g2_o21ai_1 _10813_ (.B1(_03534_),
    .Y(_04955_),
    .A1(_04954_),
    .A2(_02907_));
 sg13g2_nand2_1 _10814_ (.Y(_04956_),
    .A(_01288_),
    .B(_04955_));
 sg13g2_nor2_1 _10815_ (.A(net76),
    .B(_01419_),
    .Y(_04957_));
 sg13g2_nand3b_1 _10816_ (.B(_01494_),
    .C(_04957_),
    .Y(_04958_),
    .A_N(_04955_));
 sg13g2_a21oi_1 _10817_ (.A1(_04956_),
    .A2(_04958_),
    .Y(_00557_),
    .B1(net195));
 sg13g2_nand2_1 _10818_ (.Y(_04959_),
    .A(_01262_),
    .B(_03034_));
 sg13g2_o21ai_1 _10819_ (.B1(_04959_),
    .Y(_04960_),
    .A1(_01262_),
    .A2(_03845_));
 sg13g2_a22oi_1 _10820_ (.Y(_04961_),
    .B1(_01281_),
    .B2(_04960_),
    .A2(net74),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_o21ai_1 _10821_ (.B1(_01408_),
    .Y(_04962_),
    .A1(_01431_),
    .A2(_01433_));
 sg13g2_nand3b_1 _10822_ (.B(net65),
    .C(_04962_),
    .Y(_04963_),
    .A_N(_01434_));
 sg13g2_a21oi_1 _10823_ (.A1(_04961_),
    .A2(_04963_),
    .Y(_00558_),
    .B1(net195));
 sg13g2_mux2_1 _10824_ (.A0(_03040_),
    .A1(_03917_),
    .S(_04790_),
    .X(_04964_));
 sg13g2_a22oi_1 _10825_ (.Y(_04965_),
    .B1(net76),
    .B2(_04964_),
    .A2(net75),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_xnor2_1 _10826_ (.Y(_04966_),
    .A(_00158_),
    .B(_01434_));
 sg13g2_nand2_1 _10827_ (.Y(_04967_),
    .A(net65),
    .B(_04966_));
 sg13g2_a21oi_1 _10828_ (.A1(_04965_),
    .A2(_04967_),
    .Y(_00559_),
    .B1(net199));
 sg13g2_nand2_1 _10829_ (.Y(_04968_),
    .A(_03534_),
    .B(_02907_));
 sg13g2_a22oi_1 _10830_ (.Y(_04969_),
    .B1(_04968_),
    .B2(_04763_),
    .A2(net79),
    .A1(_04954_));
 sg13g2_nor2_1 _10831_ (.A(net194),
    .B(_04969_),
    .Y(_00561_));
 sg13g2_o21ai_1 _10832_ (.B1(_02959_),
    .Y(_04970_),
    .A1(net115),
    .A2(_02984_));
 sg13g2_a21oi_1 _10833_ (.A1(net101),
    .A2(_04970_),
    .Y(_04971_),
    .B1(_03169_));
 sg13g2_o21ai_1 _10834_ (.B1(_03199_),
    .Y(_04972_),
    .A1(net108),
    .A2(_04971_));
 sg13g2_nor3_1 _10835_ (.A(net90),
    .B(_01345_),
    .C(_02937_),
    .Y(_04973_));
 sg13g2_a21oi_1 _10836_ (.A1(net90),
    .A2(_04972_),
    .Y(_04974_),
    .B1(_04973_));
 sg13g2_nor2_1 _10837_ (.A(net56),
    .B(_04974_),
    .Y(_04975_));
 sg13g2_a21oi_1 _10838_ (.A1(\i_tinyqv.cpu.is_alu_imm ),
    .A2(net46),
    .Y(_04976_),
    .B1(_04975_));
 sg13g2_nor2_1 _10839_ (.A(net194),
    .B(_04976_),
    .Y(_00562_));
 sg13g2_nor2_1 _10840_ (.A(net90),
    .B(_02937_),
    .Y(_04977_));
 sg13g2_o21ai_1 _10841_ (.B1(_01345_),
    .Y(_04978_),
    .A1(_01468_),
    .A2(_04977_));
 sg13g2_a221oi_1 _10842_ (.B2(_02984_),
    .C1(_02971_),
    .B1(_02987_),
    .A1(_02921_),
    .Y(_04979_),
    .A2(_01468_));
 sg13g2_a21oi_1 _10843_ (.A1(_04978_),
    .A2(_04979_),
    .Y(_04980_),
    .B1(net56));
 sg13g2_a21oi_1 _10844_ (.A1(\i_tinyqv.cpu.is_alu_reg ),
    .A2(net46),
    .Y(_04981_),
    .B1(_04980_));
 sg13g2_nor2_1 _10845_ (.A(net195),
    .B(_04981_),
    .Y(_00563_));
 sg13g2_nand2_1 _10846_ (.Y(_04982_),
    .A(net88),
    .B(_02922_));
 sg13g2_nor3_1 _10847_ (.A(net56),
    .B(_02951_),
    .C(_04982_),
    .Y(_04983_));
 sg13g2_a21oi_1 _10848_ (.A1(\i_tinyqv.cpu.is_auipc ),
    .A2(net46),
    .Y(_04984_),
    .B1(_04983_));
 sg13g2_nor2_1 _10849_ (.A(net195),
    .B(_04984_),
    .Y(_00564_));
 sg13g2_nor2_1 _10850_ (.A(_00868_),
    .B(_04718_),
    .Y(_04985_));
 sg13g2_a221oi_1 _10851_ (.B2(net94),
    .C1(net46),
    .B1(_02956_),
    .A1(net88),
    .Y(_04986_),
    .A2(_02933_));
 sg13g2_nor3_1 _10852_ (.A(net196),
    .B(_04985_),
    .C(_04986_),
    .Y(_00565_));
 sg13g2_nand2_1 _10853_ (.Y(_04987_),
    .A(_01364_),
    .B(_04718_));
 sg13g2_nand2_1 _10854_ (.Y(_04988_),
    .A(\i_tinyqv.cpu.is_jal ),
    .B(net46));
 sg13g2_a21oi_1 _10855_ (.A1(_04987_),
    .A2(_04988_),
    .Y(_00566_),
    .B1(net199));
 sg13g2_nand2b_1 _10856_ (.Y(_04989_),
    .B(_01469_),
    .A_N(_03178_));
 sg13g2_nand4_1 _10857_ (.B(net130),
    .C(_02923_),
    .A(net88),
    .Y(_04990_),
    .D(_01353_));
 sg13g2_a21oi_1 _10858_ (.A1(_04989_),
    .A2(_04990_),
    .Y(_04991_),
    .B1(_02911_));
 sg13g2_a21oi_1 _10859_ (.A1(\i_tinyqv.cpu.is_jalr ),
    .A2(net46),
    .Y(_04992_),
    .B1(_04991_));
 sg13g2_nor2_1 _10860_ (.A(net195),
    .B(_04992_),
    .Y(_00567_));
 sg13g2_nor2_1 _10861_ (.A(net91),
    .B(_02932_),
    .Y(_04993_));
 sg13g2_nand3_1 _10862_ (.B(_02949_),
    .C(_03589_),
    .A(net128),
    .Y(_04994_));
 sg13g2_o21ai_1 _10863_ (.B1(_04994_),
    .Y(_04995_),
    .A1(_02959_),
    .A2(net116));
 sg13g2_a221oi_1 _10864_ (.B2(_04995_),
    .C1(net88),
    .B1(_04993_),
    .A1(net103),
    .Y(_04996_),
    .A2(_03283_));
 sg13g2_a21oi_1 _10865_ (.A1(net88),
    .A2(_01455_),
    .Y(_04997_),
    .B1(_04996_));
 sg13g2_nand2_1 _10866_ (.Y(_04998_),
    .A(_04718_),
    .B(_04997_));
 sg13g2_nand2_1 _10867_ (.Y(_04999_),
    .A(_01170_),
    .B(net46));
 sg13g2_a21oi_1 _10868_ (.A1(_04998_),
    .A2(_04999_),
    .Y(_00568_),
    .B1(net199));
 sg13g2_o21ai_1 _10869_ (.B1(_03260_),
    .Y(_05000_),
    .A1(net136),
    .A2(_03298_));
 sg13g2_mux2_1 _10870_ (.A0(\i_tinyqv.cpu.is_lui ),
    .A1(_05000_),
    .S(_04718_),
    .X(_05001_));
 sg13g2_and2_1 _10871_ (.A(net241),
    .B(_05001_),
    .X(_00569_));
 sg13g2_nor2_1 _10872_ (.A(_01196_),
    .B(_04718_),
    .Y(_05002_));
 sg13g2_or2_1 _10873_ (.X(_05003_),
    .B(_02949_),
    .A(net103));
 sg13g2_o21ai_1 _10874_ (.B1(_03186_),
    .Y(_05004_),
    .A1(_01467_),
    .A2(_05003_));
 sg13g2_a221oi_1 _10875_ (.B2(net100),
    .C1(net56),
    .B1(_05004_),
    .A1(net88),
    .Y(_05005_),
    .A2(_03159_));
 sg13g2_nor3_1 _10876_ (.A(net196),
    .B(_05002_),
    .C(_05005_),
    .Y(_00570_));
 sg13g2_nand2_1 _10877_ (.Y(_05006_),
    .A(_01451_),
    .B(net123));
 sg13g2_nor3_1 _10878_ (.A(_03242_),
    .B(_01352_),
    .C(_05006_),
    .Y(_05007_));
 sg13g2_a221oi_1 _10879_ (.B2(_03566_),
    .C1(_05007_),
    .B1(_03170_),
    .A1(_01469_),
    .Y(_05008_),
    .A2(_03178_));
 sg13g2_nor2_1 _10880_ (.A(net56),
    .B(_05008_),
    .Y(_05009_));
 sg13g2_a21oi_1 _10881_ (.A1(\i_tinyqv.cpu.is_system ),
    .A2(net46),
    .Y(_05010_),
    .B1(_05009_));
 sg13g2_nor2_1 _10882_ (.A(net195),
    .B(_05010_),
    .Y(_00571_));
 sg13g2_inv_1 _10883_ (.Y(_05011_),
    .A(\i_tinyqv.cpu.load_started ));
 sg13g2_a21oi_1 _10884_ (.A1(_05011_),
    .A2(net134),
    .Y(_00572_),
    .B1(_04315_));
 sg13g2_a21oi_1 _10885_ (.A1(_01232_),
    .A2(\i_tinyqv.cpu.data_write_n[1] ),
    .Y(_05012_),
    .B1(_01565_));
 sg13g2_nand2_1 _10886_ (.Y(_05013_),
    .A(net160),
    .B(_04732_));
 sg13g2_a21oi_1 _10887_ (.A1(\i_tinyqv.cpu.no_write_in_progress ),
    .A2(net168),
    .Y(_05014_),
    .B1(net212));
 sg13g2_o21ai_1 _10888_ (.B1(_05014_),
    .Y(_00577_),
    .A1(_05012_),
    .A2(_05013_));
 sg13g2_o21ai_1 _10889_ (.B1(net65),
    .Y(_05015_),
    .A1(_01298_),
    .A2(net82));
 sg13g2_a21o_1 _10890_ (.A2(_04961_),
    .A1(_04951_),
    .B1(_04788_),
    .X(_05016_));
 sg13g2_inv_1 _10891_ (.Y(_05017_),
    .A(net309));
 sg13g2_a221oi_1 _10892_ (.B2(_05017_),
    .C1(net199),
    .B1(_05016_),
    .A1(_04961_),
    .Y(_00578_),
    .A2(_05015_));
 sg13g2_o21ai_1 _10893_ (.B1(net65),
    .Y(_05018_),
    .A1(_01300_),
    .A2(net82));
 sg13g2_a221oi_1 _10894_ (.B2(_05018_),
    .C1(net199),
    .B1(_04965_),
    .A1(_01400_),
    .Y(_00579_),
    .A2(net66));
 sg13g2_a21oi_1 _10895_ (.A1(net240),
    .A2(_01367_),
    .Y(_05019_),
    .B1(_04945_));
 sg13g2_nor2_1 _10896_ (.A(net195),
    .B(_05019_),
    .Y(_00592_));
 sg13g2_nand3_1 _10897_ (.B(net210),
    .C(_01508_),
    .A(_04140_),
    .Y(_05020_));
 sg13g2_o21ai_1 _10898_ (.B1(_05020_),
    .Y(_05021_),
    .A1(net230),
    .A2(net210));
 sg13g2_nand2_1 _10899_ (.Y(_05022_),
    .A(_04019_),
    .B(_05021_));
 sg13g2_o21ai_1 _10900_ (.B1(_05022_),
    .Y(_05023_),
    .A1(_01508_),
    .A2(_04521_));
 sg13g2_or4_1 _10901_ (.A(_04019_),
    .B(_04140_),
    .C(_01509_),
    .D(_01563_),
    .X(_05024_));
 sg13g2_a221oi_1 _10902_ (.B2(\i_tinyqv.mem.data_stall ),
    .C1(_01560_),
    .B1(_05024_),
    .A1(_01240_),
    .Y(_05025_),
    .A2(_05023_));
 sg13g2_nor2b_1 _10903_ (.A(_05025_),
    .B_N(debug_data_continue),
    .Y(_00593_));
 sg13g2_and2_1 _10904_ (.A(net213),
    .B(_03623_),
    .X(_00595_));
 sg13g2_and2_1 _10905_ (.A(net261),
    .B(_04091_),
    .X(_00596_));
 sg13g2_nor3_1 _10906_ (.A(_04136_),
    .B(_04106_),
    .C(_04108_),
    .Y(_05026_));
 sg13g2_nor2_1 _10907_ (.A(_04126_),
    .B(_05026_),
    .Y(_05027_));
 sg13g2_nor2_1 _10908_ (.A(_04097_),
    .B(_05027_),
    .Y(_00629_));
 sg13g2_nand2b_1 _10909_ (.Y(_00638_),
    .B(net213),
    .A_N(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ));
 sg13g2_nand2b_1 _10910_ (.Y(_00639_),
    .B(net213),
    .A_N(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ));
 sg13g2_nor2_1 _10911_ (.A(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .B(_04092_),
    .Y(_05028_));
 sg13g2_and2_1 _10912_ (.A(_00596_),
    .B(_05028_),
    .X(_00659_));
 sg13g2_nor2b_1 _10913_ (.A(_04180_),
    .B_N(_04181_),
    .Y(_05029_));
 sg13g2_nor4_1 _10914_ (.A(\i_uart_rx.cycle_counter[3] ),
    .B(_04179_),
    .C(\i_uart_rx.cycle_counter[9] ),
    .D(_04559_),
    .Y(_05030_));
 sg13g2_nand4_1 _10915_ (.B(_04188_),
    .C(_05029_),
    .A(_04187_),
    .Y(_05031_),
    .D(_05030_));
 sg13g2_nor4_2 _10916_ (.A(_04184_),
    .B(_04185_),
    .C(\i_uart_rx.cycle_counter[10] ),
    .Y(_05032_),
    .D(_05031_));
 sg13g2_nand2b_1 _10917_ (.Y(_05033_),
    .B(\i_uart_rx.bit_sample ),
    .A_N(_05032_));
 sg13g2_nand2_1 _10918_ (.Y(_05034_),
    .A(\i_uart_rx.rxd_reg[0] ),
    .B(_05032_));
 sg13g2_a21oi_1 _10919_ (.A1(_05033_),
    .A2(_05034_),
    .Y(_00694_),
    .B1(net177));
 sg13g2_nand2_1 _10920_ (.Y(_05035_),
    .A(_01568_),
    .B(net150));
 sg13g2_a21oi_1 _10921_ (.A1(_01378_),
    .A2(_04536_),
    .Y(_05036_),
    .B1(net299));
 sg13g2_or2_1 _10922_ (.X(_05037_),
    .B(_05036_),
    .A(_04192_));
 sg13g2_buf_1 _10923_ (.A(_05037_),
    .X(_05038_));
 sg13g2_inv_1 _10924_ (.Y(_05039_),
    .A(_05038_));
 sg13g2_a21oi_1 _10925_ (.A1(_01381_),
    .A2(_05035_),
    .Y(_05040_),
    .B1(_05039_));
 sg13g2_nand2b_1 _10926_ (.Y(_05041_),
    .B(_01379_),
    .A_N(net300));
 sg13g2_nor2_1 _10927_ (.A(_00203_),
    .B(_05041_),
    .Y(_05042_));
 sg13g2_nor2_1 _10928_ (.A(net300),
    .B(\i_uart_rx.rxd_reg[0] ),
    .Y(_05043_));
 sg13g2_a22oi_1 _10929_ (.Y(_05044_),
    .B1(_04194_),
    .B2(_05043_),
    .A2(_00202_),
    .A1(_01377_));
 sg13g2_nor2_1 _10930_ (.A(_01377_),
    .B(_04535_),
    .Y(_05045_));
 sg13g2_o21ai_1 _10931_ (.B1(_00202_),
    .Y(_05046_),
    .A1(net299),
    .A2(_05045_));
 sg13g2_o21ai_1 _10932_ (.B1(_05046_),
    .Y(_05047_),
    .A1(net278),
    .A2(_05044_));
 sg13g2_a21oi_1 _10933_ (.A1(_05032_),
    .A2(_05042_),
    .Y(_05048_),
    .B1(_05047_));
 sg13g2_o21ai_1 _10934_ (.B1(_01598_),
    .Y(_05049_),
    .A1(net300),
    .A2(_05038_));
 sg13g2_a21oi_1 _10935_ (.A1(_05040_),
    .A2(_05048_),
    .Y(_00706_),
    .B1(_05049_));
 sg13g2_a21oi_1 _10936_ (.A1(_00203_),
    .A2(_05032_),
    .Y(_05050_),
    .B1(_05041_));
 sg13g2_nor2b_1 _10937_ (.A(_05050_),
    .B_N(_05040_),
    .Y(_05051_));
 sg13g2_inv_1 _10938_ (.Y(_05052_),
    .A(_05051_));
 sg13g2_o21ai_1 _10939_ (.B1(_05038_),
    .Y(_05053_),
    .A1(net300),
    .A2(_05052_));
 sg13g2_nand2_1 _10940_ (.Y(_05054_),
    .A(_01377_),
    .B(net300));
 sg13g2_o21ai_1 _10941_ (.B1(_05054_),
    .Y(_05055_),
    .A1(net299),
    .A2(_01378_));
 sg13g2_a221oi_1 _10942_ (.B2(_05051_),
    .C1(net178),
    .B1(_05055_),
    .A1(_04534_),
    .Y(_00707_),
    .A2(_05053_));
 sg13g2_nand3_1 _10943_ (.B(_01375_),
    .C(_04192_),
    .A(_01377_),
    .Y(_05056_));
 sg13g2_nor3_1 _10944_ (.A(net299),
    .B(_04193_),
    .C(_05056_),
    .Y(_05057_));
 sg13g2_a21o_1 _10945_ (.A2(_05056_),
    .A1(net299),
    .B1(_05057_),
    .X(_05058_));
 sg13g2_and2_1 _10946_ (.A(net213),
    .B(_05058_),
    .X(_00708_));
 sg13g2_nand2b_1 _10947_ (.Y(_05059_),
    .B(net278),
    .A_N(_01375_));
 sg13g2_o21ai_1 _10948_ (.B1(_05059_),
    .Y(_05060_),
    .A1(_04193_),
    .A2(_05054_));
 sg13g2_a22oi_1 _10949_ (.Y(_05061_),
    .B1(_05060_),
    .B2(net299),
    .A2(net278),
    .A1(_04534_));
 sg13g2_o21ai_1 _10950_ (.B1(_01598_),
    .Y(_05062_),
    .A1(net278),
    .A2(_05038_));
 sg13g2_a21oi_1 _10951_ (.A1(_05051_),
    .A2(_05061_),
    .Y(_00709_),
    .B1(_05062_));
 sg13g2_nand2b_1 _10952_ (.Y(_00718_),
    .B(net213),
    .A_N(\i_uart_rx.rxd_reg[1] ));
 sg13g2_nand2b_1 _10953_ (.Y(_00719_),
    .B(_04654_),
    .A_N(net7));
 sg13g2_nand3b_1 _10954_ (.B(net213),
    .C(_04194_),
    .Y(_00720_),
    .A_N(net278));
 sg13g2_nand3_1 _10955_ (.B(_01567_),
    .C(_02182_),
    .A(net209),
    .Y(_05063_));
 sg13g2_buf_1 _10956_ (.A(_05063_),
    .X(_05064_));
 sg13g2_inv_2 _10957_ (.Y(_05065_),
    .A(_05064_));
 sg13g2_nand2_1 _10958_ (.Y(_05066_),
    .A(_01573_),
    .B(_05065_));
 sg13g2_xnor2_1 _10959_ (.Y(_05067_),
    .A(_01386_),
    .B(_01384_));
 sg13g2_and2_1 _10960_ (.A(net179),
    .B(_05067_),
    .X(_05068_));
 sg13g2_buf_2 _10961_ (.A(_05068_),
    .X(_05069_));
 sg13g2_mux2_1 _10962_ (.A0(\i_uart_tx.data_to_send[0] ),
    .A1(\i_uart_tx.data_to_send[1] ),
    .S(_05069_),
    .X(_05070_));
 sg13g2_nand2_1 _10963_ (.Y(_05071_),
    .A(net111),
    .B(_05070_));
 sg13g2_a21oi_1 _10964_ (.A1(_05066_),
    .A2(_05071_),
    .Y(_00732_),
    .B1(_04632_));
 sg13g2_nand2_1 _10965_ (.Y(_05072_),
    .A(_01600_),
    .B(_05065_));
 sg13g2_mux2_1 _10966_ (.A0(\i_uart_tx.data_to_send[1] ),
    .A1(\i_uart_tx.data_to_send[2] ),
    .S(_05069_),
    .X(_05073_));
 sg13g2_nand2_1 _10967_ (.Y(_05074_),
    .A(net111),
    .B(_05073_));
 sg13g2_a21oi_1 _10968_ (.A1(_05072_),
    .A2(_05074_),
    .Y(_00733_),
    .B1(net177));
 sg13g2_nand2_1 _10969_ (.Y(_05075_),
    .A(_01603_),
    .B(_05065_));
 sg13g2_mux2_1 _10970_ (.A0(\i_uart_tx.data_to_send[2] ),
    .A1(\i_uart_tx.data_to_send[3] ),
    .S(_05069_),
    .X(_05076_));
 sg13g2_nand2_1 _10971_ (.Y(_05077_),
    .A(net111),
    .B(_05076_));
 sg13g2_a21oi_1 _10972_ (.A1(_05075_),
    .A2(_05077_),
    .Y(_00734_),
    .B1(net177));
 sg13g2_nand2_1 _10973_ (.Y(_05078_),
    .A(_01606_),
    .B(_05065_));
 sg13g2_mux2_1 _10974_ (.A0(\i_uart_tx.data_to_send[3] ),
    .A1(\i_uart_tx.data_to_send[4] ),
    .S(_05069_),
    .X(_05079_));
 sg13g2_nand2_1 _10975_ (.Y(_05080_),
    .A(net111),
    .B(_05079_));
 sg13g2_a21oi_1 _10976_ (.A1(_05078_),
    .A2(_05080_),
    .Y(_00735_),
    .B1(net177));
 sg13g2_nand2_1 _10977_ (.Y(_05081_),
    .A(_01609_),
    .B(_05065_));
 sg13g2_mux2_1 _10978_ (.A0(\i_uart_tx.data_to_send[4] ),
    .A1(\i_uart_tx.data_to_send[5] ),
    .S(_05069_),
    .X(_05082_));
 sg13g2_nand2_1 _10979_ (.Y(_05083_),
    .A(net111),
    .B(_05082_));
 sg13g2_a21oi_1 _10980_ (.A1(_05081_),
    .A2(_05083_),
    .Y(_00736_),
    .B1(net177));
 sg13g2_nand2_1 _10981_ (.Y(_05084_),
    .A(_01612_),
    .B(_05065_));
 sg13g2_mux2_1 _10982_ (.A0(\i_uart_tx.data_to_send[5] ),
    .A1(\i_uart_tx.data_to_send[6] ),
    .S(_05069_),
    .X(_05085_));
 sg13g2_nand2_1 _10983_ (.Y(_05086_),
    .A(_05064_),
    .B(_05085_));
 sg13g2_a21oi_1 _10984_ (.A1(_05084_),
    .A2(_05086_),
    .Y(_00737_),
    .B1(net178));
 sg13g2_nand2_1 _10985_ (.Y(_05087_),
    .A(_01616_),
    .B(_05065_));
 sg13g2_mux2_1 _10986_ (.A0(\i_uart_tx.data_to_send[6] ),
    .A1(\i_uart_tx.data_to_send[7] ),
    .S(_05069_),
    .X(_05088_));
 sg13g2_nand2_1 _10987_ (.Y(_05089_),
    .A(net111),
    .B(_05088_));
 sg13g2_a21oi_1 _10988_ (.A1(_05087_),
    .A2(_05089_),
    .Y(_00738_),
    .B1(_04601_));
 sg13g2_or2_1 _10989_ (.X(_05090_),
    .B(net111),
    .A(_00201_));
 sg13g2_nand3b_1 _10990_ (.B(\i_uart_tx.data_to_send[7] ),
    .C(net111),
    .Y(_05091_),
    .A_N(_05069_));
 sg13g2_a21oi_1 _10991_ (.A1(_05090_),
    .A2(_05091_),
    .Y(_00739_),
    .B1(net178));
 sg13g2_a21oi_1 _10992_ (.A1(_01386_),
    .A2(net179),
    .Y(_05092_),
    .B1(_05065_));
 sg13g2_inv_1 _10993_ (.Y(_05093_),
    .A(_01386_));
 sg13g2_a21oi_1 _10994_ (.A1(_01382_),
    .A2(_05093_),
    .Y(_05094_),
    .B1(_01383_));
 sg13g2_nand2b_1 _10995_ (.Y(_05095_),
    .B(net179),
    .A_N(_05094_));
 sg13g2_o21ai_1 _10996_ (.B1(_05095_),
    .Y(_05096_),
    .A1(_01382_),
    .A2(_05092_));
 sg13g2_nand2_1 _10997_ (.Y(_05097_),
    .A(_01385_),
    .B(net179));
 sg13g2_o21ai_1 _10998_ (.B1(_05097_),
    .Y(_05098_),
    .A1(_01385_),
    .A2(_05096_));
 sg13g2_nor2_1 _10999_ (.A(net176),
    .B(_05098_),
    .Y(_00740_));
 sg13g2_nor2_1 _11000_ (.A(_05093_),
    .B(_01383_),
    .Y(_05099_));
 sg13g2_o21ai_1 _11001_ (.B1(net179),
    .Y(_05100_),
    .A1(_01385_),
    .A2(_05099_));
 sg13g2_nor2_1 _11002_ (.A(_01382_),
    .B(_05097_),
    .Y(_05101_));
 sg13g2_a21oi_1 _11003_ (.A1(_01382_),
    .A2(_05100_),
    .Y(_05102_),
    .B1(_05101_));
 sg13g2_nor2_1 _11004_ (.A(_04633_),
    .B(_05102_),
    .Y(_00741_));
 sg13g2_nand3_1 _11005_ (.B(_01382_),
    .C(net179),
    .A(_01385_),
    .Y(_05103_));
 sg13g2_xor2_1 _11006_ (.B(_05103_),
    .A(_01383_),
    .X(_05104_));
 sg13g2_nor2_1 _11007_ (.A(_04633_),
    .B(_05104_),
    .Y(_00742_));
 sg13g2_nand2b_1 _11008_ (.Y(_05105_),
    .B(_01383_),
    .A_N(_01385_));
 sg13g2_nand3_1 _11009_ (.B(net179),
    .C(_05105_),
    .A(_01382_),
    .Y(_05106_));
 sg13g2_nand4_1 _11010_ (.B(_05093_),
    .C(_01383_),
    .A(_01382_),
    .Y(_05107_),
    .D(net179));
 sg13g2_nand2b_1 _11011_ (.Y(_05108_),
    .B(_05107_),
    .A_N(_05099_));
 sg13g2_a22oi_1 _11012_ (.Y(_05109_),
    .B1(_05108_),
    .B2(_01385_),
    .A2(_05106_),
    .A1(_01386_));
 sg13g2_nor2_1 _11013_ (.A(_04632_),
    .B(_05109_),
    .Y(_00743_));
 sg13g2_a21oi_1 _11014_ (.A1(_01386_),
    .A2(\i_uart_tx.data_to_send[0] ),
    .Y(_05110_),
    .B1(_01387_));
 sg13g2_nor3_1 _11015_ (.A(_01386_),
    .B(\i_uart_tx.data_to_send[0] ),
    .C(_01384_),
    .Y(_05111_));
 sg13g2_a21oi_1 _11016_ (.A1(_01384_),
    .A2(_05110_),
    .Y(_05112_),
    .B1(_05111_));
 sg13g2_nand2b_1 _11017_ (.Y(_00744_),
    .B(_04654_),
    .A_N(_05112_));
 sg13g2_and2_1 _11018_ (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .B(net1),
    .X(net17));
 sg13g2_nor2_1 _11019_ (.A(_03995_),
    .B(_04007_),
    .Y(_05113_));
 sg13g2_a22oi_1 _11020_ (.Y(_05114_),
    .B1(_04504_),
    .B2(_05113_),
    .A2(net200),
    .A1(\i_tinyqv.mem.q_ctrl.addr[20] ));
 sg13g2_nand2b_1 _11021_ (.Y(_05115_),
    .B(net238),
    .A_N(_05114_));
 sg13g2_nand2b_1 _11022_ (.Y(_05116_),
    .B(net231),
    .A_N(_03429_));
 sg13g2_nand2_1 _11023_ (.Y(_05117_),
    .A(_03633_),
    .B(net214));
 sg13g2_a21o_1 _11024_ (.A2(_05116_),
    .A1(_05115_),
    .B1(_05117_),
    .X(_05118_));
 sg13g2_o21ai_1 _11025_ (.B1(_05118_),
    .Y(net21),
    .A1(_04453_),
    .A2(_05115_));
 sg13g2_a21oi_1 _11026_ (.A1(net238),
    .A2(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .Y(_05119_),
    .B1(_04509_));
 sg13g2_nor2_1 _11027_ (.A(_01519_),
    .B(_04114_),
    .Y(_05120_));
 sg13g2_a21oi_1 _11028_ (.A1(net231),
    .A2(_03431_),
    .Y(_05121_),
    .B1(_05120_));
 sg13g2_o21ai_1 _11029_ (.B1(_04424_),
    .Y(_05122_),
    .A1(_01519_),
    .A2(_04007_));
 sg13g2_nor3_1 _11030_ (.A(net235),
    .B(_05121_),
    .C(_05122_),
    .Y(_05123_));
 sg13g2_a21oi_1 _11031_ (.A1(net235),
    .A2(_05119_),
    .Y(net22),
    .B1(_05123_));
 sg13g2_nand2_1 _11032_ (.Y(_05124_),
    .A(_03684_),
    .B(\i_tinyqv.mem.q_ctrl.addr[22] ));
 sg13g2_nand2_1 _11033_ (.Y(_05125_),
    .A(_02676_),
    .B(_04010_));
 sg13g2_o21ai_1 _11034_ (.B1(_05125_),
    .Y(net24),
    .A1(_04453_),
    .A2(_05124_));
 sg13g2_nand2_1 _11035_ (.Y(_05126_),
    .A(_03684_),
    .B(\i_tinyqv.mem.q_ctrl.addr[23] ));
 sg13g2_a22oi_1 _11036_ (.Y(_05127_),
    .B1(_05126_),
    .B2(net200),
    .A2(_04504_),
    .A1(net238));
 sg13g2_nand2_1 _11037_ (.Y(_05128_),
    .A(_03435_),
    .B(_04010_));
 sg13g2_o21ai_1 _11038_ (.B1(_05128_),
    .Y(_05129_),
    .A1(net231),
    .A2(_05127_));
 sg13g2_o21ai_1 _11039_ (.B1(_05129_),
    .Y(net25),
    .A1(_05117_),
    .A2(_05115_));
 sg13g2_dfrbp_1 _11040_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net318),
    .D(_00222_),
    .Q_N(_05521_),
    .Q(\i_tinyqv.cpu.i_core.mip[17] ));
 sg13g2_dfrbp_1 _11041_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net319),
    .D(_00223_),
    .Q_N(_05520_),
    .Q(\i_tinyqv.cpu.i_core.mip[16] ));
 sg13g2_dfrbp_1 _11042_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net320),
    .D(_00224_),
    .Q_N(_05519_),
    .Q(\i_tinyqv.cpu.i_core.mie[19] ));
 sg13g2_dfrbp_1 _11043_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net321),
    .D(_00225_),
    .Q_N(_05518_),
    .Q(\i_tinyqv.cpu.i_core.mie[18] ));
 sg13g2_dfrbp_1 _11044_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net322),
    .D(_00226_),
    .Q_N(_05517_),
    .Q(\i_tinyqv.cpu.i_core.mie[17] ));
 sg13g2_dfrbp_1 _11045_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net323),
    .D(_00227_),
    .Q_N(_05522_),
    .Q(\i_tinyqv.cpu.i_core.mie[16] ));
 sg13g2_inv_1 _08242__1 (.Y(net1354),
    .A(clknet_leaf_46_clk));
 sg13g2_buf_1 _11047_ (.A(net1),
    .X(net12));
 sg13g2_buf_1 _11048_ (.A(net17),
    .X(net13));
 sg13g2_buf_1 _11049_ (.A(net17),
    .X(net14));
 sg13g2_buf_1 _11050_ (.A(net1),
    .X(net15));
 sg13g2_buf_1 _11051_ (.A(net17),
    .X(net16));
 sg13g2_buf_1 _11052_ (.A(net1),
    .X(net18));
 sg13g2_buf_1 _11053_ (.A(net1),
    .X(net19));
 sg13g2_buf_1 _11054_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .X(net20));
 sg13g2_buf_1 _11055_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .X(net23));
 sg13g2_buf_1 _11056_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .X(net26));
 sg13g2_buf_1 _11057_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .X(net27));
 sg13g2_dfrbp_1 \debug_rd_r[0]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net324),
    .D(\debug_rd[0] ),
    .Q_N(_05523_),
    .Q(\debug_rd_r[0] ));
 sg13g2_dfrbp_1 \debug_rd_r[1]$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net325),
    .D(\debug_rd[1] ),
    .Q_N(_05524_),
    .Q(\debug_rd_r[1] ));
 sg13g2_dfrbp_1 \debug_rd_r[2]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net326),
    .D(\debug_rd[2] ),
    .Q_N(_05525_),
    .Q(\debug_rd_r[2] ));
 sg13g2_dfrbp_1 \debug_rd_r[3]$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net327),
    .D(\debug_rd[3] ),
    .Q_N(_05516_),
    .Q(\debug_rd_r[3] ));
 sg13g2_dfrbp_1 \debug_register_data$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net328),
    .D(_00228_),
    .Q_N(_05526_),
    .Q(debug_register_data));
 sg13g2_dfrbp_1 \gpio_out[0]$_DFF_P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net329),
    .D(_00000_),
    .Q_N(_05527_),
    .Q(\gpio_out[0] ));
 sg13g2_dfrbp_1 \gpio_out[1]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net330),
    .D(_00001_),
    .Q_N(_05528_),
    .Q(\gpio_out[1] ));
 sg13g2_dfrbp_1 \gpio_out[2]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net331),
    .D(_00002_),
    .Q_N(_05529_),
    .Q(\gpio_out[2] ));
 sg13g2_dfrbp_1 \gpio_out[3]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net332),
    .D(_00003_),
    .Q_N(_05530_),
    .Q(\gpio_out[3] ));
 sg13g2_dfrbp_1 \gpio_out[4]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net333),
    .D(_00004_),
    .Q_N(_05531_),
    .Q(\gpio_out[4] ));
 sg13g2_dfrbp_1 \gpio_out[5]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net334),
    .D(_00005_),
    .Q_N(_05532_),
    .Q(\gpio_out[5] ));
 sg13g2_dfrbp_1 \gpio_out[6]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net335),
    .D(_00006_),
    .Q_N(_05533_),
    .Q(\gpio_out[6] ));
 sg13g2_dfrbp_1 \gpio_out[7]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net336),
    .D(_00007_),
    .Q_N(_05534_),
    .Q(\gpio_out[7] ));
 sg13g2_dfrbp_1 \gpio_out_sel[0]$_DFF_P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net337),
    .D(_00008_),
    .Q_N(_05535_),
    .Q(\gpio_out_sel[0] ));
 sg13g2_dfrbp_1 \gpio_out_sel[1]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net338),
    .D(_00009_),
    .Q_N(_05536_),
    .Q(\gpio_out_sel[1] ));
 sg13g2_dfrbp_1 \gpio_out_sel[2]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net339),
    .D(_00010_),
    .Q_N(_05537_),
    .Q(\gpio_out_sel[2] ));
 sg13g2_dfrbp_1 \gpio_out_sel[3]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net340),
    .D(_00011_),
    .Q_N(_05538_),
    .Q(\gpio_out_sel[3] ));
 sg13g2_dfrbp_1 \gpio_out_sel[4]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net341),
    .D(_00012_),
    .Q_N(_05539_),
    .Q(\gpio_out_sel[4] ));
 sg13g2_dfrbp_1 \gpio_out_sel[5]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net342),
    .D(_00013_),
    .Q_N(_05540_),
    .Q(\gpio_out_sel[5] ));
 sg13g2_dfrbp_1 \gpio_out_sel[6]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net343),
    .D(_00014_),
    .Q_N(_05541_),
    .Q(\gpio_out_sel[6] ));
 sg13g2_dfrbp_1 \gpio_out_sel[7]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net344),
    .D(_00015_),
    .Q_N(_05515_),
    .Q(\gpio_out_sel[7] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net345),
    .D(_00229_),
    .Q_N(_00217_),
    .Q(\i_debug_uart_tx.cycle_counter[0] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net346),
    .D(_00230_),
    .Q_N(_05514_),
    .Q(\i_debug_uart_tx.cycle_counter[1] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net347),
    .D(_00231_),
    .Q_N(_05513_),
    .Q(\i_debug_uart_tx.cycle_counter[2] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net348),
    .D(_00232_),
    .Q_N(_05512_),
    .Q(\i_debug_uart_tx.cycle_counter[3] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net349),
    .D(_00233_),
    .Q_N(_00166_),
    .Q(\i_debug_uart_tx.cycle_counter[4] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net350),
    .D(_00234_),
    .Q_N(_05511_),
    .Q(\i_debug_uart_tx.data_to_send[0] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net351),
    .D(_00235_),
    .Q_N(_05510_),
    .Q(\i_debug_uart_tx.data_to_send[1] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net352),
    .D(_00236_),
    .Q_N(_05509_),
    .Q(\i_debug_uart_tx.data_to_send[2] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net353),
    .D(_00237_),
    .Q_N(_05508_),
    .Q(\i_debug_uart_tx.data_to_send[3] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net354),
    .D(_00238_),
    .Q_N(_05507_),
    .Q(\i_debug_uart_tx.data_to_send[4] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net355),
    .D(_00239_),
    .Q_N(_05506_),
    .Q(\i_debug_uart_tx.data_to_send[5] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net356),
    .D(_00240_),
    .Q_N(_05505_),
    .Q(\i_debug_uart_tx.data_to_send[6] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net357),
    .D(_00241_),
    .Q_N(_05504_),
    .Q(\i_debug_uart_tx.data_to_send[7] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.fsm_state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net358),
    .D(_00242_),
    .Q_N(_05503_),
    .Q(\i_debug_uart_tx.fsm_state[0] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.fsm_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net359),
    .D(_00243_),
    .Q_N(_05502_),
    .Q(\i_debug_uart_tx.fsm_state[1] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.fsm_state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net360),
    .D(_00244_),
    .Q_N(_05501_),
    .Q(\i_debug_uart_tx.fsm_state[2] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.fsm_state[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net361),
    .D(_00245_),
    .Q_N(_05500_),
    .Q(\i_debug_uart_tx.fsm_state[3] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.txd_reg$_SDFF_PN1_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net362),
    .D(_00246_),
    .Q_N(_05499_),
    .Q(debug_uart_txd));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net363),
    .D(_00247_),
    .Q_N(_05498_),
    .Q(\i_spi.bits_remaining[0] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net364),
    .D(_00248_),
    .Q_N(_05497_),
    .Q(\i_spi.bits_remaining[1] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net365),
    .D(_00249_),
    .Q_N(_05496_),
    .Q(\i_spi.bits_remaining[2] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net366),
    .D(_00250_),
    .Q_N(_05495_),
    .Q(\i_spi.bits_remaining[3] ));
 sg13g2_dfrbp_1 \i_spi.busy$_SDFF_PN0_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net367),
    .D(_00251_),
    .Q_N(_00167_),
    .Q(\i_spi.busy ));
 sg13g2_dfrbp_1 \i_spi.clock_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net368),
    .D(_00252_),
    .Q_N(_05494_),
    .Q(\i_spi.clock_count[0] ));
 sg13g2_dfrbp_1 \i_spi.clock_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net369),
    .D(_00253_),
    .Q_N(_05493_),
    .Q(\i_spi.clock_count[1] ));
 sg13g2_dfrbp_1 \i_spi.clock_divider[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net370),
    .D(_00254_),
    .Q_N(_05492_),
    .Q(\i_spi.clock_divider[0] ));
 sg13g2_dfrbp_1 \i_spi.clock_divider[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net371),
    .D(_00255_),
    .Q_N(_05491_),
    .Q(\i_spi.clock_divider[1] ));
 sg13g2_dfrbp_1 \i_spi.data[0]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net372),
    .D(_00256_),
    .Q_N(_05490_),
    .Q(\i_spi.data[0] ));
 sg13g2_dfrbp_1 \i_spi.data[1]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net373),
    .D(_00257_),
    .Q_N(_05489_),
    .Q(\i_spi.data[1] ));
 sg13g2_dfrbp_1 \i_spi.data[2]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net374),
    .D(_00258_),
    .Q_N(_05488_),
    .Q(\i_spi.data[2] ));
 sg13g2_dfrbp_1 \i_spi.data[3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net375),
    .D(_00259_),
    .Q_N(_05487_),
    .Q(\i_spi.data[3] ));
 sg13g2_dfrbp_1 \i_spi.data[4]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net376),
    .D(_00260_),
    .Q_N(_05486_),
    .Q(\i_spi.data[4] ));
 sg13g2_dfrbp_1 \i_spi.data[5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net377),
    .D(_00261_),
    .Q_N(_05485_),
    .Q(\i_spi.data[5] ));
 sg13g2_dfrbp_1 \i_spi.data[6]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net378),
    .D(_00262_),
    .Q_N(_05484_),
    .Q(\i_spi.data[6] ));
 sg13g2_dfrbp_1 \i_spi.data[7]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net379),
    .D(_00263_),
    .Q_N(_05483_),
    .Q(\i_spi.data[7] ));
 sg13g2_dfrbp_1 \i_spi.end_txn_reg$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net380),
    .D(_00264_),
    .Q_N(_05482_),
    .Q(\i_spi.end_txn_reg ));
 sg13g2_dfrbp_1 \i_spi.read_latency$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net381),
    .D(_00265_),
    .Q_N(_05481_),
    .Q(\i_spi.read_latency ));
 sg13g2_dfrbp_1 \i_spi.spi_clk_out$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net382),
    .D(_00266_),
    .Q_N(_05480_),
    .Q(\i_spi.spi_clk_out ));
 sg13g2_dfrbp_1 \i_spi.spi_dc$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net383),
    .D(_00267_),
    .Q_N(_05479_),
    .Q(\i_spi.spi_dc ));
 sg13g2_dfrbp_1 \i_spi.spi_select$_SDFFE_PN1P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net384),
    .D(_00268_),
    .Q_N(_05478_),
    .Q(\i_spi.spi_select ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.additional_mem_ops[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net385),
    .D(_00269_),
    .Q_N(_00212_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.additional_mem_ops[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net386),
    .D(_00270_),
    .Q_N(_05477_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.additional_mem_ops[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net387),
    .D(_00271_),
    .Q_N(_05476_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.alu_op[0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net388),
    .D(_00272_),
    .Q_N(_05475_),
    .Q(\i_tinyqv.cpu.alu_op[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.alu_op[1]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net389),
    .D(_00273_),
    .Q_N(_00089_),
    .Q(\i_tinyqv.cpu.alu_op[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.alu_op[2]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net390),
    .D(_00274_),
    .Q_N(_00094_),
    .Q(\i_tinyqv.cpu.alu_op[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.alu_op[3]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net391),
    .D(_00275_),
    .Q_N(_00085_),
    .Q(\i_tinyqv.cpu.alu_op[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.counter_hi[0]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net392),
    .D(_00276_),
    .Q_N(_00216_),
    .Q(\i_tinyqv.cpu.counter[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.counter_hi[1]$_SDFF_PN0_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net393),
    .D(_00277_),
    .Q_N(_00088_),
    .Q(\i_tinyqv.cpu.counter[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.counter_hi[2]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net394),
    .D(_00278_),
    .Q_N(_00084_),
    .Q(\i_tinyqv.cpu.counter[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net395),
    .D(_00279_),
    .Q_N(_05474_),
    .Q(\addr[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[10]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net396),
    .D(_00280_),
    .Q_N(_05473_),
    .Q(\addr[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[11]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net397),
    .D(_00281_),
    .Q_N(_05472_),
    .Q(\addr[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[12]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net398),
    .D(_00282_),
    .Q_N(_05471_),
    .Q(\addr[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[13]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net399),
    .D(_00283_),
    .Q_N(_05470_),
    .Q(\addr[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[14]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net400),
    .D(_00284_),
    .Q_N(_05469_),
    .Q(\addr[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[15]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net401),
    .D(_00285_),
    .Q_N(_05468_),
    .Q(\addr[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[16]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net402),
    .D(_00286_),
    .Q_N(_05467_),
    .Q(\addr[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[17]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net403),
    .D(_00287_),
    .Q_N(_05466_),
    .Q(\addr[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[18]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net404),
    .D(_00288_),
    .Q_N(_05465_),
    .Q(\addr[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[19]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net405),
    .D(_00289_),
    .Q_N(_05464_),
    .Q(\addr[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[1]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net406),
    .D(_00290_),
    .Q_N(_05463_),
    .Q(\addr[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[20]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net407),
    .D(_00291_),
    .Q_N(_05462_),
    .Q(\addr[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[21]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net408),
    .D(_00292_),
    .Q_N(_05461_),
    .Q(\addr[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[22]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net409),
    .D(_00293_),
    .Q_N(_05460_),
    .Q(\addr[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[23]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net410),
    .D(_00294_),
    .Q_N(_00159_),
    .Q(\addr[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net411),
    .D(_00295_),
    .Q_N(_05459_),
    .Q(\addr[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net412),
    .D(_00296_),
    .Q_N(_05458_),
    .Q(\addr[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net413),
    .D(_00297_),
    .Q_N(_05457_),
    .Q(\addr[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net414),
    .D(_00298_),
    .Q_N(_05456_),
    .Q(\addr[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[2]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net415),
    .D(_00299_),
    .Q_N(_05455_),
    .Q(\addr[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[3]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net416),
    .D(_00300_),
    .Q_N(_05454_),
    .Q(\addr[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[4]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net417),
    .D(_00301_),
    .Q_N(_05453_),
    .Q(\addr[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[5]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net418),
    .D(_00302_),
    .Q_N(_05452_),
    .Q(\addr[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[6]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net419),
    .D(_00303_),
    .Q_N(_05451_),
    .Q(\addr[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[7]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net420),
    .D(_00304_),
    .Q_N(_05450_),
    .Q(\addr[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[8]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net421),
    .D(_00305_),
    .Q_N(_05449_),
    .Q(\addr[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[9]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net422),
    .D(_00306_),
    .Q_N(_05542_),
    .Q(\addr[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_continue$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net423),
    .D(_00028_),
    .Q_N(_05448_),
    .Q(debug_data_continue));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net424),
    .D(_00307_),
    .Q_N(_05447_),
    .Q(\data_to_write[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[10]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net425),
    .D(_00308_),
    .Q_N(_05446_),
    .Q(\data_to_write[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[11]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net426),
    .D(_00309_),
    .Q_N(_05445_),
    .Q(\data_to_write[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[12]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net427),
    .D(_00310_),
    .Q_N(_05444_),
    .Q(\data_to_write[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[13]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net428),
    .D(_00311_),
    .Q_N(_05443_),
    .Q(\data_to_write[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[14]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net429),
    .D(_00312_),
    .Q_N(_05442_),
    .Q(\data_to_write[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[15]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net430),
    .D(_00313_),
    .Q_N(_05441_),
    .Q(\data_to_write[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[16]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net431),
    .D(_00314_),
    .Q_N(_05440_),
    .Q(\data_to_write[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[17]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net432),
    .D(_00315_),
    .Q_N(_05439_),
    .Q(\data_to_write[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[18]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net433),
    .D(_00316_),
    .Q_N(_05438_),
    .Q(\data_to_write[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[19]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net434),
    .D(_00317_),
    .Q_N(_05437_),
    .Q(\data_to_write[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net435),
    .D(_00318_),
    .Q_N(_05436_),
    .Q(\data_to_write[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[20]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net436),
    .D(_00319_),
    .Q_N(_05435_),
    .Q(\data_to_write[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[21]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net437),
    .D(_00320_),
    .Q_N(_05434_),
    .Q(\data_to_write[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[22]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net438),
    .D(_00321_),
    .Q_N(_05433_),
    .Q(\data_to_write[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[23]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net439),
    .D(_00322_),
    .Q_N(_05432_),
    .Q(\data_to_write[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[24]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net440),
    .D(_00323_),
    .Q_N(_05431_),
    .Q(\data_to_write[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[25]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net441),
    .D(_00324_),
    .Q_N(_05430_),
    .Q(\data_to_write[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[26]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net442),
    .D(_00325_),
    .Q_N(_05429_),
    .Q(\data_to_write[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[27]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net443),
    .D(_00326_),
    .Q_N(_05428_),
    .Q(\data_to_write[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[28]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net444),
    .D(_00327_),
    .Q_N(_05427_),
    .Q(\data_to_write[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[29]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net445),
    .D(_00328_),
    .Q_N(_05426_),
    .Q(\data_to_write[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net446),
    .D(_00329_),
    .Q_N(_05425_),
    .Q(\data_to_write[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[30]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net447),
    .D(_00330_),
    .Q_N(_05424_),
    .Q(\data_to_write[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[31]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net448),
    .D(_00331_),
    .Q_N(_05423_),
    .Q(\data_to_write[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net449),
    .D(_00332_),
    .Q_N(_05422_),
    .Q(\data_to_write[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net450),
    .D(_00333_),
    .Q_N(_05421_),
    .Q(\data_to_write[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net451),
    .D(_00334_),
    .Q_N(_05420_),
    .Q(\data_to_write[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net452),
    .D(_00335_),
    .Q_N(_05419_),
    .Q(\data_to_write[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net453),
    .D(_00336_),
    .Q_N(_00201_),
    .Q(\data_to_write[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[8]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net454),
    .D(_00337_),
    .Q_N(_05418_),
    .Q(\data_to_write[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net455),
    .D(_00338_),
    .Q_N(_05417_),
    .Q(\data_to_write[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_read_n[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net456),
    .D(_00339_),
    .Q_N(_05416_),
    .Q(\i_tinyqv.cpu.data_read_n[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_read_n[1]$_SDFFE_PP1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net457),
    .D(_00340_),
    .Q_N(_05415_),
    .Q(\i_tinyqv.cpu.data_read_n[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_ready_core$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net458),
    .D(_00341_),
    .Q_N(_05414_),
    .Q(\i_tinyqv.cpu.data_ready_core ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_ready_latch$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net459),
    .D(_00342_),
    .Q_N(_05413_),
    .Q(\i_tinyqv.cpu.data_ready_latch ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_write_n[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net460),
    .D(_00343_),
    .Q_N(_05412_),
    .Q(\i_tinyqv.cpu.data_write_n[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_write_n[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net461),
    .D(_00344_),
    .Q_N(_05543_),
    .Q(\i_tinyqv.cpu.data_write_n[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.cmp$_DFF_P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net462),
    .D(\i_tinyqv.cpu.i_core.cmp_out ),
    .Q_N(_05544_),
    .Q(\i_tinyqv.cpu.i_core.cmp ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.cy$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net463),
    .D(\i_tinyqv.cpu.i_core.cy_out ),
    .Q_N(_00092_),
    .Q(\i_tinyqv.cpu.i_core.cy ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.cycle[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net464),
    .D(_00345_),
    .Q_N(_00086_),
    .Q(\i_tinyqv.cpu.i_core.cycle[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.cycle[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net465),
    .D(_00346_),
    .Q_N(_05411_),
    .Q(\i_tinyqv.cpu.i_core.cycle[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.cy$_SDFF_PN0_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net466),
    .D(_00347_),
    .Q_N(_05410_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.cy ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[0]$_SDFF_PN0_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net467),
    .D(_00348_),
    .Q_N(_05545_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[10]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net468),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ),
    .Q_N(_05546_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[11]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net469),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ),
    .Q_N(_05547_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[12]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net470),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ),
    .Q_N(_05548_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[13]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net471),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ),
    .Q_N(_05549_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[14]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net472),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ),
    .Q_N(_05550_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[15]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net473),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ),
    .Q_N(_05551_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[16]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net474),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ),
    .Q_N(_05552_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[17]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net475),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ),
    .Q_N(_05553_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[18]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net476),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ),
    .Q_N(_05554_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[19]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net477),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ),
    .Q_N(_05409_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[1]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net478),
    .D(_00349_),
    .Q_N(_05555_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[20]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net479),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ),
    .Q_N(_05556_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[21]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net480),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ),
    .Q_N(_05557_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[22]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net481),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ),
    .Q_N(_05558_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[23]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net482),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ),
    .Q_N(_05559_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[24]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net483),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ),
    .Q_N(_05560_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[25]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net484),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ),
    .Q_N(_05561_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[26]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net485),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ),
    .Q_N(_05562_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[27]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net486),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ),
    .Q_N(_05563_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[28]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net487),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ),
    .Q_N(_05564_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[29]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net488),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ),
    .Q_N(_05408_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[2]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net489),
    .D(_00350_),
    .Q_N(_05565_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[30]$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net490),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ),
    .Q_N(_05566_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[31]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net491),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ),
    .Q_N(_05407_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[3]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net492),
    .D(_00351_),
    .Q_N(_05567_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[4]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net493),
    .D(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .Q_N(_05568_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[5]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net494),
    .D(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .Q_N(_05569_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[6]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net495),
    .D(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .Q_N(_05570_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[7]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net496),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ),
    .Q_N(_05571_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[8]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net497),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ),
    .Q_N(_05572_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[9]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net498),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ),
    .Q_N(_05406_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.cy$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net499),
    .D(_00352_),
    .Q_N(_00215_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.cy ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[0]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net500),
    .D(_00353_),
    .Q_N(_05573_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[10]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net501),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ),
    .Q_N(_05574_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[11]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net502),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ),
    .Q_N(_05575_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[12]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net503),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ),
    .Q_N(_05576_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[13]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net504),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ),
    .Q_N(_05577_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[14]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net505),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ),
    .Q_N(_05578_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[15]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net506),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ),
    .Q_N(_05579_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[16]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net507),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ),
    .Q_N(_05580_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[17]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net508),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ),
    .Q_N(_05581_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[18]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net509),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ),
    .Q_N(_05582_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[19]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net510),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ),
    .Q_N(_05405_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[1]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net511),
    .D(_00354_),
    .Q_N(_05583_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[20]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net512),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ),
    .Q_N(_05584_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[21]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net513),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ),
    .Q_N(_05585_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[22]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net514),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ),
    .Q_N(_05586_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[23]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net515),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ),
    .Q_N(_05587_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[24]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net516),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ),
    .Q_N(_05588_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[25]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net517),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ),
    .Q_N(_05589_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[26]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net518),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ),
    .Q_N(_05590_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[27]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net519),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ),
    .Q_N(_05591_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[28]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net520),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ),
    .Q_N(_05592_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[29]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net521),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ),
    .Q_N(_05404_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[2]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net522),
    .D(_00355_),
    .Q_N(_05593_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[30]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net523),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ),
    .Q_N(_05594_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[31]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net524),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ),
    .Q_N(_05403_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[3]$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net525),
    .D(_00356_),
    .Q_N(_05595_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[4]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net526),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ),
    .Q_N(_00168_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[5]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net527),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ),
    .Q_N(_05596_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[6]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net528),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ),
    .Q_N(_05597_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[7]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net529),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ),
    .Q_N(_05598_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[8]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net530),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ),
    .Q_N(_05599_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[9]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net531),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ),
    .Q_N(_05600_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][0]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net532),
    .D(_00030_),
    .Q_N(_05601_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][10]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net533),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05602_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][11]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net534),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05603_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][12]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net535),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05604_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][13]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net536),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05605_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][14]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net537),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05606_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][15]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net538),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05607_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][16]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net539),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05608_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][17]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net540),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05609_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][18]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net541),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05610_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][19]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net542),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05611_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][1]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net543),
    .D(_00031_),
    .Q_N(_05612_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][20]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net544),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05613_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][21]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net545),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05614_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][22]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net546),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05615_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][23]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net547),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05616_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][24]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net548),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05617_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][25]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net549),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05618_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][26]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net550),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05619_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][27]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net551),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05620_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][28]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net552),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05621_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][29]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net553),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05622_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][2]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net554),
    .D(_00032_),
    .Q_N(_05623_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][30]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net555),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05624_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][31]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net556),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05625_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][3]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net557),
    .D(_00033_),
    .Q_N(_05626_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][4]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net558),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05627_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][5]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net559),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05628_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][6]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net560),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05629_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][7]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net561),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05630_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][8]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net562),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05631_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][9]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net563),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05632_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][0]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net564),
    .D(_00034_),
    .Q_N(_05633_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][10]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net565),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05634_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][11]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net566),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05635_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][12]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net567),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05636_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][13]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net568),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05637_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][14]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net569),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05638_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][15]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net570),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05639_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][16]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net571),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05640_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][17]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net572),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05641_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][18]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net573),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05642_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][19]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net574),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05643_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][1]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net575),
    .D(_00035_),
    .Q_N(_05644_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][20]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net576),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05645_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][21]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net577),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05646_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][22]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net578),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05647_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][23]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net579),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05648_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][24]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net580),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05649_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][25]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net581),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05650_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][26]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net582),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05651_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][27]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net583),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05652_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][28]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net584),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05653_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][29]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net585),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05654_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][2]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net586),
    .D(_00036_),
    .Q_N(_05655_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][30]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net587),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05656_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][31]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net588),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05657_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][3]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net589),
    .D(_00037_),
    .Q_N(_05658_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][4]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net590),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05659_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][5]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net591),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05660_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][6]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net592),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05661_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][7]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net593),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05662_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][8]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net594),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05663_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][9]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net595),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05664_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][0]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net596),
    .D(_00038_),
    .Q_N(_05665_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][10]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net597),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05666_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][11]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net598),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05667_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][12]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net599),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05668_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][13]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net600),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05669_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][14]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net601),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05670_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][15]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net602),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05671_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][16]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net603),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05672_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][17]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net604),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05673_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][18]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net605),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05674_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][19]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net606),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05675_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][1]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net607),
    .D(_00039_),
    .Q_N(_05676_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][20]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net608),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05677_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][21]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net609),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05678_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][22]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net610),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05679_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][23]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net611),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05680_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][24]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net612),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05681_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][25]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net613),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05682_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][26]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net614),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05683_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][27]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net615),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05684_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][28]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net616),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05685_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][29]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net617),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05686_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][2]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net618),
    .D(_00040_),
    .Q_N(_05687_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][30]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net619),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05688_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][31]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net620),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05689_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][3]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net621),
    .D(_00041_),
    .Q_N(_05690_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][4]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net622),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05691_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][5]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net623),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05692_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][6]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net624),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05693_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][7]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net625),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05694_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][8]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net626),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05695_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][9]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net627),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05696_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][0]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net628),
    .D(_00042_),
    .Q_N(_05697_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][10]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net629),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05698_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][11]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net630),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05699_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][12]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net631),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05700_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][13]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net632),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05701_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][14]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net633),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05702_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][15]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net634),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05703_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][16]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net635),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05704_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][17]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net636),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05705_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][18]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net637),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05706_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][19]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net638),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05707_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][1]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net639),
    .D(_00043_),
    .Q_N(_05708_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][20]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net640),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05709_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][21]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net641),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05710_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][22]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net642),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05711_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][23]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net643),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05712_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][24]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net644),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05713_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][25]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net645),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05714_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][26]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net646),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05715_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][27]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net647),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05716_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][28]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net648),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05717_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][29]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net649),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05718_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][2]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net650),
    .D(_00044_),
    .Q_N(_05719_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][30]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net651),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05720_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][31]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net652),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05721_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][3]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net653),
    .D(_00045_),
    .Q_N(_05722_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][4]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net654),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05723_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][5]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net655),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05724_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][6]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net656),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05725_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][7]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net657),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05726_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][8]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net658),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05727_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][9]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net659),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05728_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][0]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net660),
    .D(_00046_),
    .Q_N(_05729_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][10]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net661),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05730_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][11]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net662),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05731_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][12]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net663),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05732_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][13]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net664),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05733_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][14]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net665),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05734_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][15]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net666),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05735_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][16]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net667),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05736_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][17]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net668),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05737_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][18]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net669),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05738_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][19]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net670),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05739_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][1]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net671),
    .D(_00047_),
    .Q_N(_05740_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][20]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net672),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05741_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][21]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net673),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05742_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][22]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net674),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05743_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][23]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net675),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05744_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][24]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net676),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05745_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][25]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net677),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05746_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][26]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net678),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05747_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][27]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net679),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05748_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][28]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net680),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05749_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][29]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net681),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05750_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][2]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net682),
    .D(_00048_),
    .Q_N(_05751_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][30]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net683),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05752_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][31]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net684),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05753_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][3]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net685),
    .D(_00049_),
    .Q_N(_05754_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][4]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net686),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05755_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][5]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net687),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05756_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][6]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net688),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05757_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][7]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net689),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05758_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][8]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net690),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05759_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][9]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net691),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05760_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][0]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net692),
    .D(_00050_),
    .Q_N(_05761_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][10]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net693),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05762_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][11]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net694),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05763_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][12]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net695),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05764_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][13]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net696),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05765_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][14]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net697),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05766_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][15]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net698),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05767_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][16]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net699),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05768_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][17]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net700),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05769_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][18]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net701),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05770_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][19]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net702),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05771_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][1]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net703),
    .D(_00051_),
    .Q_N(_05772_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][20]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net704),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05773_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][21]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net705),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05774_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][22]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net706),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05775_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][23]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net707),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05776_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][24]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net708),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05777_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][25]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net709),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05778_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][26]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net710),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05779_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][27]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net711),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05780_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][28]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net712),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05781_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][29]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net713),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05782_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][2]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net714),
    .D(_00052_),
    .Q_N(_05783_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][30]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net715),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05784_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][31]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net716),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05785_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][3]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net717),
    .D(_00053_),
    .Q_N(_05786_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][4]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net718),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05787_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][5]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net719),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_00091_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][6]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net720),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_00090_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][7]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net721),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_00087_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][8]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net722),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05788_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][9]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net723),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05789_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][0]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net724),
    .D(_00054_),
    .Q_N(_05790_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][10]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net725),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05791_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][11]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net726),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05792_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][12]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net727),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05793_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][13]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net728),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05794_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][14]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net729),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05795_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][15]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net730),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05796_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][16]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net731),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05797_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][17]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net732),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05798_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][18]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net733),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05799_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][19]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net734),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05800_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][1]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net735),
    .D(_00055_),
    .Q_N(_05801_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][20]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net736),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05802_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][21]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net737),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05803_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][22]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net738),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05804_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][23]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net739),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05805_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][24]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net740),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05806_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][25]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net741),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05807_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][26]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net742),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05808_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][27]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net743),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05809_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][28]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net744),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05810_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][29]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net745),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05811_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][2]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net746),
    .D(_00056_),
    .Q_N(_05812_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][30]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net747),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05813_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][31]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net748),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05814_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][3]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net749),
    .D(_00057_),
    .Q_N(_05815_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][4]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net750),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05816_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][5]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net751),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05817_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][6]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net752),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05818_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][7]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net753),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05819_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][8]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net754),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05820_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][9]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net755),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05821_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][0]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net756),
    .D(_00058_),
    .Q_N(_05822_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][10]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net757),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05823_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][11]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net758),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05824_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][12]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net759),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05825_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][13]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net760),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05826_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][14]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net761),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05827_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][15]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net762),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05828_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][16]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net763),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05829_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][17]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net764),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05830_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][18]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net765),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05831_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][19]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net766),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05832_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][1]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net767),
    .D(_00059_),
    .Q_N(_05833_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][20]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net768),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05834_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][21]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net769),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05835_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][22]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net770),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05836_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][23]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net771),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05837_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][24]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net772),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05838_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][25]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net773),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05839_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][26]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net774),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05840_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][27]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net775),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05841_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][28]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net776),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05842_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][29]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net777),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05843_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][2]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net778),
    .D(_00060_),
    .Q_N(_05844_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][30]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net779),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05845_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][31]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net780),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05846_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][3]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net781),
    .D(_00061_),
    .Q_N(_05847_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][4]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net782),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05848_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][5]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net783),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05849_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][6]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net784),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05850_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][7]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net785),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05851_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][8]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net786),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05852_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][9]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net787),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05853_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][0]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net788),
    .D(_00062_),
    .Q_N(_05854_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][10]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net789),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05855_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][11]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net790),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05856_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][12]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net791),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05857_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][13]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net792),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05858_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][14]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net793),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05859_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][15]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net794),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05860_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][16]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net795),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05861_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][17]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net796),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05862_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][18]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net797),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05863_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][19]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net798),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05864_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][1]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net799),
    .D(_00063_),
    .Q_N(_05865_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][20]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net800),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05866_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][21]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net801),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05867_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][22]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net802),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05868_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][23]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net803),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05869_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][24]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net804),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05870_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][25]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net805),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05871_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][26]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net806),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05872_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][27]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net807),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05873_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][28]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net808),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05874_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][29]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net809),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05875_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][2]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net810),
    .D(_00064_),
    .Q_N(_05876_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][30]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net811),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05877_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][31]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net812),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05878_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][3]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net813),
    .D(_00065_),
    .Q_N(_05879_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][4]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net814),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05880_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][5]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net815),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05881_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][6]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net816),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05882_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][7]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net817),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05883_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][8]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net818),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05884_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][9]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net819),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05885_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][0]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net820),
    .D(_00066_),
    .Q_N(_05886_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][10]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net821),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05887_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][11]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net822),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05888_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][12]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net823),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05889_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][13]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net824),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05890_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][14]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net825),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05891_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][15]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net826),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05892_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][16]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net827),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05893_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][17]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net828),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05894_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][18]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net829),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05895_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][19]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net830),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05896_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][1]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net831),
    .D(_00067_),
    .Q_N(_05897_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][20]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net832),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05898_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][21]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net833),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05899_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][22]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net834),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05900_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][23]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net835),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05901_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][24]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net836),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05902_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][25]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net837),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05903_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][26]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net838),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05904_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][27]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net839),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05905_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][28]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net840),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05906_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][29]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net841),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05907_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][2]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net842),
    .D(_00068_),
    .Q_N(_05908_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][30]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net843),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05909_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][31]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net844),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05910_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][3]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net845),
    .D(_00069_),
    .Q_N(_05911_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][4]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net846),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05912_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][5]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net847),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05913_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][6]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net848),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05914_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][7]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net849),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05915_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][8]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net850),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05916_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][9]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net851),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05917_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][0]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net852),
    .D(_00070_),
    .Q_N(_05918_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][10]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net853),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05919_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][11]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net854),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05920_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][12]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net855),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05921_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][13]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net856),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05922_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][14]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net857),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05923_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][15]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net858),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05924_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][16]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net859),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05925_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][17]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net860),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05926_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][18]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net861),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05927_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][19]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net862),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05928_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][1]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net863),
    .D(_00071_),
    .Q_N(_05929_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][20]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net864),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05930_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][21]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net865),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05931_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][22]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net866),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05932_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][23]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net867),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05933_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][24]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net868),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05934_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][25]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net869),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05935_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][26]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net870),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05936_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][27]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net871),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05937_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][28]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net872),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05938_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][29]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net873),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05939_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][2]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net874),
    .D(_00072_),
    .Q_N(_05940_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][30]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net875),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05941_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][31]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net876),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05942_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][3]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net877),
    .D(_00073_),
    .Q_N(_05943_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][4]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net878),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05944_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][5]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net879),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05945_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][6]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net880),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05946_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][7]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net881),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05947_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][8]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net882),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05948_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][9]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net883),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05949_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][0]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net884),
    .D(_00074_),
    .Q_N(_05950_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][10]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net885),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05951_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][11]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net886),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05952_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][12]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net887),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05953_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][13]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net888),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05954_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][14]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net889),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05955_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][15]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net890),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05956_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][16]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net891),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05957_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][17]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net892),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05958_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][18]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net893),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05959_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][19]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net894),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05960_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][1]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net895),
    .D(_00075_),
    .Q_N(_05961_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][20]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net896),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05962_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][21]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net897),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05963_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][22]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net898),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05964_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][23]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net899),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05965_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][24]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net900),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05966_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][25]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net901),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05967_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][26]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net902),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05968_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][27]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net903),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05969_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][28]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net904),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05970_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][29]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net905),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05971_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][2]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net906),
    .D(_00076_),
    .Q_N(_05972_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][30]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net907),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05973_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][31]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net908),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05974_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][3]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net909),
    .D(_00077_),
    .Q_N(_05975_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][4]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net910),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05976_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][5]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net911),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05977_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][6]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net912),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05978_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][7]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net913),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05979_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][8]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net914),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05980_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][9]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net915),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05981_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][0]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net916),
    .D(_00078_),
    .Q_N(_05982_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][10]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net917),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05983_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][11]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net918),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05984_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][12]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net919),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05985_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][13]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net920),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05986_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][14]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net921),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05987_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][15]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net922),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05988_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][16]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net923),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05989_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][17]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net924),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05990_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][18]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net925),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05991_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][19]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net926),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05992_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][1]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net927),
    .D(_00079_),
    .Q_N(_05993_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][20]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net928),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05994_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][21]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net929),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05995_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][22]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net930),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05996_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][23]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net931),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05997_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][24]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net932),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05998_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][25]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net933),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05999_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][26]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net934),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_06000_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][27]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net935),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_06001_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][28]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net936),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_06002_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][29]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net937),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_06003_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][2]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net938),
    .D(_00080_),
    .Q_N(_06004_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][30]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net939),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_06005_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][31]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net940),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_06006_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][3]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net941),
    .D(_00081_),
    .Q_N(_06007_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][4]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net942),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_06008_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][5]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net943),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_06009_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][6]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net944),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_06010_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][7]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net945),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_06011_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][8]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net946),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_06012_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][9]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net947),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_06013_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.instr_retired$_DFF_P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net948),
    .D(_00029_),
    .Q_N(_00214_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.add ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.is_double_fault_r$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net949),
    .D(_00357_),
    .Q_N(_05402_),
    .Q(\i_tinyqv.cpu.i_core.is_double_fault_r ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.last_interrupt_req[0]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net950),
    .D(_00358_),
    .Q_N(_05401_),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.last_interrupt_req[1]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net951),
    .D(_00359_),
    .Q_N(_05400_),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.load_done$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net952),
    .D(_00360_),
    .Q_N(_05399_),
    .Q(\i_tinyqv.cpu.i_core.load_done ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.load_top_bit$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net953),
    .D(_00361_),
    .Q_N(_05398_),
    .Q(\i_tinyqv.cpu.i_core.load_top_bit ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mcause[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net954),
    .D(_00362_),
    .Q_N(_05397_),
    .Q(\i_tinyqv.cpu.i_core.mcause[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mcause[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net955),
    .D(_00363_),
    .Q_N(_05396_),
    .Q(\i_tinyqv.cpu.i_core.mcause[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mcause[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net956),
    .D(_00364_),
    .Q_N(_05395_),
    .Q(\i_tinyqv.cpu.i_core.mcause[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mcause[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net957),
    .D(_00365_),
    .Q_N(_05394_),
    .Q(\i_tinyqv.cpu.i_core.mcause[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[0]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net958),
    .D(_00366_),
    .Q_N(_05393_),
    .Q(\i_tinyqv.cpu.i_core.mepc[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[10]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net959),
    .D(_00367_),
    .Q_N(_05392_),
    .Q(\i_tinyqv.cpu.i_core.mepc[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[11]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net960),
    .D(_00368_),
    .Q_N(_05391_),
    .Q(\i_tinyqv.cpu.i_core.mepc[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[12]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net961),
    .D(_00369_),
    .Q_N(_05390_),
    .Q(\i_tinyqv.cpu.i_core.mepc[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[13]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net962),
    .D(_00370_),
    .Q_N(_05389_),
    .Q(\i_tinyqv.cpu.i_core.mepc[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[14]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net963),
    .D(_00371_),
    .Q_N(_05388_),
    .Q(\i_tinyqv.cpu.i_core.mepc[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[15]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net964),
    .D(_00372_),
    .Q_N(_05387_),
    .Q(\i_tinyqv.cpu.i_core.mepc[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[16]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net965),
    .D(_00373_),
    .Q_N(_05386_),
    .Q(\i_tinyqv.cpu.i_core.mepc[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[17]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net966),
    .D(_00374_),
    .Q_N(_05385_),
    .Q(\i_tinyqv.cpu.i_core.mepc[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[18]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net967),
    .D(_00375_),
    .Q_N(_05384_),
    .Q(\i_tinyqv.cpu.i_core.mepc[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[19]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net968),
    .D(_00376_),
    .Q_N(_05383_),
    .Q(\i_tinyqv.cpu.i_core.mepc[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[1]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net969),
    .D(_00377_),
    .Q_N(_05382_),
    .Q(\i_tinyqv.cpu.i_core.mepc[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[20]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net970),
    .D(_00378_),
    .Q_N(_05381_),
    .Q(\i_tinyqv.cpu.i_core.mepc[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[21]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net971),
    .D(_00379_),
    .Q_N(_05380_),
    .Q(\i_tinyqv.cpu.i_core.mepc[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[22]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net972),
    .D(_00380_),
    .Q_N(_05379_),
    .Q(\i_tinyqv.cpu.i_core.mepc[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[23]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net973),
    .D(_00381_),
    .Q_N(_05378_),
    .Q(\i_tinyqv.cpu.i_core.mepc[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[2]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net974),
    .D(_00382_),
    .Q_N(_05377_),
    .Q(\i_tinyqv.cpu.i_core.mepc[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[3]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net975),
    .D(_00383_),
    .Q_N(_05376_),
    .Q(\i_tinyqv.cpu.i_core.mepc[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[4]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net976),
    .D(_00384_),
    .Q_N(_05375_),
    .Q(\i_tinyqv.cpu.i_core.mepc[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[5]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net977),
    .D(_00385_),
    .Q_N(_05374_),
    .Q(\i_tinyqv.cpu.i_core.mepc[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[6]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net978),
    .D(_00386_),
    .Q_N(_05373_),
    .Q(\i_tinyqv.cpu.i_core.mepc[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[7]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net979),
    .D(_00387_),
    .Q_N(_05372_),
    .Q(\i_tinyqv.cpu.i_core.mepc[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[8]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net980),
    .D(_00388_),
    .Q_N(_05371_),
    .Q(\i_tinyqv.cpu.i_core.mepc[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[9]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net981),
    .D(_00389_),
    .Q_N(_05370_),
    .Q(\i_tinyqv.cpu.i_core.mepc[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mstatus_mie$_SDFFE_PP1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net982),
    .D(_00390_),
    .Q_N(_05369_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mie ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mstatus_mpie$_SDFFE_PP0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net983),
    .D(_00391_),
    .Q_N(_05368_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mpie ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mstatus_mte$_SDFFE_PP1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net984),
    .D(_00392_),
    .Q_N(_06014_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mte ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[0]$_DFF_P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net985),
    .D(_00016_),
    .Q_N(_06015_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[10]$_DFF_P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net986),
    .D(_00017_),
    .Q_N(_06016_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[11]$_DFF_P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net987),
    .D(_00018_),
    .Q_N(_05367_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[12]$_SDFF_PP0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net988),
    .D(_00393_),
    .Q_N(_05366_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[13]$_SDFF_PP0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net989),
    .D(_00394_),
    .Q_N(_05365_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[14]$_SDFF_PP0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net990),
    .D(_00395_),
    .Q_N(_05364_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[15]$_SDFF_PP0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net991),
    .D(_00396_),
    .Q_N(_06017_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[1]$_DFF_P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net992),
    .D(_00019_),
    .Q_N(_06018_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[2]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net993),
    .D(_00020_),
    .Q_N(_06019_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[3]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net994),
    .D(_00021_),
    .Q_N(_06020_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[4]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net995),
    .D(_00022_),
    .Q_N(_06021_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[5]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net996),
    .D(_00023_),
    .Q_N(_06022_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[6]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net997),
    .D(_00024_),
    .Q_N(_06023_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[7]$_DFF_P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net998),
    .D(_00025_),
    .Q_N(_06024_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[8]$_DFF_P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net999),
    .D(_00026_),
    .Q_N(_06025_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[9]$_DFF_P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1000),
    .D(_00027_),
    .Q_N(_05363_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[0]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1001),
    .D(_00397_),
    .Q_N(_05362_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[1]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1002),
    .D(_00398_),
    .Q_N(_05361_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[2]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1003),
    .D(_00399_),
    .Q_N(_05360_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[3]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1004),
    .D(_00400_),
    .Q_N(_05359_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[4]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1005),
    .D(_00401_),
    .Q_N(_05358_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.time_hi[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1006),
    .D(_00402_),
    .Q_N(_00218_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.time_hi[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1007),
    .D(_00403_),
    .Q_N(_05357_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.time_hi[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1008),
    .D(_00404_),
    .Q_N(_05356_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[0]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1009),
    .D(_00405_),
    .Q_N(_00169_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[10]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1010),
    .D(_00406_),
    .Q_N(_00184_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[11]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1011),
    .D(_00407_),
    .Q_N(_00186_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[12]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1012),
    .D(_00408_),
    .Q_N(_00188_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[13]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1013),
    .D(_00409_),
    .Q_N(_00190_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[14]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1014),
    .D(_00410_),
    .Q_N(_00192_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[15]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1015),
    .D(_00411_),
    .Q_N(_00194_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[16]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1016),
    .D(_00412_),
    .Q_N(_00195_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[17]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1017),
    .D(_00413_),
    .Q_N(_00193_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[18]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1018),
    .D(_00414_),
    .Q_N(_00191_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[19]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1019),
    .D(_00415_),
    .Q_N(_00189_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[1]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1020),
    .D(_00416_),
    .Q_N(_00198_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[20]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1021),
    .D(_00417_),
    .Q_N(_00187_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[21]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1022),
    .D(_00418_),
    .Q_N(_00185_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[22]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1023),
    .D(_00419_),
    .Q_N(_00183_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[23]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1024),
    .D(_00420_),
    .Q_N(_00181_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[24]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1025),
    .D(_00421_),
    .Q_N(_00179_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[25]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1026),
    .D(_00422_),
    .Q_N(_00177_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[26]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1027),
    .D(_00423_),
    .Q_N(_00175_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[27]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1028),
    .D(_00424_),
    .Q_N(_00173_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[28]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1029),
    .D(_00425_),
    .Q_N(_00171_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[29]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1030),
    .D(_00426_),
    .Q_N(_00197_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[2]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1031),
    .D(_00427_),
    .Q_N(_00196_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[30]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1032),
    .D(_00428_),
    .Q_N(_00199_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[31]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1033),
    .D(_00429_),
    .Q_N(_00200_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[3]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1034),
    .D(_00430_),
    .Q_N(_00170_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[4]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1035),
    .D(_00431_),
    .Q_N(_00172_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[5]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1036),
    .D(_00432_),
    .Q_N(_00174_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[6]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1037),
    .D(_00433_),
    .Q_N(_00176_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[7]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1038),
    .D(_00434_),
    .Q_N(_00178_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[8]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1039),
    .D(_00435_),
    .Q_N(_00180_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[9]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1040),
    .D(_00436_),
    .Q_N(_00182_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1041),
    .D(_00437_),
    .Q_N(_05355_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1042),
    .D(_00438_),
    .Q_N(_05354_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1043),
    .D(_00439_),
    .Q_N(_05353_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1044),
    .D(_00440_),
    .Q_N(_05352_),
    .Q(\i_tinyqv.cpu.imm[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1045),
    .D(_00441_),
    .Q_N(_05351_),
    .Q(\i_tinyqv.cpu.imm[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1046),
    .D(_00442_),
    .Q_N(_05350_),
    .Q(\i_tinyqv.cpu.imm[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1047),
    .D(_00443_),
    .Q_N(_05349_),
    .Q(\i_tinyqv.cpu.imm[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[16]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1048),
    .D(_00444_),
    .Q_N(_05348_),
    .Q(\i_tinyqv.cpu.imm[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[17]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1049),
    .D(_00445_),
    .Q_N(_05347_),
    .Q(\i_tinyqv.cpu.imm[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[18]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1050),
    .D(_00446_),
    .Q_N(_05346_),
    .Q(\i_tinyqv.cpu.imm[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[19]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1051),
    .D(_00447_),
    .Q_N(_05345_),
    .Q(\i_tinyqv.cpu.imm[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1052),
    .D(_00448_),
    .Q_N(_05344_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[20]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1053),
    .D(_00449_),
    .Q_N(_05343_),
    .Q(\i_tinyqv.cpu.imm[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[21]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1054),
    .D(_00450_),
    .Q_N(_05342_),
    .Q(\i_tinyqv.cpu.imm[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[22]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1055),
    .D(_00451_),
    .Q_N(_05341_),
    .Q(\i_tinyqv.cpu.imm[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[23]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1056),
    .D(_00452_),
    .Q_N(_05340_),
    .Q(\i_tinyqv.cpu.imm[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[24]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1057),
    .D(_00453_),
    .Q_N(_05339_),
    .Q(\i_tinyqv.cpu.imm[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[25]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1058),
    .D(_00454_),
    .Q_N(_05338_),
    .Q(\i_tinyqv.cpu.imm[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[26]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1059),
    .D(_00455_),
    .Q_N(_05337_),
    .Q(\i_tinyqv.cpu.imm[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[27]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1060),
    .D(_00456_),
    .Q_N(_05336_),
    .Q(\i_tinyqv.cpu.imm[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[28]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1061),
    .D(_00457_),
    .Q_N(_05335_),
    .Q(\i_tinyqv.cpu.imm[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[29]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1062),
    .D(_00458_),
    .Q_N(_05334_),
    .Q(\i_tinyqv.cpu.imm[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1063),
    .D(_00459_),
    .Q_N(_05333_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[30]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1064),
    .D(_00460_),
    .Q_N(_05332_),
    .Q(\i_tinyqv.cpu.imm[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1065),
    .D(_00461_),
    .Q_N(_05331_),
    .Q(\i_tinyqv.cpu.imm[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1066),
    .D(_00462_),
    .Q_N(_05330_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1067),
    .D(_00463_),
    .Q_N(_05329_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1068),
    .D(_00464_),
    .Q_N(_05328_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1069),
    .D(_00465_),
    .Q_N(_05327_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1070),
    .D(_00466_),
    .Q_N(_05326_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1071),
    .D(_00467_),
    .Q_N(_05325_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1072),
    .D(_00468_),
    .Q_N(_05324_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][0]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1073),
    .D(_00469_),
    .Q_N(_05323_),
    .Q(\i_tinyqv.cpu.instr_data[0][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1074),
    .D(_00470_),
    .Q_N(_00143_),
    .Q(\i_tinyqv.cpu.instr_data[0][10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1075),
    .D(_00471_),
    .Q_N(_00151_),
    .Q(\i_tinyqv.cpu.instr_data[0][11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1076),
    .D(_00472_),
    .Q_N(_00147_),
    .Q(\i_tinyqv.cpu.instr_data[0][12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1077),
    .D(_00473_),
    .Q_N(_00119_),
    .Q(\i_tinyqv.cpu.instr_data[0][13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1078),
    .D(_00474_),
    .Q_N(_00123_),
    .Q(\i_tinyqv.cpu.instr_data[0][14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1079),
    .D(_00475_),
    .Q_N(_00127_),
    .Q(\i_tinyqv.cpu.instr_data[0][15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1080),
    .D(_00476_),
    .Q_N(_00103_),
    .Q(\i_tinyqv.cpu.instr_data[0][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1081),
    .D(_00477_),
    .Q_N(_05322_),
    .Q(\i_tinyqv.cpu.instr_data[0][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1082),
    .D(_00478_),
    .Q_N(_05321_),
    .Q(\i_tinyqv.cpu.instr_data[0][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1083),
    .D(_00479_),
    .Q_N(_00107_),
    .Q(\i_tinyqv.cpu.instr_data[0][4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1084),
    .D(_00480_),
    .Q_N(_00111_),
    .Q(\i_tinyqv.cpu.instr_data[0][5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1085),
    .D(_00481_),
    .Q_N(_00115_),
    .Q(\i_tinyqv.cpu.instr_data[0][6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1086),
    .D(_00482_),
    .Q_N(_00131_),
    .Q(\i_tinyqv.cpu.instr_data[0][7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1087),
    .D(_00483_),
    .Q_N(_00135_),
    .Q(\i_tinyqv.cpu.instr_data[0][8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1088),
    .D(_00484_),
    .Q_N(_00139_),
    .Q(\i_tinyqv.cpu.instr_data[0][9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][0]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1089),
    .D(_00485_),
    .Q_N(_05320_),
    .Q(\i_tinyqv.cpu.instr_data[1][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1090),
    .D(_00486_),
    .Q_N(_00142_),
    .Q(\i_tinyqv.cpu.instr_data[1][10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1091),
    .D(_00487_),
    .Q_N(_00150_),
    .Q(\i_tinyqv.cpu.instr_data[1][11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1092),
    .D(_00488_),
    .Q_N(_00146_),
    .Q(\i_tinyqv.cpu.instr_data[1][12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1093),
    .D(_00489_),
    .Q_N(_00118_),
    .Q(\i_tinyqv.cpu.instr_data[1][13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1094),
    .D(_00490_),
    .Q_N(_00122_),
    .Q(\i_tinyqv.cpu.instr_data[1][14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1095),
    .D(_00491_),
    .Q_N(_00126_),
    .Q(\i_tinyqv.cpu.instr_data[1][15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1096),
    .D(_00492_),
    .Q_N(_00102_),
    .Q(\i_tinyqv.cpu.instr_data[1][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1097),
    .D(_00493_),
    .Q_N(_05319_),
    .Q(\i_tinyqv.cpu.instr_data[1][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1098),
    .D(_00494_),
    .Q_N(_05318_),
    .Q(\i_tinyqv.cpu.instr_data[1][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1099),
    .D(_00495_),
    .Q_N(_00106_),
    .Q(\i_tinyqv.cpu.instr_data[1][4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1100),
    .D(_00496_),
    .Q_N(_00110_),
    .Q(\i_tinyqv.cpu.instr_data[1][5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1101),
    .D(_00497_),
    .Q_N(_00114_),
    .Q(\i_tinyqv.cpu.instr_data[1][6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1102),
    .D(_00498_),
    .Q_N(_00130_),
    .Q(\i_tinyqv.cpu.instr_data[1][7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1103),
    .D(_00499_),
    .Q_N(_00134_),
    .Q(\i_tinyqv.cpu.instr_data[1][8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1104),
    .D(_00500_),
    .Q_N(_00138_),
    .Q(\i_tinyqv.cpu.instr_data[1][9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][0]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1105),
    .D(_00501_),
    .Q_N(_05317_),
    .Q(\i_tinyqv.cpu.instr_data[2][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1106),
    .D(_00502_),
    .Q_N(_00144_),
    .Q(\i_tinyqv.cpu.instr_data[2][10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1107),
    .D(_00503_),
    .Q_N(_00152_),
    .Q(\i_tinyqv.cpu.instr_data[2][11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1108),
    .D(_00504_),
    .Q_N(_00148_),
    .Q(\i_tinyqv.cpu.instr_data[2][12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1109),
    .D(_00505_),
    .Q_N(_00120_),
    .Q(\i_tinyqv.cpu.instr_data[2][13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1110),
    .D(_00506_),
    .Q_N(_00124_),
    .Q(\i_tinyqv.cpu.instr_data[2][14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1111),
    .D(_00507_),
    .Q_N(_00128_),
    .Q(\i_tinyqv.cpu.instr_data[2][15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1112),
    .D(_00508_),
    .Q_N(_00104_),
    .Q(\i_tinyqv.cpu.instr_data[2][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1113),
    .D(_00509_),
    .Q_N(_05316_),
    .Q(\i_tinyqv.cpu.instr_data[2][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1114),
    .D(_00510_),
    .Q_N(_05315_),
    .Q(\i_tinyqv.cpu.instr_data[2][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1115),
    .D(_00511_),
    .Q_N(_00108_),
    .Q(\i_tinyqv.cpu.instr_data[2][4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1116),
    .D(_00512_),
    .Q_N(_00112_),
    .Q(\i_tinyqv.cpu.instr_data[2][5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1117),
    .D(_00513_),
    .Q_N(_00116_),
    .Q(\i_tinyqv.cpu.instr_data[2][6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1118),
    .D(_00514_),
    .Q_N(_00132_),
    .Q(\i_tinyqv.cpu.instr_data[2][7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1119),
    .D(_00515_),
    .Q_N(_00136_),
    .Q(\i_tinyqv.cpu.instr_data[2][8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1120),
    .D(_00516_),
    .Q_N(_00140_),
    .Q(\i_tinyqv.cpu.instr_data[2][9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1121),
    .D(_00517_),
    .Q_N(_05314_),
    .Q(\i_tinyqv.cpu.instr_data[3][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1122),
    .D(_00518_),
    .Q_N(_00145_),
    .Q(\i_tinyqv.cpu.instr_data[3][10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1123),
    .D(_00519_),
    .Q_N(_00153_),
    .Q(\i_tinyqv.cpu.instr_data[3][11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1124),
    .D(_00520_),
    .Q_N(_00149_),
    .Q(\i_tinyqv.cpu.instr_data[3][12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1125),
    .D(_00521_),
    .Q_N(_00121_),
    .Q(\i_tinyqv.cpu.instr_data[3][13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1126),
    .D(_00522_),
    .Q_N(_00125_),
    .Q(\i_tinyqv.cpu.instr_data[3][14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1127),
    .D(_00523_),
    .Q_N(_00129_),
    .Q(\i_tinyqv.cpu.instr_data[3][15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1128),
    .D(_00524_),
    .Q_N(_00105_),
    .Q(\i_tinyqv.cpu.instr_data[3][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1129),
    .D(_00525_),
    .Q_N(_05313_),
    .Q(\i_tinyqv.cpu.instr_data[3][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1130),
    .D(_00526_),
    .Q_N(_05312_),
    .Q(\i_tinyqv.cpu.instr_data[3][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1131),
    .D(_00527_),
    .Q_N(_00109_),
    .Q(\i_tinyqv.cpu.instr_data[3][4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1132),
    .D(_00528_),
    .Q_N(_00113_),
    .Q(\i_tinyqv.cpu.instr_data[3][5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1133),
    .D(_00529_),
    .Q_N(_00117_),
    .Q(\i_tinyqv.cpu.instr_data[3][6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1134),
    .D(_00530_),
    .Q_N(_00133_),
    .Q(\i_tinyqv.cpu.instr_data[3][7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1135),
    .D(_00531_),
    .Q_N(_00137_),
    .Q(\i_tinyqv.cpu.instr_data[3][8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1136),
    .D(_00532_),
    .Q_N(_00141_),
    .Q(\i_tinyqv.cpu.instr_data[3][9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1137),
    .D(_00533_),
    .Q_N(_05311_),
    .Q(\i_tinyqv.cpu.instr_data_start[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1138),
    .D(_00534_),
    .Q_N(_05310_),
    .Q(\i_tinyqv.cpu.instr_data_start[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1139),
    .D(_00535_),
    .Q_N(_05309_),
    .Q(\i_tinyqv.cpu.instr_data_start[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1140),
    .D(_00536_),
    .Q_N(_05308_),
    .Q(\i_tinyqv.cpu.instr_data_start[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1141),
    .D(_00537_),
    .Q_N(_05307_),
    .Q(\i_tinyqv.cpu.instr_data_start[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1142),
    .D(_00538_),
    .Q_N(_05306_),
    .Q(\i_tinyqv.cpu.instr_data_start[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1143),
    .D(_00539_),
    .Q_N(_05305_),
    .Q(\i_tinyqv.cpu.instr_data_start[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1144),
    .D(_00540_),
    .Q_N(_05304_),
    .Q(\i_tinyqv.cpu.instr_data_start[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1145),
    .D(_00541_),
    .Q_N(_05303_),
    .Q(\i_tinyqv.cpu.instr_data_start[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1146),
    .D(_00542_),
    .Q_N(_05302_),
    .Q(\i_tinyqv.cpu.instr_data_start[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1147),
    .D(_00543_),
    .Q_N(_05301_),
    .Q(\i_tinyqv.cpu.instr_data_start[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1148),
    .D(_00544_),
    .Q_N(_00161_),
    .Q(\i_tinyqv.cpu.instr_data_start[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1149),
    .D(_00545_),
    .Q_N(_00160_),
    .Q(\i_tinyqv.cpu.instr_data_start[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1150),
    .D(_00546_),
    .Q_N(_05300_),
    .Q(\i_tinyqv.cpu.instr_data_start[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1151),
    .D(_00547_),
    .Q_N(_05299_),
    .Q(\i_tinyqv.cpu.instr_data_start[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1152),
    .D(_00548_),
    .Q_N(_05298_),
    .Q(\i_tinyqv.cpu.instr_data_start[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1153),
    .D(_00549_),
    .Q_N(_05297_),
    .Q(\i_tinyqv.cpu.instr_data_start[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1154),
    .D(_00550_),
    .Q_N(_05296_),
    .Q(\i_tinyqv.cpu.instr_data_start[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1155),
    .D(_00551_),
    .Q_N(_05295_),
    .Q(\i_tinyqv.cpu.instr_data_start[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1156),
    .D(_00552_),
    .Q_N(_05294_),
    .Q(\i_tinyqv.cpu.instr_data_start[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1157),
    .D(_00553_),
    .Q_N(_05293_),
    .Q(\i_tinyqv.cpu.instr_data_start[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_fetch_running$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1158),
    .D(_00554_),
    .Q_N(_00096_),
    .Q(\i_tinyqv.cpu.instr_fetch_running ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_len[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1159),
    .D(_00555_),
    .Q_N(_05292_),
    .Q(\i_tinyqv.cpu.instr_len[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_len[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1160),
    .D(_00556_),
    .Q_N(_05291_),
    .Q(\i_tinyqv.cpu.instr_len[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_valid$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1161),
    .D(_00557_),
    .Q_N(_00099_),
    .Q(debug_instr_valid));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_write_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1162),
    .D(_00558_),
    .Q_N(_00095_),
    .Q(\i_tinyqv.cpu.instr_write_offset[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_write_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1163),
    .D(_00559_),
    .Q_N(_00158_),
    .Q(\i_tinyqv.cpu.instr_write_offset[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_write_offset[2]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1164),
    .D(_00560_),
    .Q_N(_05290_),
    .Q(\i_tinyqv.cpu.instr_write_offset[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.interrupt_core$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1165),
    .D(_00561_),
    .Q_N(_00093_),
    .Q(\i_tinyqv.cpu.i_core.is_interrupt ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_alu_imm$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1166),
    .D(_00562_),
    .Q_N(_05289_),
    .Q(\i_tinyqv.cpu.is_alu_imm ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_alu_reg$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1167),
    .D(_00563_),
    .Q_N(_05288_),
    .Q(\i_tinyqv.cpu.is_alu_reg ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_auipc$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1168),
    .D(_00564_),
    .Q_N(_05287_),
    .Q(\i_tinyqv.cpu.is_auipc ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_branch$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1169),
    .D(_00565_),
    .Q_N(_05286_),
    .Q(\i_tinyqv.cpu.is_branch ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_jal$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1170),
    .D(_00566_),
    .Q_N(_05285_),
    .Q(\i_tinyqv.cpu.is_jal ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_jalr$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1171),
    .D(_00567_),
    .Q_N(_05284_),
    .Q(\i_tinyqv.cpu.is_jalr ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_load$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1172),
    .D(_00568_),
    .Q_N(_05283_),
    .Q(\i_tinyqv.cpu.is_load ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_lui$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1173),
    .D(_00569_),
    .Q_N(_05282_),
    .Q(\i_tinyqv.cpu.is_lui ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_store$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1174),
    .D(_00570_),
    .Q_N(_05281_),
    .Q(\i_tinyqv.cpu.is_store ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_system$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1175),
    .D(_00571_),
    .Q_N(_05280_),
    .Q(\i_tinyqv.cpu.is_system ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.load_started$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1176),
    .D(_00572_),
    .Q_N(_05279_),
    .Q(\i_tinyqv.cpu.load_started ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.mem_op[0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1177),
    .D(_00573_),
    .Q_N(_05278_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.mem_op[1]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1178),
    .D(_00574_),
    .Q_N(_05277_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.mem_op[2]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1179),
    .D(_00575_),
    .Q_N(_05276_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.mem_op_increment_reg$_SDFFCE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1180),
    .D(_00576_),
    .Q_N(_05275_),
    .Q(\i_tinyqv.cpu.mem_op_increment_reg ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.no_write_in_progress$_SDFFE_PN1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1181),
    .D(_00577_),
    .Q_N(_00083_),
    .Q(\i_tinyqv.cpu.no_write_in_progress ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.pc_offset[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1182),
    .D(_00578_),
    .Q_N(_00100_),
    .Q(\i_tinyqv.cpu.pc[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.pc_offset[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1183),
    .D(_00579_),
    .Q_N(_00101_),
    .Q(\i_tinyqv.cpu.pc[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1184),
    .D(_00580_),
    .Q_N(_00213_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1185),
    .D(_00581_),
    .Q_N(_05274_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1186),
    .D(_00582_),
    .Q_N(_05273_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1187),
    .D(_00583_),
    .Q_N(_05272_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1188),
    .D(_00584_),
    .Q_N(_05271_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1189),
    .D(_00585_),
    .Q_N(_05270_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1190),
    .D(_00586_),
    .Q_N(_05269_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1191),
    .D(_00587_),
    .Q_N(_05268_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1192),
    .D(_00588_),
    .Q_N(_05267_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs2[1]$_DFFE_PP_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net1193),
    .D(_00589_),
    .Q_N(_05266_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1194),
    .D(_00590_),
    .Q_N(_05265_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1195),
    .D(_00591_),
    .Q_N(_05264_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.was_early_branch$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1196),
    .D(_00592_),
    .Q_N(_00098_),
    .Q(\i_tinyqv.cpu.was_early_branch ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.data_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1197),
    .D(_00593_),
    .Q_N(_05263_),
    .Q(\i_tinyqv.mem.data_stall ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.instr_active$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1198),
    .D(_00594_),
    .Q_N(_00097_),
    .Q(\i_tinyqv.mem.instr_active ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.instr_fetch_started$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1199),
    .D(_00595_),
    .Q_N(_05262_),
    .Q(\i_tinyqv.cpu.instr_fetch_started ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.instr_fetch_stopped$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1200),
    .D(_00596_),
    .Q_N(_05261_),
    .Q(\i_tinyqv.cpu.instr_fetch_stopped ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1201),
    .D(_00597_),
    .Q_N(_05260_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[10]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1202),
    .D(_00598_),
    .Q_N(_05259_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[11]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1203),
    .D(_00599_),
    .Q_N(_05258_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[12]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1204),
    .D(_00600_),
    .Q_N(_05257_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[13]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1205),
    .D(_00601_),
    .Q_N(_05256_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[14]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1206),
    .D(_00602_),
    .Q_N(_05255_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[15]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1207),
    .D(_00603_),
    .Q_N(_05254_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[16]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1208),
    .D(_00604_),
    .Q_N(_05253_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[17]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1209),
    .D(_00605_),
    .Q_N(_05252_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[18]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1210),
    .D(_00606_),
    .Q_N(_05251_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[19]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1211),
    .D(_00607_),
    .Q_N(_05250_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1212),
    .D(_00608_),
    .Q_N(_05249_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[20]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1213),
    .D(_00609_),
    .Q_N(_05248_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[21]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1214),
    .D(_00610_),
    .Q_N(_05247_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[22]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1215),
    .D(_00611_),
    .Q_N(_05246_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[23]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1216),
    .D(_00612_),
    .Q_N(_05245_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1217),
    .D(_00613_),
    .Q_N(_05244_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1218),
    .D(_00614_),
    .Q_N(_05243_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[4]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1219),
    .D(_00615_),
    .Q_N(_05242_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[5]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1220),
    .D(_00616_),
    .Q_N(_05241_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[6]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1221),
    .D(_00617_),
    .Q_N(_05240_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[7]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1222),
    .D(_00618_),
    .Q_N(_05239_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[8]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1223),
    .D(_00619_),
    .Q_N(_05238_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[9]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1224),
    .D(_00620_),
    .Q_N(_05237_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[0]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1225),
    .D(_00621_),
    .Q_N(_00207_),
    .Q(\i_tinyqv.cpu.instr_data_in[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1226),
    .D(_00622_),
    .Q_N(_00208_),
    .Q(\i_tinyqv.cpu.instr_data_in[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1227),
    .D(_00623_),
    .Q_N(_00209_),
    .Q(\i_tinyqv.cpu.instr_data_in[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1228),
    .D(_00624_),
    .Q_N(_00210_),
    .Q(\i_tinyqv.cpu.instr_data_in[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[4]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1229),
    .D(_00625_),
    .Q_N(_00204_),
    .Q(\i_tinyqv.cpu.instr_data_in[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[5]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1230),
    .D(_00626_),
    .Q_N(_00205_),
    .Q(\i_tinyqv.cpu.instr_data_in[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1231),
    .D(_00627_),
    .Q_N(_00211_),
    .Q(\i_tinyqv.cpu.instr_data_in[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1232),
    .D(_00628_),
    .Q_N(_00206_),
    .Q(\i_tinyqv.cpu.instr_data_in[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data_ready$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1233),
    .D(_00629_),
    .Q_N(_05236_),
    .Q(\i_tinyqv.mem.q_ctrl.data_ready ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data_req$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1234),
    .D(_00630_),
    .Q_N(_05235_),
    .Q(\i_tinyqv.mem.q_ctrl.data_req ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1235),
    .D(_00631_),
    .Q_N(_05234_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1236),
    .D(_00632_),
    .Q_N(_05233_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1237),
    .D(_00633_),
    .Q_N(_05232_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.fsm_state[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1238),
    .D(_00634_),
    .Q_N(_00163_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.fsm_state[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1239),
    .D(_00635_),
    .Q_N(_05231_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.fsm_state[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1240),
    .D(_00636_),
    .Q_N(_00155_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.is_writing$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1241),
    .D(_00637_),
    .Q_N(_00162_),
    .Q(\i_tinyqv.mem.q_ctrl.is_writing ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.last_ram_a_sel$_SDFF_PN1_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1242),
    .D(_00638_),
    .Q_N(_05230_),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.last_ram_b_sel$_SDFF_PN1_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1243),
    .D(_00639_),
    .Q_N(_05229_),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.nibbles_remaining[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1244),
    .D(_00640_),
    .Q_N(_05228_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.nibbles_remaining[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1245),
    .D(_00641_),
    .Q_N(_05227_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.nibbles_remaining[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1246),
    .D(_00642_),
    .Q_N(_05226_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.read_cycles_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1247),
    .D(_00643_),
    .Q_N(_00165_),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.read_cycles_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1248),
    .D(_00644_),
    .Q_N(_05225_),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.read_cycles_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1249),
    .D(_00645_),
    .Q_N(_05224_),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_clk_out$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1250),
    .D(_00646_),
    .Q_N(_05223_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_out ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_data_oe[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1251),
    .D(_00647_),
    .Q_N(_05222_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_flash_select$_SDFFE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1252),
    .D(_00648_),
    .Q_N(_05221_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_flash_select ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1253),
    .D(_00649_),
    .Q_N(_05220_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1254),
    .D(_00650_),
    .Q_N(_05219_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1255),
    .D(_00651_),
    .Q_N(_05218_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[3]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1256),
    .D(_00652_),
    .Q_N(_05217_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[4]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1257),
    .D(_00653_),
    .Q_N(_05216_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[5]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1258),
    .D(_00654_),
    .Q_N(_05215_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1259),
    .D(_00655_),
    .Q_N(_05214_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[7]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1260),
    .D(_00656_),
    .Q_N(_05213_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_ram_a_select$_SDFFE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1261),
    .D(_00657_),
    .Q_N(_05212_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_ram_b_select$_SDFFE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1262),
    .D(_00658_),
    .Q_N(_05211_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.stop_txn_reg$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1263),
    .D(_00659_),
    .Q_N(_05210_),
    .Q(\i_tinyqv.mem.q_ctrl.stop_txn_reg ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[0]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1264),
    .D(_00660_),
    .Q_N(_05209_),
    .Q(\i_tinyqv.cpu.instr_data_in[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1265),
    .D(_00661_),
    .Q_N(_05208_),
    .Q(\i_tinyqv.mem.qspi_data_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[11]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1266),
    .D(_00662_),
    .Q_N(_05207_),
    .Q(\i_tinyqv.mem.qspi_data_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[12]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1267),
    .D(_00663_),
    .Q_N(_05206_),
    .Q(\i_tinyqv.mem.qspi_data_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[13]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1268),
    .D(_00664_),
    .Q_N(_05205_),
    .Q(\i_tinyqv.mem.qspi_data_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[14]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1269),
    .D(_00665_),
    .Q_N(_05204_),
    .Q(\i_tinyqv.mem.qspi_data_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[15]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1270),
    .D(_00666_),
    .Q_N(_05203_),
    .Q(\i_tinyqv.mem.qspi_data_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[16]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1271),
    .D(_00667_),
    .Q_N(_05202_),
    .Q(\i_tinyqv.mem.data_from_read[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[17]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1272),
    .D(_00668_),
    .Q_N(_05201_),
    .Q(\i_tinyqv.mem.data_from_read[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[18]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1273),
    .D(_00669_),
    .Q_N(_05200_),
    .Q(\i_tinyqv.mem.data_from_read[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[19]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1274),
    .D(_00670_),
    .Q_N(_05199_),
    .Q(\i_tinyqv.mem.data_from_read[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1275),
    .D(_00671_),
    .Q_N(_05198_),
    .Q(\i_tinyqv.cpu.instr_data_in[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[20]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1276),
    .D(_00672_),
    .Q_N(_05197_),
    .Q(\i_tinyqv.mem.data_from_read[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[21]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1277),
    .D(_00673_),
    .Q_N(_05196_),
    .Q(\i_tinyqv.mem.data_from_read[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[22]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1278),
    .D(_00674_),
    .Q_N(_05195_),
    .Q(\i_tinyqv.mem.data_from_read[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[23]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1279),
    .D(_00675_),
    .Q_N(_05194_),
    .Q(\i_tinyqv.mem.data_from_read[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[24]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1280),
    .D(_00676_),
    .Q_N(_05193_),
    .Q(\i_tinyqv.mem.qspi_data_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[25]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1281),
    .D(_00677_),
    .Q_N(_05192_),
    .Q(\i_tinyqv.mem.qspi_data_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[26]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1282),
    .D(_00678_),
    .Q_N(_05191_),
    .Q(\i_tinyqv.mem.qspi_data_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[27]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1283),
    .D(_00679_),
    .Q_N(_05190_),
    .Q(\i_tinyqv.mem.qspi_data_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[28]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1284),
    .D(_00680_),
    .Q_N(_05189_),
    .Q(\i_tinyqv.mem.qspi_data_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[29]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1285),
    .D(_00681_),
    .Q_N(_05188_),
    .Q(\i_tinyqv.mem.qspi_data_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1286),
    .D(_00682_),
    .Q_N(_05187_),
    .Q(\i_tinyqv.cpu.instr_data_in[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[30]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1287),
    .D(_00683_),
    .Q_N(_05186_),
    .Q(\i_tinyqv.mem.qspi_data_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[31]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1288),
    .D(_00684_),
    .Q_N(_05185_),
    .Q(\i_tinyqv.mem.qspi_data_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1289),
    .D(_00685_),
    .Q_N(_05184_),
    .Q(\i_tinyqv.cpu.instr_data_in[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1290),
    .D(_00686_),
    .Q_N(_05183_),
    .Q(\i_tinyqv.cpu.instr_data_in[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[5]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1291),
    .D(_00687_),
    .Q_N(_05182_),
    .Q(\i_tinyqv.cpu.instr_data_in[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[6]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1292),
    .D(_00688_),
    .Q_N(_05181_),
    .Q(\i_tinyqv.cpu.instr_data_in[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[7]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1293),
    .D(_00689_),
    .Q_N(_05180_),
    .Q(\i_tinyqv.cpu.instr_data_in[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[8]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1294),
    .D(_00690_),
    .Q_N(_05179_),
    .Q(\i_tinyqv.mem.qspi_data_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1295),
    .D(_00691_),
    .Q_N(_05178_),
    .Q(\i_tinyqv.mem.qspi_data_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_byte_idx[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1296),
    .D(_00692_),
    .Q_N(_00157_),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_byte_idx[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1297),
    .D(_00693_),
    .Q_N(_06026_),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_write_done$_DFF_P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1298),
    .D(_00082_),
    .Q_N(_00154_),
    .Q(\i_tinyqv.mem.qspi_write_done ));
 sg13g2_dfrbp_1 \i_tinyqv.rst_reg_n$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1299),
    .D(\i_debug_uart_tx.resetn ),
    .Q_N(_00164_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.rstn ));
 sg13g2_dfrbp_1 \i_uart_rx.bit_sample$_SDFFE_PN0N_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1300),
    .D(_00694_),
    .Q_N(_05177_),
    .Q(\i_uart_rx.bit_sample ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1301),
    .D(_00695_),
    .Q_N(_00220_),
    .Q(\i_uart_rx.cycle_counter[0] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[10]$_SDFF_PP0_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1302),
    .D(_00696_),
    .Q_N(_05176_),
    .Q(\i_uart_rx.cycle_counter[10] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1303),
    .D(_00697_),
    .Q_N(_05175_),
    .Q(\i_uart_rx.cycle_counter[1] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1304),
    .D(_00698_),
    .Q_N(_05174_),
    .Q(\i_uart_rx.cycle_counter[2] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1305),
    .D(_00699_),
    .Q_N(_05173_),
    .Q(\i_uart_rx.cycle_counter[3] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1306),
    .D(_00700_),
    .Q_N(_05172_),
    .Q(\i_uart_rx.cycle_counter[4] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[5]$_SDFF_PP0_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1307),
    .D(_00701_),
    .Q_N(_05171_),
    .Q(\i_uart_rx.cycle_counter[5] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1308),
    .D(_00702_),
    .Q_N(_05170_),
    .Q(\i_uart_rx.cycle_counter[6] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1309),
    .D(_00703_),
    .Q_N(_05169_),
    .Q(\i_uart_rx.cycle_counter[7] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[8]$_SDFF_PP0_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1310),
    .D(_00704_),
    .Q_N(_05168_),
    .Q(\i_uart_rx.cycle_counter[8] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[9]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1311),
    .D(_00705_),
    .Q_N(_05167_),
    .Q(\i_uart_rx.cycle_counter[9] ));
 sg13g2_dfrbp_1 \i_uart_rx.fsm_state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1312),
    .D(_00706_),
    .Q_N(_00202_),
    .Q(\i_uart_rx.fsm_state[0] ));
 sg13g2_dfrbp_1 \i_uart_rx.fsm_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1313),
    .D(_00707_),
    .Q_N(_05166_),
    .Q(\i_uart_rx.fsm_state[1] ));
 sg13g2_dfrbp_1 \i_uart_rx.fsm_state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1314),
    .D(_00708_),
    .Q_N(_05165_),
    .Q(\i_uart_rx.fsm_state[2] ));
 sg13g2_dfrbp_1 \i_uart_rx.fsm_state[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1315),
    .D(_00709_),
    .Q_N(_05164_),
    .Q(\i_uart_rx.fsm_state[3] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1316),
    .D(_00710_),
    .Q_N(_05163_),
    .Q(\i_uart_rx.recieved_data[0] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[1]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1317),
    .D(_00711_),
    .Q_N(_05162_),
    .Q(\i_uart_rx.recieved_data[1] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[2]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1318),
    .D(_00712_),
    .Q_N(_05161_),
    .Q(\i_uart_rx.recieved_data[2] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[3]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1319),
    .D(_00713_),
    .Q_N(_05160_),
    .Q(\i_uart_rx.recieved_data[3] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[4]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1320),
    .D(_00714_),
    .Q_N(_05159_),
    .Q(\i_uart_rx.recieved_data[4] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[5]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1321),
    .D(_00715_),
    .Q_N(_05158_),
    .Q(\i_uart_rx.recieved_data[5] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[6]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1322),
    .D(_00716_),
    .Q_N(_05157_),
    .Q(\i_uart_rx.recieved_data[6] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[7]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1323),
    .D(_00717_),
    .Q_N(_05156_),
    .Q(\i_uart_rx.recieved_data[7] ));
 sg13g2_dfrbp_1 \i_uart_rx.rxd_reg[0]$_SDFF_PN1_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1324),
    .D(_00718_),
    .Q_N(_00203_),
    .Q(\i_uart_rx.rxd_reg[0] ));
 sg13g2_dfrbp_1 \i_uart_rx.rxd_reg[1]$_SDFF_PN1_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1325),
    .D(_00719_),
    .Q_N(_05155_),
    .Q(\i_uart_rx.rxd_reg[1] ));
 sg13g2_dfrbp_1 \i_uart_rx.uart_rts$_SDFF_PN1_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1326),
    .D(_00720_),
    .Q_N(_05154_),
    .Q(\i_uart_rx.uart_rts ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1327),
    .D(_00721_),
    .Q_N(_00219_),
    .Q(\i_uart_tx.cycle_counter[0] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1328),
    .D(_00722_),
    .Q_N(_05153_),
    .Q(\i_uart_tx.cycle_counter[10] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1329),
    .D(_00723_),
    .Q_N(_05152_),
    .Q(\i_uart_tx.cycle_counter[1] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1330),
    .D(_00724_),
    .Q_N(_05151_),
    .Q(\i_uart_tx.cycle_counter[2] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1331),
    .D(_00725_),
    .Q_N(_05150_),
    .Q(\i_uart_tx.cycle_counter[3] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1332),
    .D(_00726_),
    .Q_N(_05149_),
    .Q(\i_uart_tx.cycle_counter[4] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1333),
    .D(_00727_),
    .Q_N(_05148_),
    .Q(\i_uart_tx.cycle_counter[5] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1334),
    .D(_00728_),
    .Q_N(_05147_),
    .Q(\i_uart_tx.cycle_counter[6] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1335),
    .D(_00729_),
    .Q_N(_05146_),
    .Q(\i_uart_tx.cycle_counter[7] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1336),
    .D(_00730_),
    .Q_N(_05145_),
    .Q(\i_uart_tx.cycle_counter[8] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1337),
    .D(_00731_),
    .Q_N(_05144_),
    .Q(\i_uart_tx.cycle_counter[9] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1338),
    .D(_00732_),
    .Q_N(_05143_),
    .Q(\i_uart_tx.data_to_send[0] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1339),
    .D(_00733_),
    .Q_N(_05142_),
    .Q(\i_uart_tx.data_to_send[1] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1340),
    .D(_00734_),
    .Q_N(_05141_),
    .Q(\i_uart_tx.data_to_send[2] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1341),
    .D(_00735_),
    .Q_N(_05140_),
    .Q(\i_uart_tx.data_to_send[3] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1342),
    .D(_00736_),
    .Q_N(_05139_),
    .Q(\i_uart_tx.data_to_send[4] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1343),
    .D(_00737_),
    .Q_N(_05138_),
    .Q(\i_uart_tx.data_to_send[5] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1344),
    .D(_00738_),
    .Q_N(_05137_),
    .Q(\i_uart_tx.data_to_send[6] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1345),
    .D(_00739_),
    .Q_N(_05136_),
    .Q(\i_uart_tx.data_to_send[7] ));
 sg13g2_dfrbp_1 \i_uart_tx.fsm_state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1346),
    .D(_00740_),
    .Q_N(_05135_),
    .Q(\i_uart_tx.fsm_state[0] ));
 sg13g2_dfrbp_1 \i_uart_tx.fsm_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1347),
    .D(_00741_),
    .Q_N(_05134_),
    .Q(\i_uart_tx.fsm_state[1] ));
 sg13g2_dfrbp_1 \i_uart_tx.fsm_state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1348),
    .D(_00742_),
    .Q_N(_05133_),
    .Q(\i_uart_tx.fsm_state[2] ));
 sg13g2_dfrbp_1 \i_uart_tx.fsm_state[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1349),
    .D(_00743_),
    .Q_N(_05132_),
    .Q(\i_uart_tx.fsm_state[3] ));
 sg13g2_dfrbp_1 \i_uart_tx.txd_reg$_SDFF_PN1_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1350),
    .D(_00744_),
    .Q_N(_05131_),
    .Q(\i_uart_tx.txd_reg ));
 sg13g2_dfrbp_1 \rst_reg_n$_DFF_N_  (.CLK(net1354),
    .RESET_B(net1351),
    .D(net1),
    .Q_N(_00156_),
    .Q(\i_debug_uart_tx.resetn ));
 sg13g2_dfrbp_1 \ui_in_reg[0]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1352),
    .D(net2),
    .Q_N(_06027_),
    .Q(\i_tinyqv.cpu.i_core.interrupt_req[0] ));
 sg13g2_dfrbp_1 \ui_in_reg[1]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1353),
    .D(net3),
    .Q_N(_05130_),
    .Q(\i_tinyqv.cpu.i_core.interrupt_req[1] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[0]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[1]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[2]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[4]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[5]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[6]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[7]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[0]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[1]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[2]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[3]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[4]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_out[5]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[6]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[7]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[0]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[1]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[2]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[3]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[4]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uo_out[5]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[6]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout36 (.A(_03266_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_03237_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02964_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02916_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_02915_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_03183_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_02977_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_02914_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(\debug_rd[3] ),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_03533_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_04952_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_04422_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_03446_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_03444_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_03425_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_03422_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_03481_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_03480_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_03460_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_03458_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_02911_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(\debug_rd[2] ),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_04803_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_03818_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_03817_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_03641_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_03626_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(\debug_rd[1] ),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(\debug_rd[0] ),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_04805_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_04789_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_03832_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_03724_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_03640_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_03630_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_03625_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_04809_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_04806_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_04797_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_04796_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_04795_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_04794_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_04808_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_03534_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_03515_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_03471_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_01658_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_01281_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_03301_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_01644_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_03299_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_03241_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_03343_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_03214_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_03242_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_03213_),
    .X(net91));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(_03031_));
 sg13g2_buf_2 fanout93 (.A(_03010_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_02982_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_02959_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_02956_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_02945_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_01758_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_01324_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_03329_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_03212_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_03209_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_03205_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_03191_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_03129_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_02968_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_02954_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_02932_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_01958_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_01596_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_05064_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_04015_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_03208_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_03204_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_02988_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_02967_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_02931_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_02083_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_02081_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_02046_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_01756_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_01483_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_01339_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_01310_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_01052_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_04605_),
    .X(net126));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_02990_));
 sg13g2_buf_2 fanout128 (.A(_02966_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_02935_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_02927_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_02186_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_01814_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_01709_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_01655_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_01625_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_01450_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_01221_),
    .X(net137));
 sg13g2_buf_1 fanout138 (.A(_04604_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_04575_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_04541_),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(_04233_));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(_04231_));
 sg13g2_buf_2 fanout143 (.A(_04229_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_04228_),
    .X(net144));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(_04201_));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(_04200_));
 sg13g2_buf_2 fanout147 (.A(_03021_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_03014_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_03013_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_02182_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_01699_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_01481_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_01136_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_00856_),
    .X(net154));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(_03781_));
 sg13g2_buf_2 fanout156 (.A(_03638_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_02381_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_01407_),
    .X(net158));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(_01397_));
 sg13g2_buf_2 fanout160 (.A(_01166_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_04811_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_04791_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_02603_),
    .X(net163));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(_02425_));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(_02420_));
 sg13g2_buf_2 fanout166 (.A(_02220_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_01622_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_01367_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_01304_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_01297_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_01167_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_01165_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_01060_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_04810_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_04790_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_04633_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_04632_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_04601_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_04572_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_04299_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_04168_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_04157_),
    .X(net182));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(_03000_));
 sg13g2_buf_2 fanout184 (.A(_02386_),
    .X(net184));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(_02233_));
 sg13g2_buf_2 fanout186 (.A(_02232_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_02223_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_02178_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_01532_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_01512_),
    .X(net190));
 sg13g2_buf_4 fanout191 (.X(net191),
    .A(_01303_));
 sg13g2_buf_2 fanout192 (.A(_01296_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_00827_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_04822_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_04778_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_04773_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_04747_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_04716_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_04698_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_03635_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_02264_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_02247_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_02231_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_02225_),
    .X(net204));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(_02222_));
 sg13g2_buf_2 fanout206 (.A(_02202_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_02193_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_01567_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_01389_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_01229_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_00757_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_04697_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_04654_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_04424_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_02862_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_01614_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_01598_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_01288_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_01220_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_01141_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_00887_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_00885_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_00882_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_00874_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_00790_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_00770_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_00766_),
    .X(net227));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(_00763_));
 sg13g2_buf_2 fanout229 (.A(_04145_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_04140_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_04114_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_04085_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_04019_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_04016_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_03999_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_03715_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_03711_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_03684_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_03674_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_03643_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_03470_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_03018_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_02882_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_02867_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_02431_),
    .X(net245));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(_02430_));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(_02427_));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(_02423_));
 sg13g2_buf_2 fanout249 (.A(_02414_),
    .X(net249));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(_02413_));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(_02409_));
 sg13g2_buf_2 fanout252 (.A(_02308_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_02306_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_02292_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_02291_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_02290_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_02275_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_02266_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_01661_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_01643_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_01597_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_01183_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_01174_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_01163_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_00884_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_00879_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_00877_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_00873_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_00829_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_00787_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_00786_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_00783_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_00778_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_00776_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_00765_),
    .X(net275));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(_00762_));
 sg13g2_buf_2 fanout277 (.A(_00755_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_04193_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_04002_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_03642_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_03632_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_03066_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_02866_),
    .X(net283));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_02437_));
 sg13g2_buf_2 fanout285 (.A(_02318_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_02297_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_02276_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_02274_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_02265_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_02195_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_02162_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_02085_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_02024_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_01983_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_01579_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_01576_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_01427_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_01406_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_01376_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_01375_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_01241_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_01191_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_01146_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_01142_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_01137_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_01042_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_00990_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_00989_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_00987_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_00969_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_00919_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_00857_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_00823_),
    .X(net313));
 sg13g2_buf_1 fanout314 (.A(_00775_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_00746_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_01260_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_01257_),
    .X(net317));
 sg13g2_tiehi _11040__318 (.L_HI(net318));
 sg13g2_tiehi _11041__319 (.L_HI(net319));
 sg13g2_tiehi _11042__320 (.L_HI(net320));
 sg13g2_tiehi _11043__321 (.L_HI(net321));
 sg13g2_tiehi _11044__322 (.L_HI(net322));
 sg13g2_tiehi _11045__323 (.L_HI(net323));
 sg13g2_tiehi \debug_rd_r[0]$_DFF_P__324  (.L_HI(net324));
 sg13g2_tiehi \debug_rd_r[1]$_DFF_P__325  (.L_HI(net325));
 sg13g2_tiehi \debug_rd_r[2]$_DFF_P__326  (.L_HI(net326));
 sg13g2_tiehi \debug_rd_r[3]$_DFF_P__327  (.L_HI(net327));
 sg13g2_tiehi \debug_register_data$_DFFE_PP__328  (.L_HI(net328));
 sg13g2_tiehi \gpio_out[0]$_DFF_P__329  (.L_HI(net329));
 sg13g2_tiehi \gpio_out[1]$_DFF_P__330  (.L_HI(net330));
 sg13g2_tiehi \gpio_out[2]$_DFF_P__331  (.L_HI(net331));
 sg13g2_tiehi \gpio_out[3]$_DFF_P__332  (.L_HI(net332));
 sg13g2_tiehi \gpio_out[4]$_DFF_P__333  (.L_HI(net333));
 sg13g2_tiehi \gpio_out[5]$_DFF_P__334  (.L_HI(net334));
 sg13g2_tiehi \gpio_out[6]$_DFF_P__335  (.L_HI(net335));
 sg13g2_tiehi \gpio_out[7]$_DFF_P__336  (.L_HI(net336));
 sg13g2_tiehi \gpio_out_sel[0]$_DFF_P__337  (.L_HI(net337));
 sg13g2_tiehi \gpio_out_sel[1]$_DFF_P__338  (.L_HI(net338));
 sg13g2_tiehi \gpio_out_sel[2]$_DFF_P__339  (.L_HI(net339));
 sg13g2_tiehi \gpio_out_sel[3]$_DFF_P__340  (.L_HI(net340));
 sg13g2_tiehi \gpio_out_sel[4]$_DFF_P__341  (.L_HI(net341));
 sg13g2_tiehi \gpio_out_sel[5]$_DFF_P__342  (.L_HI(net342));
 sg13g2_tiehi \gpio_out_sel[6]$_DFF_P__343  (.L_HI(net343));
 sg13g2_tiehi \gpio_out_sel[7]$_DFF_P__344  (.L_HI(net344));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[0]$_SDFFE_PP0N__345  (.L_HI(net345));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[1]$_SDFFE_PP0N__346  (.L_HI(net346));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[2]$_SDFFE_PP0N__347  (.L_HI(net347));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[3]$_SDFFE_PP0N__348  (.L_HI(net348));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[4]$_SDFFE_PP0N__349  (.L_HI(net349));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[0]$_SDFFE_PN0P__350  (.L_HI(net350));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[1]$_SDFFE_PN0P__351  (.L_HI(net351));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[2]$_SDFFE_PN0P__352  (.L_HI(net352));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[3]$_SDFFE_PN0P__353  (.L_HI(net353));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[4]$_SDFFE_PN0P__354  (.L_HI(net354));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[5]$_SDFFE_PN0P__355  (.L_HI(net355));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[6]$_SDFFE_PN0P__356  (.L_HI(net356));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[7]$_SDFFE_PN0P__357  (.L_HI(net357));
 sg13g2_tiehi \i_debug_uart_tx.fsm_state[0]$_SDFFE_PN0P__358  (.L_HI(net358));
 sg13g2_tiehi \i_debug_uart_tx.fsm_state[1]$_SDFFE_PN0P__359  (.L_HI(net359));
 sg13g2_tiehi \i_debug_uart_tx.fsm_state[2]$_SDFFE_PN0P__360  (.L_HI(net360));
 sg13g2_tiehi \i_debug_uart_tx.fsm_state[3]$_SDFFE_PN0P__361  (.L_HI(net361));
 sg13g2_tiehi \i_debug_uart_tx.txd_reg$_SDFF_PN1__362  (.L_HI(net362));
 sg13g2_tiehi \i_spi.bits_remaining[0]$_SDFFE_PN0P__363  (.L_HI(net363));
 sg13g2_tiehi \i_spi.bits_remaining[1]$_SDFFE_PN0P__364  (.L_HI(net364));
 sg13g2_tiehi \i_spi.bits_remaining[2]$_SDFFE_PN0P__365  (.L_HI(net365));
 sg13g2_tiehi \i_spi.bits_remaining[3]$_SDFFE_PN0P__366  (.L_HI(net366));
 sg13g2_tiehi \i_spi.busy$_SDFF_PN0__367  (.L_HI(net367));
 sg13g2_tiehi \i_spi.clock_count[0]$_SDFFE_PN0P__368  (.L_HI(net368));
 sg13g2_tiehi \i_spi.clock_count[1]$_SDFFE_PN0P__369  (.L_HI(net369));
 sg13g2_tiehi \i_spi.clock_divider[0]$_SDFFE_PN1P__370  (.L_HI(net370));
 sg13g2_tiehi \i_spi.clock_divider[1]$_SDFFE_PN0P__371  (.L_HI(net371));
 sg13g2_tiehi \i_spi.data[0]$_DFFE_PP__372  (.L_HI(net372));
 sg13g2_tiehi \i_spi.data[1]$_DFFE_PP__373  (.L_HI(net373));
 sg13g2_tiehi \i_spi.data[2]$_DFFE_PP__374  (.L_HI(net374));
 sg13g2_tiehi \i_spi.data[3]$_DFFE_PP__375  (.L_HI(net375));
 sg13g2_tiehi \i_spi.data[4]$_DFFE_PP__376  (.L_HI(net376));
 sg13g2_tiehi \i_spi.data[5]$_DFFE_PP__377  (.L_HI(net377));
 sg13g2_tiehi \i_spi.data[6]$_DFFE_PP__378  (.L_HI(net378));
 sg13g2_tiehi \i_spi.data[7]$_DFFE_PP__379  (.L_HI(net379));
 sg13g2_tiehi \i_spi.end_txn_reg$_DFFE_PP__380  (.L_HI(net380));
 sg13g2_tiehi \i_spi.read_latency$_SDFFE_PN0P__381  (.L_HI(net381));
 sg13g2_tiehi \i_spi.spi_clk_out$_SDFFE_PN0P__382  (.L_HI(net382));
 sg13g2_tiehi \i_spi.spi_dc$_DFFE_PP__383  (.L_HI(net383));
 sg13g2_tiehi \i_spi.spi_select$_SDFFE_PN1P__384  (.L_HI(net384));
 sg13g2_tiehi \i_tinyqv.cpu.additional_mem_ops[0]$_SDFFE_PN0P__385  (.L_HI(net385));
 sg13g2_tiehi \i_tinyqv.cpu.additional_mem_ops[1]$_SDFFE_PN0P__386  (.L_HI(net386));
 sg13g2_tiehi \i_tinyqv.cpu.additional_mem_ops[2]$_SDFFE_PN0P__387  (.L_HI(net387));
 sg13g2_tiehi \i_tinyqv.cpu.alu_op[0]$_DFFE_PP__388  (.L_HI(net388));
 sg13g2_tiehi \i_tinyqv.cpu.alu_op[1]$_DFFE_PP__389  (.L_HI(net389));
 sg13g2_tiehi \i_tinyqv.cpu.alu_op[2]$_DFFE_PP__390  (.L_HI(net390));
 sg13g2_tiehi \i_tinyqv.cpu.alu_op[3]$_DFFE_PP__391  (.L_HI(net391));
 sg13g2_tiehi \i_tinyqv.cpu.counter_hi[0]$_SDFF_PN0__392  (.L_HI(net392));
 sg13g2_tiehi \i_tinyqv.cpu.counter_hi[1]$_SDFF_PN0__393  (.L_HI(net393));
 sg13g2_tiehi \i_tinyqv.cpu.counter_hi[2]$_SDFF_PN0__394  (.L_HI(net394));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[0]$_DFFE_PP__395  (.L_HI(net395));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[10]$_DFFE_PP__396  (.L_HI(net396));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[11]$_DFFE_PP__397  (.L_HI(net397));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[12]$_DFFE_PP__398  (.L_HI(net398));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[13]$_DFFE_PP__399  (.L_HI(net399));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[14]$_DFFE_PP__400  (.L_HI(net400));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[15]$_DFFE_PP__401  (.L_HI(net401));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[16]$_DFFE_PP__402  (.L_HI(net402));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[17]$_DFFE_PP__403  (.L_HI(net403));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[18]$_DFFE_PP__404  (.L_HI(net404));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[19]$_DFFE_PP__405  (.L_HI(net405));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[1]$_DFFE_PP__406  (.L_HI(net406));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[20]$_DFFE_PP__407  (.L_HI(net407));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[21]$_DFFE_PP__408  (.L_HI(net408));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[22]$_DFFE_PP__409  (.L_HI(net409));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[23]$_DFFE_PP__410  (.L_HI(net410));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[24]$_SDFFE_PN0P__411  (.L_HI(net411));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[25]$_SDFFE_PN0P__412  (.L_HI(net412));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[26]$_SDFFE_PN0P__413  (.L_HI(net413));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[27]$_SDFFE_PN0P__414  (.L_HI(net414));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[2]$_DFFE_PP__415  (.L_HI(net415));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[3]$_DFFE_PP__416  (.L_HI(net416));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[4]$_DFFE_PP__417  (.L_HI(net417));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[5]$_DFFE_PP__418  (.L_HI(net418));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[6]$_DFFE_PP__419  (.L_HI(net419));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[7]$_DFFE_PP__420  (.L_HI(net420));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[8]$_DFFE_PP__421  (.L_HI(net421));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[9]$_DFFE_PP__422  (.L_HI(net422));
 sg13g2_tiehi \i_tinyqv.cpu.data_continue$_DFF_P__423  (.L_HI(net423));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[0]$_DFFE_PP__424  (.L_HI(net424));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[10]$_DFFE_PP__425  (.L_HI(net425));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[11]$_DFFE_PP__426  (.L_HI(net426));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[12]$_DFFE_PP__427  (.L_HI(net427));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[13]$_DFFE_PP__428  (.L_HI(net428));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[14]$_DFFE_PP__429  (.L_HI(net429));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[15]$_DFFE_PP__430  (.L_HI(net430));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[16]$_DFFE_PP__431  (.L_HI(net431));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[17]$_DFFE_PP__432  (.L_HI(net432));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[18]$_DFFE_PP__433  (.L_HI(net433));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[19]$_DFFE_PP__434  (.L_HI(net434));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[1]$_DFFE_PP__435  (.L_HI(net435));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[20]$_DFFE_PP__436  (.L_HI(net436));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[21]$_DFFE_PP__437  (.L_HI(net437));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[22]$_DFFE_PP__438  (.L_HI(net438));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[23]$_DFFE_PP__439  (.L_HI(net439));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[24]$_DFFE_PP__440  (.L_HI(net440));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[25]$_DFFE_PP__441  (.L_HI(net441));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[26]$_DFFE_PP__442  (.L_HI(net442));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[27]$_DFFE_PP__443  (.L_HI(net443));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[28]$_DFFE_PP__444  (.L_HI(net444));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[29]$_DFFE_PP__445  (.L_HI(net445));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[2]$_DFFE_PP__446  (.L_HI(net446));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[30]$_DFFE_PP__447  (.L_HI(net447));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[31]$_DFFE_PP__448  (.L_HI(net448));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[3]$_DFFE_PP__449  (.L_HI(net449));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[4]$_DFFE_PP__450  (.L_HI(net450));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[5]$_DFFE_PP__451  (.L_HI(net451));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[6]$_DFFE_PP__452  (.L_HI(net452));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[7]$_DFFE_PP__453  (.L_HI(net453));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[8]$_DFFE_PP__454  (.L_HI(net454));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[9]$_DFFE_PP__455  (.L_HI(net455));
 sg13g2_tiehi \i_tinyqv.cpu.data_read_n[0]$_SDFFE_PP1P__456  (.L_HI(net456));
 sg13g2_tiehi \i_tinyqv.cpu.data_read_n[1]$_SDFFE_PP1P__457  (.L_HI(net457));
 sg13g2_tiehi \i_tinyqv.cpu.data_ready_core$_SDFFE_PN0P__458  (.L_HI(net458));
 sg13g2_tiehi \i_tinyqv.cpu.data_ready_latch$_SDFF_PP0__459  (.L_HI(net459));
 sg13g2_tiehi \i_tinyqv.cpu.data_write_n[0]$_SDFFE_PN1P__460  (.L_HI(net460));
 sg13g2_tiehi \i_tinyqv.cpu.data_write_n[1]$_SDFFE_PN1P__461  (.L_HI(net461));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.cmp$_DFF_P__462  (.L_HI(net462));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.cy$_DFF_P__463  (.L_HI(net463));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.cycle[0]$_SDFFE_PN0P__464  (.L_HI(net464));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.cycle[1]$_SDFFE_PN0P__465  (.L_HI(net465));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.cy$_SDFF_PN0__466  (.L_HI(net466));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[0]$_SDFF_PN0__467  (.L_HI(net467));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[10]$_DFF_P__468  (.L_HI(net468));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[11]$_DFF_P__469  (.L_HI(net469));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[12]$_DFF_P__470  (.L_HI(net470));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[13]$_DFF_P__471  (.L_HI(net471));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[14]$_DFF_P__472  (.L_HI(net472));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[15]$_DFF_P__473  (.L_HI(net473));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[16]$_DFF_P__474  (.L_HI(net474));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[17]$_DFF_P__475  (.L_HI(net475));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[18]$_DFF_P__476  (.L_HI(net476));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[19]$_DFF_P__477  (.L_HI(net477));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[1]$_SDFF_PN0__478  (.L_HI(net478));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[20]$_DFF_P__479  (.L_HI(net479));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[21]$_DFF_P__480  (.L_HI(net480));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[22]$_DFF_P__481  (.L_HI(net481));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[23]$_DFF_P__482  (.L_HI(net482));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[24]$_DFF_P__483  (.L_HI(net483));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[25]$_DFF_P__484  (.L_HI(net484));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[26]$_DFF_P__485  (.L_HI(net485));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[27]$_DFF_P__486  (.L_HI(net486));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[28]$_DFF_P__487  (.L_HI(net487));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[29]$_DFF_P__488  (.L_HI(net488));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[2]$_SDFF_PN0__489  (.L_HI(net489));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[30]$_DFF_P__490  (.L_HI(net490));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[31]$_DFF_P__491  (.L_HI(net491));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[3]$_SDFF_PN0__492  (.L_HI(net492));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[4]$_DFF_P__493  (.L_HI(net493));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[5]$_DFF_P__494  (.L_HI(net494));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[6]$_DFF_P__495  (.L_HI(net495));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[7]$_DFF_P__496  (.L_HI(net496));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[8]$_DFF_P__497  (.L_HI(net497));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[9]$_DFF_P__498  (.L_HI(net498));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.cy$_SDFF_PN0__499  (.L_HI(net499));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[0]$_SDFF_PN0__500  (.L_HI(net500));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[10]$_DFF_P__501  (.L_HI(net501));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[11]$_DFF_P__502  (.L_HI(net502));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[12]$_DFF_P__503  (.L_HI(net503));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[13]$_DFF_P__504  (.L_HI(net504));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[14]$_DFF_P__505  (.L_HI(net505));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[15]$_DFF_P__506  (.L_HI(net506));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[16]$_DFF_P__507  (.L_HI(net507));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[17]$_DFF_P__508  (.L_HI(net508));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[18]$_DFF_P__509  (.L_HI(net509));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[19]$_DFF_P__510  (.L_HI(net510));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[1]$_SDFF_PN0__511  (.L_HI(net511));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[20]$_DFF_P__512  (.L_HI(net512));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[21]$_DFF_P__513  (.L_HI(net513));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[22]$_DFF_P__514  (.L_HI(net514));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[23]$_DFF_P__515  (.L_HI(net515));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[24]$_DFF_P__516  (.L_HI(net516));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[25]$_DFF_P__517  (.L_HI(net517));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[26]$_DFF_P__518  (.L_HI(net518));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[27]$_DFF_P__519  (.L_HI(net519));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[28]$_DFF_P__520  (.L_HI(net520));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[29]$_DFF_P__521  (.L_HI(net521));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[2]$_SDFF_PN0__522  (.L_HI(net522));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[30]$_DFF_P__523  (.L_HI(net523));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[31]$_DFF_P__524  (.L_HI(net524));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[3]$_SDFF_PN0__525  (.L_HI(net525));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[4]$_DFF_P__526  (.L_HI(net526));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[5]$_DFF_P__527  (.L_HI(net527));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[6]$_DFF_P__528  (.L_HI(net528));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[7]$_DFF_P__529  (.L_HI(net529));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[8]$_DFF_P__530  (.L_HI(net530));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[9]$_DFF_P__531  (.L_HI(net531));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][0]$_DFF_P__532  (.L_HI(net532));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][10]$_DFF_P__533  (.L_HI(net533));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][11]$_DFF_P__534  (.L_HI(net534));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][12]$_DFF_P__535  (.L_HI(net535));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][13]$_DFF_P__536  (.L_HI(net536));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][14]$_DFF_P__537  (.L_HI(net537));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][15]$_DFF_P__538  (.L_HI(net538));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][16]$_DFF_P__539  (.L_HI(net539));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][17]$_DFF_P__540  (.L_HI(net540));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][18]$_DFF_P__541  (.L_HI(net541));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][19]$_DFF_P__542  (.L_HI(net542));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][1]$_DFF_P__543  (.L_HI(net543));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][20]$_DFF_P__544  (.L_HI(net544));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][21]$_DFF_P__545  (.L_HI(net545));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][22]$_DFF_P__546  (.L_HI(net546));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][23]$_DFF_P__547  (.L_HI(net547));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][24]$_DFF_P__548  (.L_HI(net548));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][25]$_DFF_P__549  (.L_HI(net549));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][26]$_DFF_P__550  (.L_HI(net550));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][27]$_DFF_P__551  (.L_HI(net551));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][28]$_DFF_P__552  (.L_HI(net552));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][29]$_DFF_P__553  (.L_HI(net553));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][2]$_DFF_P__554  (.L_HI(net554));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][30]$_DFF_P__555  (.L_HI(net555));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][31]$_DFF_P__556  (.L_HI(net556));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][3]$_DFF_P__557  (.L_HI(net557));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][4]$_DFF_P__558  (.L_HI(net558));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][5]$_DFF_P__559  (.L_HI(net559));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][6]$_DFF_P__560  (.L_HI(net560));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][7]$_DFF_P__561  (.L_HI(net561));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][8]$_DFF_P__562  (.L_HI(net562));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][9]$_DFF_P__563  (.L_HI(net563));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][0]$_DFF_P__564  (.L_HI(net564));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][10]$_DFF_P__565  (.L_HI(net565));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][11]$_DFF_P__566  (.L_HI(net566));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][12]$_DFF_P__567  (.L_HI(net567));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][13]$_DFF_P__568  (.L_HI(net568));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][14]$_DFF_P__569  (.L_HI(net569));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][15]$_DFF_P__570  (.L_HI(net570));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][16]$_DFF_P__571  (.L_HI(net571));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][17]$_DFF_P__572  (.L_HI(net572));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][18]$_DFF_P__573  (.L_HI(net573));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][19]$_DFF_P__574  (.L_HI(net574));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][1]$_DFF_P__575  (.L_HI(net575));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][20]$_DFF_P__576  (.L_HI(net576));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][21]$_DFF_P__577  (.L_HI(net577));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][22]$_DFF_P__578  (.L_HI(net578));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][23]$_DFF_P__579  (.L_HI(net579));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][24]$_DFF_P__580  (.L_HI(net580));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][25]$_DFF_P__581  (.L_HI(net581));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][26]$_DFF_P__582  (.L_HI(net582));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][27]$_DFF_P__583  (.L_HI(net583));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][28]$_DFF_P__584  (.L_HI(net584));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][29]$_DFF_P__585  (.L_HI(net585));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][2]$_DFF_P__586  (.L_HI(net586));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][30]$_DFF_P__587  (.L_HI(net587));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][31]$_DFF_P__588  (.L_HI(net588));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][3]$_DFF_P__589  (.L_HI(net589));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][4]$_DFF_P__590  (.L_HI(net590));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][5]$_DFF_P__591  (.L_HI(net591));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][6]$_DFF_P__592  (.L_HI(net592));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][7]$_DFF_P__593  (.L_HI(net593));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][8]$_DFF_P__594  (.L_HI(net594));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][9]$_DFF_P__595  (.L_HI(net595));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][0]$_DFF_P__596  (.L_HI(net596));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][10]$_DFF_P__597  (.L_HI(net597));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][11]$_DFF_P__598  (.L_HI(net598));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][12]$_DFF_P__599  (.L_HI(net599));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][13]$_DFF_P__600  (.L_HI(net600));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][14]$_DFF_P__601  (.L_HI(net601));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][15]$_DFF_P__602  (.L_HI(net602));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][16]$_DFF_P__603  (.L_HI(net603));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][17]$_DFF_P__604  (.L_HI(net604));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][18]$_DFF_P__605  (.L_HI(net605));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][19]$_DFF_P__606  (.L_HI(net606));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][1]$_DFF_P__607  (.L_HI(net607));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][20]$_DFF_P__608  (.L_HI(net608));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][21]$_DFF_P__609  (.L_HI(net609));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][22]$_DFF_P__610  (.L_HI(net610));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][23]$_DFF_P__611  (.L_HI(net611));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][24]$_DFF_P__612  (.L_HI(net612));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][25]$_DFF_P__613  (.L_HI(net613));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][26]$_DFF_P__614  (.L_HI(net614));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][27]$_DFF_P__615  (.L_HI(net615));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][28]$_DFF_P__616  (.L_HI(net616));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][29]$_DFF_P__617  (.L_HI(net617));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][2]$_DFF_P__618  (.L_HI(net618));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][30]$_DFF_P__619  (.L_HI(net619));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][31]$_DFF_P__620  (.L_HI(net620));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][3]$_DFF_P__621  (.L_HI(net621));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][4]$_DFF_P__622  (.L_HI(net622));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][5]$_DFF_P__623  (.L_HI(net623));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][6]$_DFF_P__624  (.L_HI(net624));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][7]$_DFF_P__625  (.L_HI(net625));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][8]$_DFF_P__626  (.L_HI(net626));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][9]$_DFF_P__627  (.L_HI(net627));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][0]$_DFF_P__628  (.L_HI(net628));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][10]$_DFF_P__629  (.L_HI(net629));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][11]$_DFF_P__630  (.L_HI(net630));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][12]$_DFF_P__631  (.L_HI(net631));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][13]$_DFF_P__632  (.L_HI(net632));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][14]$_DFF_P__633  (.L_HI(net633));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][15]$_DFF_P__634  (.L_HI(net634));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][16]$_DFF_P__635  (.L_HI(net635));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][17]$_DFF_P__636  (.L_HI(net636));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][18]$_DFF_P__637  (.L_HI(net637));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][19]$_DFF_P__638  (.L_HI(net638));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][1]$_DFF_P__639  (.L_HI(net639));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][20]$_DFF_P__640  (.L_HI(net640));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][21]$_DFF_P__641  (.L_HI(net641));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][22]$_DFF_P__642  (.L_HI(net642));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][23]$_DFF_P__643  (.L_HI(net643));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][24]$_DFF_P__644  (.L_HI(net644));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][25]$_DFF_P__645  (.L_HI(net645));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][26]$_DFF_P__646  (.L_HI(net646));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][27]$_DFF_P__647  (.L_HI(net647));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][28]$_DFF_P__648  (.L_HI(net648));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][29]$_DFF_P__649  (.L_HI(net649));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][2]$_DFF_P__650  (.L_HI(net650));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][30]$_DFF_P__651  (.L_HI(net651));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][31]$_DFF_P__652  (.L_HI(net652));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][3]$_DFF_P__653  (.L_HI(net653));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][4]$_DFF_P__654  (.L_HI(net654));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][5]$_DFF_P__655  (.L_HI(net655));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][6]$_DFF_P__656  (.L_HI(net656));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][7]$_DFF_P__657  (.L_HI(net657));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][8]$_DFF_P__658  (.L_HI(net658));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][9]$_DFF_P__659  (.L_HI(net659));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][0]$_DFF_P__660  (.L_HI(net660));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][10]$_DFF_P__661  (.L_HI(net661));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][11]$_DFF_P__662  (.L_HI(net662));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][12]$_DFF_P__663  (.L_HI(net663));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][13]$_DFF_P__664  (.L_HI(net664));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][14]$_DFF_P__665  (.L_HI(net665));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][15]$_DFF_P__666  (.L_HI(net666));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][16]$_DFF_P__667  (.L_HI(net667));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][17]$_DFF_P__668  (.L_HI(net668));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][18]$_DFF_P__669  (.L_HI(net669));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][19]$_DFF_P__670  (.L_HI(net670));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][1]$_DFF_P__671  (.L_HI(net671));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][20]$_DFF_P__672  (.L_HI(net672));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][21]$_DFF_P__673  (.L_HI(net673));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][22]$_DFF_P__674  (.L_HI(net674));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][23]$_DFF_P__675  (.L_HI(net675));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][24]$_DFF_P__676  (.L_HI(net676));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][25]$_DFF_P__677  (.L_HI(net677));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][26]$_DFF_P__678  (.L_HI(net678));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][27]$_DFF_P__679  (.L_HI(net679));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][28]$_DFF_P__680  (.L_HI(net680));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][29]$_DFF_P__681  (.L_HI(net681));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][2]$_DFF_P__682  (.L_HI(net682));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][30]$_DFF_P__683  (.L_HI(net683));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][31]$_DFF_P__684  (.L_HI(net684));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][3]$_DFF_P__685  (.L_HI(net685));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][4]$_DFF_P__686  (.L_HI(net686));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][5]$_DFF_P__687  (.L_HI(net687));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][6]$_DFF_P__688  (.L_HI(net688));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][7]$_DFF_P__689  (.L_HI(net689));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][8]$_DFF_P__690  (.L_HI(net690));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][9]$_DFF_P__691  (.L_HI(net691));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][0]$_DFF_P__692  (.L_HI(net692));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][10]$_DFF_P__693  (.L_HI(net693));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][11]$_DFF_P__694  (.L_HI(net694));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][12]$_DFF_P__695  (.L_HI(net695));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][13]$_DFF_P__696  (.L_HI(net696));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][14]$_DFF_P__697  (.L_HI(net697));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][15]$_DFF_P__698  (.L_HI(net698));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][16]$_DFF_P__699  (.L_HI(net699));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][17]$_DFF_P__700  (.L_HI(net700));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][18]$_DFF_P__701  (.L_HI(net701));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][19]$_DFF_P__702  (.L_HI(net702));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][1]$_DFF_P__703  (.L_HI(net703));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][20]$_DFF_P__704  (.L_HI(net704));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][21]$_DFF_P__705  (.L_HI(net705));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][22]$_DFF_P__706  (.L_HI(net706));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][23]$_DFF_P__707  (.L_HI(net707));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][24]$_DFF_P__708  (.L_HI(net708));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][25]$_DFF_P__709  (.L_HI(net709));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][26]$_DFF_P__710  (.L_HI(net710));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][27]$_DFF_P__711  (.L_HI(net711));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][28]$_DFF_P__712  (.L_HI(net712));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][29]$_DFF_P__713  (.L_HI(net713));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][2]$_DFF_P__714  (.L_HI(net714));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][30]$_DFF_P__715  (.L_HI(net715));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][31]$_DFF_P__716  (.L_HI(net716));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][3]$_DFF_P__717  (.L_HI(net717));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][4]$_DFF_P__718  (.L_HI(net718));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][5]$_DFF_P__719  (.L_HI(net719));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][6]$_DFF_P__720  (.L_HI(net720));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][7]$_DFF_P__721  (.L_HI(net721));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][8]$_DFF_P__722  (.L_HI(net722));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][9]$_DFF_P__723  (.L_HI(net723));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][0]$_DFF_P__724  (.L_HI(net724));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][10]$_DFF_P__725  (.L_HI(net725));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][11]$_DFF_P__726  (.L_HI(net726));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][12]$_DFF_P__727  (.L_HI(net727));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][13]$_DFF_P__728  (.L_HI(net728));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][14]$_DFF_P__729  (.L_HI(net729));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][15]$_DFF_P__730  (.L_HI(net730));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][16]$_DFF_P__731  (.L_HI(net731));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][17]$_DFF_P__732  (.L_HI(net732));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][18]$_DFF_P__733  (.L_HI(net733));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][19]$_DFF_P__734  (.L_HI(net734));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][1]$_DFF_P__735  (.L_HI(net735));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][20]$_DFF_P__736  (.L_HI(net736));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][21]$_DFF_P__737  (.L_HI(net737));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][22]$_DFF_P__738  (.L_HI(net738));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][23]$_DFF_P__739  (.L_HI(net739));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][24]$_DFF_P__740  (.L_HI(net740));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][25]$_DFF_P__741  (.L_HI(net741));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][26]$_DFF_P__742  (.L_HI(net742));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][27]$_DFF_P__743  (.L_HI(net743));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][28]$_DFF_P__744  (.L_HI(net744));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][29]$_DFF_P__745  (.L_HI(net745));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][2]$_DFF_P__746  (.L_HI(net746));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][30]$_DFF_P__747  (.L_HI(net747));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][31]$_DFF_P__748  (.L_HI(net748));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][3]$_DFF_P__749  (.L_HI(net749));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][4]$_DFF_P__750  (.L_HI(net750));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][5]$_DFF_P__751  (.L_HI(net751));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][6]$_DFF_P__752  (.L_HI(net752));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][7]$_DFF_P__753  (.L_HI(net753));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][8]$_DFF_P__754  (.L_HI(net754));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][9]$_DFF_P__755  (.L_HI(net755));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][0]$_DFF_P__756  (.L_HI(net756));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][10]$_DFF_P__757  (.L_HI(net757));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][11]$_DFF_P__758  (.L_HI(net758));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][12]$_DFF_P__759  (.L_HI(net759));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][13]$_DFF_P__760  (.L_HI(net760));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][14]$_DFF_P__761  (.L_HI(net761));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][15]$_DFF_P__762  (.L_HI(net762));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][16]$_DFF_P__763  (.L_HI(net763));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][17]$_DFF_P__764  (.L_HI(net764));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][18]$_DFF_P__765  (.L_HI(net765));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][19]$_DFF_P__766  (.L_HI(net766));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][1]$_DFF_P__767  (.L_HI(net767));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][20]$_DFF_P__768  (.L_HI(net768));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][21]$_DFF_P__769  (.L_HI(net769));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][22]$_DFF_P__770  (.L_HI(net770));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][23]$_DFF_P__771  (.L_HI(net771));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][24]$_DFF_P__772  (.L_HI(net772));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][25]$_DFF_P__773  (.L_HI(net773));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][26]$_DFF_P__774  (.L_HI(net774));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][27]$_DFF_P__775  (.L_HI(net775));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][28]$_DFF_P__776  (.L_HI(net776));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][29]$_DFF_P__777  (.L_HI(net777));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][2]$_DFF_P__778  (.L_HI(net778));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][30]$_DFF_P__779  (.L_HI(net779));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][31]$_DFF_P__780  (.L_HI(net780));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][3]$_DFF_P__781  (.L_HI(net781));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][4]$_DFF_P__782  (.L_HI(net782));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][5]$_DFF_P__783  (.L_HI(net783));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][6]$_DFF_P__784  (.L_HI(net784));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][7]$_DFF_P__785  (.L_HI(net785));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][8]$_DFF_P__786  (.L_HI(net786));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][9]$_DFF_P__787  (.L_HI(net787));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][0]$_DFF_P__788  (.L_HI(net788));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][10]$_DFF_P__789  (.L_HI(net789));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][11]$_DFF_P__790  (.L_HI(net790));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][12]$_DFF_P__791  (.L_HI(net791));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][13]$_DFF_P__792  (.L_HI(net792));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][14]$_DFF_P__793  (.L_HI(net793));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][15]$_DFF_P__794  (.L_HI(net794));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][16]$_DFF_P__795  (.L_HI(net795));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][17]$_DFF_P__796  (.L_HI(net796));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][18]$_DFF_P__797  (.L_HI(net797));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][19]$_DFF_P__798  (.L_HI(net798));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][1]$_DFF_P__799  (.L_HI(net799));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][20]$_DFF_P__800  (.L_HI(net800));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][21]$_DFF_P__801  (.L_HI(net801));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][22]$_DFF_P__802  (.L_HI(net802));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][23]$_DFF_P__803  (.L_HI(net803));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][24]$_DFF_P__804  (.L_HI(net804));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][25]$_DFF_P__805  (.L_HI(net805));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][26]$_DFF_P__806  (.L_HI(net806));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][27]$_DFF_P__807  (.L_HI(net807));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][28]$_DFF_P__808  (.L_HI(net808));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][29]$_DFF_P__809  (.L_HI(net809));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][2]$_DFF_P__810  (.L_HI(net810));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][30]$_DFF_P__811  (.L_HI(net811));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][31]$_DFF_P__812  (.L_HI(net812));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][3]$_DFF_P__813  (.L_HI(net813));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][4]$_DFF_P__814  (.L_HI(net814));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][5]$_DFF_P__815  (.L_HI(net815));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][6]$_DFF_P__816  (.L_HI(net816));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][7]$_DFF_P__817  (.L_HI(net817));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][8]$_DFF_P__818  (.L_HI(net818));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][9]$_DFF_P__819  (.L_HI(net819));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][0]$_DFF_P__820  (.L_HI(net820));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][10]$_DFF_P__821  (.L_HI(net821));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][11]$_DFF_P__822  (.L_HI(net822));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][12]$_DFF_P__823  (.L_HI(net823));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][13]$_DFF_P__824  (.L_HI(net824));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][14]$_DFF_P__825  (.L_HI(net825));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][15]$_DFF_P__826  (.L_HI(net826));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][16]$_DFF_P__827  (.L_HI(net827));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][17]$_DFF_P__828  (.L_HI(net828));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][18]$_DFF_P__829  (.L_HI(net829));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][19]$_DFF_P__830  (.L_HI(net830));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][1]$_DFF_P__831  (.L_HI(net831));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][20]$_DFF_P__832  (.L_HI(net832));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][21]$_DFF_P__833  (.L_HI(net833));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][22]$_DFF_P__834  (.L_HI(net834));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][23]$_DFF_P__835  (.L_HI(net835));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][24]$_DFF_P__836  (.L_HI(net836));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][25]$_DFF_P__837  (.L_HI(net837));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][26]$_DFF_P__838  (.L_HI(net838));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][27]$_DFF_P__839  (.L_HI(net839));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][28]$_DFF_P__840  (.L_HI(net840));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][29]$_DFF_P__841  (.L_HI(net841));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][2]$_DFF_P__842  (.L_HI(net842));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][30]$_DFF_P__843  (.L_HI(net843));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][31]$_DFF_P__844  (.L_HI(net844));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][3]$_DFF_P__845  (.L_HI(net845));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][4]$_DFF_P__846  (.L_HI(net846));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][5]$_DFF_P__847  (.L_HI(net847));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][6]$_DFF_P__848  (.L_HI(net848));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][7]$_DFF_P__849  (.L_HI(net849));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][8]$_DFF_P__850  (.L_HI(net850));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][9]$_DFF_P__851  (.L_HI(net851));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][0]$_DFF_P__852  (.L_HI(net852));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][10]$_DFF_P__853  (.L_HI(net853));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][11]$_DFF_P__854  (.L_HI(net854));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][12]$_DFF_P__855  (.L_HI(net855));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][13]$_DFF_P__856  (.L_HI(net856));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][14]$_DFF_P__857  (.L_HI(net857));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][15]$_DFF_P__858  (.L_HI(net858));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][16]$_DFF_P__859  (.L_HI(net859));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][17]$_DFF_P__860  (.L_HI(net860));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][18]$_DFF_P__861  (.L_HI(net861));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][19]$_DFF_P__862  (.L_HI(net862));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][1]$_DFF_P__863  (.L_HI(net863));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][20]$_DFF_P__864  (.L_HI(net864));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][21]$_DFF_P__865  (.L_HI(net865));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][22]$_DFF_P__866  (.L_HI(net866));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][23]$_DFF_P__867  (.L_HI(net867));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][24]$_DFF_P__868  (.L_HI(net868));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][25]$_DFF_P__869  (.L_HI(net869));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][26]$_DFF_P__870  (.L_HI(net870));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][27]$_DFF_P__871  (.L_HI(net871));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][28]$_DFF_P__872  (.L_HI(net872));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][29]$_DFF_P__873  (.L_HI(net873));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][2]$_DFF_P__874  (.L_HI(net874));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][30]$_DFF_P__875  (.L_HI(net875));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][31]$_DFF_P__876  (.L_HI(net876));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][3]$_DFF_P__877  (.L_HI(net877));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][4]$_DFF_P__878  (.L_HI(net878));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][5]$_DFF_P__879  (.L_HI(net879));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][6]$_DFF_P__880  (.L_HI(net880));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][7]$_DFF_P__881  (.L_HI(net881));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][8]$_DFF_P__882  (.L_HI(net882));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][9]$_DFF_P__883  (.L_HI(net883));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][0]$_DFF_P__884  (.L_HI(net884));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][10]$_DFF_P__885  (.L_HI(net885));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][11]$_DFF_P__886  (.L_HI(net886));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][12]$_DFF_P__887  (.L_HI(net887));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][13]$_DFF_P__888  (.L_HI(net888));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][14]$_DFF_P__889  (.L_HI(net889));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][15]$_DFF_P__890  (.L_HI(net890));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][16]$_DFF_P__891  (.L_HI(net891));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][17]$_DFF_P__892  (.L_HI(net892));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][18]$_DFF_P__893  (.L_HI(net893));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][19]$_DFF_P__894  (.L_HI(net894));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][1]$_DFF_P__895  (.L_HI(net895));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][20]$_DFF_P__896  (.L_HI(net896));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][21]$_DFF_P__897  (.L_HI(net897));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][22]$_DFF_P__898  (.L_HI(net898));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][23]$_DFF_P__899  (.L_HI(net899));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][24]$_DFF_P__900  (.L_HI(net900));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][25]$_DFF_P__901  (.L_HI(net901));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][26]$_DFF_P__902  (.L_HI(net902));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][27]$_DFF_P__903  (.L_HI(net903));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][28]$_DFF_P__904  (.L_HI(net904));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][29]$_DFF_P__905  (.L_HI(net905));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][2]$_DFF_P__906  (.L_HI(net906));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][30]$_DFF_P__907  (.L_HI(net907));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][31]$_DFF_P__908  (.L_HI(net908));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][3]$_DFF_P__909  (.L_HI(net909));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][4]$_DFF_P__910  (.L_HI(net910));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][5]$_DFF_P__911  (.L_HI(net911));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][6]$_DFF_P__912  (.L_HI(net912));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][7]$_DFF_P__913  (.L_HI(net913));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][8]$_DFF_P__914  (.L_HI(net914));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][9]$_DFF_P__915  (.L_HI(net915));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][0]$_DFF_P__916  (.L_HI(net916));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][10]$_DFF_P__917  (.L_HI(net917));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][11]$_DFF_P__918  (.L_HI(net918));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][12]$_DFF_P__919  (.L_HI(net919));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][13]$_DFF_P__920  (.L_HI(net920));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][14]$_DFF_P__921  (.L_HI(net921));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][15]$_DFF_P__922  (.L_HI(net922));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][16]$_DFF_P__923  (.L_HI(net923));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][17]$_DFF_P__924  (.L_HI(net924));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][18]$_DFF_P__925  (.L_HI(net925));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][19]$_DFF_P__926  (.L_HI(net926));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][1]$_DFF_P__927  (.L_HI(net927));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][20]$_DFF_P__928  (.L_HI(net928));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][21]$_DFF_P__929  (.L_HI(net929));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][22]$_DFF_P__930  (.L_HI(net930));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][23]$_DFF_P__931  (.L_HI(net931));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][24]$_DFF_P__932  (.L_HI(net932));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][25]$_DFF_P__933  (.L_HI(net933));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][26]$_DFF_P__934  (.L_HI(net934));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][27]$_DFF_P__935  (.L_HI(net935));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][28]$_DFF_P__936  (.L_HI(net936));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][29]$_DFF_P__937  (.L_HI(net937));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][2]$_DFF_P__938  (.L_HI(net938));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][30]$_DFF_P__939  (.L_HI(net939));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][31]$_DFF_P__940  (.L_HI(net940));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][3]$_DFF_P__941  (.L_HI(net941));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][4]$_DFF_P__942  (.L_HI(net942));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][5]$_DFF_P__943  (.L_HI(net943));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][6]$_DFF_P__944  (.L_HI(net944));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][7]$_DFF_P__945  (.L_HI(net945));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][8]$_DFF_P__946  (.L_HI(net946));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][9]$_DFF_P__947  (.L_HI(net947));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.instr_retired$_DFF_P__948  (.L_HI(net948));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.is_double_fault_r$_DFFE_PP__949  (.L_HI(net949));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.last_interrupt_req[0]$_DFFE_PP__950  (.L_HI(net950));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.last_interrupt_req[1]$_DFFE_PP__951  (.L_HI(net951));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.load_done$_DFFE_PP__952  (.L_HI(net952));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.load_top_bit$_SDFFCE_PN0P__953  (.L_HI(net953));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mcause[0]$_SDFFE_PN0P__954  (.L_HI(net954));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mcause[1]$_SDFFE_PN0P__955  (.L_HI(net955));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mcause[3]$_SDFFE_PN0P__956  (.L_HI(net956));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mcause[4]$_SDFFE_PN0P__957  (.L_HI(net957));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[0]$_DFFE_PN__958  (.L_HI(net958));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[10]$_DFFE_PN__959  (.L_HI(net959));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[11]$_DFFE_PN__960  (.L_HI(net960));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[12]$_DFFE_PN__961  (.L_HI(net961));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[13]$_DFFE_PN__962  (.L_HI(net962));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[14]$_DFFE_PN__963  (.L_HI(net963));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[15]$_DFFE_PN__964  (.L_HI(net964));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[16]$_DFFE_PN__965  (.L_HI(net965));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[17]$_DFFE_PN__966  (.L_HI(net966));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[18]$_DFFE_PN__967  (.L_HI(net967));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[19]$_DFFE_PN__968  (.L_HI(net968));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[1]$_DFFE_PN__969  (.L_HI(net969));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[20]$_SDFFCE_PN0N__970  (.L_HI(net970));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[21]$_SDFFCE_PN0N__971  (.L_HI(net971));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[22]$_SDFFCE_PN0N__972  (.L_HI(net972));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[23]$_SDFFCE_PN0N__973  (.L_HI(net973));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[2]$_DFFE_PN__974  (.L_HI(net974));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[3]$_DFFE_PN__975  (.L_HI(net975));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[4]$_DFFE_PN__976  (.L_HI(net976));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[5]$_DFFE_PN__977  (.L_HI(net977));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[6]$_DFFE_PN__978  (.L_HI(net978));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[7]$_DFFE_PN__979  (.L_HI(net979));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[8]$_DFFE_PN__980  (.L_HI(net980));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[9]$_DFFE_PN__981  (.L_HI(net981));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mstatus_mie$_SDFFE_PP1P__982  (.L_HI(net982));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mstatus_mpie$_SDFFE_PP0P__983  (.L_HI(net983));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mstatus_mte$_SDFFE_PP1P__984  (.L_HI(net984));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[0]$_DFF_P__985  (.L_HI(net985));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[10]$_DFF_P__986  (.L_HI(net986));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[11]$_DFF_P__987  (.L_HI(net987));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[12]$_SDFF_PP0__988  (.L_HI(net988));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[13]$_SDFF_PP0__989  (.L_HI(net989));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[14]$_SDFF_PP0__990  (.L_HI(net990));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[15]$_SDFF_PP0__991  (.L_HI(net991));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[1]$_DFF_P__992  (.L_HI(net992));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[2]$_DFF_P__993  (.L_HI(net993));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[3]$_DFF_P__994  (.L_HI(net994));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[4]$_DFF_P__995  (.L_HI(net995));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[5]$_DFF_P__996  (.L_HI(net996));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[6]$_DFF_P__997  (.L_HI(net997));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[7]$_DFF_P__998  (.L_HI(net998));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[8]$_DFF_P__999  (.L_HI(net999));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[9]$_DFF_P__1000  (.L_HI(net1000));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[0]$_DFFE_PP__1001  (.L_HI(net1001));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[1]$_DFFE_PP__1002  (.L_HI(net1002));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[2]$_DFFE_PP__1003  (.L_HI(net1003));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[3]$_DFFE_PP__1004  (.L_HI(net1004));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[4]$_DFFE_PP__1005  (.L_HI(net1005));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.time_hi[0]$_SDFFE_PN0P__1006  (.L_HI(net1006));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.time_hi[1]$_SDFFE_PN0P__1007  (.L_HI(net1007));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.time_hi[2]$_SDFFE_PN0P__1008  (.L_HI(net1008));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[0]$_DFFE_PN__1009  (.L_HI(net1009));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[10]$_DFFE_PN__1010  (.L_HI(net1010));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[11]$_DFFE_PN__1011  (.L_HI(net1011));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[12]$_DFFE_PN__1012  (.L_HI(net1012));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[13]$_DFFE_PN__1013  (.L_HI(net1013));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[14]$_DFFE_PN__1014  (.L_HI(net1014));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[15]$_DFFE_PN__1015  (.L_HI(net1015));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[16]$_DFFE_PN__1016  (.L_HI(net1016));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[17]$_DFFE_PN__1017  (.L_HI(net1017));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[18]$_DFFE_PN__1018  (.L_HI(net1018));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[19]$_DFFE_PN__1019  (.L_HI(net1019));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[1]$_DFFE_PN__1020  (.L_HI(net1020));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[20]$_DFFE_PN__1021  (.L_HI(net1021));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[21]$_DFFE_PN__1022  (.L_HI(net1022));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[22]$_DFFE_PN__1023  (.L_HI(net1023));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[23]$_DFFE_PN__1024  (.L_HI(net1024));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[24]$_DFFE_PN__1025  (.L_HI(net1025));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[25]$_DFFE_PN__1026  (.L_HI(net1026));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[26]$_DFFE_PN__1027  (.L_HI(net1027));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[27]$_DFFE_PN__1028  (.L_HI(net1028));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[28]$_SDFFCE_PN0N__1029  (.L_HI(net1029));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[29]$_SDFFCE_PN0N__1030  (.L_HI(net1030));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[2]$_DFFE_PN__1031  (.L_HI(net1031));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[30]$_DFFE_PN__1032  (.L_HI(net1032));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[31]$_DFFE_PN__1033  (.L_HI(net1033));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[3]$_DFFE_PN__1034  (.L_HI(net1034));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[4]$_DFFE_PN__1035  (.L_HI(net1035));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[5]$_DFFE_PN__1036  (.L_HI(net1036));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[6]$_DFFE_PN__1037  (.L_HI(net1037));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[7]$_DFFE_PN__1038  (.L_HI(net1038));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[8]$_DFFE_PN__1039  (.L_HI(net1039));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[9]$_DFFE_PN__1040  (.L_HI(net1040));
 sg13g2_tiehi \i_tinyqv.cpu.imm[0]$_DFFE_PP__1041  (.L_HI(net1041));
 sg13g2_tiehi \i_tinyqv.cpu.imm[10]$_DFFE_PP__1042  (.L_HI(net1042));
 sg13g2_tiehi \i_tinyqv.cpu.imm[11]$_DFFE_PP__1043  (.L_HI(net1043));
 sg13g2_tiehi \i_tinyqv.cpu.imm[12]$_DFFE_PP__1044  (.L_HI(net1044));
 sg13g2_tiehi \i_tinyqv.cpu.imm[13]$_DFFE_PP__1045  (.L_HI(net1045));
 sg13g2_tiehi \i_tinyqv.cpu.imm[14]$_DFFE_PP__1046  (.L_HI(net1046));
 sg13g2_tiehi \i_tinyqv.cpu.imm[15]$_DFFE_PP__1047  (.L_HI(net1047));
 sg13g2_tiehi \i_tinyqv.cpu.imm[16]$_DFFE_PP__1048  (.L_HI(net1048));
 sg13g2_tiehi \i_tinyqv.cpu.imm[17]$_DFFE_PP__1049  (.L_HI(net1049));
 sg13g2_tiehi \i_tinyqv.cpu.imm[18]$_DFFE_PP__1050  (.L_HI(net1050));
 sg13g2_tiehi \i_tinyqv.cpu.imm[19]$_DFFE_PP__1051  (.L_HI(net1051));
 sg13g2_tiehi \i_tinyqv.cpu.imm[1]$_DFFE_PP__1052  (.L_HI(net1052));
 sg13g2_tiehi \i_tinyqv.cpu.imm[20]$_DFFE_PP__1053  (.L_HI(net1053));
 sg13g2_tiehi \i_tinyqv.cpu.imm[21]$_DFFE_PP__1054  (.L_HI(net1054));
 sg13g2_tiehi \i_tinyqv.cpu.imm[22]$_DFFE_PP__1055  (.L_HI(net1055));
 sg13g2_tiehi \i_tinyqv.cpu.imm[23]$_DFFE_PP__1056  (.L_HI(net1056));
 sg13g2_tiehi \i_tinyqv.cpu.imm[24]$_DFFE_PP__1057  (.L_HI(net1057));
 sg13g2_tiehi \i_tinyqv.cpu.imm[25]$_DFFE_PP__1058  (.L_HI(net1058));
 sg13g2_tiehi \i_tinyqv.cpu.imm[26]$_DFFE_PP__1059  (.L_HI(net1059));
 sg13g2_tiehi \i_tinyqv.cpu.imm[27]$_DFFE_PP__1060  (.L_HI(net1060));
 sg13g2_tiehi \i_tinyqv.cpu.imm[28]$_DFFE_PP__1061  (.L_HI(net1061));
 sg13g2_tiehi \i_tinyqv.cpu.imm[29]$_DFFE_PP__1062  (.L_HI(net1062));
 sg13g2_tiehi \i_tinyqv.cpu.imm[2]$_DFFE_PP__1063  (.L_HI(net1063));
 sg13g2_tiehi \i_tinyqv.cpu.imm[30]$_DFFE_PP__1064  (.L_HI(net1064));
 sg13g2_tiehi \i_tinyqv.cpu.imm[31]$_DFFE_PP__1065  (.L_HI(net1065));
 sg13g2_tiehi \i_tinyqv.cpu.imm[3]$_DFFE_PP__1066  (.L_HI(net1066));
 sg13g2_tiehi \i_tinyqv.cpu.imm[4]$_DFFE_PP__1067  (.L_HI(net1067));
 sg13g2_tiehi \i_tinyqv.cpu.imm[5]$_DFFE_PP__1068  (.L_HI(net1068));
 sg13g2_tiehi \i_tinyqv.cpu.imm[6]$_DFFE_PP__1069  (.L_HI(net1069));
 sg13g2_tiehi \i_tinyqv.cpu.imm[7]$_DFFE_PP__1070  (.L_HI(net1070));
 sg13g2_tiehi \i_tinyqv.cpu.imm[8]$_DFFE_PP__1071  (.L_HI(net1071));
 sg13g2_tiehi \i_tinyqv.cpu.imm[9]$_DFFE_PP__1072  (.L_HI(net1072));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][0]$_SDFFCE_PN1P__1073  (.L_HI(net1073));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][10]$_DFFE_PP__1074  (.L_HI(net1074));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][11]$_DFFE_PP__1075  (.L_HI(net1075));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][12]$_DFFE_PP__1076  (.L_HI(net1076));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][13]$_DFFE_PP__1077  (.L_HI(net1077));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][14]$_DFFE_PP__1078  (.L_HI(net1078));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][15]$_DFFE_PP__1079  (.L_HI(net1079));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][1]$_SDFFCE_PN1P__1080  (.L_HI(net1080));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][2]$_DFFE_PP__1081  (.L_HI(net1081));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][3]$_DFFE_PP__1082  (.L_HI(net1082));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][4]$_DFFE_PP__1083  (.L_HI(net1083));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][5]$_DFFE_PP__1084  (.L_HI(net1084));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][6]$_DFFE_PP__1085  (.L_HI(net1085));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][7]$_DFFE_PP__1086  (.L_HI(net1086));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][8]$_DFFE_PP__1087  (.L_HI(net1087));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][9]$_DFFE_PP__1088  (.L_HI(net1088));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][0]$_SDFFCE_PN1P__1089  (.L_HI(net1089));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][10]$_DFFE_PP__1090  (.L_HI(net1090));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][11]$_DFFE_PP__1091  (.L_HI(net1091));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][12]$_DFFE_PP__1092  (.L_HI(net1092));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][13]$_DFFE_PP__1093  (.L_HI(net1093));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][14]$_DFFE_PP__1094  (.L_HI(net1094));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][15]$_DFFE_PP__1095  (.L_HI(net1095));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][1]$_SDFFCE_PN1P__1096  (.L_HI(net1096));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][2]$_DFFE_PP__1097  (.L_HI(net1097));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][3]$_DFFE_PP__1098  (.L_HI(net1098));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][4]$_DFFE_PP__1099  (.L_HI(net1099));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][5]$_DFFE_PP__1100  (.L_HI(net1100));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][6]$_DFFE_PP__1101  (.L_HI(net1101));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][7]$_DFFE_PP__1102  (.L_HI(net1102));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][8]$_DFFE_PP__1103  (.L_HI(net1103));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][9]$_DFFE_PP__1104  (.L_HI(net1104));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][0]$_SDFFCE_PN1P__1105  (.L_HI(net1105));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][10]$_DFFE_PP__1106  (.L_HI(net1106));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][11]$_DFFE_PP__1107  (.L_HI(net1107));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][12]$_DFFE_PP__1108  (.L_HI(net1108));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][13]$_DFFE_PP__1109  (.L_HI(net1109));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][14]$_DFFE_PP__1110  (.L_HI(net1110));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][15]$_DFFE_PP__1111  (.L_HI(net1111));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][1]$_SDFFCE_PN1P__1112  (.L_HI(net1112));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][2]$_DFFE_PP__1113  (.L_HI(net1113));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][3]$_DFFE_PP__1114  (.L_HI(net1114));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][4]$_DFFE_PP__1115  (.L_HI(net1115));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][5]$_DFFE_PP__1116  (.L_HI(net1116));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][6]$_DFFE_PP__1117  (.L_HI(net1117));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][7]$_DFFE_PP__1118  (.L_HI(net1118));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][8]$_DFFE_PP__1119  (.L_HI(net1119));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][9]$_DFFE_PP__1120  (.L_HI(net1120));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][0]$_DFFE_PP__1121  (.L_HI(net1121));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][10]$_DFFE_PP__1122  (.L_HI(net1122));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][11]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][12]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][13]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][14]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][15]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][1]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][2]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][3]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][4]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][5]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][6]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][7]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][8]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][9]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[0]$_SDFFE_PN0P__1137  (.L_HI(net1137));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[10]$_SDFFE_PN0P__1138  (.L_HI(net1138));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[11]$_SDFFE_PN0P__1139  (.L_HI(net1139));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[12]$_SDFFE_PN0P__1140  (.L_HI(net1140));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[13]$_SDFFE_PN0P__1141  (.L_HI(net1141));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[14]$_SDFFE_PN0P__1142  (.L_HI(net1142));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[15]$_SDFFE_PN0P__1143  (.L_HI(net1143));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[16]$_SDFFE_PN0P__1144  (.L_HI(net1144));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[17]$_SDFFE_PN0P__1145  (.L_HI(net1145));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[18]$_SDFFE_PN0P__1146  (.L_HI(net1146));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[19]$_SDFFE_PN0P__1147  (.L_HI(net1147));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[1]$_SDFFE_PN0P__1148  (.L_HI(net1148));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[20]$_SDFFE_PN0P__1149  (.L_HI(net1149));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[2]$_SDFFE_PN0P__1150  (.L_HI(net1150));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[3]$_SDFFE_PN0P__1151  (.L_HI(net1151));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[4]$_SDFFE_PN0P__1152  (.L_HI(net1152));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[5]$_SDFFE_PN0P__1153  (.L_HI(net1153));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[6]$_SDFFE_PN0P__1154  (.L_HI(net1154));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[7]$_SDFFE_PN0P__1155  (.L_HI(net1155));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[8]$_SDFFE_PN0P__1156  (.L_HI(net1156));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[9]$_SDFFE_PN0P__1157  (.L_HI(net1157));
 sg13g2_tiehi \i_tinyqv.cpu.instr_fetch_running$_SDFFE_PN0P__1158  (.L_HI(net1158));
 sg13g2_tiehi \i_tinyqv.cpu.instr_len[0]$_SDFFE_PN0P__1159  (.L_HI(net1159));
 sg13g2_tiehi \i_tinyqv.cpu.instr_len[1]$_SDFFE_PN1P__1160  (.L_HI(net1160));
 sg13g2_tiehi \i_tinyqv.cpu.instr_valid$_SDFFE_PN0P__1161  (.L_HI(net1161));
 sg13g2_tiehi \i_tinyqv.cpu.instr_write_offset[0]$_SDFF_PN0__1162  (.L_HI(net1162));
 sg13g2_tiehi \i_tinyqv.cpu.instr_write_offset[1]$_SDFF_PN0__1163  (.L_HI(net1163));
 sg13g2_tiehi \i_tinyqv.cpu.instr_write_offset[2]$_SDFF_PP0__1164  (.L_HI(net1164));
 sg13g2_tiehi \i_tinyqv.cpu.interrupt_core$_SDFFE_PN0P__1165  (.L_HI(net1165));
 sg13g2_tiehi \i_tinyqv.cpu.is_alu_imm$_SDFFE_PN0P__1166  (.L_HI(net1166));
 sg13g2_tiehi \i_tinyqv.cpu.is_alu_reg$_SDFFE_PN0P__1167  (.L_HI(net1167));
 sg13g2_tiehi \i_tinyqv.cpu.is_auipc$_SDFFE_PN0P__1168  (.L_HI(net1168));
 sg13g2_tiehi \i_tinyqv.cpu.is_branch$_SDFFE_PN0P__1169  (.L_HI(net1169));
 sg13g2_tiehi \i_tinyqv.cpu.is_jal$_SDFFE_PN0P__1170  (.L_HI(net1170));
 sg13g2_tiehi \i_tinyqv.cpu.is_jalr$_SDFFE_PN0P__1171  (.L_HI(net1171));
 sg13g2_tiehi \i_tinyqv.cpu.is_load$_SDFFE_PN0P__1172  (.L_HI(net1172));
 sg13g2_tiehi \i_tinyqv.cpu.is_lui$_SDFFE_PN0P__1173  (.L_HI(net1173));
 sg13g2_tiehi \i_tinyqv.cpu.is_store$_SDFFE_PN0P__1174  (.L_HI(net1174));
 sg13g2_tiehi \i_tinyqv.cpu.is_system$_SDFFE_PN0P__1175  (.L_HI(net1175));
 sg13g2_tiehi \i_tinyqv.cpu.load_started$_SDFFE_PN0P__1176  (.L_HI(net1176));
 sg13g2_tiehi \i_tinyqv.cpu.mem_op[0]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \i_tinyqv.cpu.mem_op[1]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \i_tinyqv.cpu.mem_op[2]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \i_tinyqv.cpu.mem_op_increment_reg$_SDFFCE_PN1P__1180  (.L_HI(net1180));
 sg13g2_tiehi \i_tinyqv.cpu.no_write_in_progress$_SDFFE_PN1P__1181  (.L_HI(net1181));
 sg13g2_tiehi \i_tinyqv.cpu.pc_offset[0]$_SDFFE_PN0P__1182  (.L_HI(net1182));
 sg13g2_tiehi \i_tinyqv.cpu.pc_offset[1]$_SDFFE_PN0P__1183  (.L_HI(net1183));
 sg13g2_tiehi \i_tinyqv.cpu.rd[0]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \i_tinyqv.cpu.rd[1]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \i_tinyqv.cpu.rd[2]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \i_tinyqv.cpu.rd[3]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \i_tinyqv.cpu.rs1[0]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \i_tinyqv.cpu.rs1[1]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \i_tinyqv.cpu.rs1[2]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \i_tinyqv.cpu.rs1[3]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \i_tinyqv.cpu.rs2[0]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \i_tinyqv.cpu.rs2[1]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \i_tinyqv.cpu.rs2[2]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \i_tinyqv.cpu.rs2[3]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \i_tinyqv.cpu.was_early_branch$_SDFFE_PN0P__1196  (.L_HI(net1196));
 sg13g2_tiehi \i_tinyqv.mem.data_stall$_SDFFE_PN0P__1197  (.L_HI(net1197));
 sg13g2_tiehi \i_tinyqv.mem.instr_active$_SDFFE_PP0P__1198  (.L_HI(net1198));
 sg13g2_tiehi \i_tinyqv.mem.instr_fetch_started$_SDFF_PN0__1199  (.L_HI(net1199));
 sg13g2_tiehi \i_tinyqv.mem.instr_fetch_stopped$_SDFF_PN0__1200  (.L_HI(net1200));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[0]$_SDFFCE_PP0P__1201  (.L_HI(net1201));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[10]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[11]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[12]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[13]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[14]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[15]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[16]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[17]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[18]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[19]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[1]$_SDFFCE_PN0P__1212  (.L_HI(net1212));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[20]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[21]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[22]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[23]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[2]$_SDFFCE_PN0P__1217  (.L_HI(net1217));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[3]$_SDFFCE_PN0P__1218  (.L_HI(net1218));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[4]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[5]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[6]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[7]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[8]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[9]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[0]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[1]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[2]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[3]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[4]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[5]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[6]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[7]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data_ready$_SDFF_PN0__1233  (.L_HI(net1233));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data_req$_SDFF_PP0__1234  (.L_HI(net1234));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0]$_DFFE_PN__1235  (.L_HI(net1235));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1]$_DFFE_PN__1236  (.L_HI(net1236));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2]$_DFFE_PN__1237  (.L_HI(net1237));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.fsm_state[0]$_SDFFE_PP0P__1238  (.L_HI(net1238));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.fsm_state[1]$_SDFFE_PP0P__1239  (.L_HI(net1239));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.fsm_state[2]$_SDFFE_PP0P__1240  (.L_HI(net1240));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.is_writing$_SDFFE_PP0P__1241  (.L_HI(net1241));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.last_ram_a_sel$_SDFF_PN1__1242  (.L_HI(net1242));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.last_ram_b_sel$_SDFF_PN1__1243  (.L_HI(net1243));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.nibbles_remaining[0]$_SDFFE_PP0P__1244  (.L_HI(net1244));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.nibbles_remaining[1]$_SDFFE_PP0P__1245  (.L_HI(net1245));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.nibbles_remaining[2]$_SDFFE_PP0P__1246  (.L_HI(net1246));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.read_cycles_count[0]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.read_cycles_count[1]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.read_cycles_count[2]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_clk_out$_SDFFE_PP0P__1250  (.L_HI(net1250));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_data_oe[2]$_SDFFE_PP0P__1251  (.L_HI(net1251));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_flash_select$_SDFFE_PP1P__1252  (.L_HI(net1252));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[0]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[1]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[2]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[3]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[4]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[5]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[6]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[7]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_ram_a_select$_SDFFE_PP1P__1261  (.L_HI(net1261));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_ram_b_select$_SDFFE_PP1P__1262  (.L_HI(net1262));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.stop_txn_reg$_SDFF_PN0__1263  (.L_HI(net1263));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[0]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[10]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[11]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[12]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[13]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[14]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[15]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[16]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[17]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[18]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[19]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[1]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[20]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[21]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[22]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[23]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[24]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[25]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[26]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[27]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[28]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[29]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[2]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[30]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[31]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[3]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[4]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[5]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[6]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[7]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[8]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[9]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_byte_idx[0]$_SDFFE_PP0N__1296  (.L_HI(net1296));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_byte_idx[1]$_SDFFE_PP0N__1297  (.L_HI(net1297));
 sg13g2_tiehi \i_tinyqv.mem.qspi_write_done$_DFF_P__1298  (.L_HI(net1298));
 sg13g2_tiehi \i_tinyqv.rst_reg_n$_DFF_P__1299  (.L_HI(net1299));
 sg13g2_tiehi \i_uart_rx.bit_sample$_SDFFE_PN0N__1300  (.L_HI(net1300));
 sg13g2_tiehi \i_uart_rx.cycle_counter[0]$_SDFF_PP0__1301  (.L_HI(net1301));
 sg13g2_tiehi \i_uart_rx.cycle_counter[10]$_SDFF_PP0__1302  (.L_HI(net1302));
 sg13g2_tiehi \i_uart_rx.cycle_counter[1]$_SDFF_PP0__1303  (.L_HI(net1303));
 sg13g2_tiehi \i_uart_rx.cycle_counter[2]$_SDFF_PP0__1304  (.L_HI(net1304));
 sg13g2_tiehi \i_uart_rx.cycle_counter[3]$_SDFF_PP0__1305  (.L_HI(net1305));
 sg13g2_tiehi \i_uart_rx.cycle_counter[4]$_SDFF_PP0__1306  (.L_HI(net1306));
 sg13g2_tiehi \i_uart_rx.cycle_counter[5]$_SDFF_PP0__1307  (.L_HI(net1307));
 sg13g2_tiehi \i_uart_rx.cycle_counter[6]$_SDFF_PP0__1308  (.L_HI(net1308));
 sg13g2_tiehi \i_uart_rx.cycle_counter[7]$_SDFF_PP0__1309  (.L_HI(net1309));
 sg13g2_tiehi \i_uart_rx.cycle_counter[8]$_SDFF_PP0__1310  (.L_HI(net1310));
 sg13g2_tiehi \i_uart_rx.cycle_counter[9]$_SDFF_PP0__1311  (.L_HI(net1311));
 sg13g2_tiehi \i_uart_rx.fsm_state[0]$_SDFFE_PN0P__1312  (.L_HI(net1312));
 sg13g2_tiehi \i_uart_rx.fsm_state[1]$_SDFFE_PN0P__1313  (.L_HI(net1313));
 sg13g2_tiehi \i_uart_rx.fsm_state[2]$_SDFFE_PN0P__1314  (.L_HI(net1314));
 sg13g2_tiehi \i_uart_rx.fsm_state[3]$_SDFFE_PN0P__1315  (.L_HI(net1315));
 sg13g2_tiehi \i_uart_rx.recieved_data[0]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \i_uart_rx.recieved_data[1]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \i_uart_rx.recieved_data[2]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \i_uart_rx.recieved_data[3]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \i_uart_rx.recieved_data[4]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \i_uart_rx.recieved_data[5]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \i_uart_rx.recieved_data[6]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \i_uart_rx.recieved_data[7]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \i_uart_rx.rxd_reg[0]$_SDFF_PN1__1324  (.L_HI(net1324));
 sg13g2_tiehi \i_uart_rx.rxd_reg[1]$_SDFF_PN1__1325  (.L_HI(net1325));
 sg13g2_tiehi \i_uart_rx.uart_rts$_SDFF_PN1__1326  (.L_HI(net1326));
 sg13g2_tiehi \i_uart_tx.cycle_counter[0]$_SDFFE_PP0N__1327  (.L_HI(net1327));
 sg13g2_tiehi \i_uart_tx.cycle_counter[10]$_SDFFE_PP0N__1328  (.L_HI(net1328));
 sg13g2_tiehi \i_uart_tx.cycle_counter[1]$_SDFFE_PP0N__1329  (.L_HI(net1329));
 sg13g2_tiehi \i_uart_tx.cycle_counter[2]$_SDFFE_PP0N__1330  (.L_HI(net1330));
 sg13g2_tiehi \i_uart_tx.cycle_counter[3]$_SDFFE_PP0N__1331  (.L_HI(net1331));
 sg13g2_tiehi \i_uart_tx.cycle_counter[4]$_SDFFE_PP0N__1332  (.L_HI(net1332));
 sg13g2_tiehi \i_uart_tx.cycle_counter[5]$_SDFFE_PP0N__1333  (.L_HI(net1333));
 sg13g2_tiehi \i_uart_tx.cycle_counter[6]$_SDFFE_PP0N__1334  (.L_HI(net1334));
 sg13g2_tiehi \i_uart_tx.cycle_counter[7]$_SDFFE_PP0N__1335  (.L_HI(net1335));
 sg13g2_tiehi \i_uart_tx.cycle_counter[8]$_SDFFE_PP0N__1336  (.L_HI(net1336));
 sg13g2_tiehi \i_uart_tx.cycle_counter[9]$_SDFFE_PP0N__1337  (.L_HI(net1337));
 sg13g2_tiehi \i_uart_tx.data_to_send[0]$_SDFFE_PN0P__1338  (.L_HI(net1338));
 sg13g2_tiehi \i_uart_tx.data_to_send[1]$_SDFFE_PN0P__1339  (.L_HI(net1339));
 sg13g2_tiehi \i_uart_tx.data_to_send[2]$_SDFFE_PN0P__1340  (.L_HI(net1340));
 sg13g2_tiehi \i_uart_tx.data_to_send[3]$_SDFFE_PN0P__1341  (.L_HI(net1341));
 sg13g2_tiehi \i_uart_tx.data_to_send[4]$_SDFFE_PN0P__1342  (.L_HI(net1342));
 sg13g2_tiehi \i_uart_tx.data_to_send[5]$_SDFFE_PN0P__1343  (.L_HI(net1343));
 sg13g2_tiehi \i_uart_tx.data_to_send[6]$_SDFFE_PN0P__1344  (.L_HI(net1344));
 sg13g2_tiehi \i_uart_tx.data_to_send[7]$_SDFFE_PN0P__1345  (.L_HI(net1345));
 sg13g2_tiehi \i_uart_tx.fsm_state[0]$_SDFFE_PN0P__1346  (.L_HI(net1346));
 sg13g2_tiehi \i_uart_tx.fsm_state[1]$_SDFFE_PN0P__1347  (.L_HI(net1347));
 sg13g2_tiehi \i_uart_tx.fsm_state[2]$_SDFFE_PN0P__1348  (.L_HI(net1348));
 sg13g2_tiehi \i_uart_tx.fsm_state[3]$_SDFFE_PN0P__1349  (.L_HI(net1349));
 sg13g2_tiehi \i_uart_tx.txd_reg$_SDFF_PN1__1350  (.L_HI(net1350));
 sg13g2_tiehi \rst_reg_n$_DFF_N__1351  (.L_HI(net1351));
 sg13g2_tiehi \ui_in_reg[0]$_DFF_P__1352  (.L_HI(net1352));
 sg13g2_tiehi \ui_in_reg[1]$_DFF_P__1353  (.L_HI(net1353));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_62_clk (.X(clknet_leaf_62_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_63_clk (.X(clknet_leaf_63_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_64_clk (.X(clknet_leaf_64_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_65_clk (.X(clknet_leaf_65_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_66_clk (.X(clknet_leaf_66_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_67_clk (.X(clknet_leaf_67_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_68_clk (.X(clknet_leaf_68_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_69_clk (.X(clknet_leaf_69_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_70_clk (.X(clknet_leaf_70_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_71_clk (.X(clknet_leaf_71_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_72_clk (.X(clknet_leaf_72_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_73_clk (.X(clknet_leaf_73_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_74_clk (.X(clknet_leaf_74_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_75_clk (.X(clknet_leaf_75_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_76_clk (.X(clknet_leaf_76_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_77_clk (.X(clknet_leaf_77_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_78_clk (.X(clknet_leaf_78_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_79_clk (.X(clknet_leaf_79_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_80_clk (.X(clknet_leaf_80_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_81_clk (.X(clknet_leaf_81_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_82_clk (.X(clknet_leaf_82_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_83_clk (.X(clknet_leaf_83_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_84_clk (.X(clknet_leaf_84_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_85_clk (.X(clknet_leaf_85_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_86_clk (.X(clknet_leaf_86_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_87_clk (.X(clknet_leaf_87_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_88_clk (.X(clknet_leaf_88_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_89_clk (.X(clknet_leaf_89_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_90_clk (.X(clknet_leaf_90_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_91_clk (.X(clknet_leaf_91_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_92_clk (.X(clknet_leaf_92_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_93_clk (.X(clknet_leaf_93_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_94_clk (.X(clknet_leaf_94_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_95_clk (.X(clknet_leaf_95_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_96_clk (.X(clknet_leaf_96_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_97_clk (.X(clknet_leaf_97_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_98_clk (.X(clknet_leaf_98_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_99_clk (.X(clknet_leaf_99_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_100_clk (.X(clknet_leaf_100_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_101_clk (.X(clknet_leaf_101_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_102_clk (.X(clknet_leaf_102_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_103_clk (.X(clknet_leaf_103_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_104_clk (.X(clknet_leaf_104_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_105_clk (.X(clknet_leaf_105_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_106_clk (.X(clknet_leaf_106_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_107_clk (.X(clknet_leaf_107_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_108_clk (.X(clknet_leaf_108_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_109_clk (.X(clknet_leaf_109_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_110_clk (.X(clknet_leaf_110_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_111_clk (.X(clknet_leaf_111_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_112_clk (.X(clknet_leaf_112_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_113_clk (.X(clknet_leaf_113_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_114_clk (.X(clknet_leaf_114_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_115_clk (.X(clknet_leaf_115_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_116_clk (.X(clknet_leaf_116_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_117_clk (.X(clknet_leaf_117_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_119_clk (.X(clknet_leaf_119_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_120_clk (.X(clknet_leaf_120_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_121_clk (.X(clknet_leaf_121_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_122_clk (.X(clknet_leaf_122_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_123_clk (.X(clknet_leaf_123_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_124_clk (.X(clknet_leaf_124_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_125_clk (.X(clknet_leaf_125_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_126_clk (.X(clknet_leaf_126_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_127_clk (.X(clknet_leaf_127_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_128_clk (.X(clknet_leaf_128_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_129_clk (.X(clknet_leaf_129_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_130_clk (.X(clknet_leaf_130_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_131_clk (.X(clknet_leaf_131_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_132_clk (.X(clknet_leaf_132_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_133_clk (.X(clknet_leaf_133_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_134_clk (.X(clknet_leaf_134_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_135_clk (.X(clknet_leaf_135_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_136_clk (.X(clknet_leaf_136_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_137_clk (.X(clknet_leaf_137_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkload6 (.A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkload8 (.A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkload9 (.A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkload10 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_137_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_39_clk));
 sg13g2_buf_16 clkload14 (.A(clknet_leaf_22_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_51_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_114_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_88_clk));
 sg13g2_buf_16 clkload18 (.A(clknet_leaf_91_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_93_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_leaf_94_clk));
 sg13g2_buf_8 clkload21 (.A(clknet_leaf_95_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_54_clk));
 sg13g2_buf_8 clkload23 (.A(clknet_leaf_57_clk));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_56_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_82_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_84_clk));
 sg13g2_buf_16 clkload27 (.A(clknet_leaf_50_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_75_clk));
 sg13g2_buf_16 clkload29 (.A(clknet_leaf_81_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_86_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00035_));
 sg13g2_antennanp ANTENNA_2 (.A(_00035_));
 sg13g2_antennanp ANTENNA_3 (.A(_00641_));
 sg13g2_antennanp ANTENNA_4 (.A(_03685_));
 sg13g2_antennanp ANTENNA_5 (.A(_04121_));
 sg13g2_antennanp ANTENNA_6 (.A(_04452_));
 sg13g2_antennanp ANTENNA_7 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_antennanp ANTENNA_8 (.A(net18));
 sg13g2_antennanp ANTENNA_9 (.A(net22));
 sg13g2_antennanp ANTENNA_10 (.A(_00035_));
 sg13g2_antennanp ANTENNA_11 (.A(_00035_));
 sg13g2_antennanp ANTENNA_12 (.A(_00037_));
 sg13g2_antennanp ANTENNA_13 (.A(_00043_));
 sg13g2_antennanp ANTENNA_14 (.A(_00045_));
 sg13g2_antennanp ANTENNA_15 (.A(_00045_));
 sg13g2_antennanp ANTENNA_16 (.A(_00053_));
 sg13g2_antennanp ANTENNA_17 (.A(_00641_));
 sg13g2_antennanp ANTENNA_18 (.A(_03685_));
 sg13g2_antennanp ANTENNA_19 (.A(_04121_));
 sg13g2_antennanp ANTENNA_20 (.A(_04452_));
 sg13g2_antennanp ANTENNA_21 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_antennanp ANTENNA_22 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_antennanp ANTENNA_23 (.A(net18));
 sg13g2_antennanp ANTENNA_24 (.A(net22));
 sg13g2_antennanp ANTENNA_25 (.A(net23));
 sg13g2_antennanp ANTENNA_26 (.A(_00035_));
 sg13g2_antennanp ANTENNA_27 (.A(_00035_));
 sg13g2_antennanp ANTENNA_28 (.A(_00037_));
 sg13g2_antennanp ANTENNA_29 (.A(_00039_));
 sg13g2_antennanp ANTENNA_30 (.A(_00043_));
 sg13g2_antennanp ANTENNA_31 (.A(_00053_));
 sg13g2_antennanp ANTENNA_32 (.A(_00061_));
 sg13g2_antennanp ANTENNA_33 (.A(_00641_));
 sg13g2_antennanp ANTENNA_34 (.A(_04121_));
 sg13g2_antennanp ANTENNA_35 (.A(_04452_));
 sg13g2_antennanp ANTENNA_36 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_antennanp ANTENNA_37 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_antennanp ANTENNA_38 (.A(net18));
 sg13g2_antennanp ANTENNA_39 (.A(net22));
 sg13g2_antennanp ANTENNA_40 (.A(net23));
 sg13g2_antennanp ANTENNA_41 (.A(_00035_));
 sg13g2_antennanp ANTENNA_42 (.A(_00035_));
 sg13g2_antennanp ANTENNA_43 (.A(_00037_));
 sg13g2_antennanp ANTENNA_44 (.A(_00641_));
 sg13g2_antennanp ANTENNA_45 (.A(_04121_));
 sg13g2_antennanp ANTENNA_46 (.A(_04452_));
 sg13g2_antennanp ANTENNA_47 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_antennanp ANTENNA_48 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_antennanp ANTENNA_49 (.A(net18));
 sg13g2_antennanp ANTENNA_50 (.A(net22));
 sg13g2_antennanp ANTENNA_51 (.A(net23));
 sg13g2_antennanp ANTENNA_52 (.A(_00035_));
 sg13g2_antennanp ANTENNA_53 (.A(_00035_));
 sg13g2_antennanp ANTENNA_54 (.A(_00641_));
 sg13g2_antennanp ANTENNA_55 (.A(_04121_));
 sg13g2_antennanp ANTENNA_56 (.A(_04452_));
 sg13g2_antennanp ANTENNA_57 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_antennanp ANTENNA_58 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_antennanp ANTENNA_59 (.A(net18));
 sg13g2_antennanp ANTENNA_60 (.A(net22));
 sg13g2_antennanp ANTENNA_61 (.A(net23));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_4 FILLER_0_140 ();
 sg13g2_fill_2 FILLER_0_210 ();
 sg13g2_fill_1 FILLER_0_212 ();
 sg13g2_fill_2 FILLER_0_311 ();
 sg13g2_decap_4 FILLER_0_469 ();
 sg13g2_fill_1 FILLER_0_503 ();
 sg13g2_fill_2 FILLER_0_530 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_fill_2 FILLER_0_875 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_4 FILLER_1_126 ();
 sg13g2_fill_1 FILLER_1_130 ();
 sg13g2_fill_2 FILLER_1_135 ();
 sg13g2_fill_1 FILLER_1_153 ();
 sg13g2_fill_2 FILLER_1_158 ();
 sg13g2_fill_1 FILLER_1_224 ();
 sg13g2_fill_1 FILLER_1_433 ();
 sg13g2_fill_1 FILLER_1_438 ();
 sg13g2_fill_2 FILLER_1_443 ();
 sg13g2_fill_2 FILLER_1_579 ();
 sg13g2_decap_8 FILLER_1_633 ();
 sg13g2_decap_8 FILLER_1_640 ();
 sg13g2_decap_8 FILLER_1_647 ();
 sg13g2_decap_8 FILLER_1_654 ();
 sg13g2_decap_8 FILLER_1_661 ();
 sg13g2_decap_8 FILLER_1_668 ();
 sg13g2_decap_8 FILLER_1_675 ();
 sg13g2_decap_8 FILLER_1_682 ();
 sg13g2_decap_8 FILLER_1_689 ();
 sg13g2_decap_8 FILLER_1_696 ();
 sg13g2_decap_8 FILLER_1_703 ();
 sg13g2_decap_8 FILLER_1_710 ();
 sg13g2_decap_8 FILLER_1_717 ();
 sg13g2_decap_8 FILLER_1_724 ();
 sg13g2_decap_8 FILLER_1_731 ();
 sg13g2_decap_8 FILLER_1_738 ();
 sg13g2_decap_8 FILLER_1_745 ();
 sg13g2_decap_8 FILLER_1_752 ();
 sg13g2_decap_8 FILLER_1_759 ();
 sg13g2_decap_8 FILLER_1_766 ();
 sg13g2_decap_8 FILLER_1_773 ();
 sg13g2_decap_8 FILLER_1_780 ();
 sg13g2_decap_8 FILLER_1_787 ();
 sg13g2_decap_8 FILLER_1_794 ();
 sg13g2_decap_8 FILLER_1_801 ();
 sg13g2_decap_8 FILLER_1_808 ();
 sg13g2_decap_8 FILLER_1_815 ();
 sg13g2_decap_8 FILLER_1_822 ();
 sg13g2_decap_8 FILLER_1_829 ();
 sg13g2_decap_8 FILLER_1_836 ();
 sg13g2_decap_8 FILLER_1_843 ();
 sg13g2_decap_8 FILLER_1_850 ();
 sg13g2_decap_8 FILLER_1_857 ();
 sg13g2_decap_8 FILLER_1_864 ();
 sg13g2_decap_8 FILLER_1_871 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_4 FILLER_2_119 ();
 sg13g2_fill_1 FILLER_2_123 ();
 sg13g2_fill_2 FILLER_2_184 ();
 sg13g2_fill_2 FILLER_2_294 ();
 sg13g2_fill_1 FILLER_2_296 ();
 sg13g2_fill_2 FILLER_2_335 ();
 sg13g2_fill_2 FILLER_2_363 ();
 sg13g2_fill_1 FILLER_2_365 ();
 sg13g2_fill_1 FILLER_2_392 ();
 sg13g2_fill_2 FILLER_2_397 ();
 sg13g2_fill_2 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_427 ();
 sg13g2_fill_2 FILLER_2_454 ();
 sg13g2_fill_1 FILLER_2_456 ();
 sg13g2_fill_2 FILLER_2_461 ();
 sg13g2_fill_1 FILLER_2_463 ();
 sg13g2_fill_1 FILLER_2_490 ();
 sg13g2_fill_1 FILLER_2_517 ();
 sg13g2_fill_2 FILLER_2_552 ();
 sg13g2_decap_8 FILLER_2_638 ();
 sg13g2_decap_8 FILLER_2_645 ();
 sg13g2_decap_8 FILLER_2_652 ();
 sg13g2_decap_8 FILLER_2_659 ();
 sg13g2_decap_8 FILLER_2_666 ();
 sg13g2_decap_8 FILLER_2_673 ();
 sg13g2_decap_8 FILLER_2_680 ();
 sg13g2_decap_8 FILLER_2_687 ();
 sg13g2_decap_8 FILLER_2_694 ();
 sg13g2_decap_8 FILLER_2_701 ();
 sg13g2_decap_8 FILLER_2_708 ();
 sg13g2_decap_8 FILLER_2_715 ();
 sg13g2_decap_8 FILLER_2_722 ();
 sg13g2_decap_8 FILLER_2_729 ();
 sg13g2_decap_8 FILLER_2_736 ();
 sg13g2_decap_8 FILLER_2_743 ();
 sg13g2_decap_8 FILLER_2_750 ();
 sg13g2_decap_8 FILLER_2_757 ();
 sg13g2_decap_8 FILLER_2_764 ();
 sg13g2_decap_8 FILLER_2_771 ();
 sg13g2_decap_8 FILLER_2_778 ();
 sg13g2_decap_8 FILLER_2_785 ();
 sg13g2_decap_8 FILLER_2_792 ();
 sg13g2_decap_8 FILLER_2_799 ();
 sg13g2_decap_8 FILLER_2_806 ();
 sg13g2_decap_8 FILLER_2_813 ();
 sg13g2_decap_8 FILLER_2_820 ();
 sg13g2_decap_8 FILLER_2_827 ();
 sg13g2_decap_8 FILLER_2_834 ();
 sg13g2_decap_8 FILLER_2_841 ();
 sg13g2_decap_8 FILLER_2_848 ();
 sg13g2_decap_8 FILLER_2_855 ();
 sg13g2_decap_8 FILLER_2_862 ();
 sg13g2_decap_8 FILLER_2_869 ();
 sg13g2_fill_2 FILLER_2_876 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_fill_2 FILLER_3_105 ();
 sg13g2_fill_1 FILLER_3_111 ();
 sg13g2_fill_2 FILLER_3_154 ();
 sg13g2_fill_1 FILLER_3_156 ();
 sg13g2_fill_2 FILLER_3_307 ();
 sg13g2_decap_8 FILLER_3_633 ();
 sg13g2_decap_8 FILLER_3_640 ();
 sg13g2_decap_8 FILLER_3_647 ();
 sg13g2_decap_8 FILLER_3_654 ();
 sg13g2_decap_8 FILLER_3_661 ();
 sg13g2_decap_8 FILLER_3_668 ();
 sg13g2_decap_8 FILLER_3_675 ();
 sg13g2_decap_8 FILLER_3_682 ();
 sg13g2_decap_8 FILLER_3_689 ();
 sg13g2_decap_8 FILLER_3_696 ();
 sg13g2_decap_8 FILLER_3_703 ();
 sg13g2_decap_8 FILLER_3_710 ();
 sg13g2_decap_8 FILLER_3_717 ();
 sg13g2_decap_8 FILLER_3_724 ();
 sg13g2_decap_8 FILLER_3_731 ();
 sg13g2_decap_8 FILLER_3_738 ();
 sg13g2_decap_8 FILLER_3_745 ();
 sg13g2_decap_8 FILLER_3_752 ();
 sg13g2_decap_8 FILLER_3_759 ();
 sg13g2_decap_8 FILLER_3_766 ();
 sg13g2_decap_8 FILLER_3_773 ();
 sg13g2_decap_8 FILLER_3_780 ();
 sg13g2_decap_8 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_794 ();
 sg13g2_decap_8 FILLER_3_801 ();
 sg13g2_decap_8 FILLER_3_808 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_decap_8 FILLER_3_829 ();
 sg13g2_decap_8 FILLER_3_836 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_850 ();
 sg13g2_decap_8 FILLER_3_857 ();
 sg13g2_decap_8 FILLER_3_864 ();
 sg13g2_decap_8 FILLER_3_871 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_fill_2 FILLER_4_92 ();
 sg13g2_fill_1 FILLER_4_94 ();
 sg13g2_fill_2 FILLER_4_103 ();
 sg13g2_fill_2 FILLER_4_147 ();
 sg13g2_fill_1 FILLER_4_149 ();
 sg13g2_fill_1 FILLER_4_176 ();
 sg13g2_fill_2 FILLER_4_231 ();
 sg13g2_fill_2 FILLER_4_327 ();
 sg13g2_fill_1 FILLER_4_329 ();
 sg13g2_fill_1 FILLER_4_486 ();
 sg13g2_fill_2 FILLER_4_491 ();
 sg13g2_fill_1 FILLER_4_493 ();
 sg13g2_fill_2 FILLER_4_502 ();
 sg13g2_fill_1 FILLER_4_504 ();
 sg13g2_fill_1 FILLER_4_517 ();
 sg13g2_fill_2 FILLER_4_526 ();
 sg13g2_fill_2 FILLER_4_566 ();
 sg13g2_fill_1 FILLER_4_568 ();
 sg13g2_decap_8 FILLER_4_647 ();
 sg13g2_decap_8 FILLER_4_654 ();
 sg13g2_decap_8 FILLER_4_661 ();
 sg13g2_decap_8 FILLER_4_668 ();
 sg13g2_decap_8 FILLER_4_675 ();
 sg13g2_decap_8 FILLER_4_682 ();
 sg13g2_decap_8 FILLER_4_689 ();
 sg13g2_decap_8 FILLER_4_696 ();
 sg13g2_decap_8 FILLER_4_703 ();
 sg13g2_decap_8 FILLER_4_710 ();
 sg13g2_decap_8 FILLER_4_717 ();
 sg13g2_decap_8 FILLER_4_724 ();
 sg13g2_decap_8 FILLER_4_731 ();
 sg13g2_decap_8 FILLER_4_738 ();
 sg13g2_decap_8 FILLER_4_745 ();
 sg13g2_decap_8 FILLER_4_752 ();
 sg13g2_decap_8 FILLER_4_759 ();
 sg13g2_decap_8 FILLER_4_766 ();
 sg13g2_decap_8 FILLER_4_773 ();
 sg13g2_decap_8 FILLER_4_780 ();
 sg13g2_decap_8 FILLER_4_787 ();
 sg13g2_decap_8 FILLER_4_794 ();
 sg13g2_decap_8 FILLER_4_801 ();
 sg13g2_decap_8 FILLER_4_808 ();
 sg13g2_decap_8 FILLER_4_815 ();
 sg13g2_decap_8 FILLER_4_822 ();
 sg13g2_decap_8 FILLER_4_829 ();
 sg13g2_decap_8 FILLER_4_836 ();
 sg13g2_decap_8 FILLER_4_843 ();
 sg13g2_decap_8 FILLER_4_850 ();
 sg13g2_decap_8 FILLER_4_857 ();
 sg13g2_decap_8 FILLER_4_864 ();
 sg13g2_decap_8 FILLER_4_871 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_4 FILLER_5_77 ();
 sg13g2_fill_1 FILLER_5_185 ();
 sg13g2_fill_1 FILLER_5_243 ();
 sg13g2_fill_2 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_271 ();
 sg13g2_fill_1 FILLER_5_287 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_fill_1 FILLER_5_316 ();
 sg13g2_fill_1 FILLER_5_377 ();
 sg13g2_fill_1 FILLER_5_382 ();
 sg13g2_fill_1 FILLER_5_387 ();
 sg13g2_fill_1 FILLER_5_459 ();
 sg13g2_fill_2 FILLER_5_550 ();
 sg13g2_fill_1 FILLER_5_552 ();
 sg13g2_decap_8 FILLER_5_649 ();
 sg13g2_decap_8 FILLER_5_656 ();
 sg13g2_decap_8 FILLER_5_663 ();
 sg13g2_decap_8 FILLER_5_670 ();
 sg13g2_decap_8 FILLER_5_677 ();
 sg13g2_decap_8 FILLER_5_684 ();
 sg13g2_decap_8 FILLER_5_691 ();
 sg13g2_decap_8 FILLER_5_698 ();
 sg13g2_decap_8 FILLER_5_705 ();
 sg13g2_decap_8 FILLER_5_712 ();
 sg13g2_decap_8 FILLER_5_719 ();
 sg13g2_decap_8 FILLER_5_726 ();
 sg13g2_decap_8 FILLER_5_733 ();
 sg13g2_decap_8 FILLER_5_740 ();
 sg13g2_decap_8 FILLER_5_747 ();
 sg13g2_decap_8 FILLER_5_754 ();
 sg13g2_decap_8 FILLER_5_761 ();
 sg13g2_decap_8 FILLER_5_768 ();
 sg13g2_decap_8 FILLER_5_775 ();
 sg13g2_decap_8 FILLER_5_782 ();
 sg13g2_decap_8 FILLER_5_789 ();
 sg13g2_decap_8 FILLER_5_796 ();
 sg13g2_decap_8 FILLER_5_803 ();
 sg13g2_decap_8 FILLER_5_810 ();
 sg13g2_decap_8 FILLER_5_817 ();
 sg13g2_decap_8 FILLER_5_824 ();
 sg13g2_decap_8 FILLER_5_831 ();
 sg13g2_decap_8 FILLER_5_838 ();
 sg13g2_decap_8 FILLER_5_845 ();
 sg13g2_decap_8 FILLER_5_852 ();
 sg13g2_decap_8 FILLER_5_859 ();
 sg13g2_decap_8 FILLER_5_866 ();
 sg13g2_decap_4 FILLER_5_873 ();
 sg13g2_fill_1 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_4 FILLER_6_56 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_fill_2 FILLER_6_287 ();
 sg13g2_fill_1 FILLER_6_353 ();
 sg13g2_fill_1 FILLER_6_380 ();
 sg13g2_fill_1 FILLER_6_385 ();
 sg13g2_fill_2 FILLER_6_412 ();
 sg13g2_decap_8 FILLER_6_638 ();
 sg13g2_decap_8 FILLER_6_645 ();
 sg13g2_decap_8 FILLER_6_652 ();
 sg13g2_decap_8 FILLER_6_659 ();
 sg13g2_decap_8 FILLER_6_666 ();
 sg13g2_decap_8 FILLER_6_673 ();
 sg13g2_decap_8 FILLER_6_680 ();
 sg13g2_decap_8 FILLER_6_687 ();
 sg13g2_decap_8 FILLER_6_694 ();
 sg13g2_decap_8 FILLER_6_701 ();
 sg13g2_decap_8 FILLER_6_708 ();
 sg13g2_decap_8 FILLER_6_715 ();
 sg13g2_decap_8 FILLER_6_722 ();
 sg13g2_decap_8 FILLER_6_729 ();
 sg13g2_decap_8 FILLER_6_736 ();
 sg13g2_decap_8 FILLER_6_743 ();
 sg13g2_decap_8 FILLER_6_750 ();
 sg13g2_decap_8 FILLER_6_757 ();
 sg13g2_decap_8 FILLER_6_764 ();
 sg13g2_decap_8 FILLER_6_771 ();
 sg13g2_decap_8 FILLER_6_778 ();
 sg13g2_decap_8 FILLER_6_785 ();
 sg13g2_decap_8 FILLER_6_792 ();
 sg13g2_decap_8 FILLER_6_799 ();
 sg13g2_decap_8 FILLER_6_806 ();
 sg13g2_decap_8 FILLER_6_813 ();
 sg13g2_decap_8 FILLER_6_820 ();
 sg13g2_decap_8 FILLER_6_827 ();
 sg13g2_decap_8 FILLER_6_834 ();
 sg13g2_decap_8 FILLER_6_841 ();
 sg13g2_decap_8 FILLER_6_848 ();
 sg13g2_decap_8 FILLER_6_855 ();
 sg13g2_decap_8 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_869 ();
 sg13g2_fill_2 FILLER_6_876 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_4 FILLER_7_28 ();
 sg13g2_decap_4 FILLER_7_36 ();
 sg13g2_fill_2 FILLER_7_40 ();
 sg13g2_fill_2 FILLER_7_68 ();
 sg13g2_fill_2 FILLER_7_184 ();
 sg13g2_fill_1 FILLER_7_230 ();
 sg13g2_fill_1 FILLER_7_241 ();
 sg13g2_fill_1 FILLER_7_296 ();
 sg13g2_fill_2 FILLER_7_302 ();
 sg13g2_fill_1 FILLER_7_360 ();
 sg13g2_fill_2 FILLER_7_425 ();
 sg13g2_fill_1 FILLER_7_503 ();
 sg13g2_fill_2 FILLER_7_520 ();
 sg13g2_fill_2 FILLER_7_552 ();
 sg13g2_fill_2 FILLER_7_622 ();
 sg13g2_fill_1 FILLER_7_624 ();
 sg13g2_decap_8 FILLER_7_649 ();
 sg13g2_decap_8 FILLER_7_656 ();
 sg13g2_decap_8 FILLER_7_663 ();
 sg13g2_decap_8 FILLER_7_670 ();
 sg13g2_decap_8 FILLER_7_677 ();
 sg13g2_decap_8 FILLER_7_684 ();
 sg13g2_decap_8 FILLER_7_691 ();
 sg13g2_decap_8 FILLER_7_698 ();
 sg13g2_decap_8 FILLER_7_705 ();
 sg13g2_decap_8 FILLER_7_712 ();
 sg13g2_decap_8 FILLER_7_719 ();
 sg13g2_decap_8 FILLER_7_726 ();
 sg13g2_decap_8 FILLER_7_733 ();
 sg13g2_decap_8 FILLER_7_740 ();
 sg13g2_decap_8 FILLER_7_747 ();
 sg13g2_decap_8 FILLER_7_754 ();
 sg13g2_decap_8 FILLER_7_761 ();
 sg13g2_decap_8 FILLER_7_768 ();
 sg13g2_decap_8 FILLER_7_775 ();
 sg13g2_decap_8 FILLER_7_782 ();
 sg13g2_decap_8 FILLER_7_789 ();
 sg13g2_decap_8 FILLER_7_796 ();
 sg13g2_decap_8 FILLER_7_803 ();
 sg13g2_decap_8 FILLER_7_810 ();
 sg13g2_decap_8 FILLER_7_817 ();
 sg13g2_decap_8 FILLER_7_824 ();
 sg13g2_decap_8 FILLER_7_831 ();
 sg13g2_decap_8 FILLER_7_838 ();
 sg13g2_decap_8 FILLER_7_845 ();
 sg13g2_decap_8 FILLER_7_852 ();
 sg13g2_decap_8 FILLER_7_859 ();
 sg13g2_decap_8 FILLER_7_866 ();
 sg13g2_decap_4 FILLER_7_873 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_23 ();
 sg13g2_fill_2 FILLER_8_90 ();
 sg13g2_fill_2 FILLER_8_164 ();
 sg13g2_fill_2 FILLER_8_343 ();
 sg13g2_fill_2 FILLER_8_349 ();
 sg13g2_fill_1 FILLER_8_377 ();
 sg13g2_fill_2 FILLER_8_404 ();
 sg13g2_fill_2 FILLER_8_604 ();
 sg13g2_fill_1 FILLER_8_606 ();
 sg13g2_decap_8 FILLER_8_659 ();
 sg13g2_decap_8 FILLER_8_666 ();
 sg13g2_decap_8 FILLER_8_673 ();
 sg13g2_decap_8 FILLER_8_680 ();
 sg13g2_decap_8 FILLER_8_687 ();
 sg13g2_decap_8 FILLER_8_694 ();
 sg13g2_decap_8 FILLER_8_701 ();
 sg13g2_decap_8 FILLER_8_708 ();
 sg13g2_decap_8 FILLER_8_715 ();
 sg13g2_decap_8 FILLER_8_722 ();
 sg13g2_decap_8 FILLER_8_729 ();
 sg13g2_decap_8 FILLER_8_736 ();
 sg13g2_decap_8 FILLER_8_743 ();
 sg13g2_decap_8 FILLER_8_750 ();
 sg13g2_decap_8 FILLER_8_757 ();
 sg13g2_decap_8 FILLER_8_764 ();
 sg13g2_decap_8 FILLER_8_771 ();
 sg13g2_decap_8 FILLER_8_778 ();
 sg13g2_decap_8 FILLER_8_785 ();
 sg13g2_decap_8 FILLER_8_792 ();
 sg13g2_decap_8 FILLER_8_799 ();
 sg13g2_decap_8 FILLER_8_806 ();
 sg13g2_decap_8 FILLER_8_813 ();
 sg13g2_decap_8 FILLER_8_820 ();
 sg13g2_decap_8 FILLER_8_827 ();
 sg13g2_decap_8 FILLER_8_834 ();
 sg13g2_decap_8 FILLER_8_841 ();
 sg13g2_decap_8 FILLER_8_848 ();
 sg13g2_decap_8 FILLER_8_855 ();
 sg13g2_decap_8 FILLER_8_862 ();
 sg13g2_decap_8 FILLER_8_869 ();
 sg13g2_fill_2 FILLER_8_876 ();
 sg13g2_fill_2 FILLER_9_30 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_fill_1 FILLER_9_97 ();
 sg13g2_fill_1 FILLER_9_124 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_fill_1 FILLER_9_204 ();
 sg13g2_fill_1 FILLER_9_215 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_fill_1 FILLER_9_353 ();
 sg13g2_fill_1 FILLER_9_384 ();
 sg13g2_fill_2 FILLER_9_389 ();
 sg13g2_fill_1 FILLER_9_417 ();
 sg13g2_fill_2 FILLER_9_444 ();
 sg13g2_fill_1 FILLER_9_588 ();
 sg13g2_fill_2 FILLER_9_619 ();
 sg13g2_fill_2 FILLER_9_647 ();
 sg13g2_decap_8 FILLER_9_675 ();
 sg13g2_decap_8 FILLER_9_682 ();
 sg13g2_decap_8 FILLER_9_689 ();
 sg13g2_decap_8 FILLER_9_696 ();
 sg13g2_decap_8 FILLER_9_703 ();
 sg13g2_decap_8 FILLER_9_718 ();
 sg13g2_decap_8 FILLER_9_733 ();
 sg13g2_decap_8 FILLER_9_740 ();
 sg13g2_decap_8 FILLER_9_747 ();
 sg13g2_decap_8 FILLER_9_754 ();
 sg13g2_decap_8 FILLER_9_761 ();
 sg13g2_decap_8 FILLER_9_768 ();
 sg13g2_decap_8 FILLER_9_775 ();
 sg13g2_decap_8 FILLER_9_782 ();
 sg13g2_decap_8 FILLER_9_789 ();
 sg13g2_decap_8 FILLER_9_796 ();
 sg13g2_decap_8 FILLER_9_803 ();
 sg13g2_decap_8 FILLER_9_810 ();
 sg13g2_decap_8 FILLER_9_817 ();
 sg13g2_decap_8 FILLER_9_824 ();
 sg13g2_decap_8 FILLER_9_831 ();
 sg13g2_decap_8 FILLER_9_838 ();
 sg13g2_decap_8 FILLER_9_845 ();
 sg13g2_decap_8 FILLER_9_852 ();
 sg13g2_decap_8 FILLER_9_859 ();
 sg13g2_decap_8 FILLER_9_866 ();
 sg13g2_decap_4 FILLER_9_873 ();
 sg13g2_fill_1 FILLER_9_877 ();
 sg13g2_fill_2 FILLER_10_34 ();
 sg13g2_fill_1 FILLER_10_36 ();
 sg13g2_fill_2 FILLER_10_45 ();
 sg13g2_fill_1 FILLER_10_99 ();
 sg13g2_fill_2 FILLER_10_108 ();
 sg13g2_fill_2 FILLER_10_188 ();
 sg13g2_fill_1 FILLER_10_190 ();
 sg13g2_fill_2 FILLER_10_261 ();
 sg13g2_fill_1 FILLER_10_263 ();
 sg13g2_fill_1 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_decap_4 FILLER_10_426 ();
 sg13g2_fill_2 FILLER_10_434 ();
 sg13g2_fill_1 FILLER_10_446 ();
 sg13g2_fill_1 FILLER_10_451 ();
 sg13g2_fill_1 FILLER_10_456 ();
 sg13g2_fill_1 FILLER_10_483 ();
 sg13g2_fill_2 FILLER_10_488 ();
 sg13g2_fill_1 FILLER_10_494 ();
 sg13g2_fill_2 FILLER_10_525 ();
 sg13g2_fill_1 FILLER_10_639 ();
 sg13g2_decap_8 FILLER_10_670 ();
 sg13g2_decap_4 FILLER_10_677 ();
 sg13g2_fill_1 FILLER_10_685 ();
 sg13g2_decap_8 FILLER_10_694 ();
 sg13g2_decap_8 FILLER_10_701 ();
 sg13g2_fill_2 FILLER_10_708 ();
 sg13g2_fill_2 FILLER_10_715 ();
 sg13g2_fill_1 FILLER_10_717 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_4 FILLER_10_770 ();
 sg13g2_fill_1 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_decap_8 FILLER_10_786 ();
 sg13g2_decap_8 FILLER_10_793 ();
 sg13g2_decap_8 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_10_835 ();
 sg13g2_decap_8 FILLER_10_842 ();
 sg13g2_decap_8 FILLER_10_849 ();
 sg13g2_decap_8 FILLER_10_856 ();
 sg13g2_decap_8 FILLER_10_863 ();
 sg13g2_decap_8 FILLER_10_870 ();
 sg13g2_fill_1 FILLER_10_877 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_9 ();
 sg13g2_fill_2 FILLER_11_74 ();
 sg13g2_fill_1 FILLER_11_76 ();
 sg13g2_fill_2 FILLER_11_150 ();
 sg13g2_fill_2 FILLER_11_160 ();
 sg13g2_fill_1 FILLER_11_234 ();
 sg13g2_fill_1 FILLER_11_295 ();
 sg13g2_fill_2 FILLER_11_390 ();
 sg13g2_fill_1 FILLER_11_418 ();
 sg13g2_fill_2 FILLER_11_531 ();
 sg13g2_fill_2 FILLER_11_563 ();
 sg13g2_fill_2 FILLER_11_651 ();
 sg13g2_decap_4 FILLER_11_662 ();
 sg13g2_fill_2 FILLER_11_666 ();
 sg13g2_fill_1 FILLER_11_685 ();
 sg13g2_fill_1 FILLER_11_709 ();
 sg13g2_fill_1 FILLER_11_720 ();
 sg13g2_fill_1 FILLER_11_751 ();
 sg13g2_fill_2 FILLER_11_757 ();
 sg13g2_fill_1 FILLER_11_759 ();
 sg13g2_decap_8 FILLER_11_794 ();
 sg13g2_decap_8 FILLER_11_801 ();
 sg13g2_decap_8 FILLER_11_808 ();
 sg13g2_decap_8 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_822 ();
 sg13g2_decap_8 FILLER_11_829 ();
 sg13g2_decap_8 FILLER_11_836 ();
 sg13g2_decap_8 FILLER_11_843 ();
 sg13g2_decap_8 FILLER_11_850 ();
 sg13g2_decap_8 FILLER_11_857 ();
 sg13g2_decap_8 FILLER_11_864 ();
 sg13g2_decap_8 FILLER_11_871 ();
 sg13g2_fill_2 FILLER_12_32 ();
 sg13g2_fill_2 FILLER_12_121 ();
 sg13g2_fill_1 FILLER_12_123 ();
 sg13g2_fill_1 FILLER_12_210 ();
 sg13g2_fill_2 FILLER_12_275 ();
 sg13g2_fill_1 FILLER_12_311 ();
 sg13g2_fill_2 FILLER_12_325 ();
 sg13g2_fill_1 FILLER_12_327 ();
 sg13g2_decap_4 FILLER_12_436 ();
 sg13g2_fill_1 FILLER_12_440 ();
 sg13g2_decap_4 FILLER_12_445 ();
 sg13g2_fill_2 FILLER_12_449 ();
 sg13g2_fill_1 FILLER_12_459 ();
 sg13g2_fill_2 FILLER_12_464 ();
 sg13g2_fill_1 FILLER_12_504 ();
 sg13g2_fill_2 FILLER_12_656 ();
 sg13g2_fill_2 FILLER_12_671 ();
 sg13g2_fill_1 FILLER_12_698 ();
 sg13g2_fill_1 FILLER_12_707 ();
 sg13g2_fill_2 FILLER_12_737 ();
 sg13g2_fill_1 FILLER_12_739 ();
 sg13g2_fill_2 FILLER_12_752 ();
 sg13g2_decap_8 FILLER_12_800 ();
 sg13g2_decap_8 FILLER_12_811 ();
 sg13g2_decap_8 FILLER_12_818 ();
 sg13g2_fill_2 FILLER_12_825 ();
 sg13g2_fill_1 FILLER_12_827 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_decap_8 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_12_868 ();
 sg13g2_fill_2 FILLER_12_875 ();
 sg13g2_fill_1 FILLER_12_877 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_1 FILLER_13_113 ();
 sg13g2_fill_1 FILLER_13_140 ();
 sg13g2_fill_2 FILLER_13_193 ();
 sg13g2_fill_2 FILLER_13_225 ();
 sg13g2_fill_1 FILLER_13_241 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_fill_2 FILLER_13_379 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_fill_2 FILLER_13_413 ();
 sg13g2_fill_1 FILLER_13_415 ();
 sg13g2_fill_2 FILLER_13_546 ();
 sg13g2_fill_1 FILLER_13_556 ();
 sg13g2_fill_1 FILLER_13_630 ();
 sg13g2_fill_1 FILLER_13_652 ();
 sg13g2_fill_2 FILLER_13_671 ();
 sg13g2_fill_2 FILLER_13_689 ();
 sg13g2_decap_4 FILLER_13_696 ();
 sg13g2_fill_1 FILLER_13_708 ();
 sg13g2_fill_1 FILLER_13_716 ();
 sg13g2_fill_2 FILLER_13_741 ();
 sg13g2_fill_1 FILLER_13_764 ();
 sg13g2_fill_2 FILLER_13_811 ();
 sg13g2_fill_1 FILLER_13_818 ();
 sg13g2_decap_8 FILLER_13_848 ();
 sg13g2_decap_8 FILLER_13_855 ();
 sg13g2_decap_8 FILLER_13_862 ();
 sg13g2_decap_8 FILLER_13_869 ();
 sg13g2_fill_2 FILLER_13_876 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_187 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_fill_1 FILLER_14_229 ();
 sg13g2_fill_1 FILLER_14_240 ();
 sg13g2_fill_2 FILLER_14_267 ();
 sg13g2_fill_2 FILLER_14_325 ();
 sg13g2_fill_2 FILLER_14_339 ();
 sg13g2_fill_1 FILLER_14_341 ();
 sg13g2_fill_2 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_492 ();
 sg13g2_fill_1 FILLER_14_494 ();
 sg13g2_fill_2 FILLER_14_521 ();
 sg13g2_fill_1 FILLER_14_549 ();
 sg13g2_fill_2 FILLER_14_580 ();
 sg13g2_fill_1 FILLER_14_582 ();
 sg13g2_fill_1 FILLER_14_609 ();
 sg13g2_fill_1 FILLER_14_615 ();
 sg13g2_fill_1 FILLER_14_634 ();
 sg13g2_fill_1 FILLER_14_654 ();
 sg13g2_fill_2 FILLER_14_673 ();
 sg13g2_fill_1 FILLER_14_675 ();
 sg13g2_fill_2 FILLER_14_692 ();
 sg13g2_fill_2 FILLER_14_705 ();
 sg13g2_fill_1 FILLER_14_712 ();
 sg13g2_fill_2 FILLER_14_724 ();
 sg13g2_fill_2 FILLER_14_742 ();
 sg13g2_fill_1 FILLER_14_744 ();
 sg13g2_fill_1 FILLER_14_766 ();
 sg13g2_fill_2 FILLER_14_776 ();
 sg13g2_fill_2 FILLER_14_820 ();
 sg13g2_fill_1 FILLER_14_836 ();
 sg13g2_decap_8 FILLER_14_845 ();
 sg13g2_decap_8 FILLER_14_852 ();
 sg13g2_decap_8 FILLER_14_863 ();
 sg13g2_decap_8 FILLER_14_870 ();
 sg13g2_fill_1 FILLER_14_877 ();
 sg13g2_fill_1 FILLER_15_85 ();
 sg13g2_fill_1 FILLER_15_112 ();
 sg13g2_fill_1 FILLER_15_139 ();
 sg13g2_fill_2 FILLER_15_166 ();
 sg13g2_fill_2 FILLER_15_194 ();
 sg13g2_fill_2 FILLER_15_222 ();
 sg13g2_fill_1 FILLER_15_250 ();
 sg13g2_fill_1 FILLER_15_277 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_fill_1 FILLER_15_328 ();
 sg13g2_fill_2 FILLER_15_333 ();
 sg13g2_fill_2 FILLER_15_345 ();
 sg13g2_fill_2 FILLER_15_374 ();
 sg13g2_fill_2 FILLER_15_426 ();
 sg13g2_fill_1 FILLER_15_480 ();
 sg13g2_fill_1 FILLER_15_507 ();
 sg13g2_fill_2 FILLER_15_600 ();
 sg13g2_fill_1 FILLER_15_602 ();
 sg13g2_fill_1 FILLER_15_664 ();
 sg13g2_decap_4 FILLER_15_669 ();
 sg13g2_fill_1 FILLER_15_673 ();
 sg13g2_fill_2 FILLER_15_696 ();
 sg13g2_fill_1 FILLER_15_703 ();
 sg13g2_fill_2 FILLER_15_731 ();
 sg13g2_fill_1 FILLER_15_737 ();
 sg13g2_fill_1 FILLER_15_745 ();
 sg13g2_decap_4 FILLER_15_763 ();
 sg13g2_fill_2 FILLER_15_791 ();
 sg13g2_fill_1 FILLER_15_793 ();
 sg13g2_fill_2 FILLER_15_802 ();
 sg13g2_fill_2 FILLER_15_812 ();
 sg13g2_fill_1 FILLER_15_814 ();
 sg13g2_fill_2 FILLER_15_842 ();
 sg13g2_decap_4 FILLER_15_870 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_fill_1 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_24 ();
 sg13g2_fill_2 FILLER_16_52 ();
 sg13g2_fill_1 FILLER_16_54 ();
 sg13g2_fill_1 FILLER_16_59 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_fill_1 FILLER_16_178 ();
 sg13g2_fill_1 FILLER_16_205 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_fill_2 FILLER_16_299 ();
 sg13g2_fill_2 FILLER_16_320 ();
 sg13g2_fill_1 FILLER_16_327 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_fill_1 FILLER_16_349 ();
 sg13g2_fill_2 FILLER_16_355 ();
 sg13g2_fill_2 FILLER_16_364 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_fill_1 FILLER_16_388 ();
 sg13g2_fill_2 FILLER_16_426 ();
 sg13g2_fill_2 FILLER_16_438 ();
 sg13g2_fill_1 FILLER_16_440 ();
 sg13g2_fill_1 FILLER_16_445 ();
 sg13g2_decap_8 FILLER_16_450 ();
 sg13g2_fill_2 FILLER_16_457 ();
 sg13g2_decap_4 FILLER_16_463 ();
 sg13g2_fill_1 FILLER_16_467 ();
 sg13g2_fill_2 FILLER_16_498 ();
 sg13g2_fill_2 FILLER_16_526 ();
 sg13g2_fill_1 FILLER_16_528 ();
 sg13g2_decap_8 FILLER_16_593 ();
 sg13g2_fill_2 FILLER_16_600 ();
 sg13g2_fill_1 FILLER_16_602 ();
 sg13g2_fill_2 FILLER_16_606 ();
 sg13g2_fill_1 FILLER_16_608 ();
 sg13g2_fill_2 FILLER_16_618 ();
 sg13g2_fill_2 FILLER_16_654 ();
 sg13g2_fill_1 FILLER_16_656 ();
 sg13g2_decap_8 FILLER_16_681 ();
 sg13g2_fill_1 FILLER_16_693 ();
 sg13g2_decap_4 FILLER_16_707 ();
 sg13g2_fill_1 FILLER_16_711 ();
 sg13g2_fill_2 FILLER_16_731 ();
 sg13g2_fill_2 FILLER_16_762 ();
 sg13g2_fill_2 FILLER_16_790 ();
 sg13g2_fill_1 FILLER_16_818 ();
 sg13g2_fill_1 FILLER_16_877 ();
 sg13g2_fill_1 FILLER_17_26 ();
 sg13g2_fill_2 FILLER_17_35 ();
 sg13g2_fill_1 FILLER_17_37 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_262 ();
 sg13g2_fill_2 FILLER_17_287 ();
 sg13g2_fill_2 FILLER_17_570 ();
 sg13g2_decap_8 FILLER_17_576 ();
 sg13g2_decap_4 FILLER_17_583 ();
 sg13g2_fill_2 FILLER_17_609 ();
 sg13g2_fill_1 FILLER_17_637 ();
 sg13g2_fill_1 FILLER_17_646 ();
 sg13g2_fill_1 FILLER_17_655 ();
 sg13g2_fill_2 FILLER_17_704 ();
 sg13g2_fill_1 FILLER_17_749 ();
 sg13g2_fill_1 FILLER_17_755 ();
 sg13g2_fill_1 FILLER_17_769 ();
 sg13g2_fill_1 FILLER_17_775 ();
 sg13g2_fill_2 FILLER_17_781 ();
 sg13g2_fill_2 FILLER_17_793 ();
 sg13g2_fill_2 FILLER_17_804 ();
 sg13g2_fill_2 FILLER_17_810 ();
 sg13g2_fill_2 FILLER_17_817 ();
 sg13g2_fill_1 FILLER_17_819 ();
 sg13g2_fill_1 FILLER_17_824 ();
 sg13g2_fill_2 FILLER_17_846 ();
 sg13g2_fill_2 FILLER_18_8 ();
 sg13g2_fill_2 FILLER_18_51 ();
 sg13g2_fill_1 FILLER_18_53 ();
 sg13g2_fill_2 FILLER_18_62 ();
 sg13g2_fill_2 FILLER_18_76 ();
 sg13g2_fill_2 FILLER_18_120 ();
 sg13g2_fill_1 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_181 ();
 sg13g2_fill_1 FILLER_18_183 ();
 sg13g2_fill_1 FILLER_18_218 ();
 sg13g2_fill_1 FILLER_18_237 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_fill_2 FILLER_18_405 ();
 sg13g2_fill_1 FILLER_18_412 ();
 sg13g2_fill_2 FILLER_18_435 ();
 sg13g2_decap_4 FILLER_18_442 ();
 sg13g2_fill_1 FILLER_18_446 ();
 sg13g2_fill_2 FILLER_18_455 ();
 sg13g2_fill_1 FILLER_18_457 ();
 sg13g2_fill_1 FILLER_18_512 ();
 sg13g2_fill_2 FILLER_18_525 ();
 sg13g2_fill_2 FILLER_18_531 ();
 sg13g2_fill_2 FILLER_18_563 ();
 sg13g2_decap_8 FILLER_18_569 ();
 sg13g2_decap_8 FILLER_18_576 ();
 sg13g2_decap_4 FILLER_18_583 ();
 sg13g2_fill_2 FILLER_18_587 ();
 sg13g2_fill_1 FILLER_18_602 ();
 sg13g2_fill_1 FILLER_18_616 ();
 sg13g2_fill_1 FILLER_18_625 ();
 sg13g2_fill_2 FILLER_18_642 ();
 sg13g2_fill_1 FILLER_18_644 ();
 sg13g2_fill_1 FILLER_18_674 ();
 sg13g2_decap_8 FILLER_18_685 ();
 sg13g2_decap_4 FILLER_18_692 ();
 sg13g2_fill_1 FILLER_18_696 ();
 sg13g2_fill_1 FILLER_18_750 ();
 sg13g2_fill_1 FILLER_18_755 ();
 sg13g2_decap_4 FILLER_18_775 ();
 sg13g2_fill_2 FILLER_18_795 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_4 FILLER_18_815 ();
 sg13g2_fill_1 FILLER_18_819 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_6 ();
 sg13g2_fill_2 FILLER_19_12 ();
 sg13g2_fill_2 FILLER_19_44 ();
 sg13g2_fill_1 FILLER_19_46 ();
 sg13g2_fill_2 FILLER_19_103 ();
 sg13g2_fill_1 FILLER_19_131 ();
 sg13g2_fill_1 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_260 ();
 sg13g2_fill_1 FILLER_19_271 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_fill_1 FILLER_19_311 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_fill_1 FILLER_19_350 ();
 sg13g2_fill_1 FILLER_19_380 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_491 ();
 sg13g2_fill_2 FILLER_19_523 ();
 sg13g2_decap_4 FILLER_19_529 ();
 sg13g2_decap_4 FILLER_19_559 ();
 sg13g2_fill_1 FILLER_19_589 ();
 sg13g2_fill_1 FILLER_19_598 ();
 sg13g2_fill_2 FILLER_19_705 ();
 sg13g2_fill_1 FILLER_19_748 ();
 sg13g2_fill_2 FILLER_19_753 ();
 sg13g2_fill_1 FILLER_19_771 ();
 sg13g2_fill_2 FILLER_19_777 ();
 sg13g2_decap_4 FILLER_19_803 ();
 sg13g2_fill_1 FILLER_19_819 ();
 sg13g2_fill_1 FILLER_19_859 ();
 sg13g2_fill_2 FILLER_19_868 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_237 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_fill_2 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_358 ();
 sg13g2_fill_1 FILLER_20_363 ();
 sg13g2_decap_4 FILLER_20_391 ();
 sg13g2_fill_1 FILLER_20_400 ();
 sg13g2_fill_1 FILLER_20_405 ();
 sg13g2_fill_1 FILLER_20_412 ();
 sg13g2_fill_1 FILLER_20_419 ();
 sg13g2_fill_1 FILLER_20_433 ();
 sg13g2_fill_1 FILLER_20_439 ();
 sg13g2_decap_4 FILLER_20_444 ();
 sg13g2_decap_8 FILLER_20_452 ();
 sg13g2_decap_4 FILLER_20_459 ();
 sg13g2_fill_2 FILLER_20_463 ();
 sg13g2_fill_1 FILLER_20_473 ();
 sg13g2_fill_1 FILLER_20_512 ();
 sg13g2_fill_1 FILLER_20_517 ();
 sg13g2_fill_1 FILLER_20_544 ();
 sg13g2_fill_1 FILLER_20_596 ();
 sg13g2_fill_2 FILLER_20_630 ();
 sg13g2_fill_2 FILLER_20_658 ();
 sg13g2_fill_2 FILLER_20_674 ();
 sg13g2_fill_1 FILLER_20_676 ();
 sg13g2_fill_1 FILLER_20_730 ();
 sg13g2_fill_1 FILLER_20_747 ();
 sg13g2_fill_1 FILLER_20_752 ();
 sg13g2_fill_2 FILLER_20_774 ();
 sg13g2_fill_1 FILLER_20_796 ();
 sg13g2_fill_2 FILLER_20_828 ();
 sg13g2_fill_1 FILLER_20_842 ();
 sg13g2_fill_2 FILLER_20_875 ();
 sg13g2_fill_1 FILLER_20_877 ();
 sg13g2_fill_1 FILLER_21_26 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_fill_2 FILLER_21_108 ();
 sg13g2_fill_2 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_246 ();
 sg13g2_fill_2 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_fill_1 FILLER_21_291 ();
 sg13g2_fill_2 FILLER_21_310 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_329 ();
 sg13g2_decap_4 FILLER_21_360 ();
 sg13g2_fill_1 FILLER_21_364 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_499 ();
 sg13g2_fill_1 FILLER_21_501 ();
 sg13g2_decap_4 FILLER_21_506 ();
 sg13g2_fill_1 FILLER_21_510 ();
 sg13g2_decap_4 FILLER_21_546 ();
 sg13g2_fill_2 FILLER_21_550 ();
 sg13g2_fill_2 FILLER_21_556 ();
 sg13g2_decap_4 FILLER_21_562 ();
 sg13g2_fill_2 FILLER_21_629 ();
 sg13g2_fill_2 FILLER_21_661 ();
 sg13g2_fill_1 FILLER_21_737 ();
 sg13g2_fill_1 FILLER_21_754 ();
 sg13g2_fill_2 FILLER_21_763 ();
 sg13g2_fill_1 FILLER_21_771 ();
 sg13g2_fill_2 FILLER_21_788 ();
 sg13g2_fill_1 FILLER_21_803 ();
 sg13g2_fill_1 FILLER_21_824 ();
 sg13g2_fill_2 FILLER_21_846 ();
 sg13g2_fill_2 FILLER_21_870 ();
 sg13g2_fill_1 FILLER_21_877 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_239 ();
 sg13g2_fill_2 FILLER_22_253 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_319 ();
 sg13g2_fill_1 FILLER_22_328 ();
 sg13g2_fill_2 FILLER_22_333 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_353 ();
 sg13g2_decap_4 FILLER_22_360 ();
 sg13g2_fill_1 FILLER_22_405 ();
 sg13g2_fill_1 FILLER_22_410 ();
 sg13g2_fill_1 FILLER_22_415 ();
 sg13g2_fill_1 FILLER_22_434 ();
 sg13g2_fill_1 FILLER_22_439 ();
 sg13g2_fill_1 FILLER_22_444 ();
 sg13g2_fill_1 FILLER_22_450 ();
 sg13g2_fill_2 FILLER_22_455 ();
 sg13g2_fill_1 FILLER_22_457 ();
 sg13g2_fill_2 FILLER_22_462 ();
 sg13g2_fill_1 FILLER_22_464 ();
 sg13g2_decap_8 FILLER_22_662 ();
 sg13g2_fill_1 FILLER_22_669 ();
 sg13g2_fill_1 FILLER_22_679 ();
 sg13g2_fill_2 FILLER_22_730 ();
 sg13g2_fill_2 FILLER_22_748 ();
 sg13g2_fill_1 FILLER_22_759 ();
 sg13g2_fill_2 FILLER_22_765 ();
 sg13g2_fill_2 FILLER_22_816 ();
 sg13g2_fill_1 FILLER_22_818 ();
 sg13g2_fill_2 FILLER_22_846 ();
 sg13g2_fill_2 FILLER_22_858 ();
 sg13g2_fill_2 FILLER_22_875 ();
 sg13g2_fill_1 FILLER_22_877 ();
 sg13g2_fill_1 FILLER_23_44 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_304 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_decap_4 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_fill_1 FILLER_23_375 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_2 FILLER_23_387 ();
 sg13g2_fill_2 FILLER_23_393 ();
 sg13g2_decap_4 FILLER_23_411 ();
 sg13g2_fill_2 FILLER_23_420 ();
 sg13g2_fill_1 FILLER_23_422 ();
 sg13g2_fill_2 FILLER_23_426 ();
 sg13g2_fill_2 FILLER_23_448 ();
 sg13g2_fill_1 FILLER_23_450 ();
 sg13g2_fill_2 FILLER_23_507 ();
 sg13g2_decap_8 FILLER_23_521 ();
 sg13g2_fill_1 FILLER_23_528 ();
 sg13g2_fill_1 FILLER_23_537 ();
 sg13g2_fill_2 FILLER_23_542 ();
 sg13g2_fill_2 FILLER_23_570 ();
 sg13g2_fill_1 FILLER_23_572 ();
 sg13g2_fill_1 FILLER_23_627 ();
 sg13g2_fill_2 FILLER_23_634 ();
 sg13g2_fill_2 FILLER_23_669 ();
 sg13g2_fill_1 FILLER_23_717 ();
 sg13g2_fill_2 FILLER_23_741 ();
 sg13g2_fill_1 FILLER_23_781 ();
 sg13g2_fill_1 FILLER_23_804 ();
 sg13g2_fill_2 FILLER_23_841 ();
 sg13g2_fill_1 FILLER_23_843 ();
 sg13g2_fill_2 FILLER_23_849 ();
 sg13g2_fill_1 FILLER_23_851 ();
 sg13g2_fill_2 FILLER_24_26 ();
 sg13g2_decap_4 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_decap_4 FILLER_24_335 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_fill_1 FILLER_24_368 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_fill_1 FILLER_24_388 ();
 sg13g2_fill_2 FILLER_24_394 ();
 sg13g2_fill_1 FILLER_24_419 ();
 sg13g2_fill_2 FILLER_24_430 ();
 sg13g2_fill_1 FILLER_24_432 ();
 sg13g2_fill_2 FILLER_24_596 ();
 sg13g2_fill_1 FILLER_24_598 ();
 sg13g2_fill_2 FILLER_24_618 ();
 sg13g2_fill_2 FILLER_24_649 ();
 sg13g2_fill_2 FILLER_24_674 ();
 sg13g2_fill_2 FILLER_24_693 ();
 sg13g2_fill_1 FILLER_24_700 ();
 sg13g2_fill_2 FILLER_24_706 ();
 sg13g2_fill_1 FILLER_24_729 ();
 sg13g2_fill_1 FILLER_24_759 ();
 sg13g2_fill_1 FILLER_24_777 ();
 sg13g2_fill_1 FILLER_24_800 ();
 sg13g2_fill_1 FILLER_24_811 ();
 sg13g2_fill_2 FILLER_24_839 ();
 sg13g2_fill_1 FILLER_24_841 ();
 sg13g2_fill_1 FILLER_24_850 ();
 sg13g2_decap_4 FILLER_24_863 ();
 sg13g2_fill_2 FILLER_24_871 ();
 sg13g2_fill_1 FILLER_24_873 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_2 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_341 ();
 sg13g2_decap_4 FILLER_25_348 ();
 sg13g2_fill_1 FILLER_25_378 ();
 sg13g2_fill_2 FILLER_25_392 ();
 sg13g2_fill_2 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_431 ();
 sg13g2_fill_2 FILLER_25_459 ();
 sg13g2_fill_1 FILLER_25_545 ();
 sg13g2_fill_2 FILLER_25_575 ();
 sg13g2_fill_2 FILLER_25_581 ();
 sg13g2_fill_2 FILLER_25_587 ();
 sg13g2_fill_2 FILLER_25_638 ();
 sg13g2_decap_8 FILLER_25_645 ();
 sg13g2_fill_1 FILLER_25_652 ();
 sg13g2_fill_2 FILLER_25_687 ();
 sg13g2_fill_1 FILLER_25_707 ();
 sg13g2_fill_2 FILLER_25_718 ();
 sg13g2_fill_2 FILLER_25_775 ();
 sg13g2_decap_8 FILLER_25_817 ();
 sg13g2_decap_4 FILLER_25_824 ();
 sg13g2_fill_1 FILLER_25_846 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_50 ();
 sg13g2_fill_2 FILLER_26_96 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_fill_1 FILLER_26_269 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_fill_1 FILLER_26_318 ();
 sg13g2_fill_2 FILLER_26_323 ();
 sg13g2_decap_4 FILLER_26_329 ();
 sg13g2_decap_4 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_fill_1 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_486 ();
 sg13g2_fill_1 FILLER_26_569 ();
 sg13g2_fill_1 FILLER_26_579 ();
 sg13g2_fill_1 FILLER_26_586 ();
 sg13g2_decap_4 FILLER_26_592 ();
 sg13g2_fill_1 FILLER_26_596 ();
 sg13g2_fill_1 FILLER_26_603 ();
 sg13g2_fill_2 FILLER_26_612 ();
 sg13g2_fill_1 FILLER_26_622 ();
 sg13g2_fill_2 FILLER_26_675 ();
 sg13g2_fill_2 FILLER_26_689 ();
 sg13g2_fill_1 FILLER_26_691 ();
 sg13g2_fill_2 FILLER_26_795 ();
 sg13g2_fill_2 FILLER_26_817 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_fill_2 FILLER_27_69 ();
 sg13g2_fill_1 FILLER_27_71 ();
 sg13g2_fill_1 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_fill_1 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_229 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_305 ();
 sg13g2_fill_2 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_413 ();
 sg13g2_fill_1 FILLER_27_483 ();
 sg13g2_fill_1 FILLER_27_509 ();
 sg13g2_fill_1 FILLER_27_530 ();
 sg13g2_fill_2 FILLER_27_536 ();
 sg13g2_fill_1 FILLER_27_546 ();
 sg13g2_fill_1 FILLER_27_565 ();
 sg13g2_fill_1 FILLER_27_571 ();
 sg13g2_fill_1 FILLER_27_582 ();
 sg13g2_fill_2 FILLER_27_597 ();
 sg13g2_fill_1 FILLER_27_599 ();
 sg13g2_fill_1 FILLER_27_605 ();
 sg13g2_fill_2 FILLER_27_616 ();
 sg13g2_fill_1 FILLER_27_618 ();
 sg13g2_fill_2 FILLER_27_635 ();
 sg13g2_fill_2 FILLER_27_641 ();
 sg13g2_fill_1 FILLER_27_643 ();
 sg13g2_fill_2 FILLER_27_648 ();
 sg13g2_fill_1 FILLER_27_650 ();
 sg13g2_fill_2 FILLER_27_707 ();
 sg13g2_fill_2 FILLER_27_729 ();
 sg13g2_fill_1 FILLER_27_731 ();
 sg13g2_fill_1 FILLER_27_785 ();
 sg13g2_fill_2 FILLER_27_812 ();
 sg13g2_fill_1 FILLER_27_814 ();
 sg13g2_fill_1 FILLER_27_845 ();
 sg13g2_fill_2 FILLER_28_153 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_decap_4 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_186 ();
 sg13g2_fill_2 FILLER_28_266 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_fill_2 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_28_438 ();
 sg13g2_decap_4 FILLER_28_470 ();
 sg13g2_fill_2 FILLER_28_474 ();
 sg13g2_fill_2 FILLER_28_519 ();
 sg13g2_fill_1 FILLER_28_547 ();
 sg13g2_fill_2 FILLER_28_573 ();
 sg13g2_fill_1 FILLER_28_579 ();
 sg13g2_decap_4 FILLER_28_585 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_fill_2 FILLER_28_609 ();
 sg13g2_fill_2 FILLER_28_624 ();
 sg13g2_fill_1 FILLER_28_662 ();
 sg13g2_fill_1 FILLER_28_694 ();
 sg13g2_fill_1 FILLER_28_721 ();
 sg13g2_fill_1 FILLER_28_766 ();
 sg13g2_fill_2 FILLER_28_814 ();
 sg13g2_fill_2 FILLER_28_826 ();
 sg13g2_fill_1 FILLER_28_867 ();
 sg13g2_decap_4 FILLER_28_873 ();
 sg13g2_fill_1 FILLER_28_877 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_134 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_29_395 ();
 sg13g2_fill_2 FILLER_29_423 ();
 sg13g2_fill_1 FILLER_29_425 ();
 sg13g2_fill_2 FILLER_29_513 ();
 sg13g2_fill_1 FILLER_29_560 ();
 sg13g2_decap_4 FILLER_29_613 ();
 sg13g2_fill_1 FILLER_29_635 ();
 sg13g2_fill_2 FILLER_29_649 ();
 sg13g2_fill_1 FILLER_29_661 ();
 sg13g2_fill_2 FILLER_29_681 ();
 sg13g2_fill_1 FILLER_29_683 ();
 sg13g2_fill_2 FILLER_29_718 ();
 sg13g2_fill_1 FILLER_29_720 ();
 sg13g2_fill_1 FILLER_29_814 ();
 sg13g2_fill_1 FILLER_29_867 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_fill_1 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_173 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_384 ();
 sg13g2_fill_2 FILLER_30_452 ();
 sg13g2_fill_1 FILLER_30_459 ();
 sg13g2_fill_2 FILLER_30_486 ();
 sg13g2_fill_1 FILLER_30_518 ();
 sg13g2_fill_1 FILLER_30_577 ();
 sg13g2_fill_2 FILLER_30_596 ();
 sg13g2_fill_1 FILLER_30_598 ();
 sg13g2_fill_1 FILLER_30_608 ();
 sg13g2_fill_1 FILLER_30_618 ();
 sg13g2_fill_2 FILLER_30_623 ();
 sg13g2_fill_1 FILLER_30_630 ();
 sg13g2_fill_2 FILLER_30_636 ();
 sg13g2_fill_2 FILLER_30_666 ();
 sg13g2_fill_2 FILLER_30_678 ();
 sg13g2_fill_1 FILLER_30_680 ();
 sg13g2_fill_2 FILLER_30_690 ();
 sg13g2_fill_1 FILLER_30_734 ();
 sg13g2_fill_1 FILLER_30_798 ();
 sg13g2_fill_2 FILLER_30_809 ();
 sg13g2_fill_1 FILLER_30_821 ();
 sg13g2_fill_1 FILLER_30_832 ();
 sg13g2_fill_1 FILLER_30_843 ();
 sg13g2_fill_1 FILLER_30_865 ();
 sg13g2_fill_2 FILLER_30_870 ();
 sg13g2_fill_1 FILLER_30_872 ();
 sg13g2_fill_1 FILLER_31_27 ();
 sg13g2_fill_1 FILLER_31_66 ();
 sg13g2_fill_2 FILLER_31_71 ();
 sg13g2_fill_2 FILLER_31_170 ();
 sg13g2_fill_2 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_286 ();
 sg13g2_fill_1 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_412 ();
 sg13g2_fill_2 FILLER_31_426 ();
 sg13g2_fill_2 FILLER_31_457 ();
 sg13g2_fill_2 FILLER_31_494 ();
 sg13g2_fill_1 FILLER_31_511 ();
 sg13g2_fill_1 FILLER_31_522 ();
 sg13g2_fill_1 FILLER_31_531 ();
 sg13g2_fill_1 FILLER_31_536 ();
 sg13g2_fill_2 FILLER_31_546 ();
 sg13g2_fill_2 FILLER_31_556 ();
 sg13g2_fill_2 FILLER_31_589 ();
 sg13g2_fill_1 FILLER_31_595 ();
 sg13g2_fill_2 FILLER_31_620 ();
 sg13g2_fill_1 FILLER_31_622 ();
 sg13g2_fill_2 FILLER_31_635 ();
 sg13g2_fill_1 FILLER_31_637 ();
 sg13g2_fill_1 FILLER_31_647 ();
 sg13g2_fill_2 FILLER_31_658 ();
 sg13g2_fill_1 FILLER_31_660 ();
 sg13g2_fill_2 FILLER_31_671 ();
 sg13g2_fill_1 FILLER_31_707 ();
 sg13g2_fill_2 FILLER_31_865 ();
 sg13g2_decap_4 FILLER_31_872 ();
 sg13g2_fill_2 FILLER_31_876 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_186 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_227 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_fill_1 FILLER_32_295 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_390 ();
 sg13g2_fill_2 FILLER_32_395 ();
 sg13g2_fill_1 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_432 ();
 sg13g2_fill_2 FILLER_32_437 ();
 sg13g2_fill_2 FILLER_32_465 ();
 sg13g2_fill_1 FILLER_32_471 ();
 sg13g2_decap_4 FILLER_32_498 ();
 sg13g2_fill_1 FILLER_32_502 ();
 sg13g2_fill_2 FILLER_32_521 ();
 sg13g2_fill_1 FILLER_32_523 ();
 sg13g2_fill_2 FILLER_32_529 ();
 sg13g2_fill_1 FILLER_32_531 ();
 sg13g2_fill_1 FILLER_32_544 ();
 sg13g2_fill_1 FILLER_32_550 ();
 sg13g2_fill_1 FILLER_32_565 ();
 sg13g2_fill_1 FILLER_32_571 ();
 sg13g2_fill_1 FILLER_32_576 ();
 sg13g2_fill_1 FILLER_32_582 ();
 sg13g2_fill_1 FILLER_32_588 ();
 sg13g2_fill_1 FILLER_32_603 ();
 sg13g2_fill_1 FILLER_32_609 ();
 sg13g2_fill_1 FILLER_32_614 ();
 sg13g2_fill_1 FILLER_32_620 ();
 sg13g2_fill_1 FILLER_32_626 ();
 sg13g2_fill_1 FILLER_32_632 ();
 sg13g2_fill_1 FILLER_32_638 ();
 sg13g2_fill_2 FILLER_32_643 ();
 sg13g2_fill_1 FILLER_32_645 ();
 sg13g2_fill_2 FILLER_32_658 ();
 sg13g2_fill_2 FILLER_32_709 ();
 sg13g2_fill_1 FILLER_32_711 ();
 sg13g2_fill_2 FILLER_32_741 ();
 sg13g2_fill_2 FILLER_32_764 ();
 sg13g2_fill_1 FILLER_32_766 ();
 sg13g2_fill_1 FILLER_32_863 ();
 sg13g2_decap_4 FILLER_32_874 ();
 sg13g2_fill_2 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_fill_2 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_414 ();
 sg13g2_fill_2 FILLER_33_436 ();
 sg13g2_fill_1 FILLER_33_491 ();
 sg13g2_fill_2 FILLER_33_498 ();
 sg13g2_fill_2 FILLER_33_505 ();
 sg13g2_fill_1 FILLER_33_533 ();
 sg13g2_fill_1 FILLER_33_538 ();
 sg13g2_fill_1 FILLER_33_544 ();
 sg13g2_fill_2 FILLER_33_550 ();
 sg13g2_fill_1 FILLER_33_556 ();
 sg13g2_fill_2 FILLER_33_572 ();
 sg13g2_fill_1 FILLER_33_579 ();
 sg13g2_fill_1 FILLER_33_627 ();
 sg13g2_fill_1 FILLER_33_637 ();
 sg13g2_fill_1 FILLER_33_647 ();
 sg13g2_fill_1 FILLER_33_652 ();
 sg13g2_fill_1 FILLER_33_657 ();
 sg13g2_fill_2 FILLER_33_681 ();
 sg13g2_fill_1 FILLER_33_683 ();
 sg13g2_fill_1 FILLER_33_689 ();
 sg13g2_fill_1 FILLER_33_729 ();
 sg13g2_fill_1 FILLER_33_751 ();
 sg13g2_fill_1 FILLER_33_762 ();
 sg13g2_fill_1 FILLER_33_771 ();
 sg13g2_fill_1 FILLER_33_793 ();
 sg13g2_fill_1 FILLER_33_815 ();
 sg13g2_fill_1 FILLER_33_826 ();
 sg13g2_fill_1 FILLER_33_837 ();
 sg13g2_fill_2 FILLER_33_859 ();
 sg13g2_decap_8 FILLER_33_871 ();
 sg13g2_fill_1 FILLER_34_138 ();
 sg13g2_fill_1 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_235 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_304 ();
 sg13g2_fill_1 FILLER_34_319 ();
 sg13g2_fill_1 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_423 ();
 sg13g2_fill_2 FILLER_34_446 ();
 sg13g2_fill_1 FILLER_34_452 ();
 sg13g2_fill_2 FILLER_34_457 ();
 sg13g2_fill_2 FILLER_34_485 ();
 sg13g2_fill_2 FILLER_34_496 ();
 sg13g2_fill_1 FILLER_34_502 ();
 sg13g2_fill_1 FILLER_34_529 ();
 sg13g2_fill_2 FILLER_34_534 ();
 sg13g2_fill_1 FILLER_34_544 ();
 sg13g2_fill_1 FILLER_34_572 ();
 sg13g2_fill_1 FILLER_34_581 ();
 sg13g2_decap_4 FILLER_34_587 ();
 sg13g2_fill_1 FILLER_34_614 ();
 sg13g2_decap_4 FILLER_34_624 ();
 sg13g2_fill_2 FILLER_34_706 ();
 sg13g2_fill_2 FILLER_34_831 ();
 sg13g2_fill_1 FILLER_34_868 ();
 sg13g2_fill_1 FILLER_34_877 ();
 sg13g2_fill_1 FILLER_35_11 ();
 sg13g2_fill_2 FILLER_35_38 ();
 sg13g2_fill_2 FILLER_35_100 ();
 sg13g2_fill_1 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_174 ();
 sg13g2_fill_2 FILLER_35_186 ();
 sg13g2_fill_1 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_fill_2 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_440 ();
 sg13g2_fill_1 FILLER_35_450 ();
 sg13g2_fill_2 FILLER_35_456 ();
 sg13g2_fill_2 FILLER_35_516 ();
 sg13g2_fill_2 FILLER_35_523 ();
 sg13g2_fill_1 FILLER_35_559 ();
 sg13g2_fill_2 FILLER_35_614 ();
 sg13g2_fill_1 FILLER_35_616 ();
 sg13g2_fill_2 FILLER_35_655 ();
 sg13g2_fill_1 FILLER_35_657 ();
 sg13g2_fill_1 FILLER_35_689 ();
 sg13g2_fill_2 FILLER_35_751 ();
 sg13g2_fill_1 FILLER_35_779 ();
 sg13g2_fill_1 FILLER_35_790 ();
 sg13g2_decap_8 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_35_868 ();
 sg13g2_fill_2 FILLER_35_875 ();
 sg13g2_fill_1 FILLER_35_877 ();
 sg13g2_fill_1 FILLER_36_82 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_331 ();
 sg13g2_fill_2 FILLER_36_349 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_fill_1 FILLER_36_428 ();
 sg13g2_fill_1 FILLER_36_441 ();
 sg13g2_fill_2 FILLER_36_455 ();
 sg13g2_fill_1 FILLER_36_469 ();
 sg13g2_fill_2 FILLER_36_485 ();
 sg13g2_fill_1 FILLER_36_487 ();
 sg13g2_decap_4 FILLER_36_497 ();
 sg13g2_fill_1 FILLER_36_509 ();
 sg13g2_fill_1 FILLER_36_514 ();
 sg13g2_fill_2 FILLER_36_546 ();
 sg13g2_fill_1 FILLER_36_570 ();
 sg13g2_fill_1 FILLER_36_577 ();
 sg13g2_fill_1 FILLER_36_587 ();
 sg13g2_fill_1 FILLER_36_592 ();
 sg13g2_fill_2 FILLER_36_606 ();
 sg13g2_fill_1 FILLER_36_612 ();
 sg13g2_fill_1 FILLER_36_623 ();
 sg13g2_fill_2 FILLER_36_628 ();
 sg13g2_fill_2 FILLER_36_638 ();
 sg13g2_fill_1 FILLER_36_680 ();
 sg13g2_fill_1 FILLER_36_702 ();
 sg13g2_fill_2 FILLER_36_708 ();
 sg13g2_fill_1 FILLER_36_715 ();
 sg13g2_fill_2 FILLER_36_726 ();
 sg13g2_fill_2 FILLER_36_733 ();
 sg13g2_fill_2 FILLER_36_743 ();
 sg13g2_fill_1 FILLER_36_853 ();
 sg13g2_decap_8 FILLER_36_862 ();
 sg13g2_decap_4 FILLER_36_873 ();
 sg13g2_fill_1 FILLER_36_877 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_5 ();
 sg13g2_fill_2 FILLER_37_25 ();
 sg13g2_fill_1 FILLER_37_27 ();
 sg13g2_fill_2 FILLER_37_82 ();
 sg13g2_fill_2 FILLER_37_110 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_fill_2 FILLER_37_252 ();
 sg13g2_fill_1 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_265 ();
 sg13g2_fill_2 FILLER_37_279 ();
 sg13g2_fill_1 FILLER_37_286 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_1 FILLER_37_316 ();
 sg13g2_fill_2 FILLER_37_356 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_fill_2 FILLER_37_377 ();
 sg13g2_fill_1 FILLER_37_406 ();
 sg13g2_fill_2 FILLER_37_415 ();
 sg13g2_fill_2 FILLER_37_439 ();
 sg13g2_fill_1 FILLER_37_441 ();
 sg13g2_fill_2 FILLER_37_449 ();
 sg13g2_fill_2 FILLER_37_491 ();
 sg13g2_fill_2 FILLER_37_498 ();
 sg13g2_fill_2 FILLER_37_505 ();
 sg13g2_fill_1 FILLER_37_507 ();
 sg13g2_fill_2 FILLER_37_513 ();
 sg13g2_fill_1 FILLER_37_515 ();
 sg13g2_fill_1 FILLER_37_521 ();
 sg13g2_fill_1 FILLER_37_585 ();
 sg13g2_fill_1 FILLER_37_601 ();
 sg13g2_fill_2 FILLER_37_628 ();
 sg13g2_fill_2 FILLER_37_694 ();
 sg13g2_fill_1 FILLER_37_696 ();
 sg13g2_fill_2 FILLER_37_710 ();
 sg13g2_fill_1 FILLER_37_722 ();
 sg13g2_fill_1 FILLER_37_749 ();
 sg13g2_fill_2 FILLER_37_806 ();
 sg13g2_fill_1 FILLER_37_808 ();
 sg13g2_fill_1 FILLER_37_830 ();
 sg13g2_fill_1 FILLER_37_839 ();
 sg13g2_fill_2 FILLER_37_876 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_5 ();
 sg13g2_fill_1 FILLER_38_43 ();
 sg13g2_fill_2 FILLER_38_74 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_152 ();
 sg13g2_fill_1 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_163 ();
 sg13g2_fill_2 FILLER_38_168 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_fill_1 FILLER_38_189 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_211 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_fill_2 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_2 FILLER_38_312 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_360 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_2 FILLER_38_417 ();
 sg13g2_decap_4 FILLER_38_423 ();
 sg13g2_decap_4 FILLER_38_432 ();
 sg13g2_fill_1 FILLER_38_449 ();
 sg13g2_fill_1 FILLER_38_454 ();
 sg13g2_fill_1 FILLER_38_489 ();
 sg13g2_fill_1 FILLER_38_525 ();
 sg13g2_fill_1 FILLER_38_531 ();
 sg13g2_fill_2 FILLER_38_549 ();
 sg13g2_fill_2 FILLER_38_556 ();
 sg13g2_fill_2 FILLER_38_569 ();
 sg13g2_fill_2 FILLER_38_674 ();
 sg13g2_fill_1 FILLER_38_756 ();
 sg13g2_fill_2 FILLER_38_834 ();
 sg13g2_fill_2 FILLER_38_876 ();
 sg13g2_fill_2 FILLER_39_70 ();
 sg13g2_fill_1 FILLER_39_72 ();
 sg13g2_fill_1 FILLER_39_103 ();
 sg13g2_fill_1 FILLER_39_108 ();
 sg13g2_fill_2 FILLER_39_133 ();
 sg13g2_fill_1 FILLER_39_163 ();
 sg13g2_fill_1 FILLER_39_169 ();
 sg13g2_fill_1 FILLER_39_246 ();
 sg13g2_fill_1 FILLER_39_302 ();
 sg13g2_fill_2 FILLER_39_311 ();
 sg13g2_fill_2 FILLER_39_328 ();
 sg13g2_fill_2 FILLER_39_335 ();
 sg13g2_fill_1 FILLER_39_337 ();
 sg13g2_fill_1 FILLER_39_385 ();
 sg13g2_fill_2 FILLER_39_396 ();
 sg13g2_fill_1 FILLER_39_433 ();
 sg13g2_fill_1 FILLER_39_465 ();
 sg13g2_fill_2 FILLER_39_487 ();
 sg13g2_fill_1 FILLER_39_501 ();
 sg13g2_fill_1 FILLER_39_507 ();
 sg13g2_fill_1 FILLER_39_534 ();
 sg13g2_fill_1 FILLER_39_540 ();
 sg13g2_fill_1 FILLER_39_546 ();
 sg13g2_fill_1 FILLER_39_566 ();
 sg13g2_decap_4 FILLER_39_575 ();
 sg13g2_fill_1 FILLER_39_598 ();
 sg13g2_fill_1 FILLER_39_603 ();
 sg13g2_decap_4 FILLER_39_651 ();
 sg13g2_decap_8 FILLER_39_659 ();
 sg13g2_decap_4 FILLER_39_666 ();
 sg13g2_fill_2 FILLER_39_670 ();
 sg13g2_fill_1 FILLER_39_676 ();
 sg13g2_fill_1 FILLER_39_682 ();
 sg13g2_fill_2 FILLER_39_688 ();
 sg13g2_fill_1 FILLER_39_699 ();
 sg13g2_fill_1 FILLER_39_718 ();
 sg13g2_fill_2 FILLER_39_727 ();
 sg13g2_decap_4 FILLER_39_874 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_1 FILLER_40_29 ();
 sg13g2_fill_1 FILLER_40_40 ();
 sg13g2_fill_2 FILLER_40_55 ();
 sg13g2_fill_2 FILLER_40_77 ();
 sg13g2_fill_1 FILLER_40_115 ();
 sg13g2_fill_1 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_141 ();
 sg13g2_fill_1 FILLER_40_143 ();
 sg13g2_fill_2 FILLER_40_158 ();
 sg13g2_fill_1 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_206 ();
 sg13g2_fill_2 FILLER_40_227 ();
 sg13g2_fill_2 FILLER_40_243 ();
 sg13g2_fill_2 FILLER_40_250 ();
 sg13g2_fill_1 FILLER_40_268 ();
 sg13g2_fill_2 FILLER_40_311 ();
 sg13g2_fill_1 FILLER_40_330 ();
 sg13g2_fill_2 FILLER_40_335 ();
 sg13g2_fill_2 FILLER_40_341 ();
 sg13g2_fill_2 FILLER_40_348 ();
 sg13g2_fill_2 FILLER_40_354 ();
 sg13g2_fill_1 FILLER_40_401 ();
 sg13g2_fill_2 FILLER_40_411 ();
 sg13g2_fill_2 FILLER_40_433 ();
 sg13g2_fill_1 FILLER_40_435 ();
 sg13g2_decap_8 FILLER_40_444 ();
 sg13g2_fill_2 FILLER_40_459 ();
 sg13g2_fill_1 FILLER_40_466 ();
 sg13g2_fill_1 FILLER_40_472 ();
 sg13g2_fill_2 FILLER_40_502 ();
 sg13g2_fill_1 FILLER_40_509 ();
 sg13g2_fill_2 FILLER_40_522 ();
 sg13g2_fill_1 FILLER_40_529 ();
 sg13g2_fill_1 FILLER_40_540 ();
 sg13g2_fill_2 FILLER_40_545 ();
 sg13g2_fill_1 FILLER_40_560 ();
 sg13g2_fill_1 FILLER_40_566 ();
 sg13g2_fill_1 FILLER_40_598 ();
 sg13g2_fill_1 FILLER_40_608 ();
 sg13g2_fill_1 FILLER_40_619 ();
 sg13g2_fill_1 FILLER_40_624 ();
 sg13g2_fill_2 FILLER_40_635 ();
 sg13g2_decap_8 FILLER_40_641 ();
 sg13g2_decap_4 FILLER_40_648 ();
 sg13g2_fill_1 FILLER_40_763 ();
 sg13g2_fill_1 FILLER_40_774 ();
 sg13g2_fill_1 FILLER_40_801 ();
 sg13g2_fill_1 FILLER_40_816 ();
 sg13g2_fill_2 FILLER_40_831 ();
 sg13g2_decap_4 FILLER_40_872 ();
 sg13g2_fill_2 FILLER_40_876 ();
 sg13g2_fill_1 FILLER_41_44 ();
 sg13g2_fill_2 FILLER_41_81 ();
 sg13g2_fill_1 FILLER_41_95 ();
 sg13g2_fill_1 FILLER_41_104 ();
 sg13g2_fill_1 FILLER_41_109 ();
 sg13g2_fill_1 FILLER_41_125 ();
 sg13g2_fill_1 FILLER_41_136 ();
 sg13g2_fill_1 FILLER_41_141 ();
 sg13g2_fill_1 FILLER_41_165 ();
 sg13g2_fill_2 FILLER_41_186 ();
 sg13g2_fill_1 FILLER_41_212 ();
 sg13g2_fill_1 FILLER_41_231 ();
 sg13g2_fill_1 FILLER_41_265 ();
 sg13g2_fill_1 FILLER_41_272 ();
 sg13g2_fill_1 FILLER_41_288 ();
 sg13g2_decap_8 FILLER_41_307 ();
 sg13g2_fill_1 FILLER_41_314 ();
 sg13g2_fill_1 FILLER_41_354 ();
 sg13g2_fill_2 FILLER_41_378 ();
 sg13g2_fill_1 FILLER_41_385 ();
 sg13g2_fill_1 FILLER_41_394 ();
 sg13g2_fill_2 FILLER_41_416 ();
 sg13g2_fill_1 FILLER_41_422 ();
 sg13g2_fill_1 FILLER_41_443 ();
 sg13g2_fill_1 FILLER_41_449 ();
 sg13g2_fill_1 FILLER_41_468 ();
 sg13g2_fill_1 FILLER_41_473 ();
 sg13g2_fill_1 FILLER_41_483 ();
 sg13g2_fill_1 FILLER_41_490 ();
 sg13g2_fill_1 FILLER_41_497 ();
 sg13g2_fill_1 FILLER_41_509 ();
 sg13g2_decap_4 FILLER_41_526 ();
 sg13g2_decap_4 FILLER_41_536 ();
 sg13g2_fill_2 FILLER_41_540 ();
 sg13g2_fill_2 FILLER_41_546 ();
 sg13g2_fill_2 FILLER_41_561 ();
 sg13g2_fill_1 FILLER_41_609 ();
 sg13g2_fill_1 FILLER_41_642 ();
 sg13g2_fill_1 FILLER_41_648 ();
 sg13g2_fill_1 FILLER_41_675 ();
 sg13g2_fill_1 FILLER_41_680 ();
 sg13g2_fill_2 FILLER_41_695 ();
 sg13g2_fill_1 FILLER_41_707 ();
 sg13g2_fill_1 FILLER_41_748 ();
 sg13g2_fill_1 FILLER_41_759 ();
 sg13g2_fill_2 FILLER_41_792 ();
 sg13g2_fill_1 FILLER_41_804 ();
 sg13g2_fill_1 FILLER_41_810 ();
 sg13g2_fill_2 FILLER_41_837 ();
 sg13g2_fill_2 FILLER_41_875 ();
 sg13g2_fill_1 FILLER_41_877 ();
 sg13g2_fill_2 FILLER_42_60 ();
 sg13g2_fill_2 FILLER_42_87 ();
 sg13g2_fill_1 FILLER_42_89 ();
 sg13g2_fill_2 FILLER_42_124 ();
 sg13g2_fill_1 FILLER_42_126 ();
 sg13g2_fill_1 FILLER_42_137 ();
 sg13g2_fill_1 FILLER_42_148 ();
 sg13g2_fill_2 FILLER_42_167 ();
 sg13g2_fill_1 FILLER_42_209 ();
 sg13g2_fill_2 FILLER_42_235 ();
 sg13g2_fill_1 FILLER_42_253 ();
 sg13g2_fill_2 FILLER_42_260 ();
 sg13g2_fill_1 FILLER_42_266 ();
 sg13g2_fill_1 FILLER_42_276 ();
 sg13g2_fill_2 FILLER_42_287 ();
 sg13g2_fill_2 FILLER_42_334 ();
 sg13g2_fill_1 FILLER_42_423 ();
 sg13g2_decap_4 FILLER_42_462 ();
 sg13g2_fill_1 FILLER_42_466 ();
 sg13g2_fill_1 FILLER_42_503 ();
 sg13g2_fill_2 FILLER_42_509 ();
 sg13g2_fill_1 FILLER_42_516 ();
 sg13g2_fill_1 FILLER_42_523 ();
 sg13g2_fill_1 FILLER_42_589 ();
 sg13g2_fill_1 FILLER_42_598 ();
 sg13g2_fill_2 FILLER_42_608 ();
 sg13g2_fill_2 FILLER_42_625 ();
 sg13g2_fill_1 FILLER_42_631 ();
 sg13g2_fill_1 FILLER_42_637 ();
 sg13g2_fill_1 FILLER_42_643 ();
 sg13g2_fill_2 FILLER_42_679 ();
 sg13g2_fill_1 FILLER_42_720 ();
 sg13g2_fill_1 FILLER_42_726 ();
 sg13g2_fill_1 FILLER_42_747 ();
 sg13g2_fill_1 FILLER_42_758 ();
 sg13g2_fill_2 FILLER_42_809 ();
 sg13g2_fill_1 FILLER_42_815 ();
 sg13g2_fill_2 FILLER_43_54 ();
 sg13g2_fill_1 FILLER_43_60 ();
 sg13g2_fill_1 FILLER_43_82 ();
 sg13g2_fill_2 FILLER_43_134 ();
 sg13g2_fill_2 FILLER_43_146 ();
 sg13g2_fill_1 FILLER_43_148 ();
 sg13g2_fill_1 FILLER_43_155 ();
 sg13g2_fill_1 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_167 ();
 sg13g2_fill_1 FILLER_43_174 ();
 sg13g2_fill_2 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_187 ();
 sg13g2_fill_2 FILLER_43_193 ();
 sg13g2_fill_2 FILLER_43_200 ();
 sg13g2_fill_1 FILLER_43_231 ();
 sg13g2_fill_1 FILLER_43_236 ();
 sg13g2_fill_1 FILLER_43_242 ();
 sg13g2_fill_1 FILLER_43_248 ();
 sg13g2_fill_2 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_290 ();
 sg13g2_fill_2 FILLER_43_297 ();
 sg13g2_fill_2 FILLER_43_309 ();
 sg13g2_fill_1 FILLER_43_316 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_fill_1 FILLER_43_333 ();
 sg13g2_fill_1 FILLER_43_339 ();
 sg13g2_fill_2 FILLER_43_345 ();
 sg13g2_fill_1 FILLER_43_360 ();
 sg13g2_fill_2 FILLER_43_369 ();
 sg13g2_fill_1 FILLER_43_371 ();
 sg13g2_fill_2 FILLER_43_377 ();
 sg13g2_fill_1 FILLER_43_392 ();
 sg13g2_fill_1 FILLER_43_398 ();
 sg13g2_fill_2 FILLER_43_403 ();
 sg13g2_decap_8 FILLER_43_417 ();
 sg13g2_decap_8 FILLER_43_424 ();
 sg13g2_fill_2 FILLER_43_431 ();
 sg13g2_fill_2 FILLER_43_438 ();
 sg13g2_fill_1 FILLER_43_440 ();
 sg13g2_decap_8 FILLER_43_445 ();
 sg13g2_decap_8 FILLER_43_452 ();
 sg13g2_fill_2 FILLER_43_459 ();
 sg13g2_fill_1 FILLER_43_476 ();
 sg13g2_fill_1 FILLER_43_487 ();
 sg13g2_fill_2 FILLER_43_507 ();
 sg13g2_fill_1 FILLER_43_509 ();
 sg13g2_fill_2 FILLER_43_519 ();
 sg13g2_fill_1 FILLER_43_521 ();
 sg13g2_fill_2 FILLER_43_531 ();
 sg13g2_fill_1 FILLER_43_546 ();
 sg13g2_fill_2 FILLER_43_553 ();
 sg13g2_fill_2 FILLER_43_601 ();
 sg13g2_fill_1 FILLER_43_603 ();
 sg13g2_fill_2 FILLER_43_616 ();
 sg13g2_fill_1 FILLER_43_623 ();
 sg13g2_fill_2 FILLER_43_650 ();
 sg13g2_fill_2 FILLER_43_678 ();
 sg13g2_fill_1 FILLER_43_680 ();
 sg13g2_fill_1 FILLER_43_783 ();
 sg13g2_fill_2 FILLER_43_830 ();
 sg13g2_decap_4 FILLER_43_872 ();
 sg13g2_fill_2 FILLER_43_876 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_27 ();
 sg13g2_fill_1 FILLER_44_45 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_fill_1 FILLER_44_119 ();
 sg13g2_fill_1 FILLER_44_140 ();
 sg13g2_fill_2 FILLER_44_155 ();
 sg13g2_fill_1 FILLER_44_157 ();
 sg13g2_fill_1 FILLER_44_174 ();
 sg13g2_fill_2 FILLER_44_241 ();
 sg13g2_fill_2 FILLER_44_289 ();
 sg13g2_fill_1 FILLER_44_295 ();
 sg13g2_fill_2 FILLER_44_369 ();
 sg13g2_fill_1 FILLER_44_371 ();
 sg13g2_decap_4 FILLER_44_398 ();
 sg13g2_fill_1 FILLER_44_463 ();
 sg13g2_fill_2 FILLER_44_507 ();
 sg13g2_fill_1 FILLER_44_601 ();
 sg13g2_fill_2 FILLER_44_636 ();
 sg13g2_fill_1 FILLER_44_642 ();
 sg13g2_fill_1 FILLER_44_657 ();
 sg13g2_fill_1 FILLER_44_662 ();
 sg13g2_fill_2 FILLER_44_688 ();
 sg13g2_fill_1 FILLER_44_690 ();
 sg13g2_fill_2 FILLER_44_704 ();
 sg13g2_fill_2 FILLER_44_716 ();
 sg13g2_fill_2 FILLER_44_732 ();
 sg13g2_fill_1 FILLER_44_734 ();
 sg13g2_fill_1 FILLER_44_753 ();
 sg13g2_fill_2 FILLER_44_780 ();
 sg13g2_fill_2 FILLER_44_792 ();
 sg13g2_fill_1 FILLER_44_794 ();
 sg13g2_fill_1 FILLER_44_805 ();
 sg13g2_fill_2 FILLER_44_810 ();
 sg13g2_fill_1 FILLER_44_812 ();
 sg13g2_fill_2 FILLER_44_849 ();
 sg13g2_fill_1 FILLER_44_851 ();
 sg13g2_fill_2 FILLER_45_34 ();
 sg13g2_fill_1 FILLER_45_87 ();
 sg13g2_fill_2 FILLER_45_134 ();
 sg13g2_fill_2 FILLER_45_146 ();
 sg13g2_fill_1 FILLER_45_192 ();
 sg13g2_fill_1 FILLER_45_198 ();
 sg13g2_fill_2 FILLER_45_228 ();
 sg13g2_fill_2 FILLER_45_235 ();
 sg13g2_fill_2 FILLER_45_317 ();
 sg13g2_fill_1 FILLER_45_319 ();
 sg13g2_fill_2 FILLER_45_396 ();
 sg13g2_fill_2 FILLER_45_402 ();
 sg13g2_fill_1 FILLER_45_404 ();
 sg13g2_fill_2 FILLER_45_440 ();
 sg13g2_fill_2 FILLER_45_446 ();
 sg13g2_fill_1 FILLER_45_448 ();
 sg13g2_decap_4 FILLER_45_453 ();
 sg13g2_decap_4 FILLER_45_466 ();
 sg13g2_fill_1 FILLER_45_470 ();
 sg13g2_fill_1 FILLER_45_503 ();
 sg13g2_fill_2 FILLER_45_547 ();
 sg13g2_fill_1 FILLER_45_577 ();
 sg13g2_fill_1 FILLER_45_582 ();
 sg13g2_fill_1 FILLER_45_587 ();
 sg13g2_fill_1 FILLER_45_630 ();
 sg13g2_decap_4 FILLER_45_635 ();
 sg13g2_fill_1 FILLER_45_644 ();
 sg13g2_fill_1 FILLER_45_689 ();
 sg13g2_fill_2 FILLER_45_702 ();
 sg13g2_fill_2 FILLER_45_712 ();
 sg13g2_fill_2 FILLER_45_725 ();
 sg13g2_fill_1 FILLER_45_727 ();
 sg13g2_fill_2 FILLER_45_741 ();
 sg13g2_fill_1 FILLER_45_753 ();
 sg13g2_fill_2 FILLER_45_768 ();
 sg13g2_fill_1 FILLER_45_770 ();
 sg13g2_fill_2 FILLER_45_791 ();
 sg13g2_fill_2 FILLER_45_839 ();
 sg13g2_fill_1 FILLER_45_841 ();
 sg13g2_fill_1 FILLER_46_50 ();
 sg13g2_fill_1 FILLER_46_77 ();
 sg13g2_fill_1 FILLER_46_119 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_150 ();
 sg13g2_fill_1 FILLER_46_168 ();
 sg13g2_fill_1 FILLER_46_177 ();
 sg13g2_fill_1 FILLER_46_187 ();
 sg13g2_fill_2 FILLER_46_228 ();
 sg13g2_fill_2 FILLER_46_269 ();
 sg13g2_fill_2 FILLER_46_280 ();
 sg13g2_fill_2 FILLER_46_291 ();
 sg13g2_fill_1 FILLER_46_312 ();
 sg13g2_fill_2 FILLER_46_366 ();
 sg13g2_fill_1 FILLER_46_368 ();
 sg13g2_fill_1 FILLER_46_379 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_2 FILLER_46_434 ();
 sg13g2_fill_1 FILLER_46_436 ();
 sg13g2_fill_2 FILLER_46_442 ();
 sg13g2_fill_1 FILLER_46_444 ();
 sg13g2_fill_2 FILLER_46_450 ();
 sg13g2_fill_1 FILLER_46_460 ();
 sg13g2_decap_8 FILLER_46_465 ();
 sg13g2_fill_2 FILLER_46_485 ();
 sg13g2_fill_1 FILLER_46_496 ();
 sg13g2_fill_2 FILLER_46_566 ();
 sg13g2_fill_1 FILLER_46_642 ();
 sg13g2_fill_2 FILLER_46_652 ();
 sg13g2_fill_1 FILLER_46_662 ();
 sg13g2_fill_2 FILLER_46_667 ();
 sg13g2_fill_2 FILLER_46_682 ();
 sg13g2_fill_1 FILLER_46_684 ();
 sg13g2_fill_2 FILLER_46_705 ();
 sg13g2_fill_1 FILLER_46_747 ();
 sg13g2_fill_1 FILLER_46_778 ();
 sg13g2_fill_1 FILLER_46_805 ();
 sg13g2_fill_2 FILLER_46_816 ();
 sg13g2_fill_1 FILLER_46_828 ();
 sg13g2_fill_1 FILLER_46_833 ();
 sg13g2_fill_2 FILLER_46_864 ();
 sg13g2_fill_1 FILLER_46_866 ();
 sg13g2_decap_8 FILLER_46_871 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_38 ();
 sg13g2_fill_1 FILLER_47_111 ();
 sg13g2_fill_2 FILLER_47_126 ();
 sg13g2_fill_1 FILLER_47_128 ();
 sg13g2_fill_2 FILLER_47_151 ();
 sg13g2_fill_1 FILLER_47_153 ();
 sg13g2_fill_1 FILLER_47_235 ();
 sg13g2_fill_1 FILLER_47_251 ();
 sg13g2_fill_2 FILLER_47_352 ();
 sg13g2_fill_1 FILLER_47_354 ();
 sg13g2_fill_1 FILLER_47_370 ();
 sg13g2_fill_2 FILLER_47_381 ();
 sg13g2_fill_1 FILLER_47_383 ();
 sg13g2_fill_1 FILLER_47_397 ();
 sg13g2_fill_2 FILLER_47_403 ();
 sg13g2_fill_2 FILLER_47_417 ();
 sg13g2_fill_1 FILLER_47_440 ();
 sg13g2_fill_1 FILLER_47_446 ();
 sg13g2_fill_2 FILLER_47_452 ();
 sg13g2_fill_1 FILLER_47_488 ();
 sg13g2_fill_2 FILLER_47_515 ();
 sg13g2_fill_1 FILLER_47_529 ();
 sg13g2_fill_2 FILLER_47_534 ();
 sg13g2_fill_2 FILLER_47_570 ();
 sg13g2_fill_2 FILLER_47_672 ();
 sg13g2_fill_2 FILLER_47_679 ();
 sg13g2_fill_2 FILLER_47_718 ();
 sg13g2_fill_2 FILLER_47_753 ();
 sg13g2_fill_1 FILLER_47_755 ();
 sg13g2_fill_2 FILLER_47_790 ();
 sg13g2_fill_1 FILLER_47_792 ();
 sg13g2_fill_1 FILLER_47_803 ();
 sg13g2_fill_2 FILLER_47_830 ();
 sg13g2_fill_1 FILLER_47_832 ();
 sg13g2_decap_8 FILLER_47_859 ();
 sg13g2_decap_8 FILLER_47_866 ();
 sg13g2_decap_4 FILLER_47_873 ();
 sg13g2_fill_1 FILLER_47_877 ();
 sg13g2_fill_1 FILLER_48_34 ();
 sg13g2_fill_1 FILLER_48_45 ();
 sg13g2_fill_1 FILLER_48_119 ();
 sg13g2_fill_2 FILLER_48_148 ();
 sg13g2_fill_2 FILLER_48_155 ();
 sg13g2_fill_1 FILLER_48_220 ();
 sg13g2_fill_2 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_307 ();
 sg13g2_fill_1 FILLER_48_424 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_fill_2 FILLER_48_490 ();
 sg13g2_fill_2 FILLER_48_590 ();
 sg13g2_fill_2 FILLER_48_651 ();
 sg13g2_fill_2 FILLER_48_711 ();
 sg13g2_fill_1 FILLER_48_713 ();
 sg13g2_fill_2 FILLER_48_823 ();
 sg13g2_fill_1 FILLER_48_825 ();
 sg13g2_decap_8 FILLER_48_848 ();
 sg13g2_decap_8 FILLER_48_855 ();
 sg13g2_decap_8 FILLER_48_862 ();
 sg13g2_decap_8 FILLER_48_869 ();
 sg13g2_fill_2 FILLER_48_876 ();
 sg13g2_fill_1 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_76 ();
 sg13g2_fill_1 FILLER_49_123 ();
 sg13g2_fill_1 FILLER_49_129 ();
 sg13g2_fill_1 FILLER_49_187 ();
 sg13g2_fill_1 FILLER_49_193 ();
 sg13g2_fill_2 FILLER_49_225 ();
 sg13g2_fill_2 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_1 FILLER_49_341 ();
 sg13g2_fill_2 FILLER_49_378 ();
 sg13g2_fill_1 FILLER_49_380 ();
 sg13g2_fill_1 FILLER_49_393 ();
 sg13g2_fill_1 FILLER_49_398 ();
 sg13g2_fill_1 FILLER_49_403 ();
 sg13g2_fill_1 FILLER_49_409 ();
 sg13g2_fill_1 FILLER_49_423 ();
 sg13g2_fill_2 FILLER_49_432 ();
 sg13g2_fill_1 FILLER_49_461 ();
 sg13g2_fill_1 FILLER_49_472 ();
 sg13g2_fill_1 FILLER_49_486 ();
 sg13g2_fill_1 FILLER_49_495 ();
 sg13g2_fill_2 FILLER_49_504 ();
 sg13g2_fill_2 FILLER_49_522 ();
 sg13g2_fill_1 FILLER_49_524 ();
 sg13g2_fill_1 FILLER_49_623 ();
 sg13g2_fill_2 FILLER_49_664 ();
 sg13g2_decap_8 FILLER_49_671 ();
 sg13g2_fill_2 FILLER_49_706 ();
 sg13g2_fill_1 FILLER_49_724 ();
 sg13g2_fill_1 FILLER_49_735 ();
 sg13g2_fill_2 FILLER_49_757 ();
 sg13g2_fill_2 FILLER_49_803 ();
 sg13g2_decap_8 FILLER_49_839 ();
 sg13g2_decap_8 FILLER_49_846 ();
 sg13g2_decap_8 FILLER_49_853 ();
 sg13g2_decap_8 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_49_867 ();
 sg13g2_decap_4 FILLER_49_874 ();
 sg13g2_fill_2 FILLER_50_119 ();
 sg13g2_fill_2 FILLER_50_131 ();
 sg13g2_fill_2 FILLER_50_141 ();
 sg13g2_fill_1 FILLER_50_143 ();
 sg13g2_fill_2 FILLER_50_186 ();
 sg13g2_fill_1 FILLER_50_193 ();
 sg13g2_fill_1 FILLER_50_204 ();
 sg13g2_fill_1 FILLER_50_209 ();
 sg13g2_fill_1 FILLER_50_235 ();
 sg13g2_fill_1 FILLER_50_241 ();
 sg13g2_fill_1 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_403 ();
 sg13g2_fill_2 FILLER_50_438 ();
 sg13g2_fill_2 FILLER_50_530 ();
 sg13g2_fill_1 FILLER_50_563 ();
 sg13g2_fill_1 FILLER_50_670 ();
 sg13g2_fill_2 FILLER_50_675 ();
 sg13g2_fill_1 FILLER_50_677 ();
 sg13g2_fill_2 FILLER_50_687 ();
 sg13g2_fill_1 FILLER_50_689 ();
 sg13g2_fill_1 FILLER_50_708 ();
 sg13g2_fill_2 FILLER_50_729 ();
 sg13g2_fill_1 FILLER_50_731 ();
 sg13g2_fill_2 FILLER_50_757 ();
 sg13g2_fill_2 FILLER_50_773 ();
 sg13g2_decap_8 FILLER_50_843 ();
 sg13g2_decap_8 FILLER_50_850 ();
 sg13g2_decap_8 FILLER_50_857 ();
 sg13g2_decap_8 FILLER_50_864 ();
 sg13g2_decap_8 FILLER_50_871 ();
 sg13g2_fill_1 FILLER_51_79 ();
 sg13g2_fill_2 FILLER_51_92 ();
 sg13g2_fill_1 FILLER_51_94 ();
 sg13g2_fill_2 FILLER_51_128 ();
 sg13g2_fill_1 FILLER_51_140 ();
 sg13g2_fill_1 FILLER_51_167 ();
 sg13g2_fill_1 FILLER_51_194 ();
 sg13g2_fill_1 FILLER_51_213 ();
 sg13g2_fill_1 FILLER_51_244 ();
 sg13g2_fill_1 FILLER_51_271 ();
 sg13g2_fill_2 FILLER_51_308 ();
 sg13g2_fill_1 FILLER_51_320 ();
 sg13g2_fill_1 FILLER_51_347 ();
 sg13g2_fill_1 FILLER_51_353 ();
 sg13g2_fill_2 FILLER_51_371 ();
 sg13g2_fill_2 FILLER_51_382 ();
 sg13g2_fill_2 FILLER_51_444 ();
 sg13g2_fill_2 FILLER_51_464 ();
 sg13g2_fill_1 FILLER_51_473 ();
 sg13g2_fill_1 FILLER_51_484 ();
 sg13g2_fill_1 FILLER_51_493 ();
 sg13g2_fill_2 FILLER_51_498 ();
 sg13g2_fill_1 FILLER_51_500 ();
 sg13g2_fill_1 FILLER_51_531 ();
 sg13g2_fill_1 FILLER_51_542 ();
 sg13g2_fill_1 FILLER_51_565 ();
 sg13g2_fill_2 FILLER_51_576 ();
 sg13g2_fill_1 FILLER_51_604 ();
 sg13g2_fill_1 FILLER_51_657 ();
 sg13g2_decap_4 FILLER_51_674 ();
 sg13g2_fill_2 FILLER_51_768 ();
 sg13g2_fill_1 FILLER_51_779 ();
 sg13g2_fill_1 FILLER_51_806 ();
 sg13g2_fill_1 FILLER_51_817 ();
 sg13g2_decap_8 FILLER_51_854 ();
 sg13g2_decap_8 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_51_868 ();
 sg13g2_fill_2 FILLER_51_875 ();
 sg13g2_fill_1 FILLER_51_877 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_2 FILLER_52_52 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_2 FILLER_52_111 ();
 sg13g2_fill_1 FILLER_52_206 ();
 sg13g2_fill_1 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_243 ();
 sg13g2_fill_1 FILLER_52_271 ();
 sg13g2_fill_1 FILLER_52_277 ();
 sg13g2_fill_1 FILLER_52_282 ();
 sg13g2_fill_2 FILLER_52_288 ();
 sg13g2_fill_1 FILLER_52_423 ();
 sg13g2_fill_1 FILLER_52_428 ();
 sg13g2_fill_1 FILLER_52_437 ();
 sg13g2_fill_1 FILLER_52_442 ();
 sg13g2_fill_2 FILLER_52_447 ();
 sg13g2_fill_1 FILLER_52_455 ();
 sg13g2_fill_1 FILLER_52_489 ();
 sg13g2_fill_1 FILLER_52_495 ();
 sg13g2_fill_1 FILLER_52_501 ();
 sg13g2_fill_1 FILLER_52_506 ();
 sg13g2_decap_4 FILLER_52_516 ();
 sg13g2_fill_1 FILLER_52_530 ();
 sg13g2_fill_1 FILLER_52_536 ();
 sg13g2_fill_1 FILLER_52_542 ();
 sg13g2_fill_1 FILLER_52_562 ();
 sg13g2_fill_1 FILLER_52_576 ();
 sg13g2_fill_2 FILLER_52_633 ();
 sg13g2_fill_2 FILLER_52_643 ();
 sg13g2_decap_4 FILLER_52_677 ();
 sg13g2_decap_4 FILLER_52_685 ();
 sg13g2_fill_1 FILLER_52_707 ();
 sg13g2_fill_2 FILLER_52_713 ();
 sg13g2_fill_1 FILLER_52_724 ();
 sg13g2_fill_1 FILLER_52_730 ();
 sg13g2_fill_1 FILLER_52_735 ();
 sg13g2_fill_1 FILLER_52_743 ();
 sg13g2_fill_2 FILLER_52_753 ();
 sg13g2_fill_1 FILLER_52_755 ();
 sg13g2_fill_2 FILLER_52_798 ();
 sg13g2_fill_1 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_850 ();
 sg13g2_decap_8 FILLER_52_857 ();
 sg13g2_decap_8 FILLER_52_864 ();
 sg13g2_decap_8 FILLER_52_871 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_27 ();
 sg13g2_fill_1 FILLER_53_34 ();
 sg13g2_fill_2 FILLER_53_53 ();
 sg13g2_fill_1 FILLER_53_133 ();
 sg13g2_fill_1 FILLER_53_176 ();
 sg13g2_fill_1 FILLER_53_190 ();
 sg13g2_fill_2 FILLER_53_196 ();
 sg13g2_fill_1 FILLER_53_229 ();
 sg13g2_fill_2 FILLER_53_239 ();
 sg13g2_fill_1 FILLER_53_241 ();
 sg13g2_fill_1 FILLER_53_246 ();
 sg13g2_fill_1 FILLER_53_287 ();
 sg13g2_fill_1 FILLER_53_328 ();
 sg13g2_decap_4 FILLER_53_400 ();
 sg13g2_fill_1 FILLER_53_404 ();
 sg13g2_fill_2 FILLER_53_412 ();
 sg13g2_fill_1 FILLER_53_419 ();
 sg13g2_fill_1 FILLER_53_459 ();
 sg13g2_fill_2 FILLER_53_465 ();
 sg13g2_fill_2 FILLER_53_475 ();
 sg13g2_fill_2 FILLER_53_483 ();
 sg13g2_fill_1 FILLER_53_485 ();
 sg13g2_decap_4 FILLER_53_501 ();
 sg13g2_fill_1 FILLER_53_536 ();
 sg13g2_fill_2 FILLER_53_610 ();
 sg13g2_fill_1 FILLER_53_612 ();
 sg13g2_decap_4 FILLER_53_691 ();
 sg13g2_fill_1 FILLER_53_695 ();
 sg13g2_fill_2 FILLER_53_704 ();
 sg13g2_fill_1 FILLER_53_724 ();
 sg13g2_fill_1 FILLER_53_730 ();
 sg13g2_fill_1 FILLER_53_735 ();
 sg13g2_fill_2 FILLER_53_745 ();
 sg13g2_fill_1 FILLER_53_747 ();
 sg13g2_fill_1 FILLER_53_756 ();
 sg13g2_fill_1 FILLER_53_781 ();
 sg13g2_fill_2 FILLER_53_826 ();
 sg13g2_decap_8 FILLER_53_854 ();
 sg13g2_decap_8 FILLER_53_861 ();
 sg13g2_decap_8 FILLER_53_868 ();
 sg13g2_fill_2 FILLER_53_875 ();
 sg13g2_fill_1 FILLER_53_877 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_27 ();
 sg13g2_fill_1 FILLER_54_37 ();
 sg13g2_fill_1 FILLER_54_48 ();
 sg13g2_fill_2 FILLER_54_93 ();
 sg13g2_fill_1 FILLER_54_151 ();
 sg13g2_fill_2 FILLER_54_256 ();
 sg13g2_fill_2 FILLER_54_263 ();
 sg13g2_fill_1 FILLER_54_265 ();
 sg13g2_fill_1 FILLER_54_306 ();
 sg13g2_fill_2 FILLER_54_350 ();
 sg13g2_fill_1 FILLER_54_373 ();
 sg13g2_fill_1 FILLER_54_392 ();
 sg13g2_fill_1 FILLER_54_404 ();
 sg13g2_fill_2 FILLER_54_463 ();
 sg13g2_decap_4 FILLER_54_471 ();
 sg13g2_fill_2 FILLER_54_475 ();
 sg13g2_fill_1 FILLER_54_501 ();
 sg13g2_fill_1 FILLER_54_512 ();
 sg13g2_fill_1 FILLER_54_522 ();
 sg13g2_fill_1 FILLER_54_565 ();
 sg13g2_fill_1 FILLER_54_612 ();
 sg13g2_fill_1 FILLER_54_630 ();
 sg13g2_fill_1 FILLER_54_635 ();
 sg13g2_fill_1 FILLER_54_640 ();
 sg13g2_fill_2 FILLER_54_646 ();
 sg13g2_fill_1 FILLER_54_698 ();
 sg13g2_fill_1 FILLER_54_789 ();
 sg13g2_decap_8 FILLER_54_850 ();
 sg13g2_decap_8 FILLER_54_857 ();
 sg13g2_decap_8 FILLER_54_864 ();
 sg13g2_decap_8 FILLER_54_871 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_6 ();
 sg13g2_fill_2 FILLER_55_38 ();
 sg13g2_fill_2 FILLER_55_86 ();
 sg13g2_fill_1 FILLER_55_122 ();
 sg13g2_fill_1 FILLER_55_133 ();
 sg13g2_fill_2 FILLER_55_168 ();
 sg13g2_fill_1 FILLER_55_170 ();
 sg13g2_fill_2 FILLER_55_195 ();
 sg13g2_fill_2 FILLER_55_319 ();
 sg13g2_fill_2 FILLER_55_365 ();
 sg13g2_decap_4 FILLER_55_428 ();
 sg13g2_fill_2 FILLER_55_432 ();
 sg13g2_fill_1 FILLER_55_479 ();
 sg13g2_fill_1 FILLER_55_490 ();
 sg13g2_fill_2 FILLER_55_511 ();
 sg13g2_fill_1 FILLER_55_518 ();
 sg13g2_fill_1 FILLER_55_575 ();
 sg13g2_fill_2 FILLER_55_593 ();
 sg13g2_fill_1 FILLER_55_595 ();
 sg13g2_fill_2 FILLER_55_605 ();
 sg13g2_fill_1 FILLER_55_613 ();
 sg13g2_fill_1 FILLER_55_626 ();
 sg13g2_fill_2 FILLER_55_672 ();
 sg13g2_fill_2 FILLER_55_679 ();
 sg13g2_fill_1 FILLER_55_685 ();
 sg13g2_fill_1 FILLER_55_691 ();
 sg13g2_fill_1 FILLER_55_700 ();
 sg13g2_fill_2 FILLER_55_706 ();
 sg13g2_fill_1 FILLER_55_725 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_fill_1 FILLER_55_746 ();
 sg13g2_fill_2 FILLER_55_800 ();
 sg13g2_fill_2 FILLER_55_838 ();
 sg13g2_decap_8 FILLER_55_844 ();
 sg13g2_decap_8 FILLER_55_851 ();
 sg13g2_decap_8 FILLER_55_858 ();
 sg13g2_decap_8 FILLER_55_865 ();
 sg13g2_decap_4 FILLER_55_872 ();
 sg13g2_fill_2 FILLER_55_876 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_22 ();
 sg13g2_fill_1 FILLER_56_24 ();
 sg13g2_fill_2 FILLER_56_39 ();
 sg13g2_fill_1 FILLER_56_55 ();
 sg13g2_fill_2 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_76 ();
 sg13g2_fill_2 FILLER_56_82 ();
 sg13g2_fill_1 FILLER_56_113 ();
 sg13g2_fill_1 FILLER_56_190 ();
 sg13g2_fill_1 FILLER_56_209 ();
 sg13g2_fill_2 FILLER_56_290 ();
 sg13g2_fill_1 FILLER_56_292 ();
 sg13g2_fill_1 FILLER_56_323 ();
 sg13g2_fill_2 FILLER_56_360 ();
 sg13g2_fill_1 FILLER_56_367 ();
 sg13g2_fill_1 FILLER_56_398 ();
 sg13g2_fill_2 FILLER_56_403 ();
 sg13g2_fill_1 FILLER_56_418 ();
 sg13g2_fill_1 FILLER_56_445 ();
 sg13g2_fill_1 FILLER_56_454 ();
 sg13g2_fill_1 FILLER_56_460 ();
 sg13g2_fill_1 FILLER_56_477 ();
 sg13g2_fill_2 FILLER_56_493 ();
 sg13g2_fill_1 FILLER_56_575 ();
 sg13g2_fill_1 FILLER_56_580 ();
 sg13g2_fill_1 FILLER_56_590 ();
 sg13g2_fill_1 FILLER_56_596 ();
 sg13g2_fill_1 FILLER_56_614 ();
 sg13g2_fill_1 FILLER_56_620 ();
 sg13g2_fill_1 FILLER_56_627 ();
 sg13g2_fill_1 FILLER_56_632 ();
 sg13g2_fill_2 FILLER_56_638 ();
 sg13g2_fill_1 FILLER_56_718 ();
 sg13g2_fill_2 FILLER_56_752 ();
 sg13g2_fill_2 FILLER_56_787 ();
 sg13g2_fill_2 FILLER_56_795 ();
 sg13g2_fill_1 FILLER_56_813 ();
 sg13g2_fill_2 FILLER_56_857 ();
 sg13g2_decap_8 FILLER_56_863 ();
 sg13g2_decap_8 FILLER_56_870 ();
 sg13g2_fill_1 FILLER_56_877 ();
 sg13g2_fill_2 FILLER_57_44 ();
 sg13g2_fill_2 FILLER_57_106 ();
 sg13g2_fill_1 FILLER_57_130 ();
 sg13g2_fill_2 FILLER_57_165 ();
 sg13g2_fill_1 FILLER_57_240 ();
 sg13g2_fill_1 FILLER_57_245 ();
 sg13g2_fill_1 FILLER_57_255 ();
 sg13g2_fill_2 FILLER_57_260 ();
 sg13g2_fill_2 FILLER_57_315 ();
 sg13g2_fill_1 FILLER_57_317 ();
 sg13g2_fill_1 FILLER_57_339 ();
 sg13g2_fill_1 FILLER_57_345 ();
 sg13g2_fill_1 FILLER_57_351 ();
 sg13g2_fill_1 FILLER_57_361 ();
 sg13g2_fill_1 FILLER_57_424 ();
 sg13g2_fill_2 FILLER_57_452 ();
 sg13g2_fill_2 FILLER_57_642 ();
 sg13g2_fill_2 FILLER_57_656 ();
 sg13g2_fill_2 FILLER_57_680 ();
 sg13g2_fill_1 FILLER_57_687 ();
 sg13g2_fill_2 FILLER_57_693 ();
 sg13g2_fill_1 FILLER_57_695 ();
 sg13g2_fill_2 FILLER_57_726 ();
 sg13g2_fill_1 FILLER_57_736 ();
 sg13g2_fill_1 FILLER_57_745 ();
 sg13g2_fill_2 FILLER_57_824 ();
 sg13g2_fill_2 FILLER_57_876 ();
 sg13g2_fill_2 FILLER_58_4 ();
 sg13g2_fill_1 FILLER_58_6 ();
 sg13g2_fill_1 FILLER_58_57 ();
 sg13g2_fill_2 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_103 ();
 sg13g2_fill_2 FILLER_58_270 ();
 sg13g2_fill_2 FILLER_58_302 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_1 FILLER_58_383 ();
 sg13g2_fill_2 FILLER_58_448 ();
 sg13g2_fill_1 FILLER_58_455 ();
 sg13g2_fill_2 FILLER_58_460 ();
 sg13g2_fill_2 FILLER_58_470 ();
 sg13g2_fill_1 FILLER_58_472 ();
 sg13g2_fill_1 FILLER_58_481 ();
 sg13g2_fill_1 FILLER_58_518 ();
 sg13g2_fill_2 FILLER_58_600 ();
 sg13g2_fill_2 FILLER_58_655 ();
 sg13g2_fill_2 FILLER_58_665 ();
 sg13g2_fill_1 FILLER_58_667 ();
 sg13g2_fill_2 FILLER_58_677 ();
 sg13g2_fill_1 FILLER_58_679 ();
 sg13g2_decap_4 FILLER_58_710 ();
 sg13g2_fill_2 FILLER_58_714 ();
 sg13g2_fill_2 FILLER_58_736 ();
 sg13g2_fill_1 FILLER_58_738 ();
 sg13g2_fill_1 FILLER_58_797 ();
 sg13g2_fill_1 FILLER_58_840 ();
 sg13g2_fill_1 FILLER_58_877 ();
 sg13g2_fill_2 FILLER_59_44 ();
 sg13g2_fill_1 FILLER_59_61 ();
 sg13g2_fill_2 FILLER_59_121 ();
 sg13g2_fill_1 FILLER_59_123 ();
 sg13g2_fill_1 FILLER_59_137 ();
 sg13g2_fill_1 FILLER_59_148 ();
 sg13g2_fill_1 FILLER_59_187 ();
 sg13g2_fill_1 FILLER_59_201 ();
 sg13g2_fill_2 FILLER_59_211 ();
 sg13g2_fill_1 FILLER_59_222 ();
 sg13g2_fill_1 FILLER_59_227 ();
 sg13g2_fill_1 FILLER_59_246 ();
 sg13g2_fill_1 FILLER_59_287 ();
 sg13g2_fill_2 FILLER_59_380 ();
 sg13g2_fill_2 FILLER_59_421 ();
 sg13g2_fill_2 FILLER_59_485 ();
 sg13g2_fill_1 FILLER_59_487 ();
 sg13g2_fill_2 FILLER_59_531 ();
 sg13g2_fill_2 FILLER_59_548 ();
 sg13g2_fill_1 FILLER_59_560 ();
 sg13g2_fill_1 FILLER_59_566 ();
 sg13g2_fill_1 FILLER_59_575 ();
 sg13g2_fill_1 FILLER_59_581 ();
 sg13g2_fill_1 FILLER_59_638 ();
 sg13g2_fill_2 FILLER_59_648 ();
 sg13g2_fill_1 FILLER_59_690 ();
 sg13g2_fill_1 FILLER_59_701 ();
 sg13g2_fill_1 FILLER_59_780 ();
 sg13g2_fill_2 FILLER_59_790 ();
 sg13g2_fill_2 FILLER_60_26 ();
 sg13g2_fill_1 FILLER_60_28 ();
 sg13g2_fill_1 FILLER_60_55 ();
 sg13g2_fill_1 FILLER_60_141 ();
 sg13g2_fill_1 FILLER_60_209 ();
 sg13g2_fill_2 FILLER_60_219 ();
 sg13g2_fill_2 FILLER_60_234 ();
 sg13g2_fill_1 FILLER_60_236 ();
 sg13g2_fill_1 FILLER_60_254 ();
 sg13g2_fill_2 FILLER_60_347 ();
 sg13g2_fill_1 FILLER_60_366 ();
 sg13g2_fill_1 FILLER_60_372 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_fill_1 FILLER_60_414 ();
 sg13g2_fill_1 FILLER_60_420 ();
 sg13g2_decap_4 FILLER_60_468 ();
 sg13g2_fill_2 FILLER_60_472 ();
 sg13g2_fill_2 FILLER_60_512 ();
 sg13g2_fill_2 FILLER_60_595 ();
 sg13g2_fill_2 FILLER_60_606 ();
 sg13g2_fill_1 FILLER_60_608 ();
 sg13g2_fill_1 FILLER_60_614 ();
 sg13g2_fill_1 FILLER_60_623 ();
 sg13g2_fill_2 FILLER_60_629 ();
 sg13g2_fill_1 FILLER_60_680 ();
 sg13g2_fill_2 FILLER_60_685 ();
 sg13g2_fill_1 FILLER_60_695 ();
 sg13g2_fill_1 FILLER_60_706 ();
 sg13g2_fill_2 FILLER_60_717 ();
 sg13g2_fill_2 FILLER_60_731 ();
 sg13g2_fill_1 FILLER_60_790 ();
 sg13g2_fill_1 FILLER_60_799 ();
 sg13g2_fill_1 FILLER_60_826 ();
 sg13g2_fill_1 FILLER_60_865 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_11 ();
 sg13g2_fill_1 FILLER_61_23 ();
 sg13g2_fill_1 FILLER_61_177 ();
 sg13g2_fill_2 FILLER_61_229 ();
 sg13g2_fill_1 FILLER_61_251 ();
 sg13g2_fill_1 FILLER_61_261 ();
 sg13g2_fill_2 FILLER_61_271 ();
 sg13g2_fill_1 FILLER_61_273 ();
 sg13g2_fill_1 FILLER_61_299 ();
 sg13g2_fill_1 FILLER_61_343 ();
 sg13g2_fill_2 FILLER_61_350 ();
 sg13g2_fill_1 FILLER_61_357 ();
 sg13g2_fill_1 FILLER_61_372 ();
 sg13g2_fill_1 FILLER_61_378 ();
 sg13g2_fill_1 FILLER_61_389 ();
 sg13g2_fill_1 FILLER_61_479 ();
 sg13g2_fill_1 FILLER_61_511 ();
 sg13g2_fill_2 FILLER_61_522 ();
 sg13g2_fill_2 FILLER_61_571 ();
 sg13g2_fill_1 FILLER_61_573 ();
 sg13g2_fill_2 FILLER_61_601 ();
 sg13g2_fill_2 FILLER_61_616 ();
 sg13g2_fill_2 FILLER_61_627 ();
 sg13g2_fill_1 FILLER_61_634 ();
 sg13g2_fill_2 FILLER_61_664 ();
 sg13g2_fill_2 FILLER_61_678 ();
 sg13g2_fill_1 FILLER_61_680 ();
 sg13g2_fill_2 FILLER_61_711 ();
 sg13g2_fill_2 FILLER_61_744 ();
 sg13g2_fill_2 FILLER_61_787 ();
 sg13g2_fill_2 FILLER_61_829 ();
 sg13g2_fill_2 FILLER_61_843 ();
 sg13g2_fill_1 FILLER_61_845 ();
 sg13g2_fill_1 FILLER_61_877 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_13 ();
 sg13g2_fill_1 FILLER_62_56 ();
 sg13g2_fill_1 FILLER_62_62 ();
 sg13g2_fill_1 FILLER_62_112 ();
 sg13g2_fill_1 FILLER_62_123 ();
 sg13g2_fill_1 FILLER_62_137 ();
 sg13g2_fill_2 FILLER_62_143 ();
 sg13g2_fill_2 FILLER_62_201 ();
 sg13g2_fill_2 FILLER_62_278 ();
 sg13g2_fill_1 FILLER_62_280 ();
 sg13g2_fill_2 FILLER_62_332 ();
 sg13g2_fill_1 FILLER_62_340 ();
 sg13g2_fill_1 FILLER_62_347 ();
 sg13g2_fill_2 FILLER_62_368 ();
 sg13g2_fill_1 FILLER_62_435 ();
 sg13g2_fill_1 FILLER_62_441 ();
 sg13g2_fill_2 FILLER_62_447 ();
 sg13g2_fill_1 FILLER_62_611 ();
 sg13g2_fill_1 FILLER_62_617 ();
 sg13g2_fill_2 FILLER_62_628 ();
 sg13g2_fill_2 FILLER_62_695 ();
 sg13g2_fill_2 FILLER_62_703 ();
 sg13g2_fill_1 FILLER_62_705 ();
 sg13g2_fill_2 FILLER_62_724 ();
 sg13g2_fill_2 FILLER_62_772 ();
 sg13g2_fill_1 FILLER_62_774 ();
 sg13g2_fill_1 FILLER_62_869 ();
 sg13g2_fill_2 FILLER_63_36 ();
 sg13g2_fill_2 FILLER_63_119 ();
 sg13g2_fill_1 FILLER_63_168 ();
 sg13g2_fill_2 FILLER_63_173 ();
 sg13g2_fill_2 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_211 ();
 sg13g2_fill_1 FILLER_63_217 ();
 sg13g2_fill_1 FILLER_63_224 ();
 sg13g2_fill_2 FILLER_63_235 ();
 sg13g2_fill_2 FILLER_63_270 ();
 sg13g2_fill_1 FILLER_63_272 ();
 sg13g2_fill_1 FILLER_63_338 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_fill_2 FILLER_63_404 ();
 sg13g2_fill_1 FILLER_63_446 ();
 sg13g2_fill_2 FILLER_63_461 ();
 sg13g2_fill_2 FILLER_63_497 ();
 sg13g2_fill_2 FILLER_63_546 ();
 sg13g2_fill_2 FILLER_63_640 ();
 sg13g2_fill_1 FILLER_63_660 ();
 sg13g2_fill_1 FILLER_63_665 ();
 sg13g2_fill_1 FILLER_63_675 ();
 sg13g2_fill_1 FILLER_63_681 ();
 sg13g2_fill_1 FILLER_63_708 ();
 sg13g2_fill_2 FILLER_63_850 ();
 sg13g2_fill_1 FILLER_64_36 ();
 sg13g2_fill_1 FILLER_64_68 ();
 sg13g2_fill_1 FILLER_64_74 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_2 FILLER_64_204 ();
 sg13g2_fill_1 FILLER_64_225 ();
 sg13g2_fill_2 FILLER_64_284 ();
 sg13g2_fill_2 FILLER_64_360 ();
 sg13g2_fill_1 FILLER_64_367 ();
 sg13g2_fill_1 FILLER_64_386 ();
 sg13g2_fill_1 FILLER_64_396 ();
 sg13g2_fill_1 FILLER_64_402 ();
 sg13g2_fill_2 FILLER_64_411 ();
 sg13g2_fill_2 FILLER_64_418 ();
 sg13g2_fill_1 FILLER_64_486 ();
 sg13g2_fill_2 FILLER_64_521 ();
 sg13g2_fill_1 FILLER_64_527 ();
 sg13g2_fill_2 FILLER_64_580 ();
 sg13g2_fill_2 FILLER_64_678 ();
 sg13g2_fill_2 FILLER_64_689 ();
 sg13g2_fill_2 FILLER_64_700 ();
 sg13g2_fill_1 FILLER_64_702 ();
 sg13g2_fill_2 FILLER_64_713 ();
 sg13g2_fill_1 FILLER_64_715 ();
 sg13g2_fill_1 FILLER_64_747 ();
 sg13g2_fill_2 FILLER_64_764 ();
 sg13g2_fill_1 FILLER_64_766 ();
 sg13g2_fill_1 FILLER_64_780 ();
 sg13g2_fill_2 FILLER_64_822 ();
 sg13g2_fill_1 FILLER_64_877 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_40 ();
 sg13g2_fill_1 FILLER_65_111 ();
 sg13g2_fill_2 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_143 ();
 sg13g2_fill_2 FILLER_65_154 ();
 sg13g2_fill_1 FILLER_65_173 ();
 sg13g2_fill_2 FILLER_65_183 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_fill_2 FILLER_65_264 ();
 sg13g2_fill_1 FILLER_65_266 ();
 sg13g2_fill_2 FILLER_65_285 ();
 sg13g2_fill_1 FILLER_65_287 ();
 sg13g2_fill_1 FILLER_65_295 ();
 sg13g2_fill_2 FILLER_65_341 ();
 sg13g2_fill_1 FILLER_65_349 ();
 sg13g2_fill_1 FILLER_65_356 ();
 sg13g2_fill_1 FILLER_65_361 ();
 sg13g2_fill_2 FILLER_65_373 ();
 sg13g2_fill_1 FILLER_65_395 ();
 sg13g2_fill_1 FILLER_65_410 ();
 sg13g2_fill_2 FILLER_65_477 ();
 sg13g2_fill_2 FILLER_65_505 ();
 sg13g2_fill_1 FILLER_65_507 ();
 sg13g2_fill_1 FILLER_65_544 ();
 sg13g2_fill_2 FILLER_65_553 ();
 sg13g2_fill_1 FILLER_65_555 ();
 sg13g2_fill_1 FILLER_65_641 ();
 sg13g2_fill_2 FILLER_65_825 ();
 sg13g2_fill_1 FILLER_65_827 ();
 sg13g2_fill_2 FILLER_65_837 ();
 sg13g2_fill_1 FILLER_65_839 ();
 sg13g2_fill_2 FILLER_65_848 ();
 sg13g2_fill_1 FILLER_65_850 ();
 sg13g2_fill_2 FILLER_65_868 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_44 ();
 sg13g2_fill_2 FILLER_66_79 ();
 sg13g2_fill_1 FILLER_66_81 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_fill_1 FILLER_66_147 ();
 sg13g2_fill_1 FILLER_66_184 ();
 sg13g2_fill_2 FILLER_66_219 ();
 sg13g2_fill_2 FILLER_66_245 ();
 sg13g2_fill_1 FILLER_66_385 ();
 sg13g2_fill_2 FILLER_66_421 ();
 sg13g2_fill_2 FILLER_66_446 ();
 sg13g2_fill_1 FILLER_66_470 ();
 sg13g2_fill_2 FILLER_66_481 ();
 sg13g2_fill_1 FILLER_66_483 ();
 sg13g2_fill_2 FILLER_66_498 ();
 sg13g2_fill_2 FILLER_66_504 ();
 sg13g2_fill_1 FILLER_66_506 ();
 sg13g2_fill_1 FILLER_66_527 ();
 sg13g2_fill_1 FILLER_66_558 ();
 sg13g2_fill_1 FILLER_66_564 ();
 sg13g2_fill_1 FILLER_66_570 ();
 sg13g2_fill_1 FILLER_66_581 ();
 sg13g2_fill_1 FILLER_66_591 ();
 sg13g2_fill_2 FILLER_66_742 ();
 sg13g2_fill_1 FILLER_66_744 ();
 sg13g2_fill_1 FILLER_66_863 ();
 sg13g2_decap_8 FILLER_66_871 ();
 sg13g2_fill_2 FILLER_67_89 ();
 sg13g2_fill_2 FILLER_67_124 ();
 sg13g2_fill_1 FILLER_67_126 ();
 sg13g2_fill_2 FILLER_67_136 ();
 sg13g2_fill_1 FILLER_67_138 ();
 sg13g2_fill_2 FILLER_67_187 ();
 sg13g2_fill_2 FILLER_67_248 ();
 sg13g2_fill_2 FILLER_67_276 ();
 sg13g2_fill_1 FILLER_67_287 ();
 sg13g2_fill_1 FILLER_67_328 ();
 sg13g2_fill_1 FILLER_67_378 ();
 sg13g2_fill_1 FILLER_67_388 ();
 sg13g2_fill_2 FILLER_67_400 ();
 sg13g2_fill_1 FILLER_67_402 ();
 sg13g2_fill_2 FILLER_67_416 ();
 sg13g2_fill_1 FILLER_67_426 ();
 sg13g2_fill_1 FILLER_67_441 ();
 sg13g2_fill_2 FILLER_67_447 ();
 sg13g2_fill_1 FILLER_67_457 ();
 sg13g2_fill_2 FILLER_67_464 ();
 sg13g2_fill_2 FILLER_67_478 ();
 sg13g2_fill_1 FILLER_67_480 ();
 sg13g2_fill_1 FILLER_67_498 ();
 sg13g2_fill_1 FILLER_67_503 ();
 sg13g2_fill_1 FILLER_67_541 ();
 sg13g2_fill_1 FILLER_67_546 ();
 sg13g2_fill_1 FILLER_67_592 ();
 sg13g2_fill_2 FILLER_67_652 ();
 sg13g2_fill_1 FILLER_67_720 ();
 sg13g2_fill_1 FILLER_67_729 ();
 sg13g2_fill_1 FILLER_67_740 ();
 sg13g2_fill_1 FILLER_67_756 ();
 sg13g2_fill_2 FILLER_67_798 ();
 sg13g2_fill_2 FILLER_67_830 ();
 sg13g2_fill_1 FILLER_67_832 ();
 sg13g2_fill_2 FILLER_67_837 ();
 sg13g2_fill_1 FILLER_67_851 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_149 ();
 sg13g2_fill_2 FILLER_68_187 ();
 sg13g2_fill_1 FILLER_68_206 ();
 sg13g2_fill_1 FILLER_68_271 ();
 sg13g2_fill_1 FILLER_68_323 ();
 sg13g2_fill_2 FILLER_68_329 ();
 sg13g2_fill_1 FILLER_68_331 ();
 sg13g2_fill_1 FILLER_68_382 ();
 sg13g2_fill_1 FILLER_68_399 ();
 sg13g2_fill_1 FILLER_68_433 ();
 sg13g2_fill_1 FILLER_68_464 ();
 sg13g2_fill_2 FILLER_68_532 ();
 sg13g2_fill_1 FILLER_68_544 ();
 sg13g2_fill_2 FILLER_68_585 ();
 sg13g2_fill_1 FILLER_68_611 ();
 sg13g2_fill_2 FILLER_68_630 ();
 sg13g2_fill_2 FILLER_68_688 ();
 sg13g2_fill_1 FILLER_68_690 ();
 sg13g2_fill_2 FILLER_68_726 ();
 sg13g2_fill_2 FILLER_68_776 ();
 sg13g2_fill_1 FILLER_68_778 ();
 sg13g2_fill_1 FILLER_68_793 ();
 sg13g2_fill_1 FILLER_68_828 ();
 sg13g2_fill_2 FILLER_68_863 ();
 sg13g2_fill_1 FILLER_68_870 ();
 sg13g2_fill_2 FILLER_68_875 ();
 sg13g2_fill_1 FILLER_68_877 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_69 ();
 sg13g2_fill_1 FILLER_69_80 ();
 sg13g2_fill_2 FILLER_69_90 ();
 sg13g2_fill_1 FILLER_69_101 ();
 sg13g2_fill_2 FILLER_69_107 ();
 sg13g2_fill_1 FILLER_69_109 ();
 sg13g2_fill_2 FILLER_69_159 ();
 sg13g2_fill_1 FILLER_69_197 ();
 sg13g2_fill_1 FILLER_69_266 ();
 sg13g2_fill_2 FILLER_69_301 ();
 sg13g2_fill_1 FILLER_69_303 ();
 sg13g2_fill_1 FILLER_69_359 ();
 sg13g2_fill_2 FILLER_69_386 ();
 sg13g2_fill_1 FILLER_69_393 ();
 sg13g2_fill_2 FILLER_69_473 ();
 sg13g2_fill_1 FILLER_69_475 ();
 sg13g2_fill_2 FILLER_69_493 ();
 sg13g2_fill_1 FILLER_69_495 ();
 sg13g2_fill_2 FILLER_69_706 ();
 sg13g2_fill_1 FILLER_69_708 ();
 sg13g2_fill_1 FILLER_69_736 ();
 sg13g2_fill_1 FILLER_69_745 ();
 sg13g2_decap_4 FILLER_69_843 ();
 sg13g2_fill_2 FILLER_69_850 ();
 sg13g2_decap_8 FILLER_69_864 ();
 sg13g2_decap_8 FILLER_69_871 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_27 ();
 sg13g2_fill_1 FILLER_70_43 ();
 sg13g2_fill_1 FILLER_70_70 ();
 sg13g2_fill_2 FILLER_70_114 ();
 sg13g2_fill_1 FILLER_70_129 ();
 sg13g2_fill_2 FILLER_70_138 ();
 sg13g2_fill_1 FILLER_70_140 ();
 sg13g2_fill_2 FILLER_70_146 ();
 sg13g2_fill_2 FILLER_70_152 ();
 sg13g2_fill_1 FILLER_70_215 ();
 sg13g2_fill_1 FILLER_70_272 ();
 sg13g2_fill_1 FILLER_70_330 ();
 sg13g2_fill_2 FILLER_70_343 ();
 sg13g2_fill_1 FILLER_70_345 ();
 sg13g2_fill_2 FILLER_70_371 ();
 sg13g2_fill_2 FILLER_70_416 ();
 sg13g2_fill_1 FILLER_70_551 ();
 sg13g2_fill_2 FILLER_70_574 ();
 sg13g2_fill_1 FILLER_70_610 ();
 sg13g2_fill_1 FILLER_70_615 ();
 sg13g2_fill_2 FILLER_70_629 ();
 sg13g2_fill_1 FILLER_70_636 ();
 sg13g2_fill_1 FILLER_70_642 ();
 sg13g2_fill_1 FILLER_70_653 ();
 sg13g2_fill_2 FILLER_70_704 ();
 sg13g2_fill_2 FILLER_70_744 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_847 ();
 sg13g2_decap_8 FILLER_70_854 ();
 sg13g2_decap_8 FILLER_70_861 ();
 sg13g2_decap_8 FILLER_70_868 ();
 sg13g2_fill_2 FILLER_70_875 ();
 sg13g2_fill_1 FILLER_70_877 ();
 sg13g2_fill_1 FILLER_71_34 ();
 sg13g2_fill_1 FILLER_71_63 ();
 sg13g2_fill_1 FILLER_71_69 ();
 sg13g2_fill_2 FILLER_71_83 ();
 sg13g2_fill_1 FILLER_71_103 ();
 sg13g2_fill_2 FILLER_71_189 ();
 sg13g2_fill_1 FILLER_71_191 ();
 sg13g2_fill_1 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_279 ();
 sg13g2_fill_2 FILLER_71_324 ();
 sg13g2_fill_1 FILLER_71_326 ();
 sg13g2_fill_2 FILLER_71_353 ();
 sg13g2_fill_2 FILLER_71_385 ();
 sg13g2_fill_1 FILLER_71_417 ();
 sg13g2_fill_1 FILLER_71_437 ();
 sg13g2_fill_1 FILLER_71_468 ();
 sg13g2_fill_1 FILLER_71_473 ();
 sg13g2_fill_1 FILLER_71_484 ();
 sg13g2_fill_2 FILLER_71_490 ();
 sg13g2_fill_1 FILLER_71_497 ();
 sg13g2_fill_1 FILLER_71_503 ();
 sg13g2_fill_1 FILLER_71_509 ();
 sg13g2_fill_1 FILLER_71_521 ();
 sg13g2_fill_2 FILLER_71_545 ();
 sg13g2_fill_1 FILLER_71_571 ();
 sg13g2_fill_2 FILLER_71_581 ();
 sg13g2_fill_2 FILLER_71_657 ();
 sg13g2_fill_1 FILLER_71_704 ();
 sg13g2_fill_2 FILLER_71_734 ();
 sg13g2_fill_1 FILLER_71_767 ();
 sg13g2_fill_2 FILLER_71_801 ();
 sg13g2_fill_2 FILLER_71_817 ();
 sg13g2_decap_8 FILLER_71_839 ();
 sg13g2_decap_8 FILLER_71_846 ();
 sg13g2_decap_8 FILLER_71_853 ();
 sg13g2_decap_8 FILLER_71_860 ();
 sg13g2_decap_8 FILLER_71_867 ();
 sg13g2_decap_4 FILLER_71_874 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_5 ();
 sg13g2_fill_1 FILLER_72_31 ();
 sg13g2_fill_1 FILLER_72_47 ();
 sg13g2_fill_1 FILLER_72_91 ();
 sg13g2_fill_1 FILLER_72_181 ();
 sg13g2_fill_1 FILLER_72_213 ();
 sg13g2_fill_2 FILLER_72_274 ();
 sg13g2_fill_1 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_334 ();
 sg13g2_fill_1 FILLER_72_339 ();
 sg13g2_fill_1 FILLER_72_354 ();
 sg13g2_fill_1 FILLER_72_364 ();
 sg13g2_fill_1 FILLER_72_391 ();
 sg13g2_fill_1 FILLER_72_397 ();
 sg13g2_fill_1 FILLER_72_402 ();
 sg13g2_fill_2 FILLER_72_440 ();
 sg13g2_fill_1 FILLER_72_513 ();
 sg13g2_fill_1 FILLER_72_519 ();
 sg13g2_fill_1 FILLER_72_658 ();
 sg13g2_fill_1 FILLER_72_668 ();
 sg13g2_fill_2 FILLER_72_678 ();
 sg13g2_fill_2 FILLER_72_685 ();
 sg13g2_fill_1 FILLER_72_705 ();
 sg13g2_fill_1 FILLER_72_711 ();
 sg13g2_fill_1 FILLER_72_717 ();
 sg13g2_fill_1 FILLER_72_728 ();
 sg13g2_fill_1 FILLER_72_734 ();
 sg13g2_fill_1 FILLER_72_740 ();
 sg13g2_fill_2 FILLER_72_751 ();
 sg13g2_fill_1 FILLER_72_758 ();
 sg13g2_fill_2 FILLER_72_768 ();
 sg13g2_fill_1 FILLER_72_796 ();
 sg13g2_fill_2 FILLER_72_806 ();
 sg13g2_decap_8 FILLER_72_839 ();
 sg13g2_decap_8 FILLER_72_846 ();
 sg13g2_decap_8 FILLER_72_853 ();
 sg13g2_decap_8 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_72_867 ();
 sg13g2_decap_4 FILLER_72_874 ();
 sg13g2_fill_2 FILLER_73_31 ();
 sg13g2_fill_2 FILLER_73_83 ();
 sg13g2_fill_1 FILLER_73_98 ();
 sg13g2_fill_2 FILLER_73_144 ();
 sg13g2_fill_1 FILLER_73_180 ();
 sg13g2_fill_2 FILLER_73_221 ();
 sg13g2_fill_1 FILLER_73_386 ();
 sg13g2_fill_1 FILLER_73_392 ();
 sg13g2_fill_1 FILLER_73_423 ();
 sg13g2_fill_2 FILLER_73_485 ();
 sg13g2_fill_1 FILLER_73_504 ();
 sg13g2_fill_2 FILLER_73_577 ();
 sg13g2_fill_2 FILLER_73_662 ();
 sg13g2_fill_1 FILLER_73_789 ();
 sg13g2_fill_2 FILLER_73_802 ();
 sg13g2_fill_2 FILLER_73_813 ();
 sg13g2_fill_2 FILLER_73_823 ();
 sg13g2_decap_8 FILLER_73_851 ();
 sg13g2_decap_8 FILLER_73_858 ();
 sg13g2_decap_8 FILLER_73_865 ();
 sg13g2_decap_4 FILLER_73_872 ();
 sg13g2_fill_2 FILLER_73_876 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_10 ();
 sg13g2_fill_1 FILLER_74_27 ();
 sg13g2_fill_1 FILLER_74_83 ();
 sg13g2_fill_1 FILLER_74_133 ();
 sg13g2_fill_1 FILLER_74_182 ();
 sg13g2_fill_1 FILLER_74_231 ();
 sg13g2_fill_1 FILLER_74_258 ();
 sg13g2_fill_1 FILLER_74_285 ();
 sg13g2_fill_1 FILLER_74_296 ();
 sg13g2_fill_1 FILLER_74_307 ();
 sg13g2_fill_1 FILLER_74_336 ();
 sg13g2_fill_1 FILLER_74_341 ();
 sg13g2_fill_2 FILLER_74_414 ();
 sg13g2_fill_1 FILLER_74_421 ();
 sg13g2_fill_1 FILLER_74_432 ();
 sg13g2_fill_1 FILLER_74_438 ();
 sg13g2_fill_1 FILLER_74_485 ();
 sg13g2_fill_2 FILLER_74_571 ();
 sg13g2_fill_1 FILLER_74_660 ();
 sg13g2_fill_2 FILLER_74_695 ();
 sg13g2_fill_2 FILLER_74_766 ();
 sg13g2_fill_2 FILLER_74_807 ();
 sg13g2_decap_8 FILLER_74_851 ();
 sg13g2_decap_8 FILLER_74_858 ();
 sg13g2_decap_8 FILLER_74_865 ();
 sg13g2_decap_4 FILLER_74_872 ();
 sg13g2_fill_2 FILLER_74_876 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_11 ();
 sg13g2_fill_2 FILLER_75_27 ();
 sg13g2_fill_1 FILLER_75_70 ();
 sg13g2_fill_1 FILLER_75_76 ();
 sg13g2_fill_2 FILLER_75_82 ();
 sg13g2_fill_2 FILLER_75_93 ();
 sg13g2_fill_1 FILLER_75_100 ();
 sg13g2_fill_2 FILLER_75_106 ();
 sg13g2_fill_1 FILLER_75_140 ();
 sg13g2_fill_2 FILLER_75_181 ();
 sg13g2_fill_1 FILLER_75_183 ();
 sg13g2_fill_1 FILLER_75_192 ();
 sg13g2_fill_1 FILLER_75_223 ();
 sg13g2_fill_2 FILLER_75_228 ();
 sg13g2_fill_2 FILLER_75_235 ();
 sg13g2_fill_1 FILLER_75_245 ();
 sg13g2_fill_1 FILLER_75_256 ();
 sg13g2_fill_1 FILLER_75_288 ();
 sg13g2_fill_2 FILLER_75_320 ();
 sg13g2_fill_1 FILLER_75_332 ();
 sg13g2_fill_1 FILLER_75_343 ();
 sg13g2_fill_2 FILLER_75_377 ();
 sg13g2_fill_1 FILLER_75_387 ();
 sg13g2_fill_1 FILLER_75_436 ();
 sg13g2_fill_2 FILLER_75_451 ();
 sg13g2_fill_1 FILLER_75_496 ();
 sg13g2_fill_2 FILLER_75_566 ();
 sg13g2_fill_1 FILLER_75_581 ();
 sg13g2_fill_2 FILLER_75_640 ();
 sg13g2_fill_1 FILLER_75_697 ();
 sg13g2_fill_2 FILLER_75_716 ();
 sg13g2_fill_2 FILLER_75_761 ();
 sg13g2_decap_8 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_fill_2 FILLER_75_875 ();
 sg13g2_fill_1 FILLER_75_877 ();
 sg13g2_fill_2 FILLER_76_53 ();
 sg13g2_fill_2 FILLER_76_122 ();
 sg13g2_fill_2 FILLER_76_145 ();
 sg13g2_fill_1 FILLER_76_257 ();
 sg13g2_fill_2 FILLER_76_395 ();
 sg13g2_fill_1 FILLER_76_419 ();
 sg13g2_fill_2 FILLER_76_492 ();
 sg13g2_fill_2 FILLER_76_498 ();
 sg13g2_fill_1 FILLER_76_505 ();
 sg13g2_fill_1 FILLER_76_532 ();
 sg13g2_fill_1 FILLER_76_678 ();
 sg13g2_fill_2 FILLER_76_687 ();
 sg13g2_fill_1 FILLER_76_699 ();
 sg13g2_fill_1 FILLER_76_721 ();
 sg13g2_fill_1 FILLER_76_782 ();
 sg13g2_decap_8 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_76_868 ();
 sg13g2_fill_2 FILLER_76_875 ();
 sg13g2_fill_1 FILLER_76_877 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_4 ();
 sg13g2_fill_2 FILLER_77_45 ();
 sg13g2_fill_2 FILLER_77_94 ();
 sg13g2_fill_1 FILLER_77_144 ();
 sg13g2_fill_2 FILLER_77_150 ();
 sg13g2_fill_1 FILLER_77_208 ();
 sg13g2_fill_2 FILLER_77_283 ();
 sg13g2_fill_2 FILLER_77_314 ();
 sg13g2_fill_1 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_459 ();
 sg13g2_fill_1 FILLER_77_474 ();
 sg13g2_fill_1 FILLER_77_480 ();
 sg13g2_fill_1 FILLER_77_491 ();
 sg13g2_fill_1 FILLER_77_547 ();
 sg13g2_fill_2 FILLER_77_553 ();
 sg13g2_fill_2 FILLER_77_560 ();
 sg13g2_fill_1 FILLER_77_635 ();
 sg13g2_fill_1 FILLER_77_716 ();
 sg13g2_fill_1 FILLER_77_797 ();
 sg13g2_fill_1 FILLER_77_826 ();
 sg13g2_decap_8 FILLER_77_857 ();
 sg13g2_decap_8 FILLER_77_864 ();
 sg13g2_decap_8 FILLER_77_871 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_32 ();
 sg13g2_fill_2 FILLER_78_39 ();
 sg13g2_fill_1 FILLER_78_46 ();
 sg13g2_fill_1 FILLER_78_83 ();
 sg13g2_fill_2 FILLER_78_89 ();
 sg13g2_fill_1 FILLER_78_169 ();
 sg13g2_fill_1 FILLER_78_237 ();
 sg13g2_fill_2 FILLER_78_253 ();
 sg13g2_fill_1 FILLER_78_263 ();
 sg13g2_fill_1 FILLER_78_306 ();
 sg13g2_fill_1 FILLER_78_333 ();
 sg13g2_fill_2 FILLER_78_344 ();
 sg13g2_fill_1 FILLER_78_360 ();
 sg13g2_fill_1 FILLER_78_391 ();
 sg13g2_fill_2 FILLER_78_397 ();
 sg13g2_fill_2 FILLER_78_455 ();
 sg13g2_fill_2 FILLER_78_490 ();
 sg13g2_fill_2 FILLER_78_504 ();
 sg13g2_fill_1 FILLER_78_581 ();
 sg13g2_fill_2 FILLER_78_587 ();
 sg13g2_fill_1 FILLER_78_596 ();
 sg13g2_fill_2 FILLER_78_602 ();
 sg13g2_fill_1 FILLER_78_609 ();
 sg13g2_fill_1 FILLER_78_619 ();
 sg13g2_fill_1 FILLER_78_639 ();
 sg13g2_fill_1 FILLER_78_672 ();
 sg13g2_fill_1 FILLER_78_704 ();
 sg13g2_fill_1 FILLER_78_714 ();
 sg13g2_fill_1 FILLER_78_729 ();
 sg13g2_fill_2 FILLER_78_764 ();
 sg13g2_fill_1 FILLER_78_822 ();
 sg13g2_fill_2 FILLER_78_827 ();
 sg13g2_fill_1 FILLER_78_829 ();
 sg13g2_decap_8 FILLER_78_862 ();
 sg13g2_decap_8 FILLER_78_869 ();
 sg13g2_fill_2 FILLER_78_876 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_47 ();
 sg13g2_fill_2 FILLER_79_69 ();
 sg13g2_fill_2 FILLER_79_124 ();
 sg13g2_fill_2 FILLER_79_156 ();
 sg13g2_fill_1 FILLER_79_202 ();
 sg13g2_fill_1 FILLER_79_275 ();
 sg13g2_fill_1 FILLER_79_390 ();
 sg13g2_fill_1 FILLER_79_624 ();
 sg13g2_fill_2 FILLER_79_819 ();
 sg13g2_fill_1 FILLER_79_821 ();
 sg13g2_fill_2 FILLER_79_830 ();
 sg13g2_fill_1 FILLER_79_832 ();
 sg13g2_decap_8 FILLER_79_862 ();
 sg13g2_decap_8 FILLER_79_869 ();
 sg13g2_fill_2 FILLER_79_876 ();
 sg13g2_fill_2 FILLER_80_54 ();
 sg13g2_fill_1 FILLER_80_191 ();
 sg13g2_fill_1 FILLER_80_308 ();
 sg13g2_fill_1 FILLER_80_403 ();
 sg13g2_fill_1 FILLER_80_408 ();
 sg13g2_fill_1 FILLER_80_413 ();
 sg13g2_fill_2 FILLER_80_418 ();
 sg13g2_fill_1 FILLER_80_446 ();
 sg13g2_fill_1 FILLER_80_491 ();
 sg13g2_fill_2 FILLER_80_496 ();
 sg13g2_fill_1 FILLER_80_558 ();
 sg13g2_fill_1 FILLER_80_589 ();
 sg13g2_fill_2 FILLER_80_675 ();
 sg13g2_fill_1 FILLER_80_720 ();
 sg13g2_decap_8 FILLER_80_850 ();
 sg13g2_decap_8 FILLER_80_857 ();
 sg13g2_decap_8 FILLER_80_864 ();
 sg13g2_decap_8 FILLER_80_871 ();
endmodule
