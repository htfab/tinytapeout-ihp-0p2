module tt_um_htfab_rotfpga2 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire clknet_0_clk;
 wire net183;
 wire \g.g_y[0].g_x[0].t.out_sc ;
 wire \g.g_y[0].g_x[0].t.r_d ;
 wire \g.g_y[0].g_x[0].t.r_ghl ;
 wire \g.g_y[0].g_x[0].t.r_gnl ;
 wire \g.g_y[0].g_x[0].t.r_h ;
 wire \g.g_y[0].g_x[0].t.r_v ;
 wire \g.g_y[0].g_x[1].t.out_sc ;
 wire \g.g_y[0].g_x[1].t.r_d ;
 wire \g.g_y[0].g_x[1].t.r_h ;
 wire \g.g_y[0].g_x[1].t.r_v ;
 wire \g.g_y[0].g_x[2].t.out_sc ;
 wire \g.g_y[0].g_x[2].t.r_d ;
 wire \g.g_y[0].g_x[2].t.r_ghl ;
 wire \g.g_y[0].g_x[2].t.r_gnl ;
 wire \g.g_y[0].g_x[2].t.r_h ;
 wire \g.g_y[0].g_x[2].t.r_v ;
 wire \g.g_y[0].g_x[3].t.out_sc ;
 wire \g.g_y[0].g_x[3].t.r_d ;
 wire \g.g_y[0].g_x[3].t.r_h ;
 wire \g.g_y[0].g_x[3].t.r_v ;
 wire \g.g_y[0].g_x[4].t.out_sc ;
 wire \g.g_y[0].g_x[4].t.r_d ;
 wire \g.g_y[0].g_x[4].t.r_ghl ;
 wire \g.g_y[0].g_x[4].t.r_gnl ;
 wire \g.g_y[0].g_x[4].t.r_h ;
 wire \g.g_y[0].g_x[4].t.r_v ;
 wire \g.g_y[0].g_x[5].t.out_sc ;
 wire \g.g_y[0].g_x[5].t.r_d ;
 wire \g.g_y[0].g_x[5].t.r_h ;
 wire \g.g_y[0].g_x[5].t.r_v ;
 wire \g.g_y[0].g_x[6].t.out_sc ;
 wire \g.g_y[0].g_x[6].t.r_d ;
 wire \g.g_y[0].g_x[6].t.r_ghl ;
 wire \g.g_y[0].g_x[6].t.r_gnl ;
 wire \g.g_y[0].g_x[6].t.r_h ;
 wire \g.g_y[0].g_x[6].t.r_v ;
 wire \g.g_y[0].g_x[7].t.out_r ;
 wire \g.g_y[0].g_x[7].t.out_sc ;
 wire \g.g_y[0].g_x[7].t.r_d ;
 wire \g.g_y[0].g_x[7].t.r_h ;
 wire \g.g_y[0].g_x[7].t.r_v ;
 wire \g.g_y[1].g_x[0].t.out_sc ;
 wire \g.g_y[1].g_x[0].t.r_d ;
 wire \g.g_y[1].g_x[0].t.r_h ;
 wire \g.g_y[1].g_x[0].t.r_v ;
 wire \g.g_y[1].g_x[1].t.out_sc ;
 wire \g.g_y[1].g_x[1].t.r_d ;
 wire \g.g_y[1].g_x[1].t.r_ghl ;
 wire \g.g_y[1].g_x[1].t.r_gnl ;
 wire \g.g_y[1].g_x[1].t.r_h ;
 wire \g.g_y[1].g_x[1].t.r_v ;
 wire \g.g_y[1].g_x[2].t.out_sc ;
 wire \g.g_y[1].g_x[2].t.r_d ;
 wire \g.g_y[1].g_x[2].t.r_h ;
 wire \g.g_y[1].g_x[2].t.r_v ;
 wire \g.g_y[1].g_x[3].t.out_sc ;
 wire \g.g_y[1].g_x[3].t.r_d ;
 wire \g.g_y[1].g_x[3].t.r_ghl ;
 wire \g.g_y[1].g_x[3].t.r_gnl ;
 wire \g.g_y[1].g_x[3].t.r_h ;
 wire \g.g_y[1].g_x[3].t.r_v ;
 wire \g.g_y[1].g_x[4].t.out_sc ;
 wire \g.g_y[1].g_x[4].t.r_d ;
 wire \g.g_y[1].g_x[4].t.r_h ;
 wire \g.g_y[1].g_x[4].t.r_v ;
 wire \g.g_y[1].g_x[5].t.out_sc ;
 wire \g.g_y[1].g_x[5].t.r_d ;
 wire \g.g_y[1].g_x[5].t.r_ghl ;
 wire \g.g_y[1].g_x[5].t.r_gnl ;
 wire \g.g_y[1].g_x[5].t.r_h ;
 wire \g.g_y[1].g_x[5].t.r_v ;
 wire \g.g_y[1].g_x[6].t.out_sc ;
 wire \g.g_y[1].g_x[6].t.r_d ;
 wire \g.g_y[1].g_x[6].t.r_h ;
 wire \g.g_y[1].g_x[6].t.r_v ;
 wire \g.g_y[1].g_x[7].t.out_r ;
 wire \g.g_y[1].g_x[7].t.out_sc ;
 wire \g.g_y[1].g_x[7].t.r_d ;
 wire \g.g_y[1].g_x[7].t.r_ghl ;
 wire \g.g_y[1].g_x[7].t.r_gnl ;
 wire \g.g_y[1].g_x[7].t.r_h ;
 wire \g.g_y[1].g_x[7].t.r_v ;
 wire \g.g_y[2].g_x[0].t.out_sc ;
 wire \g.g_y[2].g_x[0].t.r_d ;
 wire \g.g_y[2].g_x[0].t.r_ghl ;
 wire \g.g_y[2].g_x[0].t.r_gnl ;
 wire \g.g_y[2].g_x[0].t.r_h ;
 wire \g.g_y[2].g_x[0].t.r_v ;
 wire \g.g_y[2].g_x[1].t.out_sc ;
 wire \g.g_y[2].g_x[1].t.r_d ;
 wire \g.g_y[2].g_x[1].t.r_h ;
 wire \g.g_y[2].g_x[1].t.r_v ;
 wire \g.g_y[2].g_x[2].t.out_sc ;
 wire \g.g_y[2].g_x[2].t.r_d ;
 wire \g.g_y[2].g_x[2].t.r_ghl ;
 wire \g.g_y[2].g_x[2].t.r_gnl ;
 wire \g.g_y[2].g_x[2].t.r_h ;
 wire \g.g_y[2].g_x[2].t.r_v ;
 wire \g.g_y[2].g_x[3].t.out_sc ;
 wire \g.g_y[2].g_x[3].t.r_d ;
 wire \g.g_y[2].g_x[3].t.r_h ;
 wire \g.g_y[2].g_x[3].t.r_v ;
 wire \g.g_y[2].g_x[4].t.out_sc ;
 wire \g.g_y[2].g_x[4].t.r_d ;
 wire \g.g_y[2].g_x[4].t.r_ghl ;
 wire \g.g_y[2].g_x[4].t.r_gnl ;
 wire \g.g_y[2].g_x[4].t.r_h ;
 wire \g.g_y[2].g_x[4].t.r_v ;
 wire \g.g_y[2].g_x[5].t.out_sc ;
 wire \g.g_y[2].g_x[5].t.r_d ;
 wire \g.g_y[2].g_x[5].t.r_h ;
 wire \g.g_y[2].g_x[5].t.r_v ;
 wire \g.g_y[2].g_x[6].t.out_sc ;
 wire \g.g_y[2].g_x[6].t.r_d ;
 wire \g.g_y[2].g_x[6].t.r_ghl ;
 wire \g.g_y[2].g_x[6].t.r_gnl ;
 wire \g.g_y[2].g_x[6].t.r_h ;
 wire \g.g_y[2].g_x[6].t.r_v ;
 wire \g.g_y[2].g_x[7].t.out_r ;
 wire \g.g_y[2].g_x[7].t.out_sc ;
 wire \g.g_y[2].g_x[7].t.r_d ;
 wire \g.g_y[2].g_x[7].t.r_h ;
 wire \g.g_y[2].g_x[7].t.r_v ;
 wire \g.g_y[3].g_x[0].t.out_sc ;
 wire \g.g_y[3].g_x[0].t.r_d ;
 wire \g.g_y[3].g_x[0].t.r_h ;
 wire \g.g_y[3].g_x[0].t.r_v ;
 wire \g.g_y[3].g_x[1].t.out_sc ;
 wire \g.g_y[3].g_x[1].t.r_d ;
 wire \g.g_y[3].g_x[1].t.r_ghl ;
 wire \g.g_y[3].g_x[1].t.r_gnl ;
 wire \g.g_y[3].g_x[1].t.r_h ;
 wire \g.g_y[3].g_x[1].t.r_v ;
 wire \g.g_y[3].g_x[2].t.out_sc ;
 wire \g.g_y[3].g_x[2].t.r_d ;
 wire \g.g_y[3].g_x[2].t.r_h ;
 wire \g.g_y[3].g_x[2].t.r_v ;
 wire \g.g_y[3].g_x[3].t.out_sc ;
 wire \g.g_y[3].g_x[3].t.r_d ;
 wire \g.g_y[3].g_x[3].t.r_ghl ;
 wire \g.g_y[3].g_x[3].t.r_gnl ;
 wire \g.g_y[3].g_x[3].t.r_h ;
 wire \g.g_y[3].g_x[3].t.r_v ;
 wire \g.g_y[3].g_x[4].t.out_sc ;
 wire \g.g_y[3].g_x[4].t.r_d ;
 wire \g.g_y[3].g_x[4].t.r_h ;
 wire \g.g_y[3].g_x[4].t.r_v ;
 wire \g.g_y[3].g_x[5].t.out_sc ;
 wire \g.g_y[3].g_x[5].t.r_d ;
 wire \g.g_y[3].g_x[5].t.r_ghl ;
 wire \g.g_y[3].g_x[5].t.r_gnl ;
 wire \g.g_y[3].g_x[5].t.r_h ;
 wire \g.g_y[3].g_x[5].t.r_v ;
 wire \g.g_y[3].g_x[6].t.out_sc ;
 wire \g.g_y[3].g_x[6].t.r_d ;
 wire \g.g_y[3].g_x[6].t.r_h ;
 wire \g.g_y[3].g_x[6].t.r_v ;
 wire \g.g_y[3].g_x[7].t.out_r ;
 wire \g.g_y[3].g_x[7].t.out_sc ;
 wire \g.g_y[3].g_x[7].t.r_d ;
 wire \g.g_y[3].g_x[7].t.r_ghl ;
 wire \g.g_y[3].g_x[7].t.r_gnl ;
 wire \g.g_y[3].g_x[7].t.r_h ;
 wire \g.g_y[3].g_x[7].t.r_v ;
 wire \g.g_y[4].g_x[0].t.out_sc ;
 wire \g.g_y[4].g_x[0].t.r_d ;
 wire \g.g_y[4].g_x[0].t.r_ghl ;
 wire \g.g_y[4].g_x[0].t.r_gnl ;
 wire \g.g_y[4].g_x[0].t.r_h ;
 wire \g.g_y[4].g_x[0].t.r_v ;
 wire \g.g_y[4].g_x[1].t.out_sc ;
 wire \g.g_y[4].g_x[1].t.r_d ;
 wire \g.g_y[4].g_x[1].t.r_h ;
 wire \g.g_y[4].g_x[1].t.r_v ;
 wire \g.g_y[4].g_x[2].t.out_sc ;
 wire \g.g_y[4].g_x[2].t.r_d ;
 wire \g.g_y[4].g_x[2].t.r_ghl ;
 wire \g.g_y[4].g_x[2].t.r_gnl ;
 wire \g.g_y[4].g_x[2].t.r_h ;
 wire \g.g_y[4].g_x[2].t.r_v ;
 wire \g.g_y[4].g_x[3].t.out_sc ;
 wire \g.g_y[4].g_x[3].t.r_d ;
 wire \g.g_y[4].g_x[3].t.r_h ;
 wire \g.g_y[4].g_x[3].t.r_v ;
 wire \g.g_y[4].g_x[4].t.out_sc ;
 wire \g.g_y[4].g_x[4].t.r_d ;
 wire \g.g_y[4].g_x[4].t.r_ghl ;
 wire \g.g_y[4].g_x[4].t.r_gnl ;
 wire \g.g_y[4].g_x[4].t.r_h ;
 wire \g.g_y[4].g_x[4].t.r_v ;
 wire \g.g_y[4].g_x[5].t.out_sc ;
 wire \g.g_y[4].g_x[5].t.r_d ;
 wire \g.g_y[4].g_x[5].t.r_h ;
 wire \g.g_y[4].g_x[5].t.r_v ;
 wire \g.g_y[4].g_x[6].t.out_sc ;
 wire \g.g_y[4].g_x[6].t.r_d ;
 wire \g.g_y[4].g_x[6].t.r_ghl ;
 wire \g.g_y[4].g_x[6].t.r_gnl ;
 wire \g.g_y[4].g_x[6].t.r_h ;
 wire \g.g_y[4].g_x[6].t.r_v ;
 wire \g.g_y[4].g_x[7].t.out_r ;
 wire \g.g_y[4].g_x[7].t.out_sc ;
 wire \g.g_y[4].g_x[7].t.r_d ;
 wire \g.g_y[4].g_x[7].t.r_h ;
 wire \g.g_y[4].g_x[7].t.r_v ;
 wire \g.g_y[5].g_x[0].t.out_sc ;
 wire \g.g_y[5].g_x[0].t.r_d ;
 wire \g.g_y[5].g_x[0].t.r_h ;
 wire \g.g_y[5].g_x[0].t.r_v ;
 wire \g.g_y[5].g_x[1].t.out_sc ;
 wire \g.g_y[5].g_x[1].t.r_d ;
 wire \g.g_y[5].g_x[1].t.r_ghl ;
 wire \g.g_y[5].g_x[1].t.r_gnl ;
 wire \g.g_y[5].g_x[1].t.r_h ;
 wire \g.g_y[5].g_x[1].t.r_v ;
 wire \g.g_y[5].g_x[2].t.out_sc ;
 wire \g.g_y[5].g_x[2].t.r_d ;
 wire \g.g_y[5].g_x[2].t.r_h ;
 wire \g.g_y[5].g_x[2].t.r_v ;
 wire \g.g_y[5].g_x[3].t.out_sc ;
 wire \g.g_y[5].g_x[3].t.r_d ;
 wire \g.g_y[5].g_x[3].t.r_ghl ;
 wire \g.g_y[5].g_x[3].t.r_gnl ;
 wire \g.g_y[5].g_x[3].t.r_h ;
 wire \g.g_y[5].g_x[3].t.r_v ;
 wire \g.g_y[5].g_x[4].t.out_sc ;
 wire \g.g_y[5].g_x[4].t.r_d ;
 wire \g.g_y[5].g_x[4].t.r_h ;
 wire \g.g_y[5].g_x[4].t.r_v ;
 wire \g.g_y[5].g_x[5].t.out_sc ;
 wire \g.g_y[5].g_x[5].t.r_d ;
 wire \g.g_y[5].g_x[5].t.r_ghl ;
 wire \g.g_y[5].g_x[5].t.r_gnl ;
 wire \g.g_y[5].g_x[5].t.r_h ;
 wire \g.g_y[5].g_x[5].t.r_v ;
 wire \g.g_y[5].g_x[6].t.out_sc ;
 wire \g.g_y[5].g_x[6].t.r_d ;
 wire \g.g_y[5].g_x[6].t.r_h ;
 wire \g.g_y[5].g_x[6].t.r_v ;
 wire \g.g_y[5].g_x[7].t.out_r ;
 wire \g.g_y[5].g_x[7].t.out_sc ;
 wire \g.g_y[5].g_x[7].t.r_d ;
 wire \g.g_y[5].g_x[7].t.r_ghl ;
 wire \g.g_y[5].g_x[7].t.r_gnl ;
 wire \g.g_y[5].g_x[7].t.r_h ;
 wire \g.g_y[5].g_x[7].t.r_v ;
 wire \g.g_y[6].g_x[0].t.out_sc ;
 wire \g.g_y[6].g_x[0].t.r_d ;
 wire \g.g_y[6].g_x[0].t.r_ghl ;
 wire \g.g_y[6].g_x[0].t.r_gnl ;
 wire \g.g_y[6].g_x[0].t.r_h ;
 wire \g.g_y[6].g_x[0].t.r_v ;
 wire \g.g_y[6].g_x[1].t.out_sc ;
 wire \g.g_y[6].g_x[1].t.r_d ;
 wire \g.g_y[6].g_x[1].t.r_h ;
 wire \g.g_y[6].g_x[1].t.r_v ;
 wire \g.g_y[6].g_x[2].t.out_sc ;
 wire \g.g_y[6].g_x[2].t.r_d ;
 wire \g.g_y[6].g_x[2].t.r_ghl ;
 wire \g.g_y[6].g_x[2].t.r_gnl ;
 wire \g.g_y[6].g_x[2].t.r_h ;
 wire \g.g_y[6].g_x[2].t.r_v ;
 wire \g.g_y[6].g_x[3].t.out_sc ;
 wire \g.g_y[6].g_x[3].t.r_d ;
 wire \g.g_y[6].g_x[3].t.r_h ;
 wire \g.g_y[6].g_x[3].t.r_v ;
 wire \g.g_y[6].g_x[4].t.out_sc ;
 wire \g.g_y[6].g_x[4].t.r_d ;
 wire \g.g_y[6].g_x[4].t.r_ghl ;
 wire \g.g_y[6].g_x[4].t.r_gnl ;
 wire \g.g_y[6].g_x[4].t.r_h ;
 wire \g.g_y[6].g_x[4].t.r_v ;
 wire \g.g_y[6].g_x[5].t.out_sc ;
 wire \g.g_y[6].g_x[5].t.r_d ;
 wire \g.g_y[6].g_x[5].t.r_h ;
 wire \g.g_y[6].g_x[5].t.r_v ;
 wire \g.g_y[6].g_x[6].t.out_sc ;
 wire \g.g_y[6].g_x[6].t.r_d ;
 wire \g.g_y[6].g_x[6].t.r_ghl ;
 wire \g.g_y[6].g_x[6].t.r_gnl ;
 wire \g.g_y[6].g_x[6].t.r_h ;
 wire \g.g_y[6].g_x[6].t.r_v ;
 wire \g.g_y[6].g_x[7].t.out_r ;
 wire \g.g_y[6].g_x[7].t.out_sc ;
 wire \g.g_y[6].g_x[7].t.r_d ;
 wire \g.g_y[6].g_x[7].t.r_h ;
 wire \g.g_y[6].g_x[7].t.r_v ;
 wire \g.g_y[7].g_x[0].t.out_sc ;
 wire \g.g_y[7].g_x[0].t.r_d ;
 wire \g.g_y[7].g_x[0].t.r_h ;
 wire \g.g_y[7].g_x[0].t.r_v ;
 wire \g.g_y[7].g_x[1].t.out_sc ;
 wire \g.g_y[7].g_x[1].t.r_d ;
 wire \g.g_y[7].g_x[1].t.r_ghl ;
 wire \g.g_y[7].g_x[1].t.r_gnl ;
 wire \g.g_y[7].g_x[1].t.r_h ;
 wire \g.g_y[7].g_x[1].t.r_v ;
 wire \g.g_y[7].g_x[2].t.out_sc ;
 wire \g.g_y[7].g_x[2].t.r_d ;
 wire \g.g_y[7].g_x[2].t.r_h ;
 wire \g.g_y[7].g_x[2].t.r_v ;
 wire \g.g_y[7].g_x[3].t.out_sc ;
 wire \g.g_y[7].g_x[3].t.r_d ;
 wire \g.g_y[7].g_x[3].t.r_ghl ;
 wire \g.g_y[7].g_x[3].t.r_gnl ;
 wire \g.g_y[7].g_x[3].t.r_h ;
 wire \g.g_y[7].g_x[3].t.r_v ;
 wire \g.g_y[7].g_x[4].t.out_sc ;
 wire \g.g_y[7].g_x[4].t.r_d ;
 wire \g.g_y[7].g_x[4].t.r_h ;
 wire \g.g_y[7].g_x[4].t.r_v ;
 wire \g.g_y[7].g_x[5].t.out_sc ;
 wire \g.g_y[7].g_x[5].t.r_d ;
 wire \g.g_y[7].g_x[5].t.r_ghl ;
 wire \g.g_y[7].g_x[5].t.r_gnl ;
 wire \g.g_y[7].g_x[5].t.r_h ;
 wire \g.g_y[7].g_x[5].t.r_v ;
 wire \g.g_y[7].g_x[6].t.out_sc ;
 wire \g.g_y[7].g_x[6].t.r_d ;
 wire \g.g_y[7].g_x[6].t.r_h ;
 wire \g.g_y[7].g_x[6].t.r_v ;
 wire \g.g_y[7].g_x[7].t.out_r ;
 wire \g.g_y[7].g_x[7].t.out_sc ;
 wire \g.g_y[7].g_x[7].t.r_d ;
 wire \g.g_y[7].g_x[7].t.r_ghl ;
 wire \g.g_y[7].g_x[7].t.r_gnl ;
 wire \g.g_y[7].g_x[7].t.r_h ;
 wire \g.g_y[7].g_x[7].t.r_v ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_2 _2862_ (.A(\g.g_y[7].g_x[7].t.r_d ),
    .X(_2348_));
 sg13g2_buf_1 _2863_ (.A(\g.g_y[7].g_x[6].t.r_h ),
    .X(_2349_));
 sg13g2_buf_1 _2864_ (.A(\g.g_y[7].g_x[6].t.r_d ),
    .X(_2350_));
 sg13g2_buf_1 _2865_ (.A(\g.g_y[6].g_x[6].t.r_ghl ),
    .X(_2351_));
 sg13g2_buf_2 _2866_ (.A(\g.g_y[6].g_x[6].t.r_d ),
    .X(_2352_));
 sg13g2_mux2_1 _2867_ (.A0(\g.g_y[6].g_x[6].t.r_gnl ),
    .A1(\g.g_y[6].g_x[6].t.out_sc ),
    .S(_2352_),
    .X(_2353_));
 sg13g2_buf_2 _2868_ (.A(\g.g_y[6].g_x[6].t.r_v ),
    .X(_2354_));
 sg13g2_mux2_1 _2869_ (.A0(_2351_),
    .A1(_2353_),
    .S(_2354_),
    .X(_2355_));
 sg13g2_buf_1 _2870_ (.A(\g.g_y[0].g_x[6].t.r_ghl ),
    .X(_2356_));
 sg13g2_buf_8 _2871_ (.A(\g.g_y[0].g_x[6].t.r_d ),
    .X(_2357_));
 sg13g2_mux2_1 _2872_ (.A0(\g.g_y[0].g_x[6].t.r_gnl ),
    .A1(\g.g_y[0].g_x[6].t.out_sc ),
    .S(_2357_),
    .X(_2358_));
 sg13g2_buf_2 _2873_ (.A(\g.g_y[0].g_x[6].t.r_v ),
    .X(_2359_));
 sg13g2_inv_1 _2874_ (.Y(_2360_),
    .A(_2359_));
 sg13g2_mux2_1 _2875_ (.A0(_2356_),
    .A1(_2358_),
    .S(_2360_),
    .X(_2361_));
 sg13g2_buf_1 _2876_ (.A(\g.g_y[7].g_x[6].t.r_v ),
    .X(_2362_));
 sg13g2_inv_1 _2877_ (.Y(_2363_),
    .A(_2362_));
 sg13g2_mux2_1 _2878_ (.A0(_2355_),
    .A1(_2361_),
    .S(_2363_),
    .X(_2364_));
 sg13g2_buf_1 _2879_ (.A(_2364_),
    .X(_2365_));
 sg13g2_buf_2 _2880_ (.A(\g.g_y[7].g_x[5].t.r_ghl ),
    .X(_2366_));
 sg13g2_buf_8 _2881_ (.A(\g.g_y[7].g_x[5].t.r_d ),
    .X(_2367_));
 sg13g2_mux2_1 _2882_ (.A0(\g.g_y[7].g_x[5].t.out_sc ),
    .A1(\g.g_y[7].g_x[5].t.r_gnl ),
    .S(_2367_),
    .X(_2368_));
 sg13g2_buf_1 _2883_ (.A(\g.g_y[7].g_x[5].t.r_h ),
    .X(_2369_));
 sg13g2_mux2_1 _2884_ (.A0(_2366_),
    .A1(_2368_),
    .S(net88),
    .X(_2370_));
 sg13g2_buf_1 _2885_ (.A(_2370_),
    .X(_2371_));
 sg13g2_nand4_1 _2886_ (.B(_2350_),
    .C(_2365_),
    .A(net90),
    .Y(_2372_),
    .D(_2371_));
 sg13g2_buf_1 _2887_ (.A(\g.g_y[7].g_x[6].t.out_sc ),
    .X(_2373_));
 sg13g2_nor2_1 _2888_ (.A(_2350_),
    .B(_2373_),
    .Y(_2374_));
 sg13g2_nand2b_1 _2889_ (.Y(_2375_),
    .B(_2360_),
    .A_N(_2358_));
 sg13g2_inv_1 _2890_ (.Y(_2376_),
    .A(_2356_));
 sg13g2_a21oi_1 _2891_ (.A1(_2376_),
    .A2(_2359_),
    .Y(_2377_),
    .B1(_2363_));
 sg13g2_a22oi_1 _2892_ (.Y(_2378_),
    .B1(_2375_),
    .B2(_2377_),
    .A2(_2355_),
    .A1(_2363_));
 sg13g2_inv_1 _2893_ (.Y(_2379_),
    .A(\g.g_y[7].g_x[6].t.r_d ));
 sg13g2_nor2_1 _2894_ (.A(net90),
    .B(_2379_),
    .Y(_2380_));
 sg13g2_nor3_1 _2895_ (.A(_2349_),
    .B(net89),
    .C(_2371_),
    .Y(_2381_));
 sg13g2_a221oi_1 _2896_ (.B2(_2380_),
    .C1(_2381_),
    .B1(_2378_),
    .A1(_2349_),
    .Y(_2382_),
    .A2(_2374_));
 sg13g2_buf_2 _2897_ (.A(\g.g_y[7].g_x[7].t.r_h ),
    .X(_2383_));
 sg13g2_a21o_1 _2898_ (.A2(_2382_),
    .A1(_2372_),
    .B1(_2383_),
    .X(_2384_));
 sg13g2_buf_2 _2899_ (.A(\g.g_y[7].g_x[1].t.r_h ),
    .X(_2385_));
 sg13g2_buf_2 _2900_ (.A(\g.g_y[7].g_x[1].t.r_d ),
    .X(_2386_));
 sg13g2_mux2_1 _2901_ (.A0(\g.g_y[7].g_x[1].t.out_sc ),
    .A1(\g.g_y[7].g_x[1].t.r_gnl ),
    .S(_2386_),
    .X(_2387_));
 sg13g2_buf_1 _2902_ (.A(\g.g_y[7].g_x[1].t.r_ghl ),
    .X(_2388_));
 sg13g2_nand2b_1 _2903_ (.Y(_2389_),
    .B(_2385_),
    .A_N(_2388_));
 sg13g2_o21ai_1 _2904_ (.B1(_2389_),
    .Y(_2390_),
    .A1(_2385_),
    .A2(_2387_));
 sg13g2_buf_2 _2905_ (.A(\g.g_y[0].g_x[0].t.r_d ),
    .X(_2391_));
 sg13g2_mux2_1 _2906_ (.A0(\g.g_y[0].g_x[0].t.r_gnl ),
    .A1(\g.g_y[0].g_x[0].t.out_sc ),
    .S(_2391_),
    .X(_2392_));
 sg13g2_buf_1 _2907_ (.A(_2392_),
    .X(_2393_));
 sg13g2_buf_2 _2908_ (.A(\g.g_y[0].g_x[0].t.r_v ),
    .X(_2394_));
 sg13g2_inv_1 _2909_ (.Y(_2395_),
    .A(_2394_));
 sg13g2_nand2b_1 _2910_ (.Y(_2396_),
    .B(_2395_),
    .A_N(_2393_));
 sg13g2_buf_1 _2911_ (.A(\g.g_y[7].g_x[0].t.r_v ),
    .X(_2397_));
 sg13g2_buf_1 _2912_ (.A(\g.g_y[7].g_x[0].t.r_d ),
    .X(_2398_));
 sg13g2_inv_1 _2913_ (.Y(_2399_),
    .A(net86));
 sg13g2_buf_1 _2914_ (.A(\g.g_y[0].g_x[0].t.r_ghl ),
    .X(_2400_));
 sg13g2_nor2b_1 _2915_ (.A(_2400_),
    .B_N(_2394_),
    .Y(_2401_));
 sg13g2_nor3_1 _2916_ (.A(net87),
    .B(_2399_),
    .C(_2401_),
    .Y(_2402_));
 sg13g2_buf_2 _2917_ (.A(\g.g_y[6].g_x[0].t.r_ghl ),
    .X(_2403_));
 sg13g2_buf_2 _2918_ (.A(\g.g_y[6].g_x[0].t.r_v ),
    .X(_2404_));
 sg13g2_nor2_1 _2919_ (.A(_2403_),
    .B(_2404_),
    .Y(_2405_));
 sg13g2_nand2_1 _2920_ (.Y(_2406_),
    .A(\g.g_y[7].g_x[0].t.r_v ),
    .B(_2398_));
 sg13g2_nor2_1 _2921_ (.A(_2405_),
    .B(_2406_),
    .Y(_2407_));
 sg13g2_inv_2 _2922_ (.Y(_2408_),
    .A(_2404_));
 sg13g2_buf_8 _2923_ (.A(\g.g_y[6].g_x[0].t.r_d ),
    .X(_2409_));
 sg13g2_mux2_1 _2924_ (.A0(\g.g_y[6].g_x[0].t.r_gnl ),
    .A1(\g.g_y[6].g_x[0].t.out_sc ),
    .S(_2409_),
    .X(_2410_));
 sg13g2_buf_1 _2925_ (.A(_2410_),
    .X(_2411_));
 sg13g2_or2_1 _2926_ (.X(_2412_),
    .B(_2411_),
    .A(_2408_));
 sg13g2_buf_2 _2927_ (.A(_2412_),
    .X(_2413_));
 sg13g2_a22oi_1 _2928_ (.Y(_2414_),
    .B1(_2407_),
    .B2(_2413_),
    .A2(_2402_),
    .A1(_2396_));
 sg13g2_buf_2 _2929_ (.A(\g.g_y[7].g_x[0].t.r_h ),
    .X(_2415_));
 sg13g2_nor2_1 _2930_ (.A(\g.g_y[7].g_x[0].t.out_sc ),
    .B(net86),
    .Y(_2416_));
 sg13g2_nor2_1 _2931_ (.A(_2415_),
    .B(_2416_),
    .Y(_2417_));
 sg13g2_o21ai_1 _2932_ (.B1(_2417_),
    .Y(_2418_),
    .A1(_2390_),
    .A2(_2414_));
 sg13g2_inv_1 _2933_ (.Y(_2419_),
    .A(_2415_));
 sg13g2_mux2_1 _2934_ (.A0(_2400_),
    .A1(_2393_),
    .S(_2395_),
    .X(_2420_));
 sg13g2_buf_2 _2935_ (.A(_2420_),
    .X(_2421_));
 sg13g2_nor2_1 _2936_ (.A(net87),
    .B(_2405_),
    .Y(_2422_));
 sg13g2_a221oi_1 _2937_ (.B2(_2413_),
    .C1(_2399_),
    .B1(_2422_),
    .A1(net87),
    .Y(_2423_),
    .A2(_2421_));
 sg13g2_buf_1 _2938_ (.A(ui_in[7]),
    .X(_2424_));
 sg13g2_nor2b_1 _2939_ (.A(_2385_),
    .B_N(_2415_),
    .Y(_2425_));
 sg13g2_and3_1 _2940_ (.X(_2426_),
    .A(_2388_),
    .B(_2385_),
    .C(_2415_));
 sg13g2_a221oi_1 _2941_ (.B2(_2425_),
    .C1(_2426_),
    .B1(_2387_),
    .A1(_2424_),
    .Y(_2427_),
    .A2(_2419_));
 sg13g2_and2_1 _2942_ (.A(_2399_),
    .B(_2427_),
    .X(_2428_));
 sg13g2_or3_1 _2943_ (.A(_2419_),
    .B(_2423_),
    .C(_2428_),
    .X(_2429_));
 sg13g2_nand3_1 _2944_ (.B(_2418_),
    .C(_2429_),
    .A(_2383_),
    .Y(_2430_));
 sg13g2_nand3b_1 _2945_ (.B(_2384_),
    .C(_2430_),
    .Y(_2431_),
    .A_N(_2348_));
 sg13g2_buf_2 _2946_ (.A(\g.g_y[6].g_x[6].t.r_h ),
    .X(_2432_));
 sg13g2_inv_1 _2947_ (.Y(_2433_),
    .A(_2432_));
 sg13g2_mux2_1 _2948_ (.A0(\g.g_y[6].g_x[6].t.out_sc ),
    .A1(\g.g_y[6].g_x[6].t.r_gnl ),
    .S(_2352_),
    .X(_2434_));
 sg13g2_buf_1 _2949_ (.A(_2434_),
    .X(_2435_));
 sg13g2_or2_1 _2950_ (.X(_2436_),
    .B(_2432_),
    .A(_2351_));
 sg13g2_o21ai_1 _2951_ (.B1(_2436_),
    .Y(_2437_),
    .A1(_2433_),
    .A2(_2435_));
 sg13g2_buf_1 _2952_ (.A(_2437_),
    .X(_2438_));
 sg13g2_buf_1 _2953_ (.A(\g.g_y[6].g_x[0].t.r_h ),
    .X(_2439_));
 sg13g2_mux2_1 _2954_ (.A0(\g.g_y[6].g_x[0].t.out_sc ),
    .A1(\g.g_y[6].g_x[0].t.r_gnl ),
    .S(_2409_),
    .X(_2440_));
 sg13g2_buf_1 _2955_ (.A(_2440_),
    .X(_2441_));
 sg13g2_nand2b_1 _2956_ (.Y(_2442_),
    .B(net85),
    .A_N(_2403_));
 sg13g2_o21ai_1 _2957_ (.B1(_2442_),
    .Y(_2443_),
    .A1(net85),
    .A2(_2441_));
 sg13g2_buf_2 _2958_ (.A(\g.g_y[5].g_x[7].t.r_v ),
    .X(_2444_));
 sg13g2_inv_1 _2959_ (.Y(_2445_),
    .A(_2444_));
 sg13g2_buf_2 _2960_ (.A(\g.g_y[5].g_x[7].t.r_d ),
    .X(_2446_));
 sg13g2_mux2_1 _2961_ (.A0(\g.g_y[5].g_x[7].t.r_gnl ),
    .A1(\g.g_y[5].g_x[7].t.out_sc ),
    .S(_2446_),
    .X(_2447_));
 sg13g2_buf_1 _2962_ (.A(_2447_),
    .X(_2448_));
 sg13g2_buf_1 _2963_ (.A(\g.g_y[5].g_x[7].t.r_ghl ),
    .X(_2449_));
 sg13g2_or2_1 _2964_ (.X(_2450_),
    .B(_2444_),
    .A(_2449_));
 sg13g2_o21ai_1 _2965_ (.B1(_2450_),
    .Y(_2451_),
    .A1(_2445_),
    .A2(_2448_));
 sg13g2_nor2_1 _2966_ (.A(_2451_),
    .B(_2443_),
    .Y(_2452_));
 sg13g2_nor2_1 _2967_ (.A(_2451_),
    .B(_2438_),
    .Y(_2453_));
 sg13g2_buf_2 _2968_ (.A(\g.g_y[6].g_x[7].t.r_h ),
    .X(_2454_));
 sg13g2_buf_1 _2969_ (.A(\g.g_y[6].g_x[7].t.r_v ),
    .X(_2455_));
 sg13g2_mux4_1 _2970_ (.S0(_2454_),
    .A0(_2438_),
    .A1(_2443_),
    .A2(_2452_),
    .A3(_2453_),
    .S1(net84),
    .X(_2456_));
 sg13g2_buf_2 _2971_ (.A(\g.g_y[7].g_x[7].t.r_v ),
    .X(_2457_));
 sg13g2_buf_1 _2972_ (.A(\g.g_y[6].g_x[7].t.r_d ),
    .X(_2458_));
 sg13g2_nor2_1 _2973_ (.A(_2457_),
    .B(net83),
    .Y(_2459_));
 sg13g2_buf_2 _2974_ (.A(\g.g_y[0].g_x[6].t.r_h ),
    .X(_2460_));
 sg13g2_inv_2 _2975_ (.Y(_2461_),
    .A(_2460_));
 sg13g2_mux2_1 _2976_ (.A0(\g.g_y[0].g_x[6].t.out_sc ),
    .A1(\g.g_y[0].g_x[6].t.r_gnl ),
    .S(_2357_),
    .X(_2462_));
 sg13g2_or2_1 _2977_ (.X(_2463_),
    .B(_2460_),
    .A(_2356_));
 sg13g2_o21ai_1 _2978_ (.B1(_2463_),
    .Y(_2464_),
    .A1(_2461_),
    .A2(_2462_));
 sg13g2_buf_1 _2979_ (.A(\g.g_y[0].g_x[0].t.r_h ),
    .X(_2465_));
 sg13g2_mux2_1 _2980_ (.A0(\g.g_y[0].g_x[0].t.out_sc ),
    .A1(\g.g_y[0].g_x[0].t.r_gnl ),
    .S(_2391_),
    .X(_2466_));
 sg13g2_buf_1 _2981_ (.A(_2466_),
    .X(_2467_));
 sg13g2_nand2b_1 _2982_ (.Y(_2468_),
    .B(net82),
    .A_N(_2400_));
 sg13g2_o21ai_1 _2983_ (.B1(_2468_),
    .Y(_2469_),
    .A1(net82),
    .A2(_2467_));
 sg13g2_buf_1 _2984_ (.A(_2469_),
    .X(_2470_));
 sg13g2_buf_2 _2985_ (.A(\g.g_y[1].g_x[7].t.r_v ),
    .X(_2471_));
 sg13g2_buf_2 _2986_ (.A(\g.g_y[1].g_x[7].t.r_d ),
    .X(_2472_));
 sg13g2_mux2_1 _2987_ (.A0(\g.g_y[1].g_x[7].t.r_gnl ),
    .A1(\g.g_y[1].g_x[7].t.out_sc ),
    .S(_2472_),
    .X(_2473_));
 sg13g2_buf_1 _2988_ (.A(_2473_),
    .X(_2474_));
 sg13g2_buf_1 _2989_ (.A(\g.g_y[1].g_x[7].t.r_ghl ),
    .X(_2475_));
 sg13g2_nand2b_1 _2990_ (.Y(_2476_),
    .B(_2471_),
    .A_N(_2475_));
 sg13g2_o21ai_1 _2991_ (.B1(_2476_),
    .Y(_2477_),
    .A1(_2471_),
    .A2(_2474_));
 sg13g2_buf_1 _2992_ (.A(_2477_),
    .X(_2478_));
 sg13g2_nor2_1 _2993_ (.A(_2478_),
    .B(_2470_),
    .Y(_2479_));
 sg13g2_nor2_1 _2994_ (.A(_2478_),
    .B(_2464_),
    .Y(_2480_));
 sg13g2_buf_2 _2995_ (.A(\g.g_y[0].g_x[7].t.r_h ),
    .X(_2481_));
 sg13g2_buf_2 _2996_ (.A(\g.g_y[0].g_x[7].t.r_v ),
    .X(_2482_));
 sg13g2_inv_2 _2997_ (.Y(_2483_),
    .A(_2482_));
 sg13g2_mux4_1 _2998_ (.S0(_2481_),
    .A0(_2464_),
    .A1(_2470_),
    .A2(_2479_),
    .A3(_2480_),
    .S1(_2483_),
    .X(_2484_));
 sg13g2_inv_1 _2999_ (.Y(_2485_),
    .A(_2457_));
 sg13g2_buf_1 _3000_ (.A(\g.g_y[0].g_x[7].t.r_d ),
    .X(_2486_));
 sg13g2_nor2_1 _3001_ (.A(_2485_),
    .B(net81),
    .Y(_2487_));
 sg13g2_o21ai_1 _3002_ (.B1(net83),
    .Y(_2488_),
    .A1(net84),
    .A2(_2451_));
 sg13g2_buf_2 _3003_ (.A(\g.g_y[6].g_x[7].t.out_sc ),
    .X(_2489_));
 sg13g2_a21o_1 _3004_ (.A2(_2489_),
    .A1(_2455_),
    .B1(_2457_),
    .X(_2490_));
 sg13g2_buf_1 _3005_ (.A(\g.g_y[0].g_x[7].t.out_sc ),
    .X(_2491_));
 sg13g2_nand2_1 _3006_ (.Y(_2492_),
    .A(_2457_),
    .B(net81));
 sg13g2_a21oi_1 _3007_ (.A1(_2483_),
    .A2(_2491_),
    .Y(_2493_),
    .B1(_2492_));
 sg13g2_o21ai_1 _3008_ (.B1(_2493_),
    .Y(_2494_),
    .A1(_2483_),
    .A2(_2478_));
 sg13g2_o21ai_1 _3009_ (.B1(_2494_),
    .Y(_2495_),
    .A1(_2488_),
    .A2(_2490_));
 sg13g2_a221oi_1 _3010_ (.B2(_2487_),
    .C1(_2495_),
    .B1(_2484_),
    .A1(_2456_),
    .Y(_2496_),
    .A2(_2459_));
 sg13g2_nand2_1 _3011_ (.Y(_2497_),
    .A(_2348_),
    .B(_2496_));
 sg13g2_buf_1 _3012_ (.A(rst_n),
    .X(_2498_));
 sg13g2_inv_2 _3013_ (.Y(_2499_),
    .A(net168));
 sg13g2_buf_1 _3014_ (.A(_2499_),
    .X(_2500_));
 sg13g2_buf_1 _3015_ (.A(net156),
    .X(_2501_));
 sg13g2_a21oi_1 _3016_ (.A1(_2431_),
    .A2(_2497_),
    .Y(_0133_),
    .B1(net139));
 sg13g2_inv_1 _3017_ (.Y(_2502_),
    .A(_2491_));
 sg13g2_inv_1 _3018_ (.Y(_2503_),
    .A(_2471_));
 sg13g2_mux2_1 _3019_ (.A0(_2475_),
    .A1(_2474_),
    .S(_2503_),
    .X(_2504_));
 sg13g2_mux2_1 _3020_ (.A0(\g.g_y[7].g_x[7].t.r_gnl ),
    .A1(\g.g_y[7].g_x[7].t.out_sc ),
    .S(_2348_),
    .X(_2505_));
 sg13g2_or2_1 _3021_ (.X(_2506_),
    .B(_2505_),
    .A(_2485_));
 sg13g2_buf_1 _3022_ (.A(_2506_),
    .X(_2507_));
 sg13g2_inv_1 _3023_ (.Y(_2508_),
    .A(\g.g_y[7].g_x[7].t.r_ghl ));
 sg13g2_a21oi_1 _3024_ (.A1(_2508_),
    .A2(_2485_),
    .Y(_2509_),
    .B1(_2483_));
 sg13g2_a22oi_1 _3025_ (.Y(_2510_),
    .B1(_2507_),
    .B2(_2509_),
    .A2(_2504_),
    .A1(_2483_));
 sg13g2_inv_1 _3026_ (.Y(_2511_),
    .A(_2481_));
 sg13g2_mux2_1 _3027_ (.A0(_2464_),
    .A1(_2470_),
    .S(_2511_),
    .X(_2512_));
 sg13g2_nor2_1 _3028_ (.A(_2510_),
    .B(_2512_),
    .Y(_2513_));
 sg13g2_mux2_1 _3029_ (.A0(_2356_),
    .A1(_2462_),
    .S(_2460_),
    .X(_2514_));
 sg13g2_inv_1 _3030_ (.Y(_2515_),
    .A(net82));
 sg13g2_nand2b_1 _3031_ (.Y(_2516_),
    .B(_2515_),
    .A_N(_2467_));
 sg13g2_and2_1 _3032_ (.A(_2481_),
    .B(_2468_),
    .X(_2517_));
 sg13g2_a22oi_1 _3033_ (.Y(_2518_),
    .B1(_2516_),
    .B2(_2517_),
    .A2(_2514_),
    .A1(_2511_));
 sg13g2_inv_1 _3034_ (.Y(_2519_),
    .A(net81));
 sg13g2_mux4_1 _3035_ (.S0(_2482_),
    .A0(_2502_),
    .A1(_2478_),
    .A2(_2513_),
    .A3(_2518_),
    .S1(_2519_),
    .X(_2520_));
 sg13g2_inv_1 _3036_ (.Y(_2521_),
    .A(_2455_));
 sg13g2_mux2_1 _3037_ (.A0(_2449_),
    .A1(_2448_),
    .S(_2444_),
    .X(_2522_));
 sg13g2_mux2_1 _3038_ (.A0(_2351_),
    .A1(_2435_),
    .S(_2432_),
    .X(_2523_));
 sg13g2_mux2_1 _3039_ (.A0(_2441_),
    .A1(_2403_),
    .S(net85),
    .X(_2524_));
 sg13g2_buf_1 _3040_ (.A(_2524_),
    .X(_2525_));
 sg13g2_mux2_1 _3041_ (.A0(_2523_),
    .A1(_2525_),
    .S(_2454_),
    .X(_2526_));
 sg13g2_inv_1 _3042_ (.Y(_2527_),
    .A(\g.g_y[6].g_x[7].t.r_d ));
 sg13g2_mux2_1 _3043_ (.A0(_2522_),
    .A1(_2526_),
    .S(_2527_),
    .X(_2528_));
 sg13g2_mux2_1 _3044_ (.A0(\g.g_y[7].g_x[7].t.r_ghl ),
    .A1(_2505_),
    .S(_2485_),
    .X(_2529_));
 sg13g2_buf_2 _3045_ (.A(_2529_),
    .X(_2530_));
 sg13g2_mux2_1 _3046_ (.A0(_2522_),
    .A1(_2530_),
    .S(_2521_),
    .X(_2531_));
 sg13g2_mux2_1 _3047_ (.A0(_2525_),
    .A1(_2523_),
    .S(_2454_),
    .X(_2532_));
 sg13g2_nand2_1 _3048_ (.Y(_2533_),
    .A(_2531_),
    .B(_2532_));
 sg13g2_nor2_1 _3049_ (.A(_2521_),
    .B(_2458_),
    .Y(_2534_));
 sg13g2_a22oi_1 _3050_ (.Y(_2535_),
    .B1(_2533_),
    .B2(_2534_),
    .A2(_2528_),
    .A1(_2521_));
 sg13g2_nand3_1 _3051_ (.B(net83),
    .C(_2489_),
    .A(net84),
    .Y(_2536_));
 sg13g2_and2_1 _3052_ (.A(_2457_),
    .B(_2536_),
    .X(_2537_));
 sg13g2_a22oi_1 _3053_ (.Y(_2538_),
    .B1(_2535_),
    .B2(_2537_),
    .A2(_2520_),
    .A1(_2485_));
 sg13g2_and2_1 _3054_ (.A(_2418_),
    .B(_2429_),
    .X(_2539_));
 sg13g2_nand3_1 _3055_ (.B(_2372_),
    .C(_2382_),
    .A(_2383_),
    .Y(_2540_));
 sg13g2_o21ai_1 _3056_ (.B1(_2540_),
    .Y(_2541_),
    .A1(_2383_),
    .A2(_2539_));
 sg13g2_a21oi_1 _3057_ (.A1(_2538_),
    .A2(_2541_),
    .Y(_0134_),
    .B1(net139));
 sg13g2_buf_1 _3058_ (.A(net168),
    .X(_2542_));
 sg13g2_buf_1 _3059_ (.A(net166),
    .X(_2543_));
 sg13g2_and2_1 _3060_ (.A(\g.g_y[7].g_x[7].t.out_sc ),
    .B(net155),
    .X(_0132_));
 sg13g2_inv_1 _3061_ (.Y(_2544_),
    .A(_2373_));
 sg13g2_buf_1 _3062_ (.A(_2499_),
    .X(_2545_));
 sg13g2_buf_1 _3063_ (.A(net154),
    .X(_2546_));
 sg13g2_nor2_1 _3064_ (.A(_2544_),
    .B(net138),
    .Y(_0131_));
 sg13g2_buf_2 _3065_ (.A(\g.g_y[0].g_x[5].t.r_v ),
    .X(_2547_));
 sg13g2_buf_2 _3066_ (.A(\g.g_y[1].g_x[5].t.r_ghl ),
    .X(_2548_));
 sg13g2_buf_8 _3067_ (.A(\g.g_y[1].g_x[5].t.r_d ),
    .X(_2549_));
 sg13g2_mux2_1 _3068_ (.A0(\g.g_y[1].g_x[5].t.r_gnl ),
    .A1(\g.g_y[1].g_x[5].t.out_sc ),
    .S(_2549_),
    .X(_2550_));
 sg13g2_buf_2 _3069_ (.A(\g.g_y[1].g_x[5].t.r_v ),
    .X(_2551_));
 sg13g2_inv_2 _3070_ (.Y(_2552_),
    .A(_2551_));
 sg13g2_mux2_1 _3071_ (.A0(_2548_),
    .A1(_2550_),
    .S(_2552_),
    .X(_2553_));
 sg13g2_inv_2 _3072_ (.Y(_2554_),
    .A(\g.g_y[7].g_x[5].t.r_v ));
 sg13g2_mux2_1 _3073_ (.A0(\g.g_y[7].g_x[5].t.r_gnl ),
    .A1(\g.g_y[7].g_x[5].t.out_sc ),
    .S(_2367_),
    .X(_2555_));
 sg13g2_or2_1 _3074_ (.X(_2556_),
    .B(_2555_),
    .A(_2554_));
 sg13g2_inv_1 _3075_ (.Y(_2557_),
    .A(_2366_));
 sg13g2_a21oi_1 _3076_ (.A1(_2557_),
    .A2(_2554_),
    .Y(_2558_),
    .B1(_2547_));
 sg13g2_buf_1 _3077_ (.A(\g.g_y[0].g_x[5].t.r_d ),
    .X(_2559_));
 sg13g2_inv_1 _3078_ (.Y(_2560_),
    .A(_2559_));
 sg13g2_a221oi_1 _3079_ (.B2(_2558_),
    .C1(_2560_),
    .B1(_2556_),
    .A1(_2547_),
    .Y(_2561_),
    .A2(_2553_));
 sg13g2_buf_2 _3080_ (.A(\g.g_y[0].g_x[4].t.r_h ),
    .X(_2562_));
 sg13g2_inv_1 _3081_ (.Y(_2563_),
    .A(_2562_));
 sg13g2_buf_8 _3082_ (.A(\g.g_y[0].g_x[4].t.r_d ),
    .X(_2564_));
 sg13g2_mux2_1 _3083_ (.A0(\g.g_y[0].g_x[4].t.out_sc ),
    .A1(\g.g_y[0].g_x[4].t.r_gnl ),
    .S(_2564_),
    .X(_2565_));
 sg13g2_or2_1 _3084_ (.X(_2566_),
    .B(_2565_),
    .A(_2563_));
 sg13g2_buf_1 _3085_ (.A(\g.g_y[0].g_x[4].t.r_ghl ),
    .X(_2567_));
 sg13g2_inv_1 _3086_ (.Y(_2568_),
    .A(_2567_));
 sg13g2_buf_1 _3087_ (.A(\g.g_y[0].g_x[5].t.r_h ),
    .X(_2569_));
 sg13g2_a21oi_1 _3088_ (.A1(_2568_),
    .A2(_2563_),
    .Y(_2570_),
    .B1(net80));
 sg13g2_mux2_1 _3089_ (.A0(_2356_),
    .A1(_2462_),
    .S(_2461_),
    .X(_2571_));
 sg13g2_a221oi_1 _3090_ (.B2(net80),
    .C1(_2559_),
    .B1(_2571_),
    .A1(_2566_),
    .Y(_2572_),
    .A2(_2570_));
 sg13g2_nor2_2 _3091_ (.A(_2561_),
    .B(_2572_),
    .Y(_2573_));
 sg13g2_mux2_1 _3092_ (.A0(_2366_),
    .A1(_2555_),
    .S(\g.g_y[7].g_x[5].t.r_v ),
    .X(_2574_));
 sg13g2_mux2_1 _3093_ (.A0(_2553_),
    .A1(_2574_),
    .S(_2547_),
    .X(_2575_));
 sg13g2_buf_1 _3094_ (.A(_2575_),
    .X(_2576_));
 sg13g2_mux2_1 _3095_ (.A0(_2567_),
    .A1(_2565_),
    .S(_2562_),
    .X(_2577_));
 sg13g2_inv_1 _3096_ (.Y(_2578_),
    .A(net80));
 sg13g2_mux2_1 _3097_ (.A0(_2577_),
    .A1(_2571_),
    .S(_2578_),
    .X(_2579_));
 sg13g2_buf_1 _3098_ (.A(_2579_),
    .X(_2580_));
 sg13g2_nand3_1 _3099_ (.B(_2576_),
    .C(_2580_),
    .A(_2560_),
    .Y(_2581_));
 sg13g2_nor2_1 _3100_ (.A(\g.g_y[0].g_x[5].t.out_sc ),
    .B(_2560_),
    .Y(_2582_));
 sg13g2_nor2_1 _3101_ (.A(_2547_),
    .B(_2582_),
    .Y(_2583_));
 sg13g2_a22oi_1 _3102_ (.Y(_2584_),
    .B1(_2581_),
    .B2(_2583_),
    .A2(_2573_),
    .A1(_2547_));
 sg13g2_buf_2 _3103_ (.A(\g.g_y[6].g_x[5].t.r_d ),
    .X(_2585_));
 sg13g2_inv_1 _3104_ (.Y(_2586_),
    .A(_2585_));
 sg13g2_buf_2 _3105_ (.A(\g.g_y[6].g_x[4].t.r_ghl ),
    .X(_2587_));
 sg13g2_buf_8 _3106_ (.A(\g.g_y[6].g_x[4].t.r_d ),
    .X(_2588_));
 sg13g2_mux2_1 _3107_ (.A0(\g.g_y[6].g_x[4].t.out_sc ),
    .A1(\g.g_y[6].g_x[4].t.r_gnl ),
    .S(_2588_),
    .X(_2589_));
 sg13g2_buf_1 _3108_ (.A(_2589_),
    .X(_2590_));
 sg13g2_buf_2 _3109_ (.A(\g.g_y[6].g_x[4].t.r_h ),
    .X(_2591_));
 sg13g2_mux2_1 _3110_ (.A0(_2587_),
    .A1(_2590_),
    .S(_2591_),
    .X(_2592_));
 sg13g2_mux2_1 _3111_ (.A0(_2351_),
    .A1(_2435_),
    .S(_2433_),
    .X(_2593_));
 sg13g2_buf_1 _3112_ (.A(_2593_),
    .X(_2594_));
 sg13g2_buf_1 _3113_ (.A(\g.g_y[6].g_x[5].t.r_h ),
    .X(_2595_));
 sg13g2_inv_2 _3114_ (.Y(_2596_),
    .A(_2595_));
 sg13g2_mux2_1 _3115_ (.A0(_2592_),
    .A1(_2594_),
    .S(_2596_),
    .X(_2597_));
 sg13g2_buf_1 _3116_ (.A(\g.g_y[5].g_x[5].t.r_ghl ),
    .X(_2598_));
 sg13g2_buf_8 _3117_ (.A(\g.g_y[5].g_x[5].t.r_d ),
    .X(_2599_));
 sg13g2_mux2_1 _3118_ (.A0(\g.g_y[5].g_x[5].t.r_gnl ),
    .A1(\g.g_y[5].g_x[5].t.out_sc ),
    .S(_2599_),
    .X(_2600_));
 sg13g2_buf_2 _3119_ (.A(\g.g_y[5].g_x[5].t.r_v ),
    .X(_2601_));
 sg13g2_mux2_1 _3120_ (.A0(_2598_),
    .A1(_2600_),
    .S(_2601_),
    .X(_2602_));
 sg13g2_mux2_1 _3121_ (.A0(_2366_),
    .A1(_2555_),
    .S(_2554_),
    .X(_2603_));
 sg13g2_buf_1 _3122_ (.A(_2603_),
    .X(_2604_));
 sg13g2_buf_1 _3123_ (.A(\g.g_y[6].g_x[5].t.r_v ),
    .X(_2605_));
 sg13g2_inv_1 _3124_ (.Y(_2606_),
    .A(_2605_));
 sg13g2_mux2_1 _3125_ (.A0(_2602_),
    .A1(_2604_),
    .S(_2606_),
    .X(_2607_));
 sg13g2_nand3_1 _3126_ (.B(_2597_),
    .C(_2607_),
    .A(_2586_),
    .Y(_2608_));
 sg13g2_nand2b_1 _3127_ (.Y(_2609_),
    .B(_2585_),
    .A_N(\g.g_y[6].g_x[5].t.out_sc ));
 sg13g2_and2_1 _3128_ (.A(_2605_),
    .B(_2609_),
    .X(_2610_));
 sg13g2_inv_1 _3129_ (.Y(_2611_),
    .A(_2598_));
 sg13g2_inv_2 _3130_ (.Y(_2612_),
    .A(_2601_));
 sg13g2_a21oi_1 _3131_ (.A1(_2611_),
    .A2(_2612_),
    .Y(_2613_),
    .B1(_2605_));
 sg13g2_or2_1 _3132_ (.X(_2614_),
    .B(_2600_),
    .A(_2612_));
 sg13g2_a221oi_1 _3133_ (.B2(_2614_),
    .C1(_2586_),
    .B1(_2613_),
    .A1(_2605_),
    .Y(_2615_),
    .A2(_2604_));
 sg13g2_inv_1 _3134_ (.Y(_2616_),
    .A(_2587_));
 sg13g2_inv_1 _3135_ (.Y(_2617_),
    .A(_2591_));
 sg13g2_a21oi_1 _3136_ (.A1(_2616_),
    .A2(_2617_),
    .Y(_2618_),
    .B1(_2595_));
 sg13g2_or2_1 _3137_ (.X(_2619_),
    .B(_2590_),
    .A(_2617_));
 sg13g2_a221oi_1 _3138_ (.B2(_2619_),
    .C1(_2585_),
    .B1(_2618_),
    .A1(_2595_),
    .Y(_2620_),
    .A2(_2594_));
 sg13g2_nor2_1 _3139_ (.A(_2615_),
    .B(_2620_),
    .Y(_2621_));
 sg13g2_a22oi_1 _3140_ (.Y(_2622_),
    .B1(_2621_),
    .B2(_2606_),
    .A2(_2610_),
    .A1(_2608_));
 sg13g2_mux2_1 _3141_ (.A0(_2584_),
    .A1(_2622_),
    .S(_2554_),
    .X(_2623_));
 sg13g2_nand2_1 _3142_ (.Y(_2624_),
    .A(_2367_),
    .B(net166));
 sg13g2_inv_1 _3143_ (.Y(_2625_),
    .A(_2367_));
 sg13g2_buf_8 _3144_ (.A(\g.g_y[7].g_x[4].t.r_h ),
    .X(_2626_));
 sg13g2_inv_4 _3145_ (.A(_2626_),
    .Y(_2627_));
 sg13g2_nor2_1 _3146_ (.A(net88),
    .B(_2627_),
    .Y(_2628_));
 sg13g2_buf_8 _3147_ (.A(\g.g_y[7].g_x[4].t.r_d ),
    .X(_2629_));
 sg13g2_inv_1 _3148_ (.Y(_2630_),
    .A(_2629_));
 sg13g2_buf_8 _3149_ (.A(\g.g_y[7].g_x[3].t.r_ghl ),
    .X(_2631_));
 sg13g2_buf_8 _3150_ (.A(\g.g_y[7].g_x[3].t.r_d ),
    .X(_2632_));
 sg13g2_mux2_1 _3151_ (.A0(\g.g_y[7].g_x[3].t.out_sc ),
    .A1(\g.g_y[7].g_x[3].t.r_gnl ),
    .S(_2632_),
    .X(_2633_));
 sg13g2_buf_1 _3152_ (.A(_2633_),
    .X(_2634_));
 sg13g2_buf_8 _3153_ (.A(\g.g_y[7].g_x[3].t.r_h ),
    .X(_2635_));
 sg13g2_mux2_1 _3154_ (.A0(_2631_),
    .A1(_2634_),
    .S(net79),
    .X(_2636_));
 sg13g2_buf_1 _3155_ (.A(_2636_),
    .X(_2637_));
 sg13g2_nand2b_1 _3156_ (.Y(_2638_),
    .B(net88),
    .A_N(_2366_));
 sg13g2_and2_1 _3157_ (.A(_2627_),
    .B(_2638_),
    .X(_2639_));
 sg13g2_or2_1 _3158_ (.X(_2640_),
    .B(_2368_),
    .A(net88));
 sg13g2_buf_1 _3159_ (.A(_2640_),
    .X(_2641_));
 sg13g2_a22oi_1 _3160_ (.Y(_2642_),
    .B1(_2639_),
    .B2(_2641_),
    .A2(_2637_),
    .A1(_2626_));
 sg13g2_buf_1 _3161_ (.A(\g.g_y[7].g_x[4].t.r_v ),
    .X(_2643_));
 sg13g2_inv_2 _3162_ (.Y(_2644_),
    .A(net78));
 sg13g2_mux2_1 _3163_ (.A0(\g.g_y[0].g_x[4].t.r_gnl ),
    .A1(\g.g_y[0].g_x[4].t.out_sc ),
    .S(_2564_),
    .X(_2645_));
 sg13g2_buf_1 _3164_ (.A(\g.g_y[0].g_x[4].t.r_v ),
    .X(_2646_));
 sg13g2_inv_1 _3165_ (.Y(_2647_),
    .A(_2646_));
 sg13g2_mux2_1 _3166_ (.A0(_2567_),
    .A1(_2645_),
    .S(_2647_),
    .X(_2648_));
 sg13g2_buf_1 _3167_ (.A(_2648_),
    .X(_2649_));
 sg13g2_buf_2 _3168_ (.A(\g.g_y[6].g_x[4].t.r_v ),
    .X(_2650_));
 sg13g2_inv_2 _3169_ (.Y(_2651_),
    .A(_2650_));
 sg13g2_mux2_1 _3170_ (.A0(\g.g_y[6].g_x[4].t.r_gnl ),
    .A1(\g.g_y[6].g_x[4].t.out_sc ),
    .S(_2588_),
    .X(_2652_));
 sg13g2_or2_1 _3171_ (.X(_2653_),
    .B(_2652_),
    .A(_2651_));
 sg13g2_buf_1 _3172_ (.A(_2653_),
    .X(_2654_));
 sg13g2_nor2_1 _3173_ (.A(_2587_),
    .B(_2650_),
    .Y(_2655_));
 sg13g2_nor2_1 _3174_ (.A(_2644_),
    .B(_2655_),
    .Y(_2656_));
 sg13g2_a22oi_1 _3175_ (.Y(_2657_),
    .B1(_2654_),
    .B2(_2656_),
    .A2(_2649_),
    .A1(_2644_));
 sg13g2_nor3_2 _3176_ (.A(_2630_),
    .B(_2642_),
    .C(_2657_),
    .Y(_2658_));
 sg13g2_and3_1 _3177_ (.X(_2659_),
    .A(net90),
    .B(net89),
    .C(_2378_));
 sg13g2_a22oi_1 _3178_ (.Y(_2660_),
    .B1(_2659_),
    .B2(net88),
    .A2(_2658_),
    .A1(_2628_));
 sg13g2_and2_1 _3179_ (.A(_2626_),
    .B(_2638_),
    .X(_2661_));
 sg13g2_buf_1 _3180_ (.A(_2661_),
    .X(_2662_));
 sg13g2_a221oi_1 _3181_ (.B2(_2627_),
    .C1(_2629_),
    .B1(_2637_),
    .A1(_2641_),
    .Y(_2663_),
    .A2(_2662_));
 sg13g2_buf_8 _3182_ (.A(_2663_),
    .X(_2664_));
 sg13g2_nor2_1 _3183_ (.A(net78),
    .B(_2655_),
    .Y(_2665_));
 sg13g2_a221oi_1 _3184_ (.B2(_2665_),
    .C1(_2630_),
    .B1(_2654_),
    .A1(net78),
    .Y(_2666_),
    .A2(_2649_));
 sg13g2_buf_8 _3185_ (.A(_2666_),
    .X(_2667_));
 sg13g2_nor2_1 _3186_ (.A(net88),
    .B(_2626_),
    .Y(_2668_));
 sg13g2_o21ai_1 _3187_ (.B1(_2668_),
    .Y(_2669_),
    .A1(_2664_),
    .A2(_2667_));
 sg13g2_mux2_1 _3188_ (.A0(\g.g_y[7].g_x[7].t.out_sc ),
    .A1(\g.g_y[7].g_x[7].t.r_gnl ),
    .S(_2348_),
    .X(_2670_));
 sg13g2_mux2_1 _3189_ (.A0(_2670_),
    .A1(\g.g_y[7].g_x[7].t.r_ghl ),
    .S(_2383_),
    .X(_2671_));
 sg13g2_buf_1 _3190_ (.A(_2671_),
    .X(_2672_));
 sg13g2_mux2_1 _3191_ (.A0(_2672_),
    .A1(_2371_),
    .S(net90),
    .X(_2673_));
 sg13g2_nor2b_1 _3192_ (.A(net90),
    .B_N(_2369_),
    .Y(_2674_));
 sg13g2_nand4_1 _3193_ (.B(_2365_),
    .C(_2673_),
    .A(net89),
    .Y(_2675_),
    .D(_2674_));
 sg13g2_buf_1 _3194_ (.A(\g.g_y[7].g_x[4].t.out_sc ),
    .X(_2676_));
 sg13g2_nor2_1 _3195_ (.A(_2629_),
    .B(_2676_),
    .Y(_2677_));
 sg13g2_o21ai_1 _3196_ (.B1(_2379_),
    .Y(_2678_),
    .A1(net90),
    .A2(_2544_));
 sg13g2_a21oi_1 _3197_ (.A1(net90),
    .A2(_2672_),
    .Y(_2679_),
    .B1(_2678_));
 sg13g2_a22oi_1 _3198_ (.Y(_2680_),
    .B1(_2679_),
    .B2(net88),
    .A2(_2628_),
    .A1(_2677_));
 sg13g2_and3_1 _3199_ (.X(_2681_),
    .A(_2669_),
    .B(_2675_),
    .C(_2680_));
 sg13g2_nand4_1 _3200_ (.B(_2542_),
    .C(_2660_),
    .A(_2625_),
    .Y(_2682_),
    .D(_2681_));
 sg13g2_o21ai_1 _3201_ (.B1(_2682_),
    .Y(_0129_),
    .A1(_2623_),
    .A2(_2624_));
 sg13g2_nand2_1 _3202_ (.Y(_2683_),
    .A(_2365_),
    .B(_2673_));
 sg13g2_mux2_1 _3203_ (.A0(_2355_),
    .A1(_2361_),
    .S(_2362_),
    .X(_2684_));
 sg13g2_mux4_1 _3204_ (.S0(net90),
    .A0(_2373_),
    .A1(_2672_),
    .A2(_2683_),
    .A3(_2684_),
    .S1(net89),
    .X(_2685_));
 sg13g2_o21ai_1 _3205_ (.B1(_2626_),
    .Y(_2686_),
    .A1(_2629_),
    .A2(_2676_));
 sg13g2_or3_1 _3206_ (.A(_2626_),
    .B(_2664_),
    .C(_2667_),
    .X(_2687_));
 sg13g2_o21ai_1 _3207_ (.B1(_2687_),
    .Y(_2688_),
    .A1(_2658_),
    .A2(_2686_));
 sg13g2_mux2_1 _3208_ (.A0(_2685_),
    .A1(_2688_),
    .S(net88),
    .X(_2689_));
 sg13g2_a221oi_1 _3209_ (.B2(_2606_),
    .C1(_2554_),
    .B1(_2621_),
    .A1(_2608_),
    .Y(_2690_),
    .A2(_2610_));
 sg13g2_a21oi_1 _3210_ (.A1(_2554_),
    .A2(_2584_),
    .Y(_2691_),
    .B1(_2690_));
 sg13g2_a21oi_1 _3211_ (.A1(_2689_),
    .A2(_2691_),
    .Y(_0130_),
    .B1(net139));
 sg13g2_buf_1 _3212_ (.A(_2542_),
    .X(_2692_));
 sg13g2_and2_1 _3213_ (.A(\g.g_y[7].g_x[5].t.out_sc ),
    .B(net153),
    .X(_0128_));
 sg13g2_and2_1 _3214_ (.A(_2676_),
    .B(net153),
    .X(_0127_));
 sg13g2_buf_1 _3215_ (.A(\g.g_y[0].g_x[3].t.r_d ),
    .X(_2693_));
 sg13g2_buf_1 _3216_ (.A(_2693_),
    .X(_2694_));
 sg13g2_buf_2 _3217_ (.A(\g.g_y[0].g_x[2].t.r_ghl ),
    .X(_2695_));
 sg13g2_buf_2 _3218_ (.A(\g.g_y[0].g_x[2].t.r_d ),
    .X(_2696_));
 sg13g2_mux2_1 _3219_ (.A0(\g.g_y[0].g_x[2].t.out_sc ),
    .A1(\g.g_y[0].g_x[2].t.r_gnl ),
    .S(_2696_),
    .X(_2697_));
 sg13g2_buf_1 _3220_ (.A(_2697_),
    .X(_2698_));
 sg13g2_buf_2 _3221_ (.A(\g.g_y[0].g_x[2].t.r_h ),
    .X(_2699_));
 sg13g2_mux2_1 _3222_ (.A0(_2695_),
    .A1(_2698_),
    .S(_2699_),
    .X(_2700_));
 sg13g2_buf_1 _3223_ (.A(_2700_),
    .X(_2701_));
 sg13g2_mux2_1 _3224_ (.A0(_2567_),
    .A1(_2565_),
    .S(_2563_),
    .X(_2702_));
 sg13g2_buf_1 _3225_ (.A(\g.g_y[0].g_x[3].t.r_h ),
    .X(_2703_));
 sg13g2_mux2_1 _3226_ (.A0(_2701_),
    .A1(_2702_),
    .S(net77),
    .X(_2704_));
 sg13g2_nand2b_1 _3227_ (.Y(_2705_),
    .B(_2704_),
    .A_N(net31));
 sg13g2_buf_1 _3228_ (.A(\g.g_y[1].g_x[3].t.r_ghl ),
    .X(_2706_));
 sg13g2_buf_8 _3229_ (.A(\g.g_y[1].g_x[3].t.r_d ),
    .X(_2707_));
 sg13g2_mux2_1 _3230_ (.A0(\g.g_y[1].g_x[3].t.r_gnl ),
    .A1(\g.g_y[1].g_x[3].t.out_sc ),
    .S(_2707_),
    .X(_2708_));
 sg13g2_buf_2 _3231_ (.A(\g.g_y[1].g_x[3].t.r_v ),
    .X(_2709_));
 sg13g2_inv_2 _3232_ (.Y(_2710_),
    .A(_2709_));
 sg13g2_mux2_1 _3233_ (.A0(_2706_),
    .A1(_2708_),
    .S(_2710_),
    .X(_2711_));
 sg13g2_buf_1 _3234_ (.A(_2711_),
    .X(_2712_));
 sg13g2_buf_1 _3235_ (.A(\g.g_y[7].g_x[3].t.r_v ),
    .X(_2713_));
 sg13g2_buf_2 _3236_ (.A(\g.g_y[0].g_x[3].t.r_v ),
    .X(_2714_));
 sg13g2_nand2_1 _3237_ (.Y(_2715_),
    .A(net76),
    .B(_2714_));
 sg13g2_a21oi_1 _3238_ (.A1(net31),
    .A2(_2712_),
    .Y(_2716_),
    .B1(_2715_));
 sg13g2_mux2_1 _3239_ (.A0(_2702_),
    .A1(_2701_),
    .S(net77),
    .X(_2717_));
 sg13g2_mux2_1 _3240_ (.A0(\g.g_y[7].g_x[3].t.r_gnl ),
    .A1(\g.g_y[7].g_x[3].t.out_sc ),
    .S(_2632_),
    .X(_2718_));
 sg13g2_buf_1 _3241_ (.A(_2718_),
    .X(_2719_));
 sg13g2_mux2_1 _3242_ (.A0(_2631_),
    .A1(_2719_),
    .S(net76),
    .X(_2720_));
 sg13g2_mux2_1 _3243_ (.A0(_2712_),
    .A1(_2720_),
    .S(_2714_),
    .X(_2721_));
 sg13g2_buf_1 _3244_ (.A(_2721_),
    .X(_2722_));
 sg13g2_and2_1 _3245_ (.A(_2717_),
    .B(_2722_),
    .X(_2723_));
 sg13g2_inv_1 _3246_ (.Y(_2724_),
    .A(_2714_));
 sg13g2_nand2_1 _3247_ (.Y(_2725_),
    .A(net76),
    .B(_2724_));
 sg13g2_nor2_1 _3248_ (.A(net31),
    .B(_2725_),
    .Y(_2726_));
 sg13g2_nand2b_1 _3249_ (.Y(_2727_),
    .B(_2693_),
    .A_N(\g.g_y[0].g_x[3].t.out_sc ));
 sg13g2_inv_1 _3250_ (.Y(_2728_),
    .A(_2713_));
 sg13g2_buf_1 _3251_ (.A(\g.g_y[6].g_x[3].t.r_v ),
    .X(_2729_));
 sg13g2_buf_2 _3252_ (.A(\g.g_y[6].g_x[3].t.r_d ),
    .X(_2730_));
 sg13g2_inv_2 _3253_ (.Y(_2731_),
    .A(_2730_));
 sg13g2_buf_2 _3254_ (.A(\g.g_y[6].g_x[3].t.out_sc ),
    .X(_2732_));
 sg13g2_nor2_1 _3255_ (.A(_2731_),
    .B(_2732_),
    .Y(_2733_));
 sg13g2_nand3_1 _3256_ (.B(_2729_),
    .C(_2733_),
    .A(_2728_),
    .Y(_2734_));
 sg13g2_o21ai_1 _3257_ (.B1(_2734_),
    .Y(_2735_),
    .A1(_2725_),
    .A2(_2727_));
 sg13g2_a221oi_1 _3258_ (.B2(_2726_),
    .C1(_2735_),
    .B1(_2723_),
    .A1(_2705_),
    .Y(_2736_),
    .A2(_2716_));
 sg13g2_nand2b_1 _3259_ (.Y(_2737_),
    .B(_2728_),
    .A_N(_2719_));
 sg13g2_nand2b_1 _3260_ (.Y(_2738_),
    .B(net76),
    .A_N(_2631_));
 sg13g2_and2_1 _3261_ (.A(_2729_),
    .B(_2738_),
    .X(_2739_));
 sg13g2_buf_1 _3262_ (.A(\g.g_y[5].g_x[3].t.r_v ),
    .X(_2740_));
 sg13g2_buf_2 _3263_ (.A(\g.g_y[5].g_x[3].t.r_d ),
    .X(_2741_));
 sg13g2_mux2_1 _3264_ (.A0(\g.g_y[5].g_x[3].t.r_gnl ),
    .A1(\g.g_y[5].g_x[3].t.out_sc ),
    .S(_2741_),
    .X(_2742_));
 sg13g2_buf_1 _3265_ (.A(\g.g_y[5].g_x[3].t.r_ghl ),
    .X(_2743_));
 sg13g2_nor2b_1 _3266_ (.A(net75),
    .B_N(_2743_),
    .Y(_2744_));
 sg13g2_a21o_1 _3267_ (.A2(_2742_),
    .A1(net75),
    .B1(_2744_),
    .X(_2745_));
 sg13g2_inv_1 _3268_ (.Y(_2746_),
    .A(_2729_));
 sg13g2_a221oi_1 _3269_ (.B2(_2746_),
    .C1(_2731_),
    .B1(_2745_),
    .A1(_2737_),
    .Y(_2747_),
    .A2(_2739_));
 sg13g2_nand2b_1 _3270_ (.Y(_2748_),
    .B(_2617_),
    .A_N(_2590_));
 sg13g2_buf_1 _3271_ (.A(\g.g_y[6].g_x[3].t.r_h ),
    .X(_2749_));
 sg13g2_nand2b_1 _3272_ (.Y(_2750_),
    .B(_2591_),
    .A_N(_2587_));
 sg13g2_and2_1 _3273_ (.A(net74),
    .B(_2750_),
    .X(_2751_));
 sg13g2_buf_2 _3274_ (.A(\g.g_y[6].g_x[2].t.r_ghl ),
    .X(_2752_));
 sg13g2_buf_8 _3275_ (.A(\g.g_y[6].g_x[2].t.r_d ),
    .X(_2753_));
 sg13g2_mux2_1 _3276_ (.A0(\g.g_y[6].g_x[2].t.out_sc ),
    .A1(\g.g_y[6].g_x[2].t.r_gnl ),
    .S(_2753_),
    .X(_2754_));
 sg13g2_mux2_1 _3277_ (.A0(_2752_),
    .A1(_2754_),
    .S(\g.g_y[6].g_x[2].t.r_h ),
    .X(_2755_));
 sg13g2_buf_2 _3278_ (.A(_2755_),
    .X(_2756_));
 sg13g2_inv_1 _3279_ (.Y(_2757_),
    .A(_2749_));
 sg13g2_a221oi_1 _3280_ (.B2(_2757_),
    .C1(_2730_),
    .B1(_2756_),
    .A1(_2748_),
    .Y(_2758_),
    .A2(_2751_));
 sg13g2_nor3_1 _3281_ (.A(_2729_),
    .B(_2747_),
    .C(_2758_),
    .Y(_2759_));
 sg13g2_mux2_1 _3282_ (.A0(_2587_),
    .A1(_2590_),
    .S(_2617_),
    .X(_2760_));
 sg13g2_mux2_1 _3283_ (.A0(_2760_),
    .A1(_2756_),
    .S(net74),
    .X(_2761_));
 sg13g2_a21oi_1 _3284_ (.A1(net75),
    .A2(_2742_),
    .Y(_2762_),
    .B1(_2744_));
 sg13g2_nor2_1 _3285_ (.A(_2730_),
    .B(_2762_),
    .Y(_2763_));
 sg13g2_a21oi_1 _3286_ (.A1(_2761_),
    .A2(_2763_),
    .Y(_2764_),
    .B1(_2746_));
 sg13g2_or3_1 _3287_ (.A(net76),
    .B(_2759_),
    .C(_2764_),
    .X(_2765_));
 sg13g2_inv_1 _3288_ (.Y(_2766_),
    .A(_2632_));
 sg13g2_a21oi_1 _3289_ (.A1(_2736_),
    .A2(_2765_),
    .Y(_2767_),
    .B1(_2766_));
 sg13g2_nand3b_1 _3290_ (.B(net79),
    .C(_2627_),
    .Y(_2768_),
    .A_N(_2677_));
 sg13g2_nand2_1 _3291_ (.Y(_2769_),
    .A(net79),
    .B(_2626_));
 sg13g2_or3_1 _3292_ (.A(_2664_),
    .B(_2667_),
    .C(_2769_),
    .X(_2770_));
 sg13g2_o21ai_1 _3293_ (.B1(_2770_),
    .Y(_2771_),
    .A1(_2658_),
    .A2(_2768_));
 sg13g2_buf_1 _3294_ (.A(\g.g_y[7].g_x[2].t.r_d ),
    .X(_2772_));
 sg13g2_inv_2 _3295_ (.Y(_2773_),
    .A(net73));
 sg13g2_or2_1 _3296_ (.X(_2774_),
    .B(_2634_),
    .A(net79));
 sg13g2_nand2b_1 _3297_ (.Y(_2775_),
    .B(net79),
    .A_N(_2631_));
 sg13g2_nor2b_1 _3298_ (.A(\g.g_y[7].g_x[2].t.r_h ),
    .B_N(_2775_),
    .Y(_2776_));
 sg13g2_mux2_1 _3299_ (.A0(_2388_),
    .A1(_2387_),
    .S(_2385_),
    .X(_2777_));
 sg13g2_buf_1 _3300_ (.A(\g.g_y[7].g_x[2].t.r_h ),
    .X(_2778_));
 sg13g2_a22oi_1 _3301_ (.Y(_2779_),
    .B1(_2777_),
    .B2(net72),
    .A2(_2776_),
    .A1(_2774_));
 sg13g2_buf_1 _3302_ (.A(_2779_),
    .X(_2780_));
 sg13g2_buf_1 _3303_ (.A(\g.g_y[6].g_x[2].t.r_v ),
    .X(_2781_));
 sg13g2_inv_1 _3304_ (.Y(_2782_),
    .A(_2781_));
 sg13g2_mux2_1 _3305_ (.A0(\g.g_y[6].g_x[2].t.r_gnl ),
    .A1(\g.g_y[6].g_x[2].t.out_sc ),
    .S(_2753_),
    .X(_2783_));
 sg13g2_buf_1 _3306_ (.A(_2783_),
    .X(_2784_));
 sg13g2_or2_1 _3307_ (.X(_2785_),
    .B(_2781_),
    .A(_2752_));
 sg13g2_o21ai_1 _3308_ (.B1(_2785_),
    .Y(_2786_),
    .A1(_2782_),
    .A2(_2784_));
 sg13g2_buf_2 _3309_ (.A(\g.g_y[0].g_x[2].t.r_v ),
    .X(_2787_));
 sg13g2_mux2_1 _3310_ (.A0(\g.g_y[0].g_x[2].t.r_gnl ),
    .A1(\g.g_y[0].g_x[2].t.out_sc ),
    .S(_2696_),
    .X(_2788_));
 sg13g2_buf_1 _3311_ (.A(_2788_),
    .X(_2789_));
 sg13g2_nand2b_1 _3312_ (.Y(_2790_),
    .B(_2787_),
    .A_N(_2695_));
 sg13g2_o21ai_1 _3313_ (.B1(_2790_),
    .Y(_2791_),
    .A1(_2787_),
    .A2(_2789_));
 sg13g2_buf_2 _3314_ (.A(\g.g_y[7].g_x[2].t.r_v ),
    .X(_2792_));
 sg13g2_inv_1 _3315_ (.Y(_2793_),
    .A(_2792_));
 sg13g2_mux2_1 _3316_ (.A0(_2786_),
    .A1(_2791_),
    .S(_2793_),
    .X(_2794_));
 sg13g2_buf_1 _3317_ (.A(_2794_),
    .X(_2795_));
 sg13g2_nor3_1 _3318_ (.A(_2773_),
    .B(_2780_),
    .C(_2795_),
    .Y(_0199_));
 sg13g2_buf_1 _3319_ (.A(\g.g_y[7].g_x[2].t.out_sc ),
    .X(_0200_));
 sg13g2_nor2b_1 _3320_ (.A(net79),
    .B_N(net72),
    .Y(_0201_));
 sg13g2_o21ai_1 _3321_ (.B1(_0201_),
    .Y(_0202_),
    .A1(net73),
    .A2(_0200_));
 sg13g2_nor2_1 _3322_ (.A(net73),
    .B(_2777_),
    .Y(_0203_));
 sg13g2_inv_1 _3323_ (.Y(_0204_),
    .A(_2787_));
 sg13g2_mux2_1 _3324_ (.A0(_2695_),
    .A1(_2789_),
    .S(_0204_),
    .X(_0205_));
 sg13g2_and2_1 _3325_ (.A(_2793_),
    .B(_2785_),
    .X(_0206_));
 sg13g2_or2_1 _3326_ (.X(_0207_),
    .B(_2784_),
    .A(_2782_));
 sg13g2_a221oi_1 _3327_ (.B2(_0207_),
    .C1(_2773_),
    .B1(_0206_),
    .A1(_2792_),
    .Y(_0208_),
    .A2(_0205_));
 sg13g2_or4_1 _3328_ (.A(net79),
    .B(net72),
    .C(_0203_),
    .D(_0208_),
    .X(_0209_));
 sg13g2_o21ai_1 _3329_ (.B1(_0209_),
    .Y(_0210_),
    .A1(_0199_),
    .A2(_0202_));
 sg13g2_nor3_1 _3330_ (.A(_2632_),
    .B(_2771_),
    .C(_0210_),
    .Y(_0211_));
 sg13g2_nor3_1 _3331_ (.A(net154),
    .B(_2767_),
    .C(_0211_),
    .Y(_0125_));
 sg13g2_nand2b_1 _3332_ (.Y(_0212_),
    .B(_2730_),
    .A_N(_2732_));
 sg13g2_a21oi_1 _3333_ (.A1(_0212_),
    .A2(_2764_),
    .Y(_0213_),
    .B1(_2759_));
 sg13g2_mux2_1 _3334_ (.A0(_2712_),
    .A1(_2720_),
    .S(_2724_),
    .X(_0214_));
 sg13g2_mux2_1 _3335_ (.A0(_2704_),
    .A1(_0214_),
    .S(_2693_),
    .X(_0215_));
 sg13g2_nand3b_1 _3336_ (.B(_2717_),
    .C(_2722_),
    .Y(_0216_),
    .A_N(net31));
 sg13g2_and2_1 _3337_ (.A(_2724_),
    .B(_2727_),
    .X(_0217_));
 sg13g2_a221oi_1 _3338_ (.B2(_0217_),
    .C1(net76),
    .B1(_0216_),
    .A1(_2714_),
    .Y(_0218_),
    .A2(_0215_));
 sg13g2_a21oi_1 _3339_ (.A1(net76),
    .A2(_0213_),
    .Y(_0219_),
    .B1(_0218_));
 sg13g2_or2_1 _3340_ (.X(_0220_),
    .B(_2677_),
    .A(_2626_));
 sg13g2_or3_1 _3341_ (.A(_2627_),
    .B(_2664_),
    .C(_2667_),
    .X(_0221_));
 sg13g2_o21ai_1 _3342_ (.B1(_0221_),
    .Y(_0222_),
    .A1(_2658_),
    .A2(_0220_));
 sg13g2_o21ai_1 _3343_ (.B1(net72),
    .Y(_0223_),
    .A1(net73),
    .A2(_0200_));
 sg13g2_or3_1 _3344_ (.A(net72),
    .B(_0203_),
    .C(_0208_),
    .X(_0224_));
 sg13g2_o21ai_1 _3345_ (.B1(_0224_),
    .Y(_0225_),
    .A1(_0199_),
    .A2(_0223_));
 sg13g2_mux2_1 _3346_ (.A0(_0222_),
    .A1(_0225_),
    .S(net79),
    .X(_0226_));
 sg13g2_a21oi_1 _3347_ (.A1(_0219_),
    .A2(_0226_),
    .Y(_0126_),
    .B1(net139));
 sg13g2_and2_1 _3348_ (.A(\g.g_y[7].g_x[3].t.out_sc ),
    .B(net153),
    .X(_0124_));
 sg13g2_inv_1 _3349_ (.Y(_0227_),
    .A(_0200_));
 sg13g2_nor2_1 _3350_ (.A(_0227_),
    .B(_2499_),
    .Y(_0123_));
 sg13g2_buf_1 _3351_ (.A(\g.g_y[7].g_x[1].t.r_v ),
    .X(_0228_));
 sg13g2_buf_2 _3352_ (.A(\g.g_y[1].g_x[1].t.r_v ),
    .X(_0229_));
 sg13g2_buf_2 _3353_ (.A(\g.g_y[1].g_x[1].t.r_d ),
    .X(_0230_));
 sg13g2_mux2_1 _3354_ (.A0(\g.g_y[1].g_x[1].t.r_gnl ),
    .A1(\g.g_y[1].g_x[1].t.out_sc ),
    .S(_0230_),
    .X(_0231_));
 sg13g2_buf_1 _3355_ (.A(_0231_),
    .X(_0232_));
 sg13g2_buf_2 _3356_ (.A(\g.g_y[1].g_x[1].t.r_ghl ),
    .X(_0233_));
 sg13g2_nand2b_1 _3357_ (.Y(_0234_),
    .B(_0229_),
    .A_N(_0233_));
 sg13g2_o21ai_1 _3358_ (.B1(_0234_),
    .Y(_0235_),
    .A1(_0229_),
    .A2(_0232_));
 sg13g2_inv_1 _3359_ (.Y(_0236_),
    .A(_2699_));
 sg13g2_nand2b_1 _3360_ (.Y(_0237_),
    .B(_0236_),
    .A_N(_2698_));
 sg13g2_buf_2 _3361_ (.A(\g.g_y[0].g_x[1].t.r_h ),
    .X(_0238_));
 sg13g2_inv_1 _3362_ (.Y(_0239_),
    .A(_0238_));
 sg13g2_buf_1 _3363_ (.A(\g.g_y[0].g_x[1].t.r_d ),
    .X(_0240_));
 sg13g2_inv_2 _3364_ (.Y(_0241_),
    .A(net70));
 sg13g2_nand2b_1 _3365_ (.Y(_0242_),
    .B(_2699_),
    .A_N(_2695_));
 sg13g2_and3_1 _3366_ (.X(_0243_),
    .A(_0239_),
    .B(_0241_),
    .C(_0242_));
 sg13g2_nor2_1 _3367_ (.A(_2400_),
    .B(net82),
    .Y(_0244_));
 sg13g2_nor3_1 _3368_ (.A(_0239_),
    .B(net70),
    .C(_0244_),
    .Y(_0245_));
 sg13g2_or2_1 _3369_ (.X(_0246_),
    .B(_2467_),
    .A(_2515_));
 sg13g2_buf_1 _3370_ (.A(_0246_),
    .X(_0247_));
 sg13g2_a22oi_1 _3371_ (.Y(_0248_),
    .B1(_0245_),
    .B2(_0247_),
    .A2(_0243_),
    .A1(_0237_));
 sg13g2_inv_1 _3372_ (.Y(_0249_),
    .A(\g.g_y[0].g_x[1].t.out_sc ));
 sg13g2_a21oi_1 _3373_ (.A1(_0249_),
    .A2(net70),
    .Y(_0250_),
    .B1(\g.g_y[0].g_x[1].t.r_v ));
 sg13g2_o21ai_1 _3374_ (.B1(_0250_),
    .Y(_0251_),
    .A1(_0235_),
    .A2(_0248_));
 sg13g2_mux2_1 _3375_ (.A0(_2695_),
    .A1(_2698_),
    .S(_0236_),
    .X(_0252_));
 sg13g2_nor2_1 _3376_ (.A(_0238_),
    .B(_0244_),
    .Y(_0253_));
 sg13g2_a221oi_1 _3377_ (.B2(_0247_),
    .C1(net70),
    .B1(_0253_),
    .A1(_0238_),
    .Y(_0254_),
    .A2(_0252_));
 sg13g2_inv_1 _3378_ (.Y(_0255_),
    .A(\g.g_y[0].g_x[1].t.r_v ));
 sg13g2_a21oi_1 _3379_ (.A1(net70),
    .A2(_0235_),
    .Y(_0256_),
    .B1(_0255_));
 sg13g2_nand2b_1 _3380_ (.Y(_0257_),
    .B(_0256_),
    .A_N(_0254_));
 sg13g2_nand3_1 _3381_ (.B(_0251_),
    .C(_0257_),
    .A(net71),
    .Y(_0258_));
 sg13g2_nor2b_1 _3382_ (.A(\g.g_y[6].g_x[0].t.r_h ),
    .B_N(_2403_),
    .Y(_0259_));
 sg13g2_a21oi_1 _3383_ (.A1(_2439_),
    .A2(_2441_),
    .Y(_0260_),
    .B1(_0259_));
 sg13g2_buf_1 _3384_ (.A(\g.g_y[6].g_x[2].t.r_h ),
    .X(_0261_));
 sg13g2_nand2b_1 _3385_ (.Y(_0262_),
    .B(net69),
    .A_N(_2752_));
 sg13g2_o21ai_1 _3386_ (.B1(_0262_),
    .Y(_0263_),
    .A1(net69),
    .A2(_2754_));
 sg13g2_buf_2 _3387_ (.A(\g.g_y[6].g_x[1].t.r_h ),
    .X(_0264_));
 sg13g2_inv_2 _3388_ (.Y(_0265_),
    .A(_0264_));
 sg13g2_mux2_1 _3389_ (.A0(_0260_),
    .A1(_0263_),
    .S(_0265_),
    .X(_0266_));
 sg13g2_buf_1 _3390_ (.A(_0266_),
    .X(_0267_));
 sg13g2_buf_1 _3391_ (.A(\g.g_y[6].g_x[1].t.r_d ),
    .X(_0268_));
 sg13g2_inv_1 _3392_ (.Y(_0269_),
    .A(_0268_));
 sg13g2_buf_2 _3393_ (.A(\g.g_y[5].g_x[1].t.r_v ),
    .X(_0270_));
 sg13g2_buf_2 _3394_ (.A(\g.g_y[5].g_x[1].t.r_d ),
    .X(_0271_));
 sg13g2_mux2_1 _3395_ (.A0(\g.g_y[5].g_x[1].t.r_gnl ),
    .A1(\g.g_y[5].g_x[1].t.out_sc ),
    .S(_0271_),
    .X(_0272_));
 sg13g2_buf_1 _3396_ (.A(_0272_),
    .X(_0273_));
 sg13g2_buf_1 _3397_ (.A(\g.g_y[5].g_x[1].t.r_ghl ),
    .X(_0274_));
 sg13g2_nor2b_1 _3398_ (.A(_0270_),
    .B_N(_0274_),
    .Y(_0275_));
 sg13g2_a21o_1 _3399_ (.A2(_0273_),
    .A1(_0270_),
    .B1(_0275_),
    .X(_0276_));
 sg13g2_nand2_1 _3400_ (.Y(_0277_),
    .A(net30),
    .B(_0276_));
 sg13g2_inv_1 _3401_ (.Y(_0278_),
    .A(\g.g_y[6].g_x[1].t.out_sc ));
 sg13g2_buf_2 _3402_ (.A(\g.g_y[6].g_x[1].t.r_v ),
    .X(_0279_));
 sg13g2_inv_1 _3403_ (.Y(_0280_),
    .A(_0279_));
 sg13g2_a21oi_1 _3404_ (.A1(net68),
    .A2(_0278_),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_o21ai_1 _3405_ (.B1(_0281_),
    .Y(_0282_),
    .A1(_0267_),
    .A2(_0277_));
 sg13g2_a21o_1 _3406_ (.A2(_2441_),
    .A1(_2439_),
    .B1(_0259_),
    .X(_0283_));
 sg13g2_buf_1 _3407_ (.A(_0283_),
    .X(_0284_));
 sg13g2_or2_1 _3408_ (.X(_0285_),
    .B(_2754_),
    .A(net69));
 sg13g2_and2_1 _3409_ (.A(_0264_),
    .B(_0262_),
    .X(_0286_));
 sg13g2_a221oi_1 _3410_ (.B2(_0286_),
    .C1(net68),
    .B1(_0285_),
    .A1(_0265_),
    .Y(_0287_),
    .A2(_0284_));
 sg13g2_a21oi_1 _3411_ (.A1(_0270_),
    .A2(_0273_),
    .Y(_0288_),
    .B1(_0275_));
 sg13g2_a21oi_1 _3412_ (.A1(net68),
    .A2(_0288_),
    .Y(_0289_),
    .B1(_0279_));
 sg13g2_nand2b_1 _3413_ (.Y(_0290_),
    .B(_0289_),
    .A_N(_0287_));
 sg13g2_nand3b_1 _3414_ (.B(_0282_),
    .C(_0290_),
    .Y(_0291_),
    .A_N(net71));
 sg13g2_nand3_1 _3415_ (.B(_0258_),
    .C(_0291_),
    .A(_2386_),
    .Y(_0292_));
 sg13g2_o21ai_1 _3416_ (.B1(_2775_),
    .Y(_0293_),
    .A1(_2635_),
    .A2(_2634_));
 sg13g2_nor4_1 _3417_ (.A(_2778_),
    .B(_2773_),
    .C(_0293_),
    .D(_2795_),
    .Y(_0294_));
 sg13g2_mux2_1 _3418_ (.A0(_2752_),
    .A1(_2784_),
    .S(_2781_),
    .X(_0295_));
 sg13g2_mux2_1 _3419_ (.A0(_0295_),
    .A1(_0205_),
    .S(_2792_),
    .X(_0296_));
 sg13g2_nand2_1 _3420_ (.Y(_0297_),
    .A(net72),
    .B(net73));
 sg13g2_nor2b_1 _3421_ (.A(net73),
    .B_N(_2778_),
    .Y(_0298_));
 sg13g2_nor3_1 _3422_ (.A(net72),
    .B(net73),
    .C(_0200_),
    .Y(_0299_));
 sg13g2_a21oi_1 _3423_ (.A1(_0293_),
    .A2(_0298_),
    .Y(_0300_),
    .B1(_0299_));
 sg13g2_o21ai_1 _3424_ (.B1(_0300_),
    .Y(_0301_),
    .A1(_0296_),
    .A2(_0297_));
 sg13g2_o21ai_1 _3425_ (.B1(_2385_),
    .Y(_0302_),
    .A1(_0294_),
    .A2(_0301_));
 sg13g2_inv_1 _3426_ (.Y(_0303_),
    .A(_2385_));
 sg13g2_nand3_1 _3427_ (.B(net86),
    .C(_2421_),
    .A(net87),
    .Y(_0304_));
 sg13g2_nor3_1 _3428_ (.A(net87),
    .B(_2399_),
    .C(_2405_),
    .Y(_0305_));
 sg13g2_a22oi_1 _3429_ (.Y(_0306_),
    .B1(_2413_),
    .B2(_0305_),
    .A2(_2399_),
    .A1(_2424_));
 sg13g2_and4_1 _3430_ (.A(_0303_),
    .B(_2419_),
    .C(_0304_),
    .D(_0306_),
    .X(_0307_));
 sg13g2_nand3_1 _3431_ (.B(_2424_),
    .C(_2415_),
    .A(_0303_),
    .Y(_0308_));
 sg13g2_nand2_1 _3432_ (.Y(_0309_),
    .A(_2416_),
    .B(_2425_));
 sg13g2_o21ai_1 _3433_ (.B1(_0309_),
    .Y(_0310_),
    .A1(_2414_),
    .A2(_0308_));
 sg13g2_nor3_1 _3434_ (.A(_2386_),
    .B(_0307_),
    .C(_0310_),
    .Y(_0311_));
 sg13g2_nand2_1 _3435_ (.Y(_0312_),
    .A(_0302_),
    .B(_0311_));
 sg13g2_buf_1 _3436_ (.A(net154),
    .X(_0313_));
 sg13g2_a21oi_1 _3437_ (.A1(_0292_),
    .A2(_0312_),
    .Y(_0121_),
    .B1(net137));
 sg13g2_nand3b_1 _3438_ (.B(_0251_),
    .C(_0257_),
    .Y(_0314_),
    .A_N(net71));
 sg13g2_nand3_1 _3439_ (.B(_0282_),
    .C(_0290_),
    .A(net71),
    .Y(_0315_));
 sg13g2_inv_1 _3440_ (.Y(_0316_),
    .A(_2424_));
 sg13g2_nor2_1 _3441_ (.A(_2419_),
    .B(_2416_),
    .Y(_0317_));
 sg13g2_o21ai_1 _3442_ (.B1(_0317_),
    .Y(_0318_),
    .A1(_0316_),
    .A2(_2414_));
 sg13g2_a21o_1 _3443_ (.A2(_0306_),
    .A1(_0304_),
    .B1(_2415_),
    .X(_0319_));
 sg13g2_nand3_1 _3444_ (.B(_0318_),
    .C(_0319_),
    .A(_2385_),
    .Y(_0320_));
 sg13g2_o21ai_1 _3445_ (.B1(_0303_),
    .Y(_0321_),
    .A1(_0294_),
    .A2(_0301_));
 sg13g2_nand4_1 _3446_ (.B(_0315_),
    .C(_0320_),
    .A(_0314_),
    .Y(_0322_),
    .D(_0321_));
 sg13g2_and2_1 _3447_ (.A(net155),
    .B(_0322_),
    .X(_0122_));
 sg13g2_and2_1 _3448_ (.A(\g.g_y[7].g_x[1].t.out_sc ),
    .B(_2692_),
    .X(_0120_));
 sg13g2_and2_1 _3449_ (.A(\g.g_y[7].g_x[0].t.out_sc ),
    .B(_2692_),
    .X(_0119_));
 sg13g2_and2_1 _3450_ (.A(_2489_),
    .B(net153),
    .X(_0118_));
 sg13g2_buf_1 _3451_ (.A(\g.g_y[5].g_x[6].t.r_d ),
    .X(_0323_));
 sg13g2_buf_1 _3452_ (.A(\g.g_y[4].g_x[6].t.r_ghl ),
    .X(_0324_));
 sg13g2_buf_2 _3453_ (.A(\g.g_y[4].g_x[6].t.r_v ),
    .X(_0325_));
 sg13g2_nor2_1 _3454_ (.A(_0324_),
    .B(_0325_),
    .Y(_0326_));
 sg13g2_inv_1 _3455_ (.Y(_0327_),
    .A(_0325_));
 sg13g2_buf_2 _3456_ (.A(\g.g_y[4].g_x[6].t.r_d ),
    .X(_0328_));
 sg13g2_mux2_1 _3457_ (.A0(\g.g_y[4].g_x[6].t.r_gnl ),
    .A1(\g.g_y[4].g_x[6].t.out_sc ),
    .S(_0328_),
    .X(_0329_));
 sg13g2_or2_1 _3458_ (.X(_0330_),
    .B(_0329_),
    .A(_0327_));
 sg13g2_buf_1 _3459_ (.A(_0330_),
    .X(_0331_));
 sg13g2_nand2b_1 _3460_ (.Y(_0332_),
    .B(_0331_),
    .A_N(_0326_));
 sg13g2_buf_1 _3461_ (.A(\g.g_y[5].g_x[6].t.r_h ),
    .X(_0333_));
 sg13g2_mux2_1 _3462_ (.A0(\g.g_y[5].g_x[7].t.out_sc ),
    .A1(\g.g_y[5].g_x[7].t.r_gnl ),
    .S(_2446_),
    .X(_0334_));
 sg13g2_buf_1 _3463_ (.A(\g.g_y[5].g_x[7].t.r_h ),
    .X(_0335_));
 sg13g2_mux2_1 _3464_ (.A0(_0334_),
    .A1(_2449_),
    .S(net65),
    .X(_0336_));
 sg13g2_buf_1 _3465_ (.A(_0336_),
    .X(_0337_));
 sg13g2_buf_2 _3466_ (.A(\g.g_y[5].g_x[5].t.r_h ),
    .X(_0338_));
 sg13g2_inv_2 _3467_ (.Y(_0339_),
    .A(_0338_));
 sg13g2_mux2_1 _3468_ (.A0(\g.g_y[5].g_x[5].t.out_sc ),
    .A1(\g.g_y[5].g_x[5].t.r_gnl ),
    .S(_2599_),
    .X(_0340_));
 sg13g2_or2_1 _3469_ (.X(_0341_),
    .B(_0340_),
    .A(_0339_));
 sg13g2_buf_1 _3470_ (.A(_0341_),
    .X(_0342_));
 sg13g2_nor2_1 _3471_ (.A(_2598_),
    .B(_0338_),
    .Y(_0343_));
 sg13g2_nor2_1 _3472_ (.A(net66),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_a221oi_1 _3473_ (.B2(_0344_),
    .C1(net67),
    .B1(_0342_),
    .A1(net66),
    .Y(_0345_),
    .A2(_0337_));
 sg13g2_a21o_1 _3474_ (.A2(_0332_),
    .A1(net67),
    .B1(_0345_),
    .X(_0346_));
 sg13g2_or2_1 _3475_ (.X(_0347_),
    .B(_0334_),
    .A(net65));
 sg13g2_inv_1 _3476_ (.Y(_0348_),
    .A(net66));
 sg13g2_inv_1 _3477_ (.Y(_0349_),
    .A(net67));
 sg13g2_nand2b_1 _3478_ (.Y(_0350_),
    .B(net65),
    .A_N(_2449_));
 sg13g2_and3_1 _3479_ (.X(_0351_),
    .A(_0348_),
    .B(_0349_),
    .C(_0350_));
 sg13g2_nor3_1 _3480_ (.A(_0348_),
    .B(net67),
    .C(_0343_),
    .Y(_0352_));
 sg13g2_a22oi_1 _3481_ (.Y(_0353_),
    .B1(_0352_),
    .B2(_0342_),
    .A2(_0351_),
    .A1(_0347_));
 sg13g2_nand2b_1 _3482_ (.Y(_0354_),
    .B(_0323_),
    .A_N(\g.g_y[5].g_x[6].t.out_sc ));
 sg13g2_o21ai_1 _3483_ (.B1(_0354_),
    .Y(_0355_),
    .A1(_0332_),
    .A2(_0353_));
 sg13g2_buf_1 _3484_ (.A(\g.g_y[5].g_x[6].t.r_v ),
    .X(_0356_));
 sg13g2_mux2_1 _3485_ (.A0(_0346_),
    .A1(_0355_),
    .S(net64),
    .X(_0357_));
 sg13g2_mux2_1 _3486_ (.A0(_2371_),
    .A1(_2672_),
    .S(\g.g_y[7].g_x[6].t.r_h ),
    .X(_0358_));
 sg13g2_mux2_1 _3487_ (.A0(_2684_),
    .A1(_0358_),
    .S(_2379_),
    .X(_0359_));
 sg13g2_buf_1 _3488_ (.A(_0359_),
    .X(_0360_));
 sg13g2_nand3_1 _3489_ (.B(_2365_),
    .C(_2673_),
    .A(_2379_),
    .Y(_0361_));
 sg13g2_buf_2 _3490_ (.A(_0361_),
    .X(_0362_));
 sg13g2_a21oi_1 _3491_ (.A1(net89),
    .A2(_2544_),
    .Y(_0363_),
    .B1(_2362_));
 sg13g2_a22oi_1 _3492_ (.Y(_0364_),
    .B1(_0362_),
    .B2(_0363_),
    .A2(_0360_),
    .A1(_2362_));
 sg13g2_mux2_1 _3493_ (.A0(_0357_),
    .A1(_0364_),
    .S(_2354_),
    .X(_0365_));
 sg13g2_nor2_1 _3494_ (.A(_2454_),
    .B(_2527_),
    .Y(_0366_));
 sg13g2_nor2_1 _3495_ (.A(_2454_),
    .B(\g.g_y[6].g_x[7].t.r_d ),
    .Y(_0367_));
 sg13g2_or2_1 _3496_ (.X(_0368_),
    .B(_2448_),
    .A(_2445_));
 sg13g2_and2_1 _3497_ (.A(_2521_),
    .B(_2450_),
    .X(_0369_));
 sg13g2_a221oi_1 _3498_ (.B2(net84),
    .C1(_2527_),
    .B1(_2530_),
    .A1(_0368_),
    .Y(_0370_),
    .A2(_0369_));
 sg13g2_o21ai_1 _3499_ (.B1(_2454_),
    .Y(_0371_),
    .A1(net83),
    .A2(_2525_));
 sg13g2_nor2_1 _3500_ (.A(_0370_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_a221oi_1 _3501_ (.B2(_2489_),
    .C1(_0372_),
    .B1(_0367_),
    .A1(_2533_),
    .Y(_0373_),
    .A2(_0366_));
 sg13g2_nand2b_1 _3502_ (.Y(_0374_),
    .B(_2432_),
    .A_N(_0373_));
 sg13g2_nand3_1 _3503_ (.B(_2597_),
    .C(_2607_),
    .A(_2585_),
    .Y(_0375_));
 sg13g2_nor2_1 _3504_ (.A(_2585_),
    .B(\g.g_y[6].g_x[5].t.out_sc ),
    .Y(_0376_));
 sg13g2_nor3_1 _3505_ (.A(_2432_),
    .B(_2596_),
    .C(_0376_),
    .Y(_0377_));
 sg13g2_nor2_1 _3506_ (.A(_2585_),
    .B(_2592_),
    .Y(_0378_));
 sg13g2_nor3_1 _3507_ (.A(_2432_),
    .B(_2595_),
    .C(_0378_),
    .Y(_0379_));
 sg13g2_a22oi_1 _3508_ (.Y(_0380_),
    .B1(_2613_),
    .B2(_2614_),
    .A2(_2604_),
    .A1(_2605_));
 sg13g2_nand2_1 _3509_ (.Y(_0381_),
    .A(_2585_),
    .B(_0380_));
 sg13g2_a221oi_1 _3510_ (.B2(_0381_),
    .C1(_2352_),
    .B1(_0379_),
    .A1(_0375_),
    .Y(_0382_),
    .A2(_0377_));
 sg13g2_a221oi_1 _3511_ (.B2(_0382_),
    .C1(net154),
    .B1(_0374_),
    .A1(_2352_),
    .Y(_0116_),
    .A2(_0365_));
 sg13g2_nor2_1 _3512_ (.A(_2596_),
    .B(_0376_),
    .Y(_0383_));
 sg13g2_a221oi_1 _3513_ (.B2(_0383_),
    .C1(_2433_),
    .B1(_0375_),
    .A1(_2596_),
    .Y(_0384_),
    .A2(_2621_));
 sg13g2_a21oi_1 _3514_ (.A1(_2433_),
    .A2(_0373_),
    .Y(_0385_),
    .B1(_0384_));
 sg13g2_a221oi_1 _3515_ (.B2(_0363_),
    .C1(_2354_),
    .B1(_0362_),
    .A1(_2362_),
    .Y(_0386_),
    .A2(_0360_));
 sg13g2_a21oi_1 _3516_ (.A1(_2354_),
    .A2(_0357_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_a21oi_1 _3517_ (.A1(_0385_),
    .A2(_0387_),
    .Y(_0117_),
    .B1(net137));
 sg13g2_and2_1 _3518_ (.A(\g.g_y[6].g_x[6].t.out_sc ),
    .B(net153),
    .X(_0115_));
 sg13g2_and2_1 _3519_ (.A(\g.g_y[6].g_x[5].t.out_sc ),
    .B(net153),
    .X(_0114_));
 sg13g2_buf_1 _3520_ (.A(\g.g_y[5].g_x[4].t.r_d ),
    .X(_0388_));
 sg13g2_inv_2 _3521_ (.Y(_0389_),
    .A(net63));
 sg13g2_buf_1 _3522_ (.A(\g.g_y[5].g_x[4].t.out_sc ),
    .X(_0390_));
 sg13g2_nor2_1 _3523_ (.A(_0389_),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_buf_1 _3524_ (.A(\g.g_y[5].g_x[4].t.r_v ),
    .X(_0392_));
 sg13g2_inv_1 _3525_ (.Y(_0393_),
    .A(_0392_));
 sg13g2_mux2_1 _3526_ (.A0(_2587_),
    .A1(_2652_),
    .S(_2651_),
    .X(_0394_));
 sg13g2_buf_1 _3527_ (.A(_0394_),
    .X(_0395_));
 sg13g2_buf_2 _3528_ (.A(\g.g_y[4].g_x[4].t.r_v ),
    .X(_0396_));
 sg13g2_inv_1 _3529_ (.Y(_0397_),
    .A(_0396_));
 sg13g2_buf_8 _3530_ (.A(\g.g_y[4].g_x[4].t.r_d ),
    .X(_0398_));
 sg13g2_mux2_1 _3531_ (.A0(\g.g_y[4].g_x[4].t.r_gnl ),
    .A1(\g.g_y[4].g_x[4].t.out_sc ),
    .S(_0398_),
    .X(_0399_));
 sg13g2_buf_1 _3532_ (.A(_0399_),
    .X(_0400_));
 sg13g2_or2_1 _3533_ (.X(_0401_),
    .B(_0400_),
    .A(_0397_));
 sg13g2_buf_1 _3534_ (.A(_0401_),
    .X(_0402_));
 sg13g2_buf_2 _3535_ (.A(\g.g_y[4].g_x[4].t.r_ghl ),
    .X(_0403_));
 sg13g2_nor2_1 _3536_ (.A(_0403_),
    .B(_0396_),
    .Y(_0404_));
 sg13g2_nor2_1 _3537_ (.A(_0393_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_a22oi_1 _3538_ (.Y(_0406_),
    .B1(_0402_),
    .B2(_0405_),
    .A2(_0395_),
    .A1(_0393_));
 sg13g2_buf_2 _3539_ (.A(\g.g_y[5].g_x[4].t.r_h ),
    .X(_0407_));
 sg13g2_inv_2 _3540_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_mux2_1 _3541_ (.A0(_2598_),
    .A1(_0340_),
    .S(_0339_),
    .X(_0409_));
 sg13g2_buf_1 _3542_ (.A(_0409_),
    .X(_0410_));
 sg13g2_buf_2 _3543_ (.A(\g.g_y[5].g_x[3].t.r_h ),
    .X(_0411_));
 sg13g2_inv_1 _3544_ (.Y(_0412_),
    .A(_0411_));
 sg13g2_mux2_1 _3545_ (.A0(\g.g_y[5].g_x[3].t.out_sc ),
    .A1(\g.g_y[5].g_x[3].t.r_gnl ),
    .S(_2741_),
    .X(_0413_));
 sg13g2_or2_1 _3546_ (.X(_0414_),
    .B(_0413_),
    .A(_0412_));
 sg13g2_nor2_1 _3547_ (.A(_2743_),
    .B(_0411_),
    .Y(_0415_));
 sg13g2_nor2_1 _3548_ (.A(_0408_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_a22oi_1 _3549_ (.Y(_0417_),
    .B1(_0414_),
    .B2(_0416_),
    .A2(_0410_),
    .A1(_0408_));
 sg13g2_buf_1 _3550_ (.A(_0417_),
    .X(_0418_));
 sg13g2_nor3_1 _3551_ (.A(net63),
    .B(_0406_),
    .C(_0418_),
    .Y(_0419_));
 sg13g2_nor2_1 _3552_ (.A(_2650_),
    .B(_0393_),
    .Y(_0420_));
 sg13g2_o21ai_1 _3553_ (.B1(_0420_),
    .Y(_0421_),
    .A1(_0391_),
    .A2(_0419_));
 sg13g2_nor2_1 _3554_ (.A(_2650_),
    .B(_0392_),
    .Y(_0422_));
 sg13g2_nor2_1 _3555_ (.A(_0407_),
    .B(_0415_),
    .Y(_0423_));
 sg13g2_a221oi_1 _3556_ (.B2(_0423_),
    .C1(_0388_),
    .B1(_0414_),
    .A1(_0407_),
    .Y(_0424_),
    .A2(_0410_));
 sg13g2_nor2_1 _3557_ (.A(net62),
    .B(_0404_),
    .Y(_0425_));
 sg13g2_a221oi_1 _3558_ (.B2(_0425_),
    .C1(_0389_),
    .B1(_0402_),
    .A1(net62),
    .Y(_0426_),
    .A2(_0395_));
 sg13g2_or2_1 _3559_ (.X(_0427_),
    .B(_0426_),
    .A(_0424_));
 sg13g2_nor3_1 _3560_ (.A(_2651_),
    .B(net78),
    .C(_2629_),
    .Y(_0428_));
 sg13g2_nor2_1 _3561_ (.A(_2642_),
    .B(_2657_),
    .Y(_0429_));
 sg13g2_nand2b_1 _3562_ (.Y(_0430_),
    .B(_2629_),
    .A_N(_2676_));
 sg13g2_nor3_1 _3563_ (.A(_2651_),
    .B(net78),
    .C(_0430_),
    .Y(_0431_));
 sg13g2_nand3_1 _3564_ (.B(_2643_),
    .C(_2630_),
    .A(_2650_),
    .Y(_0432_));
 sg13g2_a221oi_1 _3565_ (.B2(_2627_),
    .C1(_0432_),
    .B1(_2637_),
    .A1(_2641_),
    .Y(_0433_),
    .A2(_2662_));
 sg13g2_nor4_1 _3566_ (.A(_2651_),
    .B(_2644_),
    .C(_2630_),
    .D(_2649_),
    .Y(_0434_));
 sg13g2_or3_1 _3567_ (.A(_0431_),
    .B(_0433_),
    .C(_0434_),
    .X(_0435_));
 sg13g2_a221oi_1 _3568_ (.B2(_0429_),
    .C1(_0435_),
    .B1(_0428_),
    .A1(_0422_),
    .Y(_0436_),
    .A2(_0427_));
 sg13g2_nand3_1 _3569_ (.B(_0421_),
    .C(_0436_),
    .A(_2588_),
    .Y(_0437_));
 sg13g2_and2_1 _3570_ (.A(_2757_),
    .B(_2750_),
    .X(_0438_));
 sg13g2_a22oi_1 _3571_ (.Y(_0439_),
    .B1(_0438_),
    .B2(_2748_),
    .A2(_2756_),
    .A1(_2749_));
 sg13g2_buf_1 _3572_ (.A(_0439_),
    .X(_0440_));
 sg13g2_o21ai_1 _3573_ (.B1(_2738_),
    .Y(_0441_),
    .A1(net76),
    .A2(_2719_));
 sg13g2_mux2_1 _3574_ (.A0(_0441_),
    .A1(_2762_),
    .S(_2729_),
    .X(_0442_));
 sg13g2_or4_1 _3575_ (.A(_2757_),
    .B(_2731_),
    .C(_0440_),
    .D(_0442_),
    .X(_0443_));
 sg13g2_nor2_1 _3576_ (.A(_2730_),
    .B(_2732_),
    .Y(_0444_));
 sg13g2_nor2_1 _3577_ (.A(net74),
    .B(_2731_),
    .Y(_0445_));
 sg13g2_a22oi_1 _3578_ (.Y(_0446_),
    .B1(_2745_),
    .B2(_2746_),
    .A2(_2739_),
    .A1(_2737_));
 sg13g2_nor3_1 _3579_ (.A(net74),
    .B(_2730_),
    .C(_2756_),
    .Y(_0447_));
 sg13g2_a221oi_1 _3580_ (.B2(_0446_),
    .C1(_0447_),
    .B1(_0445_),
    .A1(net74),
    .Y(_0448_),
    .A2(_0444_));
 sg13g2_a21o_1 _3581_ (.A2(_0448_),
    .A1(_0443_),
    .B1(_2591_),
    .X(_0449_));
 sg13g2_and4_1 _3582_ (.A(_2596_),
    .B(_2585_),
    .C(_2594_),
    .D(_2607_),
    .X(_0450_));
 sg13g2_nor2_1 _3583_ (.A(_2596_),
    .B(_2586_),
    .Y(_0451_));
 sg13g2_nand2_1 _3584_ (.Y(_0452_),
    .A(_2595_),
    .B(_2586_));
 sg13g2_nand2_1 _3585_ (.Y(_0453_),
    .A(_2596_),
    .B(_0376_));
 sg13g2_o21ai_1 _3586_ (.B1(_0453_),
    .Y(_0454_),
    .A1(_2594_),
    .A2(_0452_));
 sg13g2_a21o_1 _3587_ (.A2(_0451_),
    .A1(_0380_),
    .B1(_0454_),
    .X(_0455_));
 sg13g2_o21ai_1 _3588_ (.B1(_2591_),
    .Y(_0456_),
    .A1(_0450_),
    .A2(_0455_));
 sg13g2_nand3b_1 _3589_ (.B(_0449_),
    .C(_0456_),
    .Y(_0457_),
    .A_N(_2588_));
 sg13g2_a21oi_1 _3590_ (.A1(_0437_),
    .A2(_0457_),
    .Y(_0112_),
    .B1(net137));
 sg13g2_a21oi_1 _3591_ (.A1(_0443_),
    .A2(_0448_),
    .Y(_0458_),
    .B1(_2617_));
 sg13g2_o21ai_1 _3592_ (.B1(_2617_),
    .Y(_0459_),
    .A1(_0450_),
    .A2(_0455_));
 sg13g2_nor2b_1 _3593_ (.A(_0458_),
    .B_N(_0459_),
    .Y(_0460_));
 sg13g2_nor2_1 _3594_ (.A(_2664_),
    .B(_2667_),
    .Y(_0461_));
 sg13g2_or3_1 _3595_ (.A(_2629_),
    .B(_2642_),
    .C(_2657_),
    .X(_0462_));
 sg13g2_buf_1 _3596_ (.A(_0462_),
    .X(_0463_));
 sg13g2_and2_1 _3597_ (.A(_2644_),
    .B(_0430_),
    .X(_0464_));
 sg13g2_a22oi_1 _3598_ (.Y(_0465_),
    .B1(_0463_),
    .B2(_0464_),
    .A2(_0461_),
    .A1(net78));
 sg13g2_or3_1 _3599_ (.A(_0393_),
    .B(_0391_),
    .C(_0419_),
    .X(_0466_));
 sg13g2_nor3_1 _3600_ (.A(net62),
    .B(_0424_),
    .C(_0426_),
    .Y(_0467_));
 sg13g2_nor2_1 _3601_ (.A(_2651_),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_a22oi_1 _3602_ (.Y(_0469_),
    .B1(_0466_),
    .B2(_0468_),
    .A2(_0465_),
    .A1(_2651_));
 sg13g2_a21oi_1 _3603_ (.A1(_0460_),
    .A2(_0469_),
    .Y(_0113_),
    .B1(net137));
 sg13g2_and2_1 _3604_ (.A(\g.g_y[6].g_x[4].t.out_sc ),
    .B(net153),
    .X(_0111_));
 sg13g2_and2_1 _3605_ (.A(_2732_),
    .B(net153),
    .X(_0110_));
 sg13g2_nor2_1 _3606_ (.A(_2780_),
    .B(_2795_),
    .Y(_0470_));
 sg13g2_mux2_1 _3607_ (.A0(_2634_),
    .A1(_2631_),
    .S(_2635_),
    .X(_0471_));
 sg13g2_mux2_1 _3608_ (.A0(_2777_),
    .A1(_0471_),
    .S(net72),
    .X(_0472_));
 sg13g2_inv_1 _3609_ (.Y(_0473_),
    .A(_0472_));
 sg13g2_mux4_1 _3610_ (.S0(_2792_),
    .A0(_0227_),
    .A1(_2791_),
    .A2(_0470_),
    .A3(_0473_),
    .S1(_2773_),
    .X(_0474_));
 sg13g2_buf_1 _3611_ (.A(\g.g_y[5].g_x[2].t.r_d ),
    .X(_0475_));
 sg13g2_inv_1 _3612_ (.Y(_0476_),
    .A(_0475_));
 sg13g2_buf_2 _3613_ (.A(\g.g_y[4].g_x[2].t.r_ghl ),
    .X(_0477_));
 sg13g2_buf_8 _3614_ (.A(\g.g_y[4].g_x[2].t.r_d ),
    .X(_0478_));
 sg13g2_mux2_1 _3615_ (.A0(\g.g_y[4].g_x[2].t.r_gnl ),
    .A1(\g.g_y[4].g_x[2].t.out_sc ),
    .S(_0478_),
    .X(_0479_));
 sg13g2_buf_2 _3616_ (.A(\g.g_y[4].g_x[2].t.r_v ),
    .X(_0480_));
 sg13g2_mux2_1 _3617_ (.A0(_0477_),
    .A1(_0479_),
    .S(_0480_),
    .X(_0481_));
 sg13g2_mux2_1 _3618_ (.A0(_2752_),
    .A1(_2784_),
    .S(_2782_),
    .X(_0482_));
 sg13g2_buf_2 _3619_ (.A(_0482_),
    .X(_0483_));
 sg13g2_buf_1 _3620_ (.A(\g.g_y[5].g_x[2].t.r_v ),
    .X(_0484_));
 sg13g2_inv_1 _3621_ (.Y(_0485_),
    .A(_0484_));
 sg13g2_mux2_1 _3622_ (.A0(_0481_),
    .A1(_0483_),
    .S(_0485_),
    .X(_0486_));
 sg13g2_mux2_1 _3623_ (.A0(\g.g_y[5].g_x[1].t.out_sc ),
    .A1(\g.g_y[5].g_x[1].t.r_gnl ),
    .S(_0271_),
    .X(_0487_));
 sg13g2_buf_1 _3624_ (.A(_0487_),
    .X(_0488_));
 sg13g2_buf_2 _3625_ (.A(\g.g_y[5].g_x[1].t.r_h ),
    .X(_0489_));
 sg13g2_mux2_1 _3626_ (.A0(_0274_),
    .A1(_0488_),
    .S(_0489_),
    .X(_0490_));
 sg13g2_mux2_1 _3627_ (.A0(_2743_),
    .A1(_0413_),
    .S(_0412_),
    .X(_0491_));
 sg13g2_buf_2 _3628_ (.A(_0491_),
    .X(_0492_));
 sg13g2_buf_2 _3629_ (.A(\g.g_y[5].g_x[2].t.r_h ),
    .X(_0493_));
 sg13g2_inv_1 _3630_ (.Y(_0494_),
    .A(_0493_));
 sg13g2_mux2_1 _3631_ (.A0(_0490_),
    .A1(_0492_),
    .S(_0494_),
    .X(_0495_));
 sg13g2_nand3_1 _3632_ (.B(_0486_),
    .C(_0495_),
    .A(_0476_),
    .Y(_0496_));
 sg13g2_nand2b_1 _3633_ (.Y(_0497_),
    .B(_0475_),
    .A_N(\g.g_y[5].g_x[2].t.out_sc ));
 sg13g2_and2_1 _3634_ (.A(_0484_),
    .B(_0497_),
    .X(_0498_));
 sg13g2_inv_1 _3635_ (.Y(_0499_),
    .A(_0477_));
 sg13g2_inv_2 _3636_ (.Y(_0500_),
    .A(_0480_));
 sg13g2_a21oi_1 _3637_ (.A1(_0499_),
    .A2(_0500_),
    .Y(_0501_),
    .B1(_0484_));
 sg13g2_or2_1 _3638_ (.X(_0502_),
    .B(_0479_),
    .A(_0500_));
 sg13g2_buf_1 _3639_ (.A(_0502_),
    .X(_0503_));
 sg13g2_a221oi_1 _3640_ (.B2(_0503_),
    .C1(_0476_),
    .B1(_0501_),
    .A1(_0484_),
    .Y(_0504_),
    .A2(_0483_));
 sg13g2_inv_1 _3641_ (.Y(_0505_),
    .A(_0274_));
 sg13g2_inv_1 _3642_ (.Y(_0506_),
    .A(_0489_));
 sg13g2_a21oi_1 _3643_ (.A1(_0505_),
    .A2(_0506_),
    .Y(_0507_),
    .B1(_0493_));
 sg13g2_or2_1 _3644_ (.X(_0508_),
    .B(_0488_),
    .A(_0506_));
 sg13g2_buf_1 _3645_ (.A(_0475_),
    .X(_0509_));
 sg13g2_a221oi_1 _3646_ (.B2(_0508_),
    .C1(net29),
    .B1(_0507_),
    .A1(_0493_),
    .Y(_0510_),
    .A2(_0492_));
 sg13g2_nor2_1 _3647_ (.A(_0504_),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_a221oi_1 _3648_ (.B2(_0485_),
    .C1(_2781_),
    .B1(_0511_),
    .A1(_0496_),
    .Y(_0512_),
    .A2(_0498_));
 sg13g2_a21o_1 _3649_ (.A2(_0474_),
    .A1(_2781_),
    .B1(_0512_),
    .X(_0513_));
 sg13g2_nand2_1 _3650_ (.Y(_0514_),
    .A(_2753_),
    .B(net168));
 sg13g2_buf_8 _3651_ (.A(net168),
    .X(_0515_));
 sg13g2_buf_1 _3652_ (.A(net165),
    .X(_0516_));
 sg13g2_mux2_1 _3653_ (.A0(\g.g_y[7].g_x[1].t.r_gnl ),
    .A1(\g.g_y[7].g_x[1].t.out_sc ),
    .S(_2386_),
    .X(_0517_));
 sg13g2_buf_1 _3654_ (.A(_0517_),
    .X(_0518_));
 sg13g2_mux2_1 _3655_ (.A0(_0518_),
    .A1(_2388_),
    .S(\g.g_y[7].g_x[1].t.r_v ),
    .X(_0519_));
 sg13g2_mux2_1 _3656_ (.A0(_0519_),
    .A1(_0276_),
    .S(_0279_),
    .X(_0520_));
 sg13g2_buf_1 _3657_ (.A(_0520_),
    .X(_0521_));
 sg13g2_nor4_1 _3658_ (.A(net69),
    .B(_0265_),
    .C(net30),
    .D(_0260_),
    .Y(_0522_));
 sg13g2_nor3_1 _3659_ (.A(_0261_),
    .B(_0264_),
    .C(net30),
    .Y(_0523_));
 sg13g2_nand2b_1 _3660_ (.Y(_0524_),
    .B(net71),
    .A_N(_2388_));
 sg13g2_o21ai_1 _3661_ (.B1(_0524_),
    .Y(_0525_),
    .A1(_0228_),
    .A2(_0518_));
 sg13g2_mux2_1 _3662_ (.A0(_0288_),
    .A1(_0525_),
    .S(_0279_),
    .X(_0526_));
 sg13g2_buf_1 _3663_ (.A(_0526_),
    .X(_0527_));
 sg13g2_a22oi_1 _3664_ (.Y(_0528_),
    .B1(_0523_),
    .B2(_0527_),
    .A2(_0522_),
    .A1(_0521_));
 sg13g2_nand2_1 _3665_ (.Y(_0529_),
    .A(_0265_),
    .B(_0284_));
 sg13g2_or2_1 _3666_ (.X(_0530_),
    .B(net68),
    .A(_0261_));
 sg13g2_a21oi_1 _3667_ (.A1(_0264_),
    .A2(\g.g_y[6].g_x[1].t.out_sc ),
    .Y(_0531_),
    .B1(_0530_));
 sg13g2_nand2_1 _3668_ (.Y(_0532_),
    .A(net69),
    .B(_2731_));
 sg13g2_a21oi_1 _3669_ (.A1(_2757_),
    .A2(_2732_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_nand2_1 _3670_ (.Y(_0534_),
    .A(net74),
    .B(_2760_));
 sg13g2_a22oi_1 _3671_ (.Y(_0535_),
    .B1(_0533_),
    .B2(_0534_),
    .A2(_0531_),
    .A1(_0529_));
 sg13g2_nand2_1 _3672_ (.Y(_0536_),
    .A(net69),
    .B(_2757_));
 sg13g2_or4_1 _3673_ (.A(_2731_),
    .B(_0440_),
    .C(_0442_),
    .D(_0536_),
    .X(_0537_));
 sg13g2_nand3_1 _3674_ (.B(net74),
    .C(_2747_),
    .A(net69),
    .Y(_0538_));
 sg13g2_and4_1 _3675_ (.A(_0528_),
    .B(_0535_),
    .C(_0537_),
    .D(_0538_),
    .X(_0539_));
 sg13g2_nand3b_1 _3676_ (.B(net152),
    .C(_0539_),
    .Y(_0540_),
    .A_N(_2753_));
 sg13g2_o21ai_1 _3677_ (.B1(_0540_),
    .Y(_0108_),
    .A1(_0513_),
    .A2(_0514_));
 sg13g2_or2_1 _3678_ (.X(_0541_),
    .B(_0442_),
    .A(_0440_));
 sg13g2_nand2_1 _3679_ (.Y(_0542_),
    .A(_2746_),
    .B(_2745_));
 sg13g2_o21ai_1 _3680_ (.B1(_0542_),
    .Y(_0543_),
    .A1(_2746_),
    .A2(_0441_));
 sg13g2_mux4_1 _3681_ (.S0(net74),
    .A0(_2732_),
    .A1(_2760_),
    .A2(_0541_),
    .A3(_0543_),
    .S1(_2730_),
    .X(_0544_));
 sg13g2_nand2b_1 _3682_ (.Y(_0545_),
    .B(_0521_),
    .A_N(_0267_));
 sg13g2_inv_1 _3683_ (.Y(_0546_),
    .A(_0527_));
 sg13g2_mux4_1 _3684_ (.S0(_0265_),
    .A0(\g.g_y[6].g_x[1].t.out_sc ),
    .A1(_0284_),
    .A2(_0545_),
    .A3(_0546_),
    .S1(net68),
    .X(_0547_));
 sg13g2_mux2_1 _3685_ (.A0(_0544_),
    .A1(_0547_),
    .S(net69),
    .X(_0548_));
 sg13g2_a221oi_1 _3686_ (.B2(_0485_),
    .C1(_2782_),
    .B1(_0511_),
    .A1(_0496_),
    .Y(_0549_),
    .A2(_0498_));
 sg13g2_a21oi_1 _3687_ (.A1(_2782_),
    .A2(_0474_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_a21oi_1 _3688_ (.A1(_0548_),
    .A2(_0550_),
    .Y(_0109_),
    .B1(net137));
 sg13g2_buf_1 _3689_ (.A(net166),
    .X(_0551_));
 sg13g2_and2_1 _3690_ (.A(\g.g_y[6].g_x[2].t.out_sc ),
    .B(net151),
    .X(_0107_));
 sg13g2_nor2_1 _3691_ (.A(_0278_),
    .B(_2499_),
    .Y(_0106_));
 sg13g2_nand2_1 _3692_ (.Y(_0552_),
    .A(_2424_),
    .B(_2415_));
 sg13g2_o21ai_1 _3693_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_2415_),
    .A2(_2390_));
 sg13g2_nor2_1 _3694_ (.A(net87),
    .B(net86),
    .Y(_0554_));
 sg13g2_and2_1 _3695_ (.A(_2421_),
    .B(_0554_),
    .X(_0555_));
 sg13g2_nor2b_1 _3696_ (.A(\g.g_y[7].g_x[0].t.out_sc ),
    .B_N(_2398_),
    .Y(_0556_));
 sg13g2_nand2b_1 _3697_ (.Y(_0557_),
    .B(_0556_),
    .A_N(net87));
 sg13g2_o21ai_1 _3698_ (.B1(_0557_),
    .Y(_0558_),
    .A1(_2421_),
    .A2(_2406_));
 sg13g2_a221oi_1 _3699_ (.B2(_0555_),
    .C1(_0558_),
    .B1(_0553_),
    .A1(_2397_),
    .Y(_0559_),
    .A2(_2428_));
 sg13g2_or2_1 _3700_ (.X(_0560_),
    .B(_0559_),
    .A(_2408_));
 sg13g2_buf_1 _3701_ (.A(\g.g_y[5].g_x[0].t.r_d ),
    .X(_0561_));
 sg13g2_inv_2 _3702_ (.Y(_0562_),
    .A(\g.g_y[5].g_x[0].t.r_h ));
 sg13g2_nand2b_1 _3703_ (.Y(_0563_),
    .B(_0489_),
    .A_N(_0274_));
 sg13g2_o21ai_1 _3704_ (.B1(_0563_),
    .Y(_0564_),
    .A1(_0489_),
    .A2(_0488_));
 sg13g2_nand2_1 _3705_ (.Y(_0565_),
    .A(net6),
    .B(_0562_));
 sg13g2_o21ai_1 _3706_ (.B1(_0565_),
    .Y(_0566_),
    .A1(_0562_),
    .A2(_0564_));
 sg13g2_buf_2 _3707_ (.A(\g.g_y[4].g_x[0].t.r_v ),
    .X(_0567_));
 sg13g2_inv_1 _3708_ (.Y(_0568_),
    .A(_0567_));
 sg13g2_buf_2 _3709_ (.A(\g.g_y[4].g_x[0].t.r_d ),
    .X(_0569_));
 sg13g2_mux2_1 _3710_ (.A0(\g.g_y[4].g_x[0].t.r_gnl ),
    .A1(\g.g_y[4].g_x[0].t.out_sc ),
    .S(_0569_),
    .X(_0570_));
 sg13g2_buf_2 _3711_ (.A(_0570_),
    .X(_0571_));
 sg13g2_buf_2 _3712_ (.A(\g.g_y[4].g_x[0].t.r_ghl ),
    .X(_0572_));
 sg13g2_or2_1 _3713_ (.X(_0573_),
    .B(_0567_),
    .A(_0572_));
 sg13g2_buf_1 _3714_ (.A(_0573_),
    .X(_0574_));
 sg13g2_o21ai_1 _3715_ (.B1(_0574_),
    .Y(_0575_),
    .A1(_0568_),
    .A2(_0571_));
 sg13g2_buf_1 _3716_ (.A(\g.g_y[5].g_x[0].t.r_v ),
    .X(_0576_));
 sg13g2_a21oi_1 _3717_ (.A1(net61),
    .A2(_0575_),
    .Y(_0577_),
    .B1(_0576_));
 sg13g2_o21ai_1 _3718_ (.B1(_0577_),
    .Y(_0578_),
    .A1(net61),
    .A2(_0566_));
 sg13g2_inv_1 _3719_ (.Y(_0579_),
    .A(\g.g_y[5].g_x[0].t.r_d ));
 sg13g2_inv_1 _3720_ (.Y(_0580_),
    .A(net6));
 sg13g2_nor2_1 _3721_ (.A(_0580_),
    .B(_0562_),
    .Y(_0581_));
 sg13g2_and3_1 _3722_ (.X(_0582_),
    .A(_0562_),
    .B(_0579_),
    .C(_0563_));
 sg13g2_nand2b_1 _3723_ (.Y(_0583_),
    .B(_0506_),
    .A_N(_0488_));
 sg13g2_a22oi_1 _3724_ (.Y(_0584_),
    .B1(_0582_),
    .B2(_0583_),
    .A2(_0581_),
    .A1(_0579_));
 sg13g2_nand2b_1 _3725_ (.Y(_0585_),
    .B(net61),
    .A_N(\g.g_y[5].g_x[0].t.out_sc ));
 sg13g2_and2_1 _3726_ (.A(_0576_),
    .B(_0585_),
    .X(_0586_));
 sg13g2_o21ai_1 _3727_ (.B1(_0586_),
    .Y(_0587_),
    .A1(_0575_),
    .A2(_0584_));
 sg13g2_nand3_1 _3728_ (.B(_0578_),
    .C(_0587_),
    .A(_2408_),
    .Y(_0588_));
 sg13g2_nand3_1 _3729_ (.B(_0560_),
    .C(_0588_),
    .A(_2409_),
    .Y(_0589_));
 sg13g2_nor2_1 _3730_ (.A(net30),
    .B(_0267_),
    .Y(_0590_));
 sg13g2_nand2_1 _3731_ (.Y(_0591_),
    .A(net85),
    .B(_0265_));
 sg13g2_a221oi_1 _3732_ (.B2(_0590_),
    .C1(_0591_),
    .B1(_0521_),
    .A1(_0269_),
    .Y(_0592_),
    .A2(_0278_));
 sg13g2_and2_1 _3733_ (.A(net68),
    .B(_0527_),
    .X(_0593_));
 sg13g2_nand3b_1 _3734_ (.B(_0264_),
    .C(net85),
    .Y(_0594_),
    .A_N(_0287_));
 sg13g2_nand2b_1 _3735_ (.Y(_0595_),
    .B(net7),
    .A_N(net85));
 sg13g2_o21ai_1 _3736_ (.B1(_0595_),
    .Y(_0596_),
    .A1(_0593_),
    .A2(_0594_));
 sg13g2_inv_1 _3737_ (.Y(_0597_),
    .A(_2409_));
 sg13g2_o21ai_1 _3738_ (.B1(_0597_),
    .Y(_0598_),
    .A1(_0592_),
    .A2(_0596_));
 sg13g2_a21oi_1 _3739_ (.A1(_0589_),
    .A2(_0598_),
    .Y(_0104_),
    .B1(_0313_));
 sg13g2_a21oi_1 _3740_ (.A1(_0578_),
    .A2(_0587_),
    .Y(_0599_),
    .B1(_2408_));
 sg13g2_a21o_1 _3741_ (.A2(_0559_),
    .A1(_2408_),
    .B1(_0599_),
    .X(_0600_));
 sg13g2_nor2b_1 _3742_ (.A(_0267_),
    .B_N(_0521_),
    .Y(_0601_));
 sg13g2_mux4_1 _3743_ (.S0(_0264_),
    .A0(_0278_),
    .A1(_0263_),
    .A2(_0601_),
    .A3(_0527_),
    .S1(net68),
    .X(_0602_));
 sg13g2_nand2_1 _3744_ (.Y(_0603_),
    .A(net85),
    .B(net7));
 sg13g2_o21ai_1 _3745_ (.B1(_0603_),
    .Y(_0604_),
    .A1(net85),
    .A2(_0602_));
 sg13g2_a21oi_1 _3746_ (.A1(_0600_),
    .A2(_0604_),
    .Y(_0105_),
    .B1(_0313_));
 sg13g2_and2_1 _3747_ (.A(\g.g_y[6].g_x[0].t.out_sc ),
    .B(net151),
    .X(_0103_));
 sg13g2_mux2_1 _3748_ (.A0(_2489_),
    .A1(_2530_),
    .S(net84),
    .X(_0605_));
 sg13g2_a21oi_1 _3749_ (.A1(net84),
    .A2(_2438_),
    .Y(_0606_),
    .B1(_2525_));
 sg13g2_or2_1 _3750_ (.X(_0607_),
    .B(_2435_),
    .A(_2433_));
 sg13g2_nand2_1 _3751_ (.Y(_0608_),
    .A(_2454_),
    .B(_2527_));
 sg13g2_a221oi_1 _3752_ (.B2(net84),
    .C1(_0608_),
    .B1(_2443_),
    .A1(_2436_),
    .Y(_0609_),
    .A2(_0607_));
 sg13g2_a221oi_1 _3753_ (.B2(_0367_),
    .C1(_0609_),
    .B1(_0606_),
    .A1(net83),
    .Y(_0610_),
    .A2(_0605_));
 sg13g2_a21oi_1 _3754_ (.A1(_2521_),
    .A2(_2530_),
    .Y(_0611_),
    .B1(net83));
 sg13g2_o21ai_1 _3755_ (.B1(_0611_),
    .Y(_0612_),
    .A1(_2521_),
    .A2(_2526_));
 sg13g2_nand3_1 _3756_ (.B(_0610_),
    .C(_0612_),
    .A(_2444_),
    .Y(_0613_));
 sg13g2_buf_1 _3757_ (.A(\g.g_y[4].g_x[7].t.r_v ),
    .X(_0614_));
 sg13g2_inv_1 _3758_ (.Y(_0615_),
    .A(net60));
 sg13g2_buf_2 _3759_ (.A(\g.g_y[3].g_x[7].t.r_d ),
    .X(_0616_));
 sg13g2_mux2_1 _3760_ (.A0(\g.g_y[3].g_x[7].t.r_gnl ),
    .A1(\g.g_y[3].g_x[7].t.out_sc ),
    .S(_0616_),
    .X(_0617_));
 sg13g2_buf_1 _3761_ (.A(_0617_),
    .X(_0618_));
 sg13g2_buf_1 _3762_ (.A(\g.g_y[3].g_x[7].t.r_v ),
    .X(_0619_));
 sg13g2_mux2_1 _3763_ (.A0(\g.g_y[3].g_x[7].t.r_ghl ),
    .A1(_0618_),
    .S(_0619_),
    .X(_0620_));
 sg13g2_buf_1 _3764_ (.A(_0620_),
    .X(_0621_));
 sg13g2_and2_1 _3765_ (.A(_0615_),
    .B(_0621_),
    .X(_0622_));
 sg13g2_inv_1 _3766_ (.Y(_0623_),
    .A(\g.g_y[4].g_x[7].t.out_sc ));
 sg13g2_nor2_1 _3767_ (.A(_0615_),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_buf_1 _3768_ (.A(\g.g_y[4].g_x[7].t.r_d ),
    .X(_0625_));
 sg13g2_o21ai_1 _3769_ (.B1(net59),
    .Y(_0626_),
    .A1(_0622_),
    .A2(_0624_));
 sg13g2_buf_2 _3770_ (.A(\g.g_y[4].g_x[0].t.r_h ),
    .X(_0627_));
 sg13g2_mux2_1 _3771_ (.A0(\g.g_y[4].g_x[0].t.out_sc ),
    .A1(\g.g_y[4].g_x[0].t.r_gnl ),
    .S(_0569_),
    .X(_0628_));
 sg13g2_buf_1 _3772_ (.A(_0628_),
    .X(_0629_));
 sg13g2_nand2b_1 _3773_ (.Y(_0630_),
    .B(_0627_),
    .A_N(_0572_));
 sg13g2_o21ai_1 _3774_ (.B1(_0630_),
    .Y(_0631_),
    .A1(_0627_),
    .A2(_0629_));
 sg13g2_buf_1 _3775_ (.A(_0631_),
    .X(_0632_));
 sg13g2_nand2_1 _3776_ (.Y(_0633_),
    .A(net60),
    .B(_0621_));
 sg13g2_buf_2 _3777_ (.A(\g.g_y[4].g_x[6].t.r_h ),
    .X(_0634_));
 sg13g2_mux2_1 _3778_ (.A0(\g.g_y[4].g_x[6].t.out_sc ),
    .A1(\g.g_y[4].g_x[6].t.r_gnl ),
    .S(_0328_),
    .X(_0635_));
 sg13g2_nor2b_1 _3779_ (.A(_0634_),
    .B_N(_0324_),
    .Y(_0636_));
 sg13g2_a21oi_1 _3780_ (.A1(_0634_),
    .A2(_0635_),
    .Y(_0637_),
    .B1(_0636_));
 sg13g2_buf_2 _3781_ (.A(_0637_),
    .X(_0638_));
 sg13g2_or2_1 _3782_ (.X(_0639_),
    .B(net59),
    .A(\g.g_y[4].g_x[7].t.r_h ));
 sg13g2_a21oi_1 _3783_ (.A1(_0615_),
    .A2(_0638_),
    .Y(_0640_),
    .B1(_0639_));
 sg13g2_o21ai_1 _3784_ (.B1(_0640_),
    .Y(_0641_),
    .A1(net23),
    .A2(_0633_));
 sg13g2_buf_1 _3785_ (.A(\g.g_y[4].g_x[7].t.r_h ),
    .X(_0642_));
 sg13g2_nor2b_1 _3786_ (.A(net59),
    .B_N(net58),
    .Y(_0643_));
 sg13g2_nand2_1 _3787_ (.Y(_0644_),
    .A(_0615_),
    .B(_0632_));
 sg13g2_nand3b_1 _3788_ (.B(net60),
    .C(_0621_),
    .Y(_0645_),
    .A_N(_0638_));
 sg13g2_nand3_1 _3789_ (.B(_0644_),
    .C(_0645_),
    .A(_0643_),
    .Y(_0646_));
 sg13g2_nand4_1 _3790_ (.B(_0626_),
    .C(_0641_),
    .A(_2445_),
    .Y(_0647_),
    .D(_0646_));
 sg13g2_nand3_1 _3791_ (.B(_0613_),
    .C(_0647_),
    .A(_2446_),
    .Y(_0648_));
 sg13g2_mux2_1 _3792_ (.A0(_2403_),
    .A1(_2411_),
    .S(_2408_),
    .X(_0649_));
 sg13g2_inv_1 _3793_ (.Y(_0650_),
    .A(_0576_));
 sg13g2_and2_1 _3794_ (.A(_0650_),
    .B(_0574_),
    .X(_0651_));
 sg13g2_or2_1 _3795_ (.X(_0652_),
    .B(_0571_),
    .A(_0568_));
 sg13g2_buf_1 _3796_ (.A(_0652_),
    .X(_0653_));
 sg13g2_a221oi_1 _3797_ (.B2(_0653_),
    .C1(_0579_),
    .B1(_0651_),
    .A1(_0576_),
    .Y(_0654_),
    .A2(_0649_));
 sg13g2_a21oi_1 _3798_ (.A1(_0579_),
    .A2(_0564_),
    .Y(_0655_),
    .B1(_0562_));
 sg13g2_nand2b_1 _3799_ (.Y(_0656_),
    .B(_0655_),
    .A_N(_0654_));
 sg13g2_nand2b_1 _3800_ (.Y(_0657_),
    .B(_2408_),
    .A_N(_2411_));
 sg13g2_nand2b_1 _3801_ (.Y(_0658_),
    .B(_2404_),
    .A_N(_2403_));
 sg13g2_and3_1 _3802_ (.X(_0659_),
    .A(_0650_),
    .B(net61),
    .C(_0658_));
 sg13g2_and3_1 _3803_ (.X(_0660_),
    .A(_0576_),
    .B(_0561_),
    .C(_0574_));
 sg13g2_a22oi_1 _3804_ (.Y(_0661_),
    .B1(_0660_),
    .B2(_0653_),
    .A2(_0659_),
    .A1(_0657_));
 sg13g2_nor2_1 _3805_ (.A(net61),
    .B(\g.g_y[5].g_x[0].t.out_sc ),
    .Y(_0662_));
 sg13g2_nor2_1 _3806_ (.A(\g.g_y[5].g_x[0].t.r_h ),
    .B(_0662_),
    .Y(_0663_));
 sg13g2_o21ai_1 _3807_ (.B1(_0663_),
    .Y(_0664_),
    .A1(_0564_),
    .A2(_0661_));
 sg13g2_nand3_1 _3808_ (.B(_0656_),
    .C(_0664_),
    .A(net65),
    .Y(_0665_));
 sg13g2_or2_1 _3809_ (.X(_0666_),
    .B(_0338_),
    .A(_2598_));
 sg13g2_o21ai_1 _3810_ (.B1(_0666_),
    .Y(_0667_),
    .A1(_0339_),
    .A2(_0340_));
 sg13g2_or2_1 _3811_ (.X(_0668_),
    .B(_2353_),
    .A(_2354_));
 sg13g2_nor2b_1 _3812_ (.A(_2351_),
    .B_N(_2354_),
    .Y(_0669_));
 sg13g2_nor3_1 _3813_ (.A(net64),
    .B(_0349_),
    .C(_0669_),
    .Y(_0670_));
 sg13g2_nand2_1 _3814_ (.Y(_0671_),
    .A(net64),
    .B(net67));
 sg13g2_nor2_1 _3815_ (.A(_0326_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_a22oi_1 _3816_ (.Y(_0673_),
    .B1(_0672_),
    .B2(_0331_),
    .A2(_0670_),
    .A1(_0668_));
 sg13g2_nor2_1 _3817_ (.A(net67),
    .B(\g.g_y[5].g_x[6].t.out_sc ),
    .Y(_0674_));
 sg13g2_nor2_1 _3818_ (.A(_0348_),
    .B(_0674_),
    .Y(_0675_));
 sg13g2_o21ai_1 _3819_ (.B1(_0675_),
    .Y(_0676_),
    .A1(_0667_),
    .A2(_0673_));
 sg13g2_mux2_1 _3820_ (.A0(_2353_),
    .A1(_2351_),
    .S(_2354_),
    .X(_0677_));
 sg13g2_buf_1 _3821_ (.A(_0677_),
    .X(_0678_));
 sg13g2_nor2_1 _3822_ (.A(net64),
    .B(_0326_),
    .Y(_0679_));
 sg13g2_a221oi_1 _3823_ (.B2(_0331_),
    .C1(_0349_),
    .B1(_0679_),
    .A1(net64),
    .Y(_0680_),
    .A2(_0678_));
 sg13g2_a21oi_1 _3824_ (.A1(_0349_),
    .A2(_0667_),
    .Y(_0681_),
    .B1(net66));
 sg13g2_nand2b_1 _3825_ (.Y(_0682_),
    .B(_0681_),
    .A_N(_0680_));
 sg13g2_nand3b_1 _3826_ (.B(_0676_),
    .C(_0682_),
    .Y(_0683_),
    .A_N(net65));
 sg13g2_nand3b_1 _3827_ (.B(_0665_),
    .C(_0683_),
    .Y(_0684_),
    .A_N(_2446_));
 sg13g2_a21oi_1 _3828_ (.A1(_0648_),
    .A2(_0684_),
    .Y(_0101_),
    .B1(net137));
 sg13g2_nand3_1 _3829_ (.B(_0676_),
    .C(_0682_),
    .A(net65),
    .Y(_0685_));
 sg13g2_nand3b_1 _3830_ (.B(_0656_),
    .C(_0664_),
    .Y(_0686_),
    .A_N(net65));
 sg13g2_nand4_1 _3831_ (.B(_0626_),
    .C(_0641_),
    .A(_2444_),
    .Y(_0687_),
    .D(_0646_));
 sg13g2_nand3_1 _3832_ (.B(_0610_),
    .C(_0612_),
    .A(_2445_),
    .Y(_0688_));
 sg13g2_nand4_1 _3833_ (.B(_0686_),
    .C(_0687_),
    .A(_0685_),
    .Y(_0689_),
    .D(_0688_));
 sg13g2_and2_1 _3834_ (.A(net155),
    .B(_0689_),
    .X(_0102_));
 sg13g2_and2_1 _3835_ (.A(\g.g_y[5].g_x[7].t.out_sc ),
    .B(_0551_),
    .X(_0100_));
 sg13g2_and2_1 _3836_ (.A(\g.g_y[5].g_x[6].t.out_sc ),
    .B(net151),
    .X(_0099_));
 sg13g2_or3_1 _3837_ (.A(_2606_),
    .B(_2615_),
    .C(_2620_),
    .X(_0690_));
 sg13g2_and2_1 _3838_ (.A(_2586_),
    .B(_2604_),
    .X(_0691_));
 sg13g2_nand2_1 _3839_ (.Y(_0692_),
    .A(_2606_),
    .B(_2609_));
 sg13g2_a21o_1 _3840_ (.A2(_0691_),
    .A1(_2597_),
    .B1(_0692_),
    .X(_0693_));
 sg13g2_nand3_1 _3841_ (.B(_0690_),
    .C(_0693_),
    .A(_2601_),
    .Y(_0694_));
 sg13g2_buf_1 _3842_ (.A(\g.g_y[4].g_x[5].t.r_v ),
    .X(_0695_));
 sg13g2_mux2_1 _3843_ (.A0(_2598_),
    .A1(_2600_),
    .S(_2612_),
    .X(_0696_));
 sg13g2_buf_1 _3844_ (.A(_0696_),
    .X(_0697_));
 sg13g2_buf_2 _3845_ (.A(\g.g_y[3].g_x[5].t.r_ghl ),
    .X(_0698_));
 sg13g2_inv_1 _3846_ (.Y(_0699_),
    .A(_0698_));
 sg13g2_buf_2 _3847_ (.A(\g.g_y[3].g_x[5].t.r_v ),
    .X(_0700_));
 sg13g2_inv_2 _3848_ (.Y(_0701_),
    .A(_0700_));
 sg13g2_a21oi_1 _3849_ (.A1(_0699_),
    .A2(_0701_),
    .Y(_0702_),
    .B1(_0695_));
 sg13g2_buf_2 _3850_ (.A(\g.g_y[3].g_x[5].t.r_d ),
    .X(_0703_));
 sg13g2_mux2_1 _3851_ (.A0(\g.g_y[3].g_x[5].t.r_gnl ),
    .A1(\g.g_y[3].g_x[5].t.out_sc ),
    .S(_0703_),
    .X(_0704_));
 sg13g2_or2_1 _3852_ (.X(_0705_),
    .B(_0704_),
    .A(_0701_));
 sg13g2_buf_1 _3853_ (.A(_0705_),
    .X(_0706_));
 sg13g2_buf_1 _3854_ (.A(\g.g_y[4].g_x[5].t.r_d ),
    .X(_0707_));
 sg13g2_inv_1 _3855_ (.Y(_0708_),
    .A(net56));
 sg13g2_a221oi_1 _3856_ (.B2(_0706_),
    .C1(_0708_),
    .B1(_0702_),
    .A1(net57),
    .Y(_0709_),
    .A2(_0697_));
 sg13g2_buf_1 _3857_ (.A(_0709_),
    .X(_0710_));
 sg13g2_buf_2 _3858_ (.A(\g.g_y[4].g_x[5].t.r_h ),
    .X(_0711_));
 sg13g2_inv_1 _3859_ (.Y(_0712_),
    .A(_0711_));
 sg13g2_mux2_1 _3860_ (.A0(\g.g_y[4].g_x[4].t.out_sc ),
    .A1(\g.g_y[4].g_x[4].t.r_gnl ),
    .S(_0398_),
    .X(_0713_));
 sg13g2_buf_1 _3861_ (.A(\g.g_y[4].g_x[4].t.r_h ),
    .X(_0714_));
 sg13g2_mux2_1 _3862_ (.A0(_0403_),
    .A1(_0713_),
    .S(net55),
    .X(_0715_));
 sg13g2_buf_1 _3863_ (.A(_0715_),
    .X(_0716_));
 sg13g2_or2_1 _3864_ (.X(_0717_),
    .B(_0635_),
    .A(_0634_));
 sg13g2_buf_1 _3865_ (.A(_0717_),
    .X(_0718_));
 sg13g2_nand2b_1 _3866_ (.Y(_0719_),
    .B(_0634_),
    .A_N(_0324_));
 sg13g2_and2_1 _3867_ (.A(_0711_),
    .B(_0719_),
    .X(_0720_));
 sg13g2_a221oi_1 _3868_ (.B2(_0720_),
    .C1(net56),
    .B1(_0718_),
    .A1(_0712_),
    .Y(_0721_),
    .A2(_0716_));
 sg13g2_buf_1 _3869_ (.A(_0721_),
    .X(_0722_));
 sg13g2_or2_1 _3870_ (.X(_0723_),
    .B(_0722_),
    .A(_0710_));
 sg13g2_nor2_1 _3871_ (.A(_2601_),
    .B(net57),
    .Y(_0724_));
 sg13g2_inv_1 _3872_ (.Y(_0725_),
    .A(net57));
 sg13g2_nor3_1 _3873_ (.A(_2601_),
    .B(_0725_),
    .C(net56),
    .Y(_0726_));
 sg13g2_o21ai_1 _3874_ (.B1(net57),
    .Y(_0727_),
    .A1(_0698_),
    .A2(_0700_));
 sg13g2_inv_1 _3875_ (.Y(_0728_),
    .A(_0727_));
 sg13g2_a22oi_1 _3876_ (.Y(_0729_),
    .B1(_0697_),
    .B2(_0725_),
    .A2(_0728_),
    .A1(_0706_));
 sg13g2_buf_1 _3877_ (.A(_0729_),
    .X(_0730_));
 sg13g2_and2_1 _3878_ (.A(net28),
    .B(_0719_),
    .X(_0731_));
 sg13g2_a22oi_1 _3879_ (.Y(_0732_),
    .B1(_0718_),
    .B2(_0731_),
    .A2(_0716_),
    .A1(_0711_));
 sg13g2_buf_1 _3880_ (.A(_0732_),
    .X(_0733_));
 sg13g2_nor2_1 _3881_ (.A(_0730_),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_nand2b_1 _3882_ (.Y(_0735_),
    .B(net56),
    .A_N(\g.g_y[4].g_x[5].t.out_sc ));
 sg13g2_nor3_1 _3883_ (.A(_2601_),
    .B(_0725_),
    .C(_0735_),
    .Y(_0736_));
 sg13g2_a221oi_1 _3884_ (.B2(_0734_),
    .C1(_0736_),
    .B1(_0726_),
    .A1(_0723_),
    .Y(_0737_),
    .A2(_0724_));
 sg13g2_nand3_1 _3885_ (.B(_0694_),
    .C(_0737_),
    .A(_2599_),
    .Y(_0738_));
 sg13g2_mux2_1 _3886_ (.A0(_2743_),
    .A1(_0413_),
    .S(_0411_),
    .X(_0739_));
 sg13g2_nor2_1 _3887_ (.A(_0338_),
    .B(_0407_),
    .Y(_0740_));
 sg13g2_o21ai_1 _3888_ (.B1(_0740_),
    .Y(_0741_),
    .A1(_0388_),
    .A2(_0739_));
 sg13g2_or2_1 _3889_ (.X(_0742_),
    .B(_0390_),
    .A(\g.g_y[5].g_x[4].t.r_d ));
 sg13g2_buf_1 _3890_ (.A(_0742_),
    .X(_0743_));
 sg13g2_nor2_1 _3891_ (.A(_0338_),
    .B(_0408_),
    .Y(_0744_));
 sg13g2_nand2_1 _3892_ (.Y(_0745_),
    .A(_0348_),
    .B(_0674_));
 sg13g2_a22oi_1 _3893_ (.Y(_0746_),
    .B1(_0745_),
    .B2(_0338_),
    .A2(_0744_),
    .A1(_0743_));
 sg13g2_o21ai_1 _3894_ (.B1(_0746_),
    .Y(_0747_),
    .A1(_0426_),
    .A2(_0741_));
 sg13g2_nand2_1 _3895_ (.Y(_0748_),
    .A(net63),
    .B(_0744_));
 sg13g2_or3_1 _3896_ (.A(_0406_),
    .B(_0418_),
    .C(_0748_),
    .X(_0749_));
 sg13g2_nand2_1 _3897_ (.Y(_0750_),
    .A(_0347_),
    .B(_0350_));
 sg13g2_or4_1 _3898_ (.A(_0339_),
    .B(net66),
    .C(_0750_),
    .D(_0673_),
    .X(_0751_));
 sg13g2_nor2_1 _3899_ (.A(net67),
    .B(_0337_),
    .Y(_0752_));
 sg13g2_nor2_1 _3900_ (.A(_0339_),
    .B(_0348_),
    .Y(_0753_));
 sg13g2_o21ai_1 _3901_ (.B1(_0753_),
    .Y(_0754_),
    .A1(_0680_),
    .A2(_0752_));
 sg13g2_and4_1 _3902_ (.A(_0747_),
    .B(_0749_),
    .C(_0751_),
    .D(_0754_),
    .X(_0755_));
 sg13g2_nand2b_1 _3903_ (.Y(_0756_),
    .B(_0755_),
    .A_N(_2599_));
 sg13g2_a21oi_1 _3904_ (.A1(_0738_),
    .A2(_0756_),
    .Y(_0097_),
    .B1(net137));
 sg13g2_nor3_1 _3905_ (.A(_0339_),
    .B(_0408_),
    .C(_0743_),
    .Y(_0757_));
 sg13g2_nor2_1 _3906_ (.A(_0345_),
    .B(_0680_),
    .Y(_0758_));
 sg13g2_nor2_1 _3907_ (.A(net66),
    .B(_0674_),
    .Y(_0759_));
 sg13g2_or2_1 _3908_ (.X(_0760_),
    .B(_0673_),
    .A(_0750_));
 sg13g2_a221oi_1 _3909_ (.B2(_0760_),
    .C1(_0338_),
    .B1(_0759_),
    .A1(net66),
    .Y(_0761_),
    .A2(_0758_));
 sg13g2_and3_1 _3910_ (.X(_0762_),
    .A(_2612_),
    .B(_0690_),
    .C(_0693_));
 sg13g2_nor3_1 _3911_ (.A(_0757_),
    .B(_0761_),
    .C(_0762_),
    .Y(_0763_));
 sg13g2_nor3_1 _3912_ (.A(net56),
    .B(_0730_),
    .C(_0733_),
    .Y(_0764_));
 sg13g2_nand3b_1 _3913_ (.B(net57),
    .C(_0735_),
    .Y(_0765_),
    .A_N(_0764_));
 sg13g2_nor2_1 _3914_ (.A(_0710_),
    .B(_0722_),
    .Y(_0766_));
 sg13g2_a21oi_1 _3915_ (.A1(_0725_),
    .A2(_0766_),
    .Y(_0767_),
    .B1(_2612_));
 sg13g2_nor3_1 _3916_ (.A(_0389_),
    .B(_0406_),
    .C(_0418_),
    .Y(_0768_));
 sg13g2_mux2_1 _3917_ (.A0(_0427_),
    .A1(_0768_),
    .S(_0407_),
    .X(_0769_));
 sg13g2_a22oi_1 _3918_ (.Y(_0770_),
    .B1(_0769_),
    .B2(_0338_),
    .A2(_0767_),
    .A1(_0765_));
 sg13g2_a21oi_1 _3919_ (.A1(_0763_),
    .A2(_0770_),
    .Y(_0098_),
    .B1(net137));
 sg13g2_and2_1 _3920_ (.A(\g.g_y[5].g_x[5].t.out_sc ),
    .B(net151),
    .X(_0096_));
 sg13g2_and2_1 _3921_ (.A(_0390_),
    .B(net151),
    .X(_0095_));
 sg13g2_or3_1 _3922_ (.A(_2746_),
    .B(_2747_),
    .C(_2758_),
    .X(_0771_));
 sg13g2_nand2b_1 _3923_ (.Y(_0772_),
    .B(_2731_),
    .A_N(_0441_));
 sg13g2_nor2_1 _3924_ (.A(_2729_),
    .B(_2733_),
    .Y(_0773_));
 sg13g2_o21ai_1 _3925_ (.B1(_0773_),
    .Y(_0774_),
    .A1(_0440_),
    .A2(_0772_));
 sg13g2_nand3_1 _3926_ (.B(_0771_),
    .C(_0774_),
    .A(_2740_),
    .Y(_0775_));
 sg13g2_buf_1 _3927_ (.A(\g.g_y[4].g_x[3].t.r_d ),
    .X(_0776_));
 sg13g2_inv_2 _3928_ (.Y(_0777_),
    .A(net54));
 sg13g2_buf_1 _3929_ (.A(\g.g_y[4].g_x[3].t.r_h ),
    .X(_0778_));
 sg13g2_inv_1 _3930_ (.Y(_0779_),
    .A(net53));
 sg13g2_mux2_1 _3931_ (.A0(\g.g_y[4].g_x[2].t.out_sc ),
    .A1(\g.g_y[4].g_x[2].t.r_gnl ),
    .S(_0478_),
    .X(_0780_));
 sg13g2_buf_2 _3932_ (.A(_0780_),
    .X(_0781_));
 sg13g2_buf_2 _3933_ (.A(\g.g_y[4].g_x[2].t.r_h ),
    .X(_0782_));
 sg13g2_mux2_1 _3934_ (.A0(_0477_),
    .A1(_0781_),
    .S(_0782_),
    .X(_0783_));
 sg13g2_or2_1 _3935_ (.X(_0784_),
    .B(_0713_),
    .A(net55));
 sg13g2_buf_1 _3936_ (.A(_0784_),
    .X(_0785_));
 sg13g2_nand2b_1 _3937_ (.Y(_0786_),
    .B(net55),
    .A_N(_0403_));
 sg13g2_and2_1 _3938_ (.A(net53),
    .B(_0786_),
    .X(_0787_));
 sg13g2_a22oi_1 _3939_ (.Y(_0788_),
    .B1(_0785_),
    .B2(_0787_),
    .A2(_0783_),
    .A1(_0779_));
 sg13g2_buf_2 _3940_ (.A(\g.g_y[4].g_x[3].t.r_v ),
    .X(_0789_));
 sg13g2_mux2_1 _3941_ (.A0(_2742_),
    .A1(_2743_),
    .S(net75),
    .X(_0790_));
 sg13g2_buf_2 _3942_ (.A(\g.g_y[3].g_x[3].t.r_ghl ),
    .X(_0791_));
 sg13g2_inv_1 _3943_ (.Y(_0792_),
    .A(_0791_));
 sg13g2_buf_2 _3944_ (.A(\g.g_y[3].g_x[3].t.r_v ),
    .X(_0793_));
 sg13g2_inv_1 _3945_ (.Y(_0794_),
    .A(_0793_));
 sg13g2_a21oi_1 _3946_ (.A1(_0792_),
    .A2(_0794_),
    .Y(_0795_),
    .B1(_0789_));
 sg13g2_buf_8 _3947_ (.A(\g.g_y[3].g_x[3].t.r_d ),
    .X(_0796_));
 sg13g2_mux2_1 _3948_ (.A0(\g.g_y[3].g_x[3].t.r_gnl ),
    .A1(\g.g_y[3].g_x[3].t.out_sc ),
    .S(_0796_),
    .X(_0797_));
 sg13g2_or2_1 _3949_ (.X(_0798_),
    .B(_0797_),
    .A(_0794_));
 sg13g2_a221oi_1 _3950_ (.B2(_0798_),
    .C1(_0777_),
    .B1(_0795_),
    .A1(_0789_),
    .Y(_0799_),
    .A2(_0790_));
 sg13g2_a21o_1 _3951_ (.A2(_0788_),
    .A1(_0777_),
    .B1(_0799_),
    .X(_0800_));
 sg13g2_nor2_1 _3952_ (.A(net75),
    .B(_0789_),
    .Y(_0801_));
 sg13g2_inv_2 _3953_ (.Y(_0802_),
    .A(_0789_));
 sg13g2_nor3_1 _3954_ (.A(net75),
    .B(_0802_),
    .C(_0776_),
    .Y(_0803_));
 sg13g2_o21ai_1 _3955_ (.B1(_0789_),
    .Y(_0804_),
    .A1(_0791_),
    .A2(_0793_));
 sg13g2_inv_1 _3956_ (.Y(_0805_),
    .A(_0804_));
 sg13g2_a22oi_1 _3957_ (.Y(_0806_),
    .B1(_0790_),
    .B2(_0802_),
    .A2(_0805_),
    .A1(_0798_));
 sg13g2_and2_1 _3958_ (.A(_0779_),
    .B(_0786_),
    .X(_0807_));
 sg13g2_a22oi_1 _3959_ (.Y(_0808_),
    .B1(_0785_),
    .B2(_0807_),
    .A2(_0783_),
    .A1(net53));
 sg13g2_nor2_1 _3960_ (.A(_0806_),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_buf_1 _3961_ (.A(\g.g_y[4].g_x[3].t.out_sc ),
    .X(_0810_));
 sg13g2_nor4_1 _3962_ (.A(net75),
    .B(_0802_),
    .C(_0777_),
    .D(net164),
    .Y(_0811_));
 sg13g2_a221oi_1 _3963_ (.B2(_0809_),
    .C1(_0811_),
    .B1(_0803_),
    .A1(_0800_),
    .Y(_0812_),
    .A2(_0801_));
 sg13g2_nand3_1 _3964_ (.B(_0775_),
    .C(_0812_),
    .A(_2741_),
    .Y(_0813_));
 sg13g2_a22oi_1 _3965_ (.Y(_0814_),
    .B1(_0402_),
    .B2(_0425_),
    .A2(_0395_),
    .A1(net62));
 sg13g2_nor2_1 _3966_ (.A(_0408_),
    .B(_0389_),
    .Y(_0815_));
 sg13g2_and3_1 _3967_ (.X(_0816_),
    .A(_0408_),
    .B(net63),
    .C(_0410_));
 sg13g2_mux2_1 _3968_ (.A0(_0403_),
    .A1(_0400_),
    .S(_0396_),
    .X(_0817_));
 sg13g2_mux2_1 _3969_ (.A0(_0395_),
    .A1(_0817_),
    .S(net62),
    .X(_0818_));
 sg13g2_nand2_1 _3970_ (.Y(_0819_),
    .A(_0407_),
    .B(_0389_));
 sg13g2_nand2b_1 _3971_ (.Y(_0820_),
    .B(_0408_),
    .A_N(_0743_));
 sg13g2_o21ai_1 _3972_ (.B1(_0820_),
    .Y(_0821_),
    .A1(_0410_),
    .A2(_0819_));
 sg13g2_a221oi_1 _3973_ (.B2(_0818_),
    .C1(_0821_),
    .B1(_0816_),
    .A1(_0814_),
    .Y(_0822_),
    .A2(_0815_));
 sg13g2_nor2_1 _3974_ (.A(net29),
    .B(\g.g_y[5].g_x[2].t.out_sc ),
    .Y(_0823_));
 sg13g2_nor3_1 _3975_ (.A(_0411_),
    .B(_0494_),
    .C(_0823_),
    .Y(_0824_));
 sg13g2_nand3_1 _3976_ (.B(_0486_),
    .C(_0495_),
    .A(_0509_),
    .Y(_0825_));
 sg13g2_nor4_1 _3977_ (.A(_0411_),
    .B(_0493_),
    .C(_0504_),
    .D(_0510_),
    .Y(_0826_));
 sg13g2_a221oi_1 _3978_ (.B2(_0825_),
    .C1(_0826_),
    .B1(_0824_),
    .A1(_0411_),
    .Y(_0827_),
    .A2(_0822_));
 sg13g2_or2_1 _3979_ (.X(_0828_),
    .B(_0827_),
    .A(_2741_));
 sg13g2_buf_1 _3980_ (.A(net154),
    .X(_0829_));
 sg13g2_a21oi_1 _3981_ (.A1(_0813_),
    .A2(_0828_),
    .Y(_0093_),
    .B1(net136));
 sg13g2_nor2_1 _3982_ (.A(_0494_),
    .B(_0823_),
    .Y(_0830_));
 sg13g2_a22oi_1 _3983_ (.Y(_0831_),
    .B1(_0825_),
    .B2(_0830_),
    .A2(_0511_),
    .A1(_0494_));
 sg13g2_nor2_1 _3984_ (.A(_0411_),
    .B(_0822_),
    .Y(_0832_));
 sg13g2_a21oi_1 _3985_ (.A1(_0411_),
    .A2(_0831_),
    .Y(_0833_),
    .B1(_0832_));
 sg13g2_or2_1 _3986_ (.X(_0834_),
    .B(_0808_),
    .A(_0806_));
 sg13g2_buf_1 _3987_ (.A(_0834_),
    .X(_0835_));
 sg13g2_mux2_1 _3988_ (.A0(_0791_),
    .A1(_0797_),
    .S(_0793_),
    .X(_0836_));
 sg13g2_mux2_1 _3989_ (.A0(_0836_),
    .A1(_0790_),
    .S(_0789_),
    .X(_0837_));
 sg13g2_buf_2 _3990_ (.A(_0837_),
    .X(_0838_));
 sg13g2_inv_2 _3991_ (.Y(_0839_),
    .A(_0782_));
 sg13g2_or2_1 _3992_ (.X(_0840_),
    .B(_0782_),
    .A(_0477_));
 sg13g2_o21ai_1 _3993_ (.B1(_0840_),
    .Y(_0841_),
    .A1(_0839_),
    .A2(_0781_));
 sg13g2_nand2_1 _3994_ (.Y(_0842_),
    .A(_0785_),
    .B(_0787_));
 sg13g2_o21ai_1 _3995_ (.B1(_0842_),
    .Y(_0843_),
    .A1(net53),
    .A2(_0841_));
 sg13g2_buf_1 _3996_ (.A(_0843_),
    .X(_0844_));
 sg13g2_mux4_1 _3997_ (.S0(_0777_),
    .A0(net164),
    .A1(_0835_),
    .A2(_0838_),
    .A3(_0844_),
    .S1(_0802_),
    .X(_0845_));
 sg13g2_a21oi_1 _3998_ (.A1(_0771_),
    .A2(_0774_),
    .Y(_0846_),
    .B1(_2740_));
 sg13g2_a21o_1 _3999_ (.A2(_0845_),
    .A1(net75),
    .B1(_0846_),
    .X(_0847_));
 sg13g2_a21oi_1 _4000_ (.A1(_0833_),
    .A2(_0847_),
    .Y(_0094_),
    .B1(net136));
 sg13g2_and2_1 _4001_ (.A(\g.g_y[5].g_x[3].t.out_sc ),
    .B(net151),
    .X(_0092_));
 sg13g2_and2_1 _4002_ (.A(\g.g_y[5].g_x[2].t.out_sc ),
    .B(net168),
    .X(_0091_));
 sg13g2_nand2_1 _4003_ (.Y(_0848_),
    .A(net30),
    .B(_0519_));
 sg13g2_a21oi_1 _4004_ (.A1(net68),
    .A2(_0278_),
    .Y(_0849_),
    .B1(_0279_));
 sg13g2_o21ai_1 _4005_ (.B1(_0849_),
    .Y(_0850_),
    .A1(_0267_),
    .A2(_0848_));
 sg13g2_o21ai_1 _4006_ (.B1(_0279_),
    .Y(_0851_),
    .A1(net30),
    .A2(_0519_));
 sg13g2_or2_1 _4007_ (.X(_0852_),
    .B(_0851_),
    .A(_0287_));
 sg13g2_nand3_1 _4008_ (.B(_0850_),
    .C(_0852_),
    .A(_0270_),
    .Y(_0853_));
 sg13g2_buf_1 _4009_ (.A(\g.g_y[4].g_x[1].t.r_v ),
    .X(_0854_));
 sg13g2_inv_1 _4010_ (.Y(_0855_),
    .A(net52));
 sg13g2_buf_1 _4011_ (.A(\g.g_y[4].g_x[1].t.r_d ),
    .X(_0856_));
 sg13g2_buf_1 _4012_ (.A(net51),
    .X(_0857_));
 sg13g2_buf_1 _4013_ (.A(\g.g_y[3].g_x[1].t.r_v ),
    .X(_0858_));
 sg13g2_buf_8 _4014_ (.A(\g.g_y[3].g_x[1].t.r_d ),
    .X(_0859_));
 sg13g2_mux2_1 _4015_ (.A0(\g.g_y[3].g_x[1].t.r_gnl ),
    .A1(\g.g_y[3].g_x[1].t.out_sc ),
    .S(_0859_),
    .X(_0860_));
 sg13g2_buf_1 _4016_ (.A(_0860_),
    .X(_0861_));
 sg13g2_buf_1 _4017_ (.A(\g.g_y[3].g_x[1].t.r_ghl ),
    .X(_0862_));
 sg13g2_nor2b_1 _4018_ (.A(net50),
    .B_N(_0862_),
    .Y(_0863_));
 sg13g2_a21oi_1 _4019_ (.A1(net50),
    .A2(_0861_),
    .Y(_0864_),
    .B1(_0863_));
 sg13g2_nand2b_1 _4020_ (.Y(_0865_),
    .B(_0782_),
    .A_N(_0477_));
 sg13g2_o21ai_1 _4021_ (.B1(_0865_),
    .Y(_0866_),
    .A1(_0782_),
    .A2(_0781_));
 sg13g2_inv_1 _4022_ (.Y(_0867_),
    .A(_0627_));
 sg13g2_or2_1 _4023_ (.X(_0868_),
    .B(_0627_),
    .A(_0572_));
 sg13g2_buf_1 _4024_ (.A(_0868_),
    .X(_0869_));
 sg13g2_o21ai_1 _4025_ (.B1(_0869_),
    .Y(_0870_),
    .A1(_0867_),
    .A2(_0629_));
 sg13g2_buf_1 _4026_ (.A(\g.g_y[4].g_x[1].t.r_h ),
    .X(_0871_));
 sg13g2_mux2_1 _4027_ (.A0(_0866_),
    .A1(_0870_),
    .S(_0871_),
    .X(_0872_));
 sg13g2_buf_1 _4028_ (.A(_0872_),
    .X(_0873_));
 sg13g2_nor4_1 _4029_ (.A(_0855_),
    .B(net27),
    .C(_0864_),
    .D(_0873_),
    .Y(_0874_));
 sg13g2_mux2_1 _4030_ (.A0(_0572_),
    .A1(_0629_),
    .S(_0627_),
    .X(_0875_));
 sg13g2_mux2_1 _4031_ (.A0(_0477_),
    .A1(_0781_),
    .S(_0839_),
    .X(_0876_));
 sg13g2_buf_1 _4032_ (.A(_0871_),
    .X(_0877_));
 sg13g2_mux2_1 _4033_ (.A0(_0875_),
    .A1(_0876_),
    .S(_0877_),
    .X(_0878_));
 sg13g2_or2_1 _4034_ (.X(_0879_),
    .B(net51),
    .A(net52));
 sg13g2_nor2b_1 _4035_ (.A(net52),
    .B_N(net51),
    .Y(_0880_));
 sg13g2_and2_1 _4036_ (.A(net52),
    .B(net51),
    .X(_0881_));
 sg13g2_buf_1 _4037_ (.A(\g.g_y[4].g_x[1].t.out_sc ),
    .X(_0882_));
 sg13g2_inv_1 _4038_ (.Y(_0883_),
    .A(_0882_));
 sg13g2_a22oi_1 _4039_ (.Y(_0884_),
    .B1(_0881_),
    .B2(_0883_),
    .A2(_0880_),
    .A1(_0864_));
 sg13g2_o21ai_1 _4040_ (.B1(_0884_),
    .Y(_0885_),
    .A1(_0878_),
    .A2(_0879_));
 sg13g2_inv_1 _4041_ (.Y(_0886_),
    .A(_0270_));
 sg13g2_o21ai_1 _4042_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0874_),
    .A2(_0885_));
 sg13g2_nand3_1 _4043_ (.B(_0853_),
    .C(_0887_),
    .A(_0271_),
    .Y(_0888_));
 sg13g2_and4_1 _4044_ (.A(_0494_),
    .B(net29),
    .C(_0486_),
    .D(_0492_),
    .X(_0889_));
 sg13g2_nand2_1 _4045_ (.Y(_0890_),
    .A(_0493_),
    .B(_0475_));
 sg13g2_a221oi_1 _4046_ (.B2(_0503_),
    .C1(_0890_),
    .B1(_0501_),
    .A1(_0484_),
    .Y(_0891_),
    .A2(_0483_));
 sg13g2_nor3_1 _4047_ (.A(_0493_),
    .B(net29),
    .C(\g.g_y[5].g_x[2].t.out_sc ),
    .Y(_0892_));
 sg13g2_nor3_1 _4048_ (.A(_0494_),
    .B(net29),
    .C(_0492_),
    .Y(_0893_));
 sg13g2_or3_1 _4049_ (.A(_0891_),
    .B(_0892_),
    .C(_0893_),
    .X(_0894_));
 sg13g2_o21ai_1 _4050_ (.B1(_0489_),
    .Y(_0895_),
    .A1(_0889_),
    .A2(_0894_));
 sg13g2_o21ai_1 _4051_ (.B1(_0562_),
    .Y(_0896_),
    .A1(net6),
    .A2(net61));
 sg13g2_or2_1 _4052_ (.X(_0897_),
    .B(_0896_),
    .A(_0654_));
 sg13g2_nor2_1 _4053_ (.A(_0562_),
    .B(_0662_),
    .Y(_0898_));
 sg13g2_o21ai_1 _4054_ (.B1(_0898_),
    .Y(_0899_),
    .A1(_0580_),
    .A2(_0661_));
 sg13g2_nand3_1 _4055_ (.B(_0897_),
    .C(_0899_),
    .A(_0506_),
    .Y(_0900_));
 sg13g2_nand3b_1 _4056_ (.B(_0895_),
    .C(_0900_),
    .Y(_0901_),
    .A_N(_0271_));
 sg13g2_a21oi_1 _4057_ (.A1(_0888_),
    .A2(_0901_),
    .Y(_0089_),
    .B1(net136));
 sg13g2_o21ai_1 _4058_ (.B1(_0506_),
    .Y(_0902_),
    .A1(_0889_),
    .A2(_0894_));
 sg13g2_nand3_1 _4059_ (.B(_0897_),
    .C(_0899_),
    .A(_0489_),
    .Y(_0903_));
 sg13g2_o21ai_1 _4060_ (.B1(_0270_),
    .Y(_0904_),
    .A1(_0874_),
    .A2(_0885_));
 sg13g2_nand3_1 _4061_ (.B(_0850_),
    .C(_0852_),
    .A(_0886_),
    .Y(_0905_));
 sg13g2_nand4_1 _4062_ (.B(_0903_),
    .C(_0904_),
    .A(_0902_),
    .Y(_0906_),
    .D(_0905_));
 sg13g2_and2_1 _4063_ (.A(net155),
    .B(_0906_),
    .X(_0090_));
 sg13g2_and2_1 _4064_ (.A(\g.g_y[5].g_x[1].t.out_sc ),
    .B(net151),
    .X(_0088_));
 sg13g2_and2_1 _4065_ (.A(\g.g_y[5].g_x[0].t.out_sc ),
    .B(_0551_),
    .X(_0087_));
 sg13g2_nor2_1 _4066_ (.A(_0623_),
    .B(net138),
    .Y(_0086_));
 sg13g2_nand2_1 _4067_ (.Y(_0907_),
    .A(net64),
    .B(_0349_));
 sg13g2_a221oi_1 _4068_ (.B2(_0344_),
    .C1(_0907_),
    .B1(_0342_),
    .A1(_0333_),
    .Y(_0908_),
    .A2(_0337_));
 sg13g2_nor2_1 _4069_ (.A(_0678_),
    .B(_0671_),
    .Y(_0909_));
 sg13g2_or2_1 _4070_ (.X(_0910_),
    .B(_0909_),
    .A(_0908_));
 sg13g2_nand2b_1 _4071_ (.Y(_0911_),
    .B(_0678_),
    .A_N(net64));
 sg13g2_or2_1 _4072_ (.X(_0912_),
    .B(_0354_),
    .A(net64));
 sg13g2_o21ai_1 _4073_ (.B1(_0912_),
    .Y(_0913_),
    .A1(_0353_),
    .A2(_0911_));
 sg13g2_o21ai_1 _4074_ (.B1(_0325_),
    .Y(_0914_),
    .A1(_0910_),
    .A2(_0913_));
 sg13g2_inv_1 _4075_ (.Y(_0915_),
    .A(\g.g_y[3].g_x[5].t.r_h ));
 sg13g2_mux2_1 _4076_ (.A0(\g.g_y[3].g_x[5].t.out_sc ),
    .A1(\g.g_y[3].g_x[5].t.r_gnl ),
    .S(_0703_),
    .X(_0916_));
 sg13g2_or2_1 _4077_ (.X(_0917_),
    .B(_0916_),
    .A(_0915_));
 sg13g2_buf_1 _4078_ (.A(_0917_),
    .X(_0918_));
 sg13g2_buf_1 _4079_ (.A(\g.g_y[3].g_x[6].t.r_h ),
    .X(_0919_));
 sg13g2_or2_1 _4080_ (.X(_0920_),
    .B(\g.g_y[3].g_x[5].t.r_h ),
    .A(_0698_));
 sg13g2_buf_1 _4081_ (.A(_0920_),
    .X(_0921_));
 sg13g2_and2_1 _4082_ (.A(_0919_),
    .B(_0921_),
    .X(_0922_));
 sg13g2_mux2_1 _4083_ (.A0(\g.g_y[3].g_x[7].t.out_sc ),
    .A1(\g.g_y[3].g_x[7].t.r_gnl ),
    .S(_0616_),
    .X(_0923_));
 sg13g2_buf_2 _4084_ (.A(\g.g_y[3].g_x[7].t.r_h ),
    .X(_0924_));
 sg13g2_inv_1 _4085_ (.Y(_0925_),
    .A(_0924_));
 sg13g2_mux2_1 _4086_ (.A0(\g.g_y[3].g_x[7].t.r_ghl ),
    .A1(_0923_),
    .S(_0925_),
    .X(_0926_));
 sg13g2_buf_1 _4087_ (.A(_0926_),
    .X(_0927_));
 sg13g2_inv_1 _4088_ (.Y(_0928_),
    .A(_0919_));
 sg13g2_a22oi_1 _4089_ (.Y(_0929_),
    .B1(_0927_),
    .B2(_0928_),
    .A2(_0922_),
    .A1(_0918_));
 sg13g2_buf_1 _4090_ (.A(_0929_),
    .X(_0930_));
 sg13g2_buf_1 _4091_ (.A(\g.g_y[3].g_x[6].t.r_d ),
    .X(_0931_));
 sg13g2_buf_2 _4092_ (.A(\g.g_y[2].g_x[6].t.r_v ),
    .X(_0932_));
 sg13g2_inv_1 _4093_ (.Y(_0933_),
    .A(_0932_));
 sg13g2_buf_1 _4094_ (.A(\g.g_y[2].g_x[6].t.r_d ),
    .X(_0934_));
 sg13g2_mux2_1 _4095_ (.A0(\g.g_y[2].g_x[6].t.r_gnl ),
    .A1(\g.g_y[2].g_x[6].t.out_sc ),
    .S(_0934_),
    .X(_0935_));
 sg13g2_buf_1 _4096_ (.A(_0935_),
    .X(_0936_));
 sg13g2_buf_2 _4097_ (.A(\g.g_y[2].g_x[6].t.r_ghl ),
    .X(_0937_));
 sg13g2_or2_1 _4098_ (.X(_0938_),
    .B(_0932_),
    .A(_0937_));
 sg13g2_buf_1 _4099_ (.A(_0938_),
    .X(_0939_));
 sg13g2_o21ai_1 _4100_ (.B1(_0939_),
    .Y(_0940_),
    .A1(_0933_),
    .A2(_0936_));
 sg13g2_or2_1 _4101_ (.X(_0941_),
    .B(_0940_),
    .A(net49));
 sg13g2_buf_1 _4102_ (.A(\g.g_y[3].g_x[6].t.r_v ),
    .X(_0942_));
 sg13g2_nand2b_1 _4103_ (.Y(_0943_),
    .B(net49),
    .A_N(\g.g_y[3].g_x[6].t.out_sc ));
 sg13g2_and2_1 _4104_ (.A(net48),
    .B(_0943_),
    .X(_0944_));
 sg13g2_o21ai_1 _4105_ (.B1(_0944_),
    .Y(_0945_),
    .A1(_0930_),
    .A2(_0941_));
 sg13g2_and2_1 _4106_ (.A(_0928_),
    .B(_0921_),
    .X(_0946_));
 sg13g2_a221oi_1 _4107_ (.B2(_0918_),
    .C1(net49),
    .B1(_0946_),
    .A1(_0919_),
    .Y(_0947_),
    .A2(_0927_));
 sg13g2_a21oi_1 _4108_ (.A1(net49),
    .A2(_0940_),
    .Y(_0948_),
    .B1(net48));
 sg13g2_nand2b_1 _4109_ (.Y(_0949_),
    .B(_0948_),
    .A_N(_0947_));
 sg13g2_nand3_1 _4110_ (.B(_0945_),
    .C(_0949_),
    .A(_0327_),
    .Y(_0950_));
 sg13g2_nand3_1 _4111_ (.B(_0914_),
    .C(_0950_),
    .A(_0328_),
    .Y(_0951_));
 sg13g2_inv_1 _4112_ (.Y(_0952_),
    .A(_0619_));
 sg13g2_or2_1 _4113_ (.X(_0953_),
    .B(_0618_),
    .A(_0952_));
 sg13g2_inv_1 _4114_ (.Y(_0954_),
    .A(\g.g_y[3].g_x[7].t.r_ghl ));
 sg13g2_a21oi_1 _4115_ (.A1(_0954_),
    .A2(_0952_),
    .Y(_0955_),
    .B1(net60));
 sg13g2_mux2_1 _4116_ (.A0(_2449_),
    .A1(_2448_),
    .S(_2445_),
    .X(_0956_));
 sg13g2_buf_2 _4117_ (.A(_0956_),
    .X(_0957_));
 sg13g2_inv_1 _4118_ (.Y(_0958_),
    .A(net59));
 sg13g2_a221oi_1 _4119_ (.B2(_0614_),
    .C1(_0958_),
    .B1(_0957_),
    .A1(_0953_),
    .Y(_0959_),
    .A2(_0955_));
 sg13g2_and2_1 _4120_ (.A(_0958_),
    .B(net23),
    .X(_0960_));
 sg13g2_o21ai_1 _4121_ (.B1(net58),
    .Y(_0961_),
    .A1(_0959_),
    .A2(_0960_));
 sg13g2_mux2_1 _4122_ (.A0(_0621_),
    .A1(_0957_),
    .S(_0615_),
    .X(_0962_));
 sg13g2_nor3_1 _4123_ (.A(net58),
    .B(_0958_),
    .C(net23),
    .Y(_0963_));
 sg13g2_o21ai_1 _4124_ (.B1(_0634_),
    .Y(_0964_),
    .A1(\g.g_y[4].g_x[7].t.out_sc ),
    .A2(_0639_));
 sg13g2_a21oi_1 _4125_ (.A1(_0962_),
    .A2(_0963_),
    .Y(_0965_),
    .B1(_0964_));
 sg13g2_or4_1 _4126_ (.A(net28),
    .B(_0708_),
    .C(_0730_),
    .D(_0733_),
    .X(_0966_));
 sg13g2_nand2_1 _4127_ (.Y(_0967_),
    .A(net28),
    .B(_0707_));
 sg13g2_a221oi_1 _4128_ (.B2(_0706_),
    .C1(_0967_),
    .B1(_0702_),
    .A1(_0695_),
    .Y(_0968_),
    .A2(_0697_));
 sg13g2_or2_1 _4129_ (.X(_0969_),
    .B(\g.g_y[4].g_x[5].t.out_sc ),
    .A(net56));
 sg13g2_buf_1 _4130_ (.A(_0969_),
    .X(_0970_));
 sg13g2_nor2_1 _4131_ (.A(net28),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_nor3_1 _4132_ (.A(_0711_),
    .B(net56),
    .C(_0716_),
    .Y(_0972_));
 sg13g2_nor4_1 _4133_ (.A(_0634_),
    .B(_0968_),
    .C(_0971_),
    .D(_0972_),
    .Y(_0973_));
 sg13g2_a22oi_1 _4134_ (.Y(_0974_),
    .B1(_0966_),
    .B2(_0973_),
    .A2(_0965_),
    .A1(_0961_));
 sg13g2_or2_1 _4135_ (.X(_0975_),
    .B(_0974_),
    .A(_0328_));
 sg13g2_a21oi_1 _4136_ (.A1(_0951_),
    .A2(_0975_),
    .Y(_0084_),
    .B1(net136));
 sg13g2_inv_1 _4137_ (.Y(_0976_),
    .A(net23));
 sg13g2_nor2b_1 _4138_ (.A(_0638_),
    .B_N(net58),
    .Y(_0977_));
 sg13g2_nor2_1 _4139_ (.A(net58),
    .B(net23),
    .Y(_0978_));
 sg13g2_o21ai_1 _4140_ (.B1(_0962_),
    .Y(_0979_),
    .A1(_0977_),
    .A2(_0978_));
 sg13g2_a21o_1 _4141_ (.A2(_0957_),
    .A1(net60),
    .B1(_0622_),
    .X(_0980_));
 sg13g2_mux4_1 _4142_ (.S0(net58),
    .A0(\g.g_y[4].g_x[7].t.out_sc ),
    .A1(_0976_),
    .A2(_0979_),
    .A3(_0980_),
    .S1(net59),
    .X(_0981_));
 sg13g2_nor3_1 _4143_ (.A(_0708_),
    .B(_0730_),
    .C(_0733_),
    .Y(_0982_));
 sg13g2_nand2_1 _4144_ (.Y(_0983_),
    .A(_0711_),
    .B(_0970_));
 sg13g2_or3_1 _4145_ (.A(_0711_),
    .B(_0710_),
    .C(_0722_),
    .X(_0984_));
 sg13g2_o21ai_1 _4146_ (.B1(_0984_),
    .Y(_0985_),
    .A1(_0982_),
    .A2(_0983_));
 sg13g2_mux2_1 _4147_ (.A0(_0981_),
    .A1(_0985_),
    .S(_0634_),
    .X(_0986_));
 sg13g2_a21oi_1 _4148_ (.A1(_0945_),
    .A2(_0949_),
    .Y(_0987_),
    .B1(_0327_));
 sg13g2_nor3_1 _4149_ (.A(_0325_),
    .B(_0910_),
    .C(_0913_),
    .Y(_0988_));
 sg13g2_or2_1 _4150_ (.X(_0989_),
    .B(_0988_),
    .A(_0987_));
 sg13g2_a21oi_1 _4151_ (.A1(_0986_),
    .A2(_0989_),
    .Y(_0085_),
    .B1(net136));
 sg13g2_and2_1 _4152_ (.A(\g.g_y[4].g_x[6].t.out_sc ),
    .B(net151),
    .X(_0083_));
 sg13g2_and2_1 _4153_ (.A(\g.g_y[4].g_x[5].t.out_sc ),
    .B(net168),
    .X(_0082_));
 sg13g2_buf_2 _4154_ (.A(\g.g_y[3].g_x[4].t.r_d ),
    .X(_0990_));
 sg13g2_inv_1 _4155_ (.Y(_0991_),
    .A(_0990_));
 sg13g2_buf_2 _4156_ (.A(\g.g_y[2].g_x[4].t.r_ghl ),
    .X(_0992_));
 sg13g2_buf_2 _4157_ (.A(\g.g_y[2].g_x[4].t.r_d ),
    .X(_0993_));
 sg13g2_mux2_1 _4158_ (.A0(\g.g_y[2].g_x[4].t.r_gnl ),
    .A1(\g.g_y[2].g_x[4].t.out_sc ),
    .S(_0993_),
    .X(_0994_));
 sg13g2_buf_1 _4159_ (.A(_0994_),
    .X(_0995_));
 sg13g2_buf_2 _4160_ (.A(\g.g_y[2].g_x[4].t.r_v ),
    .X(_0996_));
 sg13g2_mux2_1 _4161_ (.A0(_0992_),
    .A1(_0995_),
    .S(_0996_),
    .X(_0997_));
 sg13g2_buf_2 _4162_ (.A(_0997_),
    .X(_0998_));
 sg13g2_nor2_1 _4163_ (.A(net25),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_buf_1 _4164_ (.A(\g.g_y[3].g_x[4].t.r_h ),
    .X(_1000_));
 sg13g2_mux2_1 _4165_ (.A0(_0698_),
    .A1(_0916_),
    .S(_0915_),
    .X(_1001_));
 sg13g2_buf_1 _4166_ (.A(_1001_),
    .X(_1002_));
 sg13g2_buf_2 _4167_ (.A(\g.g_y[3].g_x[3].t.r_h ),
    .X(_1003_));
 sg13g2_nor2_1 _4168_ (.A(_0791_),
    .B(_1003_),
    .Y(_1004_));
 sg13g2_nor2_1 _4169_ (.A(net47),
    .B(_1004_),
    .Y(_1005_));
 sg13g2_inv_1 _4170_ (.Y(_1006_),
    .A(_1003_));
 sg13g2_mux2_1 _4171_ (.A0(\g.g_y[3].g_x[3].t.out_sc ),
    .A1(\g.g_y[3].g_x[3].t.r_gnl ),
    .S(_0796_),
    .X(_1007_));
 sg13g2_buf_1 _4172_ (.A(_1007_),
    .X(_1008_));
 sg13g2_or2_1 _4173_ (.X(_1009_),
    .B(_1008_),
    .A(_1006_));
 sg13g2_buf_1 _4174_ (.A(_1009_),
    .X(_1010_));
 sg13g2_a221oi_1 _4175_ (.B2(_1010_),
    .C1(_0990_),
    .B1(_1005_),
    .A1(net47),
    .Y(_1011_),
    .A2(_1002_));
 sg13g2_buf_1 _4176_ (.A(_1011_),
    .X(_1012_));
 sg13g2_buf_1 _4177_ (.A(\g.g_y[3].g_x[4].t.r_v ),
    .X(_1013_));
 sg13g2_inv_1 _4178_ (.Y(_1014_),
    .A(net46));
 sg13g2_o21ai_1 _4179_ (.B1(_1014_),
    .Y(_1015_),
    .A1(_0999_),
    .A2(_1012_));
 sg13g2_mux2_1 _4180_ (.A0(_0791_),
    .A1(_1008_),
    .S(_1003_),
    .X(_1016_));
 sg13g2_inv_1 _4181_ (.Y(_1017_),
    .A(net47));
 sg13g2_mux2_1 _4182_ (.A0(_1016_),
    .A1(_1002_),
    .S(_1017_),
    .X(_1018_));
 sg13g2_nand4_1 _4183_ (.B(net25),
    .C(_0998_),
    .A(net46),
    .Y(_1019_),
    .D(_1018_));
 sg13g2_nor2_1 _4184_ (.A(net25),
    .B(\g.g_y[3].g_x[4].t.out_sc ),
    .Y(_1020_));
 sg13g2_a21oi_1 _4185_ (.A1(net46),
    .A2(_1020_),
    .Y(_1021_),
    .B1(_0396_));
 sg13g2_and3_1 _4186_ (.X(_1022_),
    .A(_1015_),
    .B(_1019_),
    .C(_1021_));
 sg13g2_nand2b_1 _4187_ (.Y(_1023_),
    .B(_2650_),
    .A_N(_2587_));
 sg13g2_o21ai_1 _4188_ (.B1(_1023_),
    .Y(_1024_),
    .A1(_2650_),
    .A2(_2652_));
 sg13g2_nor4_1 _4189_ (.A(net62),
    .B(net63),
    .C(_1024_),
    .D(_0418_),
    .Y(_1025_));
 sg13g2_mux2_1 _4190_ (.A0(_0410_),
    .A1(_0739_),
    .S(_0408_),
    .X(_1026_));
 sg13g2_nand2_1 _4191_ (.Y(_1027_),
    .A(net62),
    .B(_0389_));
 sg13g2_nor2_1 _4192_ (.A(_0393_),
    .B(_0389_),
    .Y(_1028_));
 sg13g2_nor2_1 _4193_ (.A(net62),
    .B(_0390_),
    .Y(_1029_));
 sg13g2_a22oi_1 _4194_ (.Y(_1030_),
    .B1(_1029_),
    .B2(net63),
    .A2(_1028_),
    .A1(_1024_));
 sg13g2_o21ai_1 _4195_ (.B1(_1030_),
    .Y(_1031_),
    .A1(_1026_),
    .A2(_1027_));
 sg13g2_nor3_1 _4196_ (.A(_0397_),
    .B(_1025_),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_o21ai_1 _4197_ (.B1(_0398_),
    .Y(_1033_),
    .A1(_1022_),
    .A2(_1032_));
 sg13g2_nand3_1 _4198_ (.B(net28),
    .C(_0970_),
    .A(net55),
    .Y(_1034_));
 sg13g2_nand2_1 _4199_ (.Y(_1035_),
    .A(net55),
    .B(_0711_));
 sg13g2_or3_1 _4200_ (.A(_0710_),
    .B(_0722_),
    .C(_1035_),
    .X(_1036_));
 sg13g2_o21ai_1 _4201_ (.B1(_1036_),
    .Y(_1037_),
    .A1(_0982_),
    .A2(_1034_));
 sg13g2_nor4_1 _4202_ (.A(_0779_),
    .B(_0777_),
    .C(_0806_),
    .D(_0841_),
    .Y(_1038_));
 sg13g2_nand2_1 _4203_ (.Y(_1039_),
    .A(_0779_),
    .B(net54));
 sg13g2_nor2_1 _4204_ (.A(net54),
    .B(net164),
    .Y(_1040_));
 sg13g2_nor2_1 _4205_ (.A(net53),
    .B(net54),
    .Y(_1041_));
 sg13g2_a22oi_1 _4206_ (.Y(_1042_),
    .B1(_1041_),
    .B2(_0841_),
    .A2(_1040_),
    .A1(net53));
 sg13g2_o21ai_1 _4207_ (.B1(_1042_),
    .Y(_1043_),
    .A1(_0838_),
    .A2(_1039_));
 sg13g2_nor3_1 _4208_ (.A(net55),
    .B(_1038_),
    .C(_1043_),
    .Y(_1044_));
 sg13g2_inv_1 _4209_ (.Y(_1045_),
    .A(_0398_));
 sg13g2_o21ai_1 _4210_ (.B1(_1045_),
    .Y(_1046_),
    .A1(_1037_),
    .A2(_1044_));
 sg13g2_a21oi_1 _4211_ (.A1(_1033_),
    .A2(_1046_),
    .Y(_0080_),
    .B1(net136));
 sg13g2_nor2_1 _4212_ (.A(_1038_),
    .B(_1043_),
    .Y(_1047_));
 sg13g2_nand3b_1 _4213_ (.B(net28),
    .C(_0970_),
    .Y(_1048_),
    .A_N(net55));
 sg13g2_or4_1 _4214_ (.A(net55),
    .B(net28),
    .C(_0710_),
    .D(_0722_),
    .X(_1049_));
 sg13g2_o21ai_1 _4215_ (.B1(_1049_),
    .Y(_1050_),
    .A1(_0982_),
    .A2(_1048_));
 sg13g2_a21o_1 _4216_ (.A2(_1047_),
    .A1(_0714_),
    .B1(_1050_),
    .X(_1051_));
 sg13g2_o21ai_1 _4217_ (.B1(_0397_),
    .Y(_1052_),
    .A1(_1025_),
    .A2(_1031_));
 sg13g2_mux2_1 _4218_ (.A0(_0403_),
    .A1(_0400_),
    .S(_0397_),
    .X(_1053_));
 sg13g2_mux2_1 _4219_ (.A0(_0998_),
    .A1(_1053_),
    .S(_1014_),
    .X(_1054_));
 sg13g2_nand3_1 _4220_ (.B(_1054_),
    .C(_1018_),
    .A(net25),
    .Y(_1055_));
 sg13g2_buf_1 _4221_ (.A(_1055_),
    .X(_1056_));
 sg13g2_nor2_1 _4222_ (.A(_1014_),
    .B(_1020_),
    .Y(_1057_));
 sg13g2_o21ai_1 _4223_ (.B1(_1014_),
    .Y(_1058_),
    .A1(net25),
    .A2(_0998_));
 sg13g2_o21ai_1 _4224_ (.B1(_0396_),
    .Y(_1059_),
    .A1(_1012_),
    .A2(_1058_));
 sg13g2_a21o_1 _4225_ (.A2(_1057_),
    .A1(_1056_),
    .B1(_1059_),
    .X(_1060_));
 sg13g2_and2_1 _4226_ (.A(_1052_),
    .B(_1060_),
    .X(_1061_));
 sg13g2_a21oi_1 _4227_ (.A1(_1051_),
    .A2(_1061_),
    .Y(_0081_),
    .B1(net136));
 sg13g2_buf_1 _4228_ (.A(net165),
    .X(_1062_));
 sg13g2_and2_1 _4229_ (.A(\g.g_y[4].g_x[4].t.out_sc ),
    .B(net150),
    .X(_0079_));
 sg13g2_and2_1 _4230_ (.A(net164),
    .B(net150),
    .X(_0078_));
 sg13g2_buf_1 _4231_ (.A(\g.g_y[3].g_x[2].t.r_d ),
    .X(_1063_));
 sg13g2_buf_2 _4232_ (.A(\g.g_y[3].g_x[2].t.r_h ),
    .X(_1064_));
 sg13g2_inv_2 _4233_ (.Y(_1065_),
    .A(_1064_));
 sg13g2_mux2_1 _4234_ (.A0(_0791_),
    .A1(_1008_),
    .S(_1006_),
    .X(_1066_));
 sg13g2_buf_2 _4235_ (.A(\g.g_y[3].g_x[1].t.r_h ),
    .X(_1067_));
 sg13g2_inv_1 _4236_ (.Y(_1068_),
    .A(_1067_));
 sg13g2_mux2_1 _4237_ (.A0(\g.g_y[3].g_x[1].t.out_sc ),
    .A1(\g.g_y[3].g_x[1].t.r_gnl ),
    .S(_0859_),
    .X(_1069_));
 sg13g2_or2_1 _4238_ (.X(_1070_),
    .B(_1069_),
    .A(_1068_));
 sg13g2_buf_1 _4239_ (.A(_1070_),
    .X(_1071_));
 sg13g2_nor2_1 _4240_ (.A(_0862_),
    .B(_1067_),
    .Y(_1072_));
 sg13g2_nor2_1 _4241_ (.A(_1065_),
    .B(_1072_),
    .Y(_1073_));
 sg13g2_a22oi_1 _4242_ (.Y(_1074_),
    .B1(_1071_),
    .B2(_1073_),
    .A2(_1066_),
    .A1(_1065_));
 sg13g2_buf_1 _4243_ (.A(\g.g_y[3].g_x[2].t.r_v ),
    .X(_1075_));
 sg13g2_inv_1 _4244_ (.Y(_1076_),
    .A(net44));
 sg13g2_mux2_1 _4245_ (.A0(_0477_),
    .A1(_0479_),
    .S(_0500_),
    .X(_1077_));
 sg13g2_buf_2 _4246_ (.A(_1077_),
    .X(_1078_));
 sg13g2_buf_2 _4247_ (.A(\g.g_y[2].g_x[2].t.r_v ),
    .X(_1079_));
 sg13g2_inv_1 _4248_ (.Y(_1080_),
    .A(_1079_));
 sg13g2_buf_8 _4249_ (.A(\g.g_y[2].g_x[2].t.r_d ),
    .X(_1081_));
 sg13g2_mux2_1 _4250_ (.A0(\g.g_y[2].g_x[2].t.r_gnl ),
    .A1(\g.g_y[2].g_x[2].t.out_sc ),
    .S(_1081_),
    .X(_1082_));
 sg13g2_or2_1 _4251_ (.X(_1083_),
    .B(_1082_),
    .A(_1080_));
 sg13g2_buf_1 _4252_ (.A(_1083_),
    .X(_1084_));
 sg13g2_buf_1 _4253_ (.A(\g.g_y[2].g_x[2].t.r_ghl ),
    .X(_1085_));
 sg13g2_nor2_1 _4254_ (.A(_1085_),
    .B(_1079_),
    .Y(_1086_));
 sg13g2_nor2_1 _4255_ (.A(_1076_),
    .B(_1086_),
    .Y(_1087_));
 sg13g2_a22oi_1 _4256_ (.Y(_1088_),
    .B1(_1084_),
    .B2(_1087_),
    .A2(_1078_),
    .A1(_1076_));
 sg13g2_nor3_1 _4257_ (.A(net45),
    .B(_1074_),
    .C(_1088_),
    .Y(_1089_));
 sg13g2_inv_1 _4258_ (.Y(_1090_),
    .A(\g.g_y[3].g_x[2].t.out_sc ));
 sg13g2_nand2_1 _4259_ (.Y(_1091_),
    .A(net45),
    .B(_1090_));
 sg13g2_nand3_1 _4260_ (.B(net44),
    .C(_1091_),
    .A(_0500_),
    .Y(_1092_));
 sg13g2_nor2_1 _4261_ (.A(_1064_),
    .B(_1072_),
    .Y(_1093_));
 sg13g2_a221oi_1 _4262_ (.B2(_1093_),
    .C1(net45),
    .B1(_1071_),
    .A1(_1064_),
    .Y(_1094_),
    .A2(_1066_));
 sg13g2_buf_1 _4263_ (.A(_1094_),
    .X(_1095_));
 sg13g2_nor2_1 _4264_ (.A(net44),
    .B(_1086_),
    .Y(_1096_));
 sg13g2_inv_1 _4265_ (.Y(_1097_),
    .A(_1063_));
 sg13g2_a221oi_1 _4266_ (.B2(_1096_),
    .C1(_1097_),
    .B1(_1084_),
    .A1(net44),
    .Y(_1098_),
    .A2(_1078_));
 sg13g2_or4_1 _4267_ (.A(_0480_),
    .B(net44),
    .C(_1095_),
    .D(_1098_),
    .X(_1099_));
 sg13g2_o21ai_1 _4268_ (.B1(_1099_),
    .Y(_1100_),
    .A1(_1089_),
    .A2(_1092_));
 sg13g2_and4_1 _4269_ (.A(_0485_),
    .B(_0476_),
    .C(_0483_),
    .D(_0495_),
    .X(_1101_));
 sg13g2_a22oi_1 _4270_ (.Y(_1102_),
    .B1(_0507_),
    .B2(_0508_),
    .A2(_0492_),
    .A1(_0493_));
 sg13g2_nor2_1 _4271_ (.A(_0485_),
    .B(net29),
    .Y(_1103_));
 sg13g2_nand2_1 _4272_ (.Y(_1104_),
    .A(_0484_),
    .B(net29));
 sg13g2_nand2b_1 _4273_ (.Y(_1105_),
    .B(_0485_),
    .A_N(_0497_));
 sg13g2_o21ai_1 _4274_ (.B1(_1105_),
    .Y(_1106_),
    .A1(_0483_),
    .A2(_1104_));
 sg13g2_a21o_1 _4275_ (.A2(_1103_),
    .A1(_1102_),
    .B1(_1106_),
    .X(_1107_));
 sg13g2_nor3_1 _4276_ (.A(_0500_),
    .B(_1101_),
    .C(_1107_),
    .Y(_1108_));
 sg13g2_o21ai_1 _4277_ (.B1(_0478_),
    .Y(_1109_),
    .A1(_1100_),
    .A2(_1108_));
 sg13g2_nand2b_1 _4278_ (.Y(_1110_),
    .B(_0270_),
    .A_N(_0274_));
 sg13g2_o21ai_1 _4279_ (.B1(_1110_),
    .Y(_1111_),
    .A1(_0270_),
    .A2(_0273_));
 sg13g2_mux2_1 _4280_ (.A0(_0864_),
    .A1(_1111_),
    .S(net52),
    .X(_1112_));
 sg13g2_buf_1 _4281_ (.A(_1112_),
    .X(_1113_));
 sg13g2_or2_1 _4282_ (.X(_1114_),
    .B(_0629_),
    .A(_0867_));
 sg13g2_nor2b_1 _4283_ (.A(_0871_),
    .B_N(_0869_),
    .Y(_1115_));
 sg13g2_a221oi_1 _4284_ (.B2(_1115_),
    .C1(net51),
    .B1(_1114_),
    .A1(net26),
    .Y(_1116_),
    .A2(_0876_));
 sg13g2_a21o_1 _4285_ (.A2(_1113_),
    .A1(net27),
    .B1(_1116_),
    .X(_1117_));
 sg13g2_nor2_1 _4286_ (.A(_0782_),
    .B(net26),
    .Y(_1118_));
 sg13g2_and3_1 _4287_ (.X(_1119_),
    .A(_0839_),
    .B(net26),
    .C(net27));
 sg13g2_a21o_1 _4288_ (.A2(_0861_),
    .A1(net50),
    .B1(_0863_),
    .X(_1120_));
 sg13g2_nand2_1 _4289_ (.Y(_1121_),
    .A(_0854_),
    .B(_1120_));
 sg13g2_mux2_1 _4290_ (.A0(_0274_),
    .A1(_0273_),
    .S(_0886_),
    .X(_1122_));
 sg13g2_nand2_1 _4291_ (.Y(_1123_),
    .A(_0855_),
    .B(_1122_));
 sg13g2_a21oi_1 _4292_ (.A1(_1121_),
    .A2(_1123_),
    .Y(_1124_),
    .B1(_0873_));
 sg13g2_nand2b_1 _4293_ (.Y(_1125_),
    .B(net26),
    .A_N(net51));
 sg13g2_nor3_1 _4294_ (.A(_0782_),
    .B(_0882_),
    .C(_1125_),
    .Y(_1126_));
 sg13g2_a221oi_1 _4295_ (.B2(_1124_),
    .C1(_1126_),
    .B1(_1119_),
    .A1(_1117_),
    .Y(_1127_),
    .A2(_1118_));
 sg13g2_nor2_1 _4296_ (.A(_0839_),
    .B(_0779_),
    .Y(_1128_));
 sg13g2_nor3_1 _4297_ (.A(_0839_),
    .B(net53),
    .C(_0777_),
    .Y(_1129_));
 sg13g2_nor4_1 _4298_ (.A(_0839_),
    .B(net53),
    .C(net54),
    .D(net164),
    .Y(_1130_));
 sg13g2_a221oi_1 _4299_ (.B2(_0809_),
    .C1(_1130_),
    .B1(_1129_),
    .A1(_0800_),
    .Y(_1131_),
    .A2(_1128_));
 sg13g2_nand3b_1 _4300_ (.B(_1127_),
    .C(_1131_),
    .Y(_1132_),
    .A_N(_0478_));
 sg13g2_a21oi_1 _4301_ (.A1(_1109_),
    .A2(_1132_),
    .Y(_0076_),
    .B1(_0829_));
 sg13g2_inv_1 _4302_ (.Y(_1133_),
    .A(_1113_));
 sg13g2_a21o_1 _4303_ (.A2(_1123_),
    .A1(_1121_),
    .B1(_0873_),
    .X(_1134_));
 sg13g2_mux4_1 _4304_ (.S0(net27),
    .A0(_0878_),
    .A1(_1133_),
    .A2(_0882_),
    .A3(_1134_),
    .S1(net26),
    .X(_1135_));
 sg13g2_mux4_1 _4305_ (.S0(net54),
    .A0(_0810_),
    .A1(_0835_),
    .A2(_0844_),
    .A3(_0838_),
    .S1(_0778_),
    .X(_1136_));
 sg13g2_mux2_1 _4306_ (.A0(_1135_),
    .A1(_1136_),
    .S(_0839_),
    .X(_1137_));
 sg13g2_nand2_1 _4307_ (.Y(_1138_),
    .A(_1075_),
    .B(_1091_));
 sg13g2_or3_1 _4308_ (.A(_1075_),
    .B(_1095_),
    .C(_1098_),
    .X(_1139_));
 sg13g2_o21ai_1 _4309_ (.B1(_1139_),
    .Y(_1140_),
    .A1(_1089_),
    .A2(_1138_));
 sg13g2_nor3_1 _4310_ (.A(_0480_),
    .B(_1101_),
    .C(_1107_),
    .Y(_1141_));
 sg13g2_a21o_1 _4311_ (.A2(_1140_),
    .A1(_0480_),
    .B1(_1141_),
    .X(_1142_));
 sg13g2_a21oi_1 _4312_ (.A1(_1137_),
    .A2(_1142_),
    .Y(_0077_),
    .B1(net136));
 sg13g2_and2_1 _4313_ (.A(\g.g_y[4].g_x[2].t.out_sc ),
    .B(_1062_),
    .X(_0075_));
 sg13g2_nor2_1 _4314_ (.A(_0883_),
    .B(net138),
    .Y(_0074_));
 sg13g2_o21ai_1 _4315_ (.B1(_0658_),
    .Y(_1143_),
    .A1(_2404_),
    .A2(_2411_));
 sg13g2_and2_1 _4316_ (.A(_0650_),
    .B(_0585_),
    .X(_1144_));
 sg13g2_o21ai_1 _4317_ (.B1(_1144_),
    .Y(_1145_),
    .A1(_0584_),
    .A2(_1143_));
 sg13g2_a21oi_1 _4318_ (.A1(_0561_),
    .A2(_1143_),
    .Y(_1146_),
    .B1(_0650_));
 sg13g2_o21ai_1 _4319_ (.B1(_1146_),
    .Y(_1147_),
    .A1(net61),
    .A2(_0566_));
 sg13g2_nand3_1 _4320_ (.B(_1145_),
    .C(_1147_),
    .A(_0567_),
    .Y(_1148_));
 sg13g2_inv_1 _4321_ (.Y(_1149_),
    .A(\g.g_y[3].g_x[0].t.r_h ));
 sg13g2_nor3_1 _4322_ (.A(_1067_),
    .B(_1149_),
    .C(_1069_),
    .Y(_1150_));
 sg13g2_nand2b_1 _4323_ (.Y(_1151_),
    .B(_1067_),
    .A_N(_0862_));
 sg13g2_or2_1 _4324_ (.X(_1152_),
    .B(\g.g_y[3].g_x[0].t.r_h ),
    .A(net4));
 sg13g2_o21ai_1 _4325_ (.B1(_1152_),
    .Y(_1153_),
    .A1(_1149_),
    .A2(_1151_));
 sg13g2_buf_1 _4326_ (.A(\g.g_y[3].g_x[0].t.r_d ),
    .X(_1154_));
 sg13g2_inv_1 _4327_ (.Y(_1155_),
    .A(net43));
 sg13g2_o21ai_1 _4328_ (.B1(_1155_),
    .Y(_1156_),
    .A1(_1150_),
    .A2(_1153_));
 sg13g2_buf_2 _4329_ (.A(\g.g_y[2].g_x[0].t.r_v ),
    .X(_1157_));
 sg13g2_inv_1 _4330_ (.Y(_1158_),
    .A(_1157_));
 sg13g2_buf_8 _4331_ (.A(\g.g_y[2].g_x[0].t.r_d ),
    .X(_1159_));
 sg13g2_mux2_1 _4332_ (.A0(\g.g_y[2].g_x[0].t.r_gnl ),
    .A1(\g.g_y[2].g_x[0].t.out_sc ),
    .S(_1159_),
    .X(_1160_));
 sg13g2_buf_2 _4333_ (.A(_1160_),
    .X(_1161_));
 sg13g2_buf_2 _4334_ (.A(\g.g_y[2].g_x[0].t.r_ghl ),
    .X(_1162_));
 sg13g2_or2_1 _4335_ (.X(_1163_),
    .B(_1157_),
    .A(_1162_));
 sg13g2_buf_1 _4336_ (.A(_1163_),
    .X(_1164_));
 sg13g2_o21ai_1 _4337_ (.B1(_1164_),
    .Y(_1165_),
    .A1(_1158_),
    .A2(_1161_));
 sg13g2_buf_1 _4338_ (.A(\g.g_y[3].g_x[0].t.r_v ),
    .X(_1166_));
 sg13g2_a21oi_1 _4339_ (.A1(net43),
    .A2(_1165_),
    .Y(_1167_),
    .B1(net42));
 sg13g2_nand2_1 _4340_ (.Y(_1168_),
    .A(_1156_),
    .B(_1167_));
 sg13g2_inv_1 _4341_ (.Y(_1169_),
    .A(net4));
 sg13g2_nor2_1 _4342_ (.A(_1169_),
    .B(_1149_),
    .Y(_1170_));
 sg13g2_and3_1 _4343_ (.X(_1171_),
    .A(_1149_),
    .B(_1155_),
    .C(_1151_));
 sg13g2_nand2b_1 _4344_ (.Y(_1172_),
    .B(_1068_),
    .A_N(_1069_));
 sg13g2_a22oi_1 _4345_ (.Y(_1173_),
    .B1(_1171_),
    .B2(_1172_),
    .A2(_1170_),
    .A1(_1155_));
 sg13g2_nand2b_1 _4346_ (.Y(_1174_),
    .B(_1154_),
    .A_N(\g.g_y[3].g_x[0].t.out_sc ));
 sg13g2_and2_1 _4347_ (.A(net42),
    .B(_1174_),
    .X(_1175_));
 sg13g2_o21ai_1 _4348_ (.B1(_1175_),
    .Y(_1176_),
    .A1(_1165_),
    .A2(_1173_));
 sg13g2_nand3_1 _4349_ (.B(_1168_),
    .C(_1176_),
    .A(_0568_),
    .Y(_1177_));
 sg13g2_nand3_1 _4350_ (.B(_1148_),
    .C(_1177_),
    .A(_0569_),
    .Y(_1178_));
 sg13g2_mux2_1 _4351_ (.A0(_1120_),
    .A1(_1122_),
    .S(_0855_),
    .X(_1179_));
 sg13g2_nand3b_1 _4352_ (.B(net27),
    .C(_1179_),
    .Y(_1180_),
    .A_N(_0873_));
 sg13g2_or2_1 _4353_ (.X(_1181_),
    .B(_0882_),
    .A(net27));
 sg13g2_nand3b_1 _4354_ (.B(_1180_),
    .C(_1181_),
    .Y(_1182_),
    .A_N(net26));
 sg13g2_a21oi_1 _4355_ (.A1(net27),
    .A2(_1113_),
    .Y(_1183_),
    .B1(_1116_));
 sg13g2_a21oi_1 _4356_ (.A1(_0877_),
    .A2(_1183_),
    .Y(_1184_),
    .B1(_0867_));
 sg13g2_inv_1 _4357_ (.Y(_1185_),
    .A(net5));
 sg13g2_a21o_1 _4358_ (.A2(_1185_),
    .A1(_0867_),
    .B1(_0569_),
    .X(_1186_));
 sg13g2_a21o_1 _4359_ (.A2(_1184_),
    .A1(_1182_),
    .B1(_1186_),
    .X(_1187_));
 sg13g2_a21oi_1 _4360_ (.A1(_1178_),
    .A2(_1187_),
    .Y(_0072_),
    .B1(_0829_));
 sg13g2_nand2_1 _4361_ (.Y(_1188_),
    .A(_0627_),
    .B(_1185_));
 sg13g2_a21o_1 _4362_ (.A2(_1176_),
    .A1(_1168_),
    .B1(_0568_),
    .X(_1189_));
 sg13g2_a21o_1 _4363_ (.A2(_1147_),
    .A1(_1145_),
    .B1(_0567_),
    .X(_1190_));
 sg13g2_a21oi_1 _4364_ (.A1(net26),
    .A2(_1183_),
    .Y(_1191_),
    .B1(_0627_));
 sg13g2_a22oi_1 _4365_ (.Y(_1192_),
    .B1(_1191_),
    .B2(_1182_),
    .A2(_1190_),
    .A1(_1189_));
 sg13g2_buf_1 _4366_ (.A(net154),
    .X(_1193_));
 sg13g2_a21oi_1 _4367_ (.A1(_1188_),
    .A2(_1192_),
    .Y(_0073_),
    .B1(net135));
 sg13g2_and2_1 _4368_ (.A(\g.g_y[4].g_x[0].t.out_sc ),
    .B(_1062_),
    .X(_0071_));
 sg13g2_buf_2 _4369_ (.A(\g.g_y[2].g_x[7].t.r_v ),
    .X(_1194_));
 sg13g2_inv_2 _4370_ (.Y(_1195_),
    .A(_1194_));
 sg13g2_buf_1 _4371_ (.A(\g.g_y[2].g_x[7].t.r_d ),
    .X(_1196_));
 sg13g2_or2_1 _4372_ (.X(_1197_),
    .B(_2471_),
    .A(_2475_));
 sg13g2_o21ai_1 _4373_ (.B1(_1197_),
    .Y(_1198_),
    .A1(_2503_),
    .A2(_2474_));
 sg13g2_buf_2 _4374_ (.A(\g.g_y[2].g_x[0].t.r_h ),
    .X(_1199_));
 sg13g2_mux2_1 _4375_ (.A0(\g.g_y[2].g_x[0].t.out_sc ),
    .A1(\g.g_y[2].g_x[0].t.r_gnl ),
    .S(_1159_),
    .X(_1200_));
 sg13g2_nand2b_1 _4376_ (.Y(_1201_),
    .B(_1199_),
    .A_N(_1162_));
 sg13g2_o21ai_1 _4377_ (.B1(_1201_),
    .Y(_1202_),
    .A1(_1199_),
    .A2(_1200_));
 sg13g2_buf_2 _4378_ (.A(\g.g_y[2].g_x[6].t.r_h ),
    .X(_1203_));
 sg13g2_inv_2 _4379_ (.Y(_1204_),
    .A(_1203_));
 sg13g2_mux2_1 _4380_ (.A0(\g.g_y[2].g_x[6].t.out_sc ),
    .A1(\g.g_y[2].g_x[6].t.r_gnl ),
    .S(_0934_),
    .X(_1205_));
 sg13g2_buf_2 _4381_ (.A(_1205_),
    .X(_1206_));
 sg13g2_or2_1 _4382_ (.X(_1207_),
    .B(_1203_),
    .A(_0937_));
 sg13g2_buf_1 _4383_ (.A(_1207_),
    .X(_1208_));
 sg13g2_o21ai_1 _4384_ (.B1(_1208_),
    .Y(_1209_),
    .A1(_1204_),
    .A2(_1206_));
 sg13g2_mux2_1 _4385_ (.A0(_1202_),
    .A1(_1209_),
    .S(\g.g_y[2].g_x[7].t.r_h ),
    .X(_1210_));
 sg13g2_nor4_1 _4386_ (.A(_1195_),
    .B(net41),
    .C(_1198_),
    .D(_1210_),
    .Y(_1211_));
 sg13g2_mux2_1 _4387_ (.A0(_0937_),
    .A1(_1206_),
    .S(_1203_),
    .X(_1212_));
 sg13g2_inv_1 _4388_ (.Y(_1213_),
    .A(_1199_));
 sg13g2_mux2_1 _4389_ (.A0(_1162_),
    .A1(_1200_),
    .S(_1213_),
    .X(_1214_));
 sg13g2_buf_1 _4390_ (.A(_1214_),
    .X(_1215_));
 sg13g2_buf_1 _4391_ (.A(\g.g_y[2].g_x[7].t.r_h ),
    .X(_1216_));
 sg13g2_mux2_1 _4392_ (.A0(_1212_),
    .A1(_1215_),
    .S(net40),
    .X(_1217_));
 sg13g2_nor3_1 _4393_ (.A(_1194_),
    .B(net41),
    .C(_1217_),
    .Y(_1218_));
 sg13g2_mux2_1 _4394_ (.A0(_2475_),
    .A1(_2474_),
    .S(_2471_),
    .X(_1219_));
 sg13g2_nand2_1 _4395_ (.Y(_1220_),
    .A(_1195_),
    .B(net41));
 sg13g2_buf_1 _4396_ (.A(\g.g_y[2].g_x[7].t.out_sc ),
    .X(_1221_));
 sg13g2_nand3b_1 _4397_ (.B(net41),
    .C(_1194_),
    .Y(_1222_),
    .A_N(_1221_));
 sg13g2_o21ai_1 _4398_ (.B1(_1222_),
    .Y(_1223_),
    .A1(_1219_),
    .A2(_1220_));
 sg13g2_nor4_1 _4399_ (.A(_0619_),
    .B(_1211_),
    .C(_1218_),
    .D(_1223_),
    .Y(_1224_));
 sg13g2_nand2_1 _4400_ (.Y(_1225_),
    .A(_0615_),
    .B(_0957_));
 sg13g2_nand2_1 _4401_ (.Y(_1226_),
    .A(_0614_),
    .B(net23));
 sg13g2_o21ai_1 _4402_ (.B1(_1226_),
    .Y(_1227_),
    .A1(_0638_),
    .A2(_1225_));
 sg13g2_nand2_1 _4403_ (.Y(_1228_),
    .A(net60),
    .B(_0638_));
 sg13g2_o21ai_1 _4404_ (.B1(_1228_),
    .Y(_1229_),
    .A1(net23),
    .A2(_1225_));
 sg13g2_nor2_1 _4405_ (.A(_0642_),
    .B(_0625_),
    .Y(_1230_));
 sg13g2_o21ai_1 _4406_ (.B1(_0625_),
    .Y(_1231_),
    .A1(net60),
    .A2(_0623_));
 sg13g2_a21oi_1 _4407_ (.A1(net60),
    .A2(_0957_),
    .Y(_1232_),
    .B1(_1231_));
 sg13g2_nand2b_1 _4408_ (.Y(_1233_),
    .B(_0619_),
    .A_N(_1232_));
 sg13g2_a221oi_1 _4409_ (.B2(_1230_),
    .C1(_1233_),
    .B1(_1229_),
    .A1(_0643_),
    .Y(_1234_),
    .A2(_1227_));
 sg13g2_o21ai_1 _4410_ (.B1(_0616_),
    .Y(_1235_),
    .A1(_1224_),
    .A2(_1234_));
 sg13g2_nand2_1 _4411_ (.Y(_1236_),
    .A(_1151_),
    .B(_1172_));
 sg13g2_nand2b_1 _4412_ (.Y(_1237_),
    .B(_0568_),
    .A_N(_0571_));
 sg13g2_nand2b_1 _4413_ (.Y(_1238_),
    .B(_0567_),
    .A_N(_0572_));
 sg13g2_nor2b_1 _4414_ (.A(_1166_),
    .B_N(net43),
    .Y(_1239_));
 sg13g2_and2_1 _4415_ (.A(_1238_),
    .B(_1239_),
    .X(_1240_));
 sg13g2_and3_1 _4416_ (.X(_1241_),
    .A(net42),
    .B(net43),
    .C(_1164_));
 sg13g2_or2_1 _4417_ (.X(_1242_),
    .B(_1161_),
    .A(_1158_));
 sg13g2_buf_1 _4418_ (.A(_1242_),
    .X(_1243_));
 sg13g2_a22oi_1 _4419_ (.Y(_1244_),
    .B1(_1241_),
    .B2(_1243_),
    .A2(_1240_),
    .A1(_1237_));
 sg13g2_nor2_1 _4420_ (.A(net43),
    .B(\g.g_y[3].g_x[0].t.out_sc ),
    .Y(_1245_));
 sg13g2_nor2_1 _4421_ (.A(\g.g_y[3].g_x[0].t.r_h ),
    .B(_1245_),
    .Y(_1246_));
 sg13g2_o21ai_1 _4422_ (.B1(_1246_),
    .Y(_1247_),
    .A1(_1236_),
    .A2(_1244_));
 sg13g2_mux2_1 _4423_ (.A0(_0572_),
    .A1(_0571_),
    .S(_0568_),
    .X(_1248_));
 sg13g2_nor2b_1 _4424_ (.A(net42),
    .B_N(_1164_),
    .Y(_1249_));
 sg13g2_a221oi_1 _4425_ (.B2(_1243_),
    .C1(_1155_),
    .B1(_1249_),
    .A1(net42),
    .Y(_1250_),
    .A2(_1248_));
 sg13g2_nand3b_1 _4426_ (.B(\g.g_y[3].g_x[0].t.r_h ),
    .C(_1156_),
    .Y(_1251_),
    .A_N(_1250_));
 sg13g2_nand3_1 _4427_ (.B(_1247_),
    .C(_1251_),
    .A(_0924_),
    .Y(_1252_));
 sg13g2_mux2_1 _4428_ (.A0(_0324_),
    .A1(_0329_),
    .S(_0327_),
    .X(_1253_));
 sg13g2_buf_1 _4429_ (.A(_1253_),
    .X(_1254_));
 sg13g2_nor2b_1 _4430_ (.A(net48),
    .B_N(_0939_),
    .Y(_1255_));
 sg13g2_or2_1 _4431_ (.X(_1256_),
    .B(_0936_),
    .A(_0933_));
 sg13g2_buf_1 _4432_ (.A(_1256_),
    .X(_1257_));
 sg13g2_inv_1 _4433_ (.Y(_1258_),
    .A(net49));
 sg13g2_a221oi_1 _4434_ (.B2(_1257_),
    .C1(_1258_),
    .B1(_1255_),
    .A1(net48),
    .Y(_1259_),
    .A2(_1254_));
 sg13g2_o21ai_1 _4435_ (.B1(_0921_),
    .Y(_1260_),
    .A1(_0915_),
    .A2(_0916_));
 sg13g2_a21oi_1 _4436_ (.A1(_1258_),
    .A2(_1260_),
    .Y(_1261_),
    .B1(_0919_));
 sg13g2_nand2b_1 _4437_ (.Y(_1262_),
    .B(_1261_),
    .A_N(_1259_));
 sg13g2_nand2b_1 _4438_ (.Y(_1263_),
    .B(_0327_),
    .A_N(_0329_));
 sg13g2_nor2b_1 _4439_ (.A(_0324_),
    .B_N(_0325_),
    .Y(_1264_));
 sg13g2_nor3_1 _4440_ (.A(net48),
    .B(_1258_),
    .C(_1264_),
    .Y(_1265_));
 sg13g2_and3_1 _4441_ (.X(_1266_),
    .A(net48),
    .B(net49),
    .C(_0939_));
 sg13g2_a22oi_1 _4442_ (.Y(_1267_),
    .B1(_1266_),
    .B2(_1257_),
    .A2(_1265_),
    .A1(_1263_));
 sg13g2_nor2_1 _4443_ (.A(net49),
    .B(\g.g_y[3].g_x[6].t.out_sc ),
    .Y(_1268_));
 sg13g2_nor2_1 _4444_ (.A(_0928_),
    .B(_1268_),
    .Y(_1269_));
 sg13g2_o21ai_1 _4445_ (.B1(_1269_),
    .Y(_1270_),
    .A1(_0930_),
    .A2(_1267_));
 sg13g2_nand3_1 _4446_ (.B(_1262_),
    .C(_1270_),
    .A(_0925_),
    .Y(_1271_));
 sg13g2_nand3b_1 _4447_ (.B(_1252_),
    .C(_1271_),
    .Y(_1272_),
    .A_N(_0616_));
 sg13g2_a21oi_1 _4448_ (.A1(_1235_),
    .A2(_1272_),
    .Y(_0069_),
    .B1(net135));
 sg13g2_a21oi_1 _4449_ (.A1(_1262_),
    .A2(_1270_),
    .Y(_1273_),
    .B1(_0925_));
 sg13g2_a21oi_1 _4450_ (.A1(_1247_),
    .A2(_1251_),
    .Y(_1274_),
    .B1(_0924_));
 sg13g2_or2_1 _4451_ (.X(_1275_),
    .B(_1274_),
    .A(_1273_));
 sg13g2_a221oi_1 _4452_ (.B2(_1230_),
    .C1(_1232_),
    .B1(_1229_),
    .A1(_0643_),
    .Y(_1276_),
    .A2(_1227_));
 sg13g2_nor4_1 _4453_ (.A(_0952_),
    .B(_1211_),
    .C(_1218_),
    .D(_1223_),
    .Y(_1277_));
 sg13g2_a21o_1 _4454_ (.A2(_1276_),
    .A1(_0952_),
    .B1(_1277_),
    .X(_1278_));
 sg13g2_a21oi_1 _4455_ (.A1(_1275_),
    .A2(_1278_),
    .Y(_0070_),
    .B1(net135));
 sg13g2_and2_1 _4456_ (.A(\g.g_y[3].g_x[7].t.out_sc ),
    .B(_2498_),
    .X(_0068_));
 sg13g2_and2_1 _4457_ (.A(\g.g_y[3].g_x[6].t.out_sc ),
    .B(net150),
    .X(_0067_));
 sg13g2_buf_1 _4458_ (.A(\g.g_y[2].g_x[5].t.r_v ),
    .X(_1279_));
 sg13g2_inv_1 _4459_ (.Y(_1280_),
    .A(net39));
 sg13g2_mux2_1 _4460_ (.A0(_0698_),
    .A1(_0704_),
    .S(_0701_),
    .X(_1281_));
 sg13g2_buf_1 _4461_ (.A(_1281_),
    .X(_1282_));
 sg13g2_or2_1 _4462_ (.X(_1283_),
    .B(_2550_),
    .A(_2552_));
 sg13g2_buf_1 _4463_ (.A(_1283_),
    .X(_1284_));
 sg13g2_o21ai_1 _4464_ (.B1(\g.g_y[2].g_x[5].t.r_v ),
    .Y(_1285_),
    .A1(_2548_),
    .A2(_2551_));
 sg13g2_inv_1 _4465_ (.Y(_1286_),
    .A(_1285_));
 sg13g2_a22oi_1 _4466_ (.Y(_1287_),
    .B1(_1284_),
    .B2(_1286_),
    .A2(_1282_),
    .A1(_1280_));
 sg13g2_buf_1 _4467_ (.A(_1287_),
    .X(_1288_));
 sg13g2_nand2b_1 _4468_ (.Y(_1289_),
    .B(_1204_),
    .A_N(_1206_));
 sg13g2_buf_1 _4469_ (.A(\g.g_y[2].g_x[5].t.r_h ),
    .X(_1290_));
 sg13g2_buf_1 _4470_ (.A(\g.g_y[2].g_x[5].t.r_d ),
    .X(_1291_));
 sg13g2_nor2b_1 _4471_ (.A(_0937_),
    .B_N(_1203_),
    .Y(_1292_));
 sg13g2_nor3_1 _4472_ (.A(_1290_),
    .B(net38),
    .C(_1292_),
    .Y(_1293_));
 sg13g2_inv_1 _4473_ (.Y(_1294_),
    .A(_1290_));
 sg13g2_buf_2 _4474_ (.A(\g.g_y[2].g_x[4].t.r_h ),
    .X(_1295_));
 sg13g2_nor2_1 _4475_ (.A(_0992_),
    .B(_1295_),
    .Y(_1296_));
 sg13g2_nor3_1 _4476_ (.A(_1294_),
    .B(net38),
    .C(_1296_),
    .Y(_1297_));
 sg13g2_inv_1 _4477_ (.Y(_1298_),
    .A(_1295_));
 sg13g2_mux2_1 _4478_ (.A0(\g.g_y[2].g_x[4].t.out_sc ),
    .A1(\g.g_y[2].g_x[4].t.r_gnl ),
    .S(_0993_),
    .X(_1299_));
 sg13g2_or2_1 _4479_ (.X(_1300_),
    .B(_1299_),
    .A(_1298_));
 sg13g2_a22oi_1 _4480_ (.Y(_1301_),
    .B1(_1297_),
    .B2(_1300_),
    .A2(_1293_),
    .A1(_1289_));
 sg13g2_nand2b_1 _4481_ (.Y(_1302_),
    .B(net38),
    .A_N(\g.g_y[2].g_x[5].t.out_sc ));
 sg13g2_o21ai_1 _4482_ (.B1(_1302_),
    .Y(_1303_),
    .A1(_1288_),
    .A2(_1301_));
 sg13g2_nor2_1 _4483_ (.A(_0700_),
    .B(_1280_),
    .Y(_1304_));
 sg13g2_nand2_1 _4484_ (.Y(_1305_),
    .A(_1303_),
    .B(_1304_));
 sg13g2_nand2_1 _4485_ (.Y(_1306_),
    .A(_0700_),
    .B(_0725_));
 sg13g2_nor2_1 _4486_ (.A(net56),
    .B(_1306_),
    .Y(_1307_));
 sg13g2_nor2_1 _4487_ (.A(_0701_),
    .B(_0725_),
    .Y(_1308_));
 sg13g2_nor2_1 _4488_ (.A(_0735_),
    .B(_1306_),
    .Y(_1309_));
 sg13g2_inv_1 _4489_ (.Y(_1310_),
    .A(\g.g_y[2].g_x[5].t.r_d ));
 sg13g2_mux2_1 _4490_ (.A0(_2548_),
    .A1(_2550_),
    .S(_2551_),
    .X(_1311_));
 sg13g2_nor4_1 _4491_ (.A(_0700_),
    .B(net39),
    .C(_1310_),
    .D(_1311_),
    .Y(_1312_));
 sg13g2_mux2_1 _4492_ (.A0(_0992_),
    .A1(_1299_),
    .S(_1295_),
    .X(_1313_));
 sg13g2_buf_1 _4493_ (.A(_1313_),
    .X(_1314_));
 sg13g2_nor2_1 _4494_ (.A(_1294_),
    .B(_1292_),
    .Y(_1315_));
 sg13g2_nand3_1 _4495_ (.B(_1280_),
    .C(_1310_),
    .A(_0701_),
    .Y(_1316_));
 sg13g2_a221oi_1 _4496_ (.B2(_1315_),
    .C1(_1316_),
    .B1(_1289_),
    .A1(_1294_),
    .Y(_1317_),
    .A2(_1314_));
 sg13g2_or3_1 _4497_ (.A(_1309_),
    .B(_1312_),
    .C(_1317_),
    .X(_1318_));
 sg13g2_a221oi_1 _4498_ (.B2(_0723_),
    .C1(_1318_),
    .B1(_1308_),
    .A1(_0734_),
    .Y(_1319_),
    .A2(_1307_));
 sg13g2_nand3_1 _4499_ (.B(_1305_),
    .C(_1319_),
    .A(_0703_),
    .Y(_1320_));
 sg13g2_nor2_1 _4500_ (.A(_0990_),
    .B(\g.g_y[3].g_x[4].t.out_sc ),
    .Y(_1321_));
 sg13g2_and2_1 _4501_ (.A(net47),
    .B(_1321_),
    .X(_1322_));
 sg13g2_mux2_1 _4502_ (.A0(_0998_),
    .A1(_1053_),
    .S(net46),
    .X(_1323_));
 sg13g2_nor2_1 _4503_ (.A(_0990_),
    .B(_1004_),
    .Y(_1324_));
 sg13g2_a221oi_1 _4504_ (.B2(_1010_),
    .C1(net47),
    .B1(_1324_),
    .A1(_0990_),
    .Y(_1325_),
    .A2(_1323_));
 sg13g2_inv_1 _4505_ (.Y(_1326_),
    .A(_0996_));
 sg13g2_or2_1 _4506_ (.X(_1327_),
    .B(_0996_),
    .A(_0992_));
 sg13g2_o21ai_1 _4507_ (.B1(_1327_),
    .Y(_1328_),
    .A1(_1326_),
    .A2(_0995_));
 sg13g2_nand2b_1 _4508_ (.Y(_1329_),
    .B(_0396_),
    .A_N(_0403_));
 sg13g2_o21ai_1 _4509_ (.B1(_1329_),
    .Y(_1330_),
    .A1(_0396_),
    .A2(_0400_));
 sg13g2_mux2_1 _4510_ (.A0(_1328_),
    .A1(_1330_),
    .S(_1014_),
    .X(_1331_));
 sg13g2_nor2_1 _4511_ (.A(_1017_),
    .B(_1004_),
    .Y(_1332_));
 sg13g2_a22oi_1 _4512_ (.Y(_1333_),
    .B1(_1002_),
    .B2(_1017_),
    .A2(_1332_),
    .A1(_1010_));
 sg13g2_nor4_1 _4513_ (.A(_1017_),
    .B(net25),
    .C(_1331_),
    .D(_1333_),
    .Y(_1334_));
 sg13g2_nor4_1 _4514_ (.A(\g.g_y[3].g_x[5].t.r_h ),
    .B(_1322_),
    .C(_1325_),
    .D(_1334_),
    .Y(_1335_));
 sg13g2_o21ai_1 _4515_ (.B1(_0919_),
    .Y(_1336_),
    .A1(net49),
    .A2(_0927_));
 sg13g2_or2_1 _4516_ (.X(_1337_),
    .B(_1336_),
    .A(_1259_));
 sg13g2_nor2_1 _4517_ (.A(_0919_),
    .B(_1268_),
    .Y(_1338_));
 sg13g2_o21ai_1 _4518_ (.B1(_1338_),
    .Y(_1339_),
    .A1(_0930_),
    .A2(_1267_));
 sg13g2_a21oi_1 _4519_ (.A1(_1337_),
    .A2(_1339_),
    .Y(_1340_),
    .B1(_0915_));
 sg13g2_inv_1 _4520_ (.Y(_1341_),
    .A(_0703_));
 sg13g2_o21ai_1 _4521_ (.B1(_1341_),
    .Y(_1342_),
    .A1(_1335_),
    .A2(_1340_));
 sg13g2_a21oi_1 _4522_ (.A1(_1320_),
    .A2(_1342_),
    .Y(_0065_),
    .B1(net135));
 sg13g2_nor3_1 _4523_ (.A(_1322_),
    .B(_1325_),
    .C(_1334_),
    .Y(_1343_));
 sg13g2_nand2_1 _4524_ (.Y(_1344_),
    .A(_1337_),
    .B(_1339_));
 sg13g2_mux2_1 _4525_ (.A0(_1343_),
    .A1(_1344_),
    .S(_0915_),
    .X(_1345_));
 sg13g2_a22oi_1 _4526_ (.Y(_1346_),
    .B1(_1289_),
    .B2(_1315_),
    .A2(_1314_),
    .A1(_1294_));
 sg13g2_inv_1 _4527_ (.Y(_1347_),
    .A(_2548_));
 sg13g2_a21oi_1 _4528_ (.A1(_1347_),
    .A2(_2552_),
    .Y(_1348_),
    .B1(net39));
 sg13g2_a221oi_1 _4529_ (.B2(_1348_),
    .C1(_1310_),
    .B1(_1284_),
    .A1(net39),
    .Y(_1349_),
    .A2(_1282_));
 sg13g2_a21o_1 _4530_ (.A2(_1346_),
    .A1(_1310_),
    .B1(_1349_),
    .X(_1350_));
 sg13g2_mux2_1 _4531_ (.A0(_1303_),
    .A1(_1350_),
    .S(_1280_),
    .X(_1351_));
 sg13g2_inv_1 _4532_ (.Y(_1352_),
    .A(_0735_));
 sg13g2_or3_1 _4533_ (.A(net57),
    .B(_1352_),
    .C(_0764_),
    .X(_1353_));
 sg13g2_a21oi_1 _4534_ (.A1(net57),
    .A2(_0766_),
    .Y(_1354_),
    .B1(_0700_));
 sg13g2_a22oi_1 _4535_ (.Y(_1355_),
    .B1(_1353_),
    .B2(_1354_),
    .A2(_1351_),
    .A1(_0700_));
 sg13g2_a21oi_1 _4536_ (.A1(_1345_),
    .A2(_1355_),
    .Y(_0066_),
    .B1(net135));
 sg13g2_and2_1 _4537_ (.A(\g.g_y[3].g_x[5].t.out_sc ),
    .B(net150),
    .X(_0064_));
 sg13g2_and2_1 _4538_ (.A(\g.g_y[3].g_x[4].t.out_sc ),
    .B(net150),
    .X(_0063_));
 sg13g2_buf_1 _4539_ (.A(\g.g_y[2].g_x[3].t.r_v ),
    .X(_1356_));
 sg13g2_mux2_1 _4540_ (.A0(_0791_),
    .A1(_0797_),
    .S(_0794_),
    .X(_1357_));
 sg13g2_or2_1 _4541_ (.X(_1358_),
    .B(_2708_),
    .A(_2710_));
 sg13g2_nor2_1 _4542_ (.A(_2706_),
    .B(_2709_),
    .Y(_1359_));
 sg13g2_nor2_1 _4543_ (.A(net37),
    .B(_1359_),
    .Y(_1360_));
 sg13g2_buf_1 _4544_ (.A(\g.g_y[2].g_x[3].t.r_d ),
    .X(_1361_));
 sg13g2_inv_1 _4545_ (.Y(_1362_),
    .A(net36));
 sg13g2_a221oi_1 _4546_ (.B2(_1360_),
    .C1(_1362_),
    .B1(_1358_),
    .A1(net37),
    .Y(_1363_),
    .A2(_1357_));
 sg13g2_buf_1 _4547_ (.A(\g.g_y[2].g_x[3].t.r_h ),
    .X(_1364_));
 sg13g2_mux2_1 _4548_ (.A0(_0992_),
    .A1(_1299_),
    .S(_1298_),
    .X(_1365_));
 sg13g2_buf_1 _4549_ (.A(_1365_),
    .X(_1366_));
 sg13g2_inv_1 _4550_ (.Y(_1367_),
    .A(\g.g_y[2].g_x[2].t.r_h ));
 sg13g2_mux2_1 _4551_ (.A0(\g.g_y[2].g_x[2].t.out_sc ),
    .A1(\g.g_y[2].g_x[2].t.r_gnl ),
    .S(_1081_),
    .X(_1368_));
 sg13g2_or2_1 _4552_ (.X(_1369_),
    .B(_1368_),
    .A(_1367_));
 sg13g2_buf_1 _4553_ (.A(_1369_),
    .X(_1370_));
 sg13g2_nor2_1 _4554_ (.A(_1085_),
    .B(\g.g_y[2].g_x[2].t.r_h ),
    .Y(_1371_));
 sg13g2_nor2_1 _4555_ (.A(_1364_),
    .B(_1371_),
    .Y(_1372_));
 sg13g2_a221oi_1 _4556_ (.B2(_1372_),
    .C1(net36),
    .B1(_1370_),
    .A1(_1364_),
    .Y(_1373_),
    .A2(_1366_));
 sg13g2_or2_1 _4557_ (.X(_1374_),
    .B(_1373_),
    .A(_1363_));
 sg13g2_nor2_1 _4558_ (.A(_0793_),
    .B(net37),
    .Y(_1375_));
 sg13g2_nand2_1 _4559_ (.Y(_1376_),
    .A(_0794_),
    .B(net37));
 sg13g2_nor2_1 _4560_ (.A(net36),
    .B(_1376_),
    .Y(_1377_));
 sg13g2_inv_1 _4561_ (.Y(_1378_),
    .A(_1356_));
 sg13g2_nor2_1 _4562_ (.A(_1378_),
    .B(_1359_),
    .Y(_1379_));
 sg13g2_a22oi_1 _4563_ (.Y(_1380_),
    .B1(_1358_),
    .B2(_1379_),
    .A2(_1357_),
    .A1(_1378_));
 sg13g2_buf_1 _4564_ (.A(_1380_),
    .X(_1381_));
 sg13g2_inv_1 _4565_ (.Y(_1382_),
    .A(_1364_));
 sg13g2_nor2_1 _4566_ (.A(_1382_),
    .B(_1371_),
    .Y(_1383_));
 sg13g2_a22oi_1 _4567_ (.Y(_1384_),
    .B1(_1370_),
    .B2(_1383_),
    .A2(_1366_),
    .A1(_1382_));
 sg13g2_buf_1 _4568_ (.A(_1384_),
    .X(_1385_));
 sg13g2_nor2_1 _4569_ (.A(_1381_),
    .B(_1385_),
    .Y(_1386_));
 sg13g2_nand2b_1 _4570_ (.Y(_1387_),
    .B(net36),
    .A_N(\g.g_y[2].g_x[3].t.out_sc ));
 sg13g2_nor2_1 _4571_ (.A(_1387_),
    .B(_1376_),
    .Y(_1388_));
 sg13g2_a221oi_1 _4572_ (.B2(_1386_),
    .C1(_1388_),
    .B1(_1377_),
    .A1(_1374_),
    .Y(_1389_),
    .A2(_1375_));
 sg13g2_nand2_1 _4573_ (.Y(_1390_),
    .A(_0793_),
    .B(_0802_));
 sg13g2_nor2_1 _4574_ (.A(net54),
    .B(_1390_),
    .Y(_1391_));
 sg13g2_nor2_1 _4575_ (.A(_0794_),
    .B(_0802_),
    .Y(_1392_));
 sg13g2_nor3_1 _4576_ (.A(_0777_),
    .B(net164),
    .C(_1390_),
    .Y(_1393_));
 sg13g2_a221oi_1 _4577_ (.B2(_0800_),
    .C1(_1393_),
    .B1(_1392_),
    .A1(_0809_),
    .Y(_1394_),
    .A2(_1391_));
 sg13g2_inv_1 _4578_ (.Y(_1395_),
    .A(_0796_));
 sg13g2_a21oi_1 _4579_ (.A1(_1389_),
    .A2(_1394_),
    .Y(_1396_),
    .B1(_1395_));
 sg13g2_o21ai_1 _4580_ (.B1(_1065_),
    .Y(_1397_),
    .A1(_1095_),
    .A2(_1098_));
 sg13g2_nor2_1 _4581_ (.A(net45),
    .B(\g.g_y[3].g_x[2].t.out_sc ),
    .Y(_1398_));
 sg13g2_nor2_1 _4582_ (.A(_1065_),
    .B(_1097_),
    .Y(_1399_));
 sg13g2_nor2_1 _4583_ (.A(_1074_),
    .B(_1088_),
    .Y(_1400_));
 sg13g2_a221oi_1 _4584_ (.B2(_1400_),
    .C1(_1003_),
    .B1(_1399_),
    .A1(_1064_),
    .Y(_1401_),
    .A2(_1398_));
 sg13g2_nor3_1 _4585_ (.A(net25),
    .B(_1331_),
    .C(_1333_),
    .Y(_1402_));
 sg13g2_a21oi_1 _4586_ (.A1(_1017_),
    .A2(_1402_),
    .Y(_1403_),
    .B1(_1006_));
 sg13g2_mux2_1 _4587_ (.A0(_1328_),
    .A1(_1330_),
    .S(net46),
    .X(_1404_));
 sg13g2_a21oi_2 _4588_ (.B1(_1012_),
    .Y(_1405_),
    .A2(_1404_),
    .A1(_0990_));
 sg13g2_nor2_1 _4589_ (.A(net47),
    .B(_1321_),
    .Y(_1406_));
 sg13g2_a21o_1 _4590_ (.A2(_1405_),
    .A1(net47),
    .B1(_1406_),
    .X(_1407_));
 sg13g2_a221oi_1 _4591_ (.B2(_1407_),
    .C1(_0796_),
    .B1(_1403_),
    .A1(_1397_),
    .Y(_1408_),
    .A2(_1401_));
 sg13g2_nor3_1 _4592_ (.A(net154),
    .B(_1396_),
    .C(_1408_),
    .Y(_0061_));
 sg13g2_o21ai_1 _4593_ (.B1(_1071_),
    .Y(_1409_),
    .A1(_0862_),
    .A2(_1067_));
 sg13g2_a22oi_1 _4594_ (.Y(_1410_),
    .B1(_1084_),
    .B2(_1096_),
    .A2(_1078_),
    .A1(net44));
 sg13g2_mux4_1 _4595_ (.S0(_1065_),
    .A0(_1090_),
    .A1(_1409_),
    .A2(_1400_),
    .A3(_1410_),
    .S1(net45),
    .X(_1411_));
 sg13g2_nand3_1 _4596_ (.B(_1054_),
    .C(_1018_),
    .A(_0990_),
    .Y(_1412_));
 sg13g2_a221oi_1 _4597_ (.B2(_1412_),
    .C1(_1003_),
    .B1(_1406_),
    .A1(_1000_),
    .Y(_1413_),
    .A2(_1405_));
 sg13g2_a21oi_1 _4598_ (.A1(_1003_),
    .A2(_1411_),
    .Y(_1414_),
    .B1(_1413_));
 sg13g2_mux4_1 _4599_ (.S0(_0777_),
    .A0(net164),
    .A1(_0835_),
    .A2(_0838_),
    .A3(_0844_),
    .S1(_0789_),
    .X(_1415_));
 sg13g2_or3_1 _4600_ (.A(net36),
    .B(_1381_),
    .C(_1385_),
    .X(_1416_));
 sg13g2_and2_1 _4601_ (.A(net37),
    .B(_1387_),
    .X(_1417_));
 sg13g2_nor3_1 _4602_ (.A(net37),
    .B(_1363_),
    .C(_1373_),
    .Y(_1418_));
 sg13g2_a21o_1 _4603_ (.A2(_1417_),
    .A1(_1416_),
    .B1(_1418_),
    .X(_1419_));
 sg13g2_mux2_1 _4604_ (.A0(_1415_),
    .A1(_1419_),
    .S(_0793_),
    .X(_1420_));
 sg13g2_a21oi_1 _4605_ (.A1(_1414_),
    .A2(_1420_),
    .Y(_0062_),
    .B1(net135));
 sg13g2_and2_1 _4606_ (.A(\g.g_y[3].g_x[3].t.out_sc ),
    .B(net150),
    .X(_0060_));
 sg13g2_nor2_1 _4607_ (.A(_1090_),
    .B(net138),
    .Y(_0059_));
 sg13g2_nand2b_1 _4608_ (.Y(_1421_),
    .B(_1122_),
    .A_N(_0856_));
 sg13g2_a21oi_1 _4609_ (.A1(net51),
    .A2(_0883_),
    .Y(_1422_),
    .B1(net52));
 sg13g2_nor2_1 _4610_ (.A(net26),
    .B(net51),
    .Y(_1423_));
 sg13g2_a21oi_1 _4611_ (.A1(net52),
    .A2(_0870_),
    .Y(_1424_),
    .B1(_0876_));
 sg13g2_a221oi_1 _4612_ (.B2(_0869_),
    .C1(_1125_),
    .B1(_1114_),
    .A1(net52),
    .Y(_1425_),
    .A2(_0866_));
 sg13g2_a221oi_1 _4613_ (.B2(_1424_),
    .C1(_1425_),
    .B1(_1423_),
    .A1(_1421_),
    .Y(_1426_),
    .A2(_1422_));
 sg13g2_nand2_1 _4614_ (.Y(_1427_),
    .A(net27),
    .B(_1111_));
 sg13g2_nand3b_1 _4615_ (.B(_1123_),
    .C(_1427_),
    .Y(_1428_),
    .A_N(_1116_));
 sg13g2_nand3_1 _4616_ (.B(_1426_),
    .C(_1428_),
    .A(net50),
    .Y(_1429_));
 sg13g2_or2_1 _4617_ (.X(_1430_),
    .B(_1200_),
    .A(_1213_));
 sg13g2_buf_1 _4618_ (.A(_1430_),
    .X(_1431_));
 sg13g2_buf_1 _4619_ (.A(\g.g_y[2].g_x[1].t.r_h ),
    .X(_1432_));
 sg13g2_or2_1 _4620_ (.X(_1433_),
    .B(_1199_),
    .A(_1162_));
 sg13g2_buf_1 _4621_ (.A(_1433_),
    .X(_1434_));
 sg13g2_and2_1 _4622_ (.A(_1432_),
    .B(_1434_),
    .X(_1435_));
 sg13g2_mux2_1 _4623_ (.A0(_1085_),
    .A1(_1368_),
    .S(_1367_),
    .X(_1436_));
 sg13g2_buf_1 _4624_ (.A(_1436_),
    .X(_1437_));
 sg13g2_inv_1 _4625_ (.Y(_1438_),
    .A(_1432_));
 sg13g2_a22oi_1 _4626_ (.Y(_1439_),
    .B1(_1437_),
    .B2(_1438_),
    .A2(_1435_),
    .A1(_1431_));
 sg13g2_buf_1 _4627_ (.A(_1439_),
    .X(_1440_));
 sg13g2_buf_1 _4628_ (.A(\g.g_y[2].g_x[1].t.r_d ),
    .X(_1441_));
 sg13g2_inv_1 _4629_ (.Y(_1442_),
    .A(_1441_));
 sg13g2_mux2_1 _4630_ (.A0(_0233_),
    .A1(_0232_),
    .S(_0229_),
    .X(_1443_));
 sg13g2_nand2_1 _4631_ (.Y(_1444_),
    .A(_1442_),
    .B(_1443_));
 sg13g2_nor2_1 _4632_ (.A(_1442_),
    .B(\g.g_y[2].g_x[1].t.out_sc ),
    .Y(_1445_));
 sg13g2_buf_2 _4633_ (.A(\g.g_y[2].g_x[1].t.r_v ),
    .X(_1446_));
 sg13g2_nor2b_1 _4634_ (.A(_1445_),
    .B_N(_1446_),
    .Y(_1447_));
 sg13g2_o21ai_1 _4635_ (.B1(_1447_),
    .Y(_1448_),
    .A1(_1440_),
    .A2(_1444_));
 sg13g2_and2_1 _4636_ (.A(_1438_),
    .B(_1434_),
    .X(_1449_));
 sg13g2_a221oi_1 _4637_ (.B2(_1431_),
    .C1(_1441_),
    .B1(_1449_),
    .A1(_1432_),
    .Y(_1450_),
    .A2(_1437_));
 sg13g2_inv_1 _4638_ (.Y(_1451_),
    .A(_0229_));
 sg13g2_or2_1 _4639_ (.X(_1452_),
    .B(_0229_),
    .A(_0233_));
 sg13g2_o21ai_1 _4640_ (.B1(_1452_),
    .Y(_1453_),
    .A1(_1451_),
    .A2(_0232_));
 sg13g2_a21oi_1 _4641_ (.A1(_1441_),
    .A2(_1453_),
    .Y(_1454_),
    .B1(_1446_));
 sg13g2_nand2b_1 _4642_ (.Y(_1455_),
    .B(_1454_),
    .A_N(_1450_));
 sg13g2_nand3b_1 _4643_ (.B(_1448_),
    .C(_1455_),
    .Y(_1456_),
    .A_N(net50));
 sg13g2_nand3_1 _4644_ (.B(_1429_),
    .C(_1456_),
    .A(_0859_),
    .Y(_1457_));
 sg13g2_nand2b_1 _4645_ (.Y(_1458_),
    .B(_1003_),
    .A_N(_0791_));
 sg13g2_o21ai_1 _4646_ (.B1(_1458_),
    .Y(_1459_),
    .A1(_1003_),
    .A2(_1008_));
 sg13g2_nor4_2 _4647_ (.A(_1064_),
    .B(_1097_),
    .C(_1459_),
    .Y(_1460_),
    .D(_1088_));
 sg13g2_mux2_1 _4648_ (.A0(_1085_),
    .A1(_1082_),
    .S(_1079_),
    .X(_1461_));
 sg13g2_mux2_1 _4649_ (.A0(_1078_),
    .A1(_1461_),
    .S(_1076_),
    .X(_1462_));
 sg13g2_nand2_1 _4650_ (.Y(_1463_),
    .A(_1064_),
    .B(net45));
 sg13g2_nor2_1 _4651_ (.A(_1065_),
    .B(net45),
    .Y(_1464_));
 sg13g2_a22oi_1 _4652_ (.Y(_1465_),
    .B1(_1464_),
    .B2(_1459_),
    .A2(_1398_),
    .A1(_1065_));
 sg13g2_o21ai_1 _4653_ (.B1(_1465_),
    .Y(_1466_),
    .A1(_1462_),
    .A2(_1463_));
 sg13g2_o21ai_1 _4654_ (.B1(_1067_),
    .Y(_1467_),
    .A1(_1460_),
    .A2(_1466_));
 sg13g2_o21ai_1 _4655_ (.B1(_1149_),
    .Y(_1468_),
    .A1(net4),
    .A2(net43));
 sg13g2_or2_1 _4656_ (.X(_1469_),
    .B(_1468_),
    .A(_1250_));
 sg13g2_nor2_1 _4657_ (.A(_1149_),
    .B(_1245_),
    .Y(_1470_));
 sg13g2_o21ai_1 _4658_ (.B1(_1470_),
    .Y(_1471_),
    .A1(_1169_),
    .A2(_1244_));
 sg13g2_nand3_1 _4659_ (.B(_1469_),
    .C(_1471_),
    .A(_1068_),
    .Y(_1472_));
 sg13g2_nand3b_1 _4660_ (.B(_1467_),
    .C(_1472_),
    .Y(_1473_),
    .A_N(_0859_));
 sg13g2_a21oi_1 _4661_ (.A1(_1457_),
    .A2(_1473_),
    .Y(_0057_),
    .B1(_1193_));
 sg13g2_o21ai_1 _4662_ (.B1(_1068_),
    .Y(_1474_),
    .A1(_1460_),
    .A2(_1466_));
 sg13g2_nand3_1 _4663_ (.B(_1469_),
    .C(_1471_),
    .A(_1067_),
    .Y(_1475_));
 sg13g2_nand3b_1 _4664_ (.B(_1426_),
    .C(_1428_),
    .Y(_1476_),
    .A_N(net50));
 sg13g2_nand3_1 _4665_ (.B(_1448_),
    .C(_1455_),
    .A(net50),
    .Y(_1477_));
 sg13g2_nand4_1 _4666_ (.B(_1475_),
    .C(_1476_),
    .A(_1474_),
    .Y(_1478_),
    .D(_1477_));
 sg13g2_and2_1 _4667_ (.A(net155),
    .B(_1478_),
    .X(_0058_));
 sg13g2_and2_1 _4668_ (.A(\g.g_y[3].g_x[1].t.out_sc ),
    .B(net150),
    .X(_0056_));
 sg13g2_and2_1 _4669_ (.A(\g.g_y[3].g_x[0].t.out_sc ),
    .B(net150),
    .X(_0055_));
 sg13g2_buf_1 _4670_ (.A(net165),
    .X(_1479_));
 sg13g2_and2_1 _4671_ (.A(_1221_),
    .B(net149),
    .X(_0054_));
 sg13g2_nand2_1 _4672_ (.Y(_1480_),
    .A(_1258_),
    .B(_1254_));
 sg13g2_nor2b_1 _4673_ (.A(net48),
    .B_N(_0943_),
    .Y(_1481_));
 sg13g2_o21ai_1 _4674_ (.B1(_1481_),
    .Y(_1482_),
    .A1(_0930_),
    .A2(_1480_));
 sg13g2_o21ai_1 _4675_ (.B1(net48),
    .Y(_1483_),
    .A1(_1258_),
    .A2(_1254_));
 sg13g2_or2_1 _4676_ (.X(_1484_),
    .B(_1483_),
    .A(_0947_));
 sg13g2_nand3_1 _4677_ (.B(_1482_),
    .C(_1484_),
    .A(_0932_),
    .Y(_1485_));
 sg13g2_buf_1 _4678_ (.A(\g.g_y[1].g_x[6].t.r_v ),
    .X(_1486_));
 sg13g2_mux2_1 _4679_ (.A0(_2356_),
    .A1(_2358_),
    .S(_2359_),
    .X(_1487_));
 sg13g2_nand2b_1 _4680_ (.Y(_1488_),
    .B(_0933_),
    .A_N(_0936_));
 sg13g2_inv_1 _4681_ (.Y(_1489_),
    .A(_0937_));
 sg13g2_a21oi_1 _4682_ (.A1(_1489_),
    .A2(_0932_),
    .Y(_1490_),
    .B1(_1486_));
 sg13g2_a22oi_1 _4683_ (.Y(_1491_),
    .B1(_1488_),
    .B2(_1490_),
    .A2(_1487_),
    .A1(_1486_));
 sg13g2_buf_2 _4684_ (.A(\g.g_y[1].g_x[7].t.r_h ),
    .X(_1492_));
 sg13g2_mux2_1 _4685_ (.A0(\g.g_y[1].g_x[7].t.out_sc ),
    .A1(\g.g_y[1].g_x[7].t.r_gnl ),
    .S(_2472_),
    .X(_1493_));
 sg13g2_nand2b_1 _4686_ (.Y(_1494_),
    .B(_1492_),
    .A_N(_2475_));
 sg13g2_o21ai_1 _4687_ (.B1(_1494_),
    .Y(_1495_),
    .A1(_1492_),
    .A2(_1493_));
 sg13g2_buf_1 _4688_ (.A(_1495_),
    .X(_1496_));
 sg13g2_buf_2 _4689_ (.A(\g.g_y[1].g_x[5].t.r_h ),
    .X(_1497_));
 sg13g2_inv_1 _4690_ (.Y(_1498_),
    .A(_1497_));
 sg13g2_mux2_1 _4691_ (.A0(\g.g_y[1].g_x[5].t.out_sc ),
    .A1(\g.g_y[1].g_x[5].t.r_gnl ),
    .S(_2549_),
    .X(_1499_));
 sg13g2_buf_1 _4692_ (.A(_1499_),
    .X(_1500_));
 sg13g2_or2_1 _4693_ (.X(_1501_),
    .B(_1497_),
    .A(_2548_));
 sg13g2_o21ai_1 _4694_ (.B1(_1501_),
    .Y(_1502_),
    .A1(_1498_),
    .A2(_1500_));
 sg13g2_buf_2 _4695_ (.A(\g.g_y[1].g_x[6].t.r_h ),
    .X(_1503_));
 sg13g2_mux2_1 _4696_ (.A0(_1496_),
    .A1(_1502_),
    .S(_1503_),
    .X(_1504_));
 sg13g2_buf_1 _4697_ (.A(\g.g_y[1].g_x[6].t.r_d ),
    .X(_1505_));
 sg13g2_buf_1 _4698_ (.A(_1486_),
    .X(_1506_));
 sg13g2_nor2b_1 _4699_ (.A(net35),
    .B_N(net24),
    .Y(_1507_));
 sg13g2_o21ai_1 _4700_ (.B1(_1507_),
    .Y(_1508_),
    .A1(_1491_),
    .A2(_1504_));
 sg13g2_mux2_1 _4701_ (.A0(_2548_),
    .A1(_1500_),
    .S(_1497_),
    .X(_1509_));
 sg13g2_mux2_1 _4702_ (.A0(_1493_),
    .A1(_2475_),
    .S(_1492_),
    .X(_1510_));
 sg13g2_mux2_1 _4703_ (.A0(_1509_),
    .A1(_1510_),
    .S(_1503_),
    .X(_1511_));
 sg13g2_nor2_1 _4704_ (.A(net24),
    .B(net35),
    .Y(_1512_));
 sg13g2_nor2b_1 _4705_ (.A(net24),
    .B_N(net35),
    .Y(_1513_));
 sg13g2_buf_1 _4706_ (.A(\g.g_y[1].g_x[6].t.out_sc ),
    .X(_1514_));
 sg13g2_and3_1 _4707_ (.X(_1515_),
    .A(net24),
    .B(net35),
    .C(_1514_));
 sg13g2_a221oi_1 _4708_ (.B2(_1487_),
    .C1(_1515_),
    .B1(_1513_),
    .A1(_1511_),
    .Y(_1516_),
    .A2(_1512_));
 sg13g2_nand3_1 _4709_ (.B(_1508_),
    .C(_1516_),
    .A(_0933_),
    .Y(_1517_));
 sg13g2_nand3_1 _4710_ (.B(_1485_),
    .C(_1517_),
    .A(_0934_),
    .Y(_1518_));
 sg13g2_inv_1 _4711_ (.Y(_1519_),
    .A(\g.g_y[2].g_x[7].t.r_d ));
 sg13g2_nand2b_1 _4712_ (.Y(_1520_),
    .B(_0619_),
    .A_N(\g.g_y[3].g_x[7].t.r_ghl ));
 sg13g2_o21ai_1 _4713_ (.B1(_1520_),
    .Y(_1521_),
    .A1(_0619_),
    .A2(_0618_));
 sg13g2_buf_1 _4714_ (.A(_1521_),
    .X(_1522_));
 sg13g2_mux2_1 _4715_ (.A0(_1198_),
    .A1(_1522_),
    .S(_1195_),
    .X(_1523_));
 sg13g2_nor3_1 _4716_ (.A(_1519_),
    .B(_1523_),
    .C(_1210_),
    .Y(_1524_));
 sg13g2_nor2_1 _4717_ (.A(net41),
    .B(_1221_),
    .Y(_1525_));
 sg13g2_or3_1 _4718_ (.A(_1204_),
    .B(net40),
    .C(_1525_),
    .X(_1526_));
 sg13g2_or2_1 _4719_ (.X(_1527_),
    .B(_1206_),
    .A(_1204_));
 sg13g2_nor2b_1 _4720_ (.A(net40),
    .B_N(_1208_),
    .Y(_1528_));
 sg13g2_a221oi_1 _4721_ (.B2(_1528_),
    .C1(net41),
    .B1(_1527_),
    .A1(net40),
    .Y(_1529_),
    .A2(_1215_));
 sg13g2_nand2b_1 _4722_ (.Y(_1530_),
    .B(_0952_),
    .A_N(_0618_));
 sg13g2_and2_1 _4723_ (.A(_1194_),
    .B(_1520_),
    .X(_1531_));
 sg13g2_a221oi_1 _4724_ (.B2(_1531_),
    .C1(_1519_),
    .B1(_1530_),
    .A1(_1195_),
    .Y(_1532_),
    .A2(_1219_));
 sg13g2_nand2_1 _4725_ (.Y(_1533_),
    .A(_1203_),
    .B(net40));
 sg13g2_or3_1 _4726_ (.A(_1529_),
    .B(_1532_),
    .C(_1533_),
    .X(_1534_));
 sg13g2_o21ai_1 _4727_ (.B1(_1534_),
    .Y(_1535_),
    .A1(_1524_),
    .A2(_1526_));
 sg13g2_o21ai_1 _4728_ (.B1(_1294_),
    .Y(_1536_),
    .A1(net38),
    .A2(_1314_));
 sg13g2_or2_1 _4729_ (.X(_1537_),
    .B(_1536_),
    .A(_1349_));
 sg13g2_nand2_1 _4730_ (.Y(_1538_),
    .A(net38),
    .B(_1314_));
 sg13g2_nor2_1 _4731_ (.A(net38),
    .B(\g.g_y[2].g_x[5].t.out_sc ),
    .Y(_1539_));
 sg13g2_nor2_1 _4732_ (.A(_1294_),
    .B(_1539_),
    .Y(_1540_));
 sg13g2_o21ai_1 _4733_ (.B1(_1540_),
    .Y(_1541_),
    .A1(_1288_),
    .A2(_1538_));
 sg13g2_a21oi_1 _4734_ (.A1(_1537_),
    .A2(_1541_),
    .Y(_1542_),
    .B1(_1203_));
 sg13g2_inv_1 _4735_ (.Y(_1543_),
    .A(_0934_));
 sg13g2_o21ai_1 _4736_ (.B1(_1543_),
    .Y(_1544_),
    .A1(_1535_),
    .A2(_1542_));
 sg13g2_a21oi_1 _4737_ (.A1(_1518_),
    .A2(_1544_),
    .Y(_0052_),
    .B1(net135));
 sg13g2_or2_1 _4738_ (.X(_1545_),
    .B(_1210_),
    .A(_1523_));
 sg13g2_nand2_1 _4739_ (.Y(_1546_),
    .A(_1195_),
    .B(_1219_));
 sg13g2_o21ai_1 _4740_ (.B1(_1546_),
    .Y(_1547_),
    .A1(_1195_),
    .A2(_1522_));
 sg13g2_mux4_1 _4741_ (.S0(net40),
    .A0(_1221_),
    .A1(_1215_),
    .A2(_1545_),
    .A3(_1547_),
    .S1(_1196_),
    .X(_1548_));
 sg13g2_nand2b_1 _4742_ (.Y(_1549_),
    .B(_1204_),
    .A_N(_1548_));
 sg13g2_nand3_1 _4743_ (.B(_1537_),
    .C(_1541_),
    .A(_1203_),
    .Y(_1550_));
 sg13g2_nand3_1 _4744_ (.B(_1482_),
    .C(_1484_),
    .A(_0933_),
    .Y(_1551_));
 sg13g2_nand3_1 _4745_ (.B(_1508_),
    .C(_1516_),
    .A(_0932_),
    .Y(_1552_));
 sg13g2_and3_1 _4746_ (.X(_1553_),
    .A(_1550_),
    .B(_1551_),
    .C(_1552_));
 sg13g2_a21oi_1 _4747_ (.A1(_1549_),
    .A2(_1553_),
    .Y(_0053_),
    .B1(_1193_));
 sg13g2_and2_1 _4748_ (.A(\g.g_y[2].g_x[6].t.out_sc ),
    .B(net149),
    .X(_0051_));
 sg13g2_and2_1 _4749_ (.A(\g.g_y[2].g_x[5].t.out_sc ),
    .B(net149),
    .X(_0050_));
 sg13g2_inv_1 _4750_ (.Y(_1554_),
    .A(_0993_));
 sg13g2_nor2_1 _4751_ (.A(net46),
    .B(_1020_),
    .Y(_1555_));
 sg13g2_a221oi_1 _4752_ (.B2(_1056_),
    .C1(_1326_),
    .B1(_1555_),
    .A1(net46),
    .Y(_1556_),
    .A2(_1405_));
 sg13g2_buf_2 _4753_ (.A(\g.g_y[1].g_x[4].t.r_v ),
    .X(_1557_));
 sg13g2_inv_2 _4754_ (.Y(_1558_),
    .A(_1557_));
 sg13g2_mux2_1 _4755_ (.A0(_2567_),
    .A1(_2645_),
    .S(_2646_),
    .X(_1559_));
 sg13g2_buf_1 _4756_ (.A(_1559_),
    .X(_1560_));
 sg13g2_mux2_1 _4757_ (.A0(_2548_),
    .A1(_1500_),
    .S(_1498_),
    .X(_1561_));
 sg13g2_mux2_1 _4758_ (.A0(\g.g_y[1].g_x[3].t.out_sc ),
    .A1(\g.g_y[1].g_x[3].t.r_gnl ),
    .S(_2707_),
    .X(_1562_));
 sg13g2_buf_1 _4759_ (.A(_1562_),
    .X(_1563_));
 sg13g2_buf_1 _4760_ (.A(\g.g_y[1].g_x[3].t.r_h ),
    .X(_1564_));
 sg13g2_mux2_1 _4761_ (.A0(_2706_),
    .A1(_1563_),
    .S(_1564_),
    .X(_1565_));
 sg13g2_buf_2 _4762_ (.A(\g.g_y[1].g_x[4].t.r_h ),
    .X(_1566_));
 sg13g2_inv_1 _4763_ (.Y(_1567_),
    .A(_1566_));
 sg13g2_mux2_1 _4764_ (.A0(_1561_),
    .A1(_1565_),
    .S(_1567_),
    .X(_1568_));
 sg13g2_buf_1 _4765_ (.A(\g.g_y[1].g_x[4].t.r_d ),
    .X(_1569_));
 sg13g2_inv_2 _4766_ (.Y(_1570_),
    .A(net34));
 sg13g2_mux2_1 _4767_ (.A0(_1560_),
    .A1(_1568_),
    .S(_1570_),
    .X(_1571_));
 sg13g2_mux2_1 _4768_ (.A0(_0992_),
    .A1(_0995_),
    .S(_1326_),
    .X(_1572_));
 sg13g2_buf_2 _4769_ (.A(_1572_),
    .X(_1573_));
 sg13g2_mux2_1 _4770_ (.A0(_1560_),
    .A1(_1573_),
    .S(_1558_),
    .X(_1574_));
 sg13g2_mux2_1 _4771_ (.A0(_1561_),
    .A1(_1565_),
    .S(_1566_),
    .X(_1575_));
 sg13g2_nand3_1 _4772_ (.B(_1574_),
    .C(_1575_),
    .A(_1570_),
    .Y(_1576_));
 sg13g2_buf_1 _4773_ (.A(\g.g_y[1].g_x[4].t.out_sc ),
    .X(_1577_));
 sg13g2_inv_1 _4774_ (.Y(_1578_),
    .A(_1577_));
 sg13g2_a21oi_1 _4775_ (.A1(net34),
    .A2(_1578_),
    .Y(_1579_),
    .B1(_1558_));
 sg13g2_a221oi_1 _4776_ (.B2(_1579_),
    .C1(_0996_),
    .B1(_1576_),
    .A1(_1558_),
    .Y(_1580_),
    .A2(_1571_));
 sg13g2_or3_1 _4777_ (.A(_1554_),
    .B(_1556_),
    .C(_1580_),
    .X(_1581_));
 sg13g2_nor2_1 _4778_ (.A(_1382_),
    .B(_1362_),
    .Y(_1582_));
 sg13g2_o21ai_1 _4779_ (.B1(_1582_),
    .Y(_1583_),
    .A1(_1381_),
    .A2(_1385_));
 sg13g2_mux2_1 _4780_ (.A0(_2706_),
    .A1(_2708_),
    .S(_2709_),
    .X(_1584_));
 sg13g2_mux2_1 _4781_ (.A0(_1357_),
    .A1(_1584_),
    .S(_1378_),
    .X(_1585_));
 sg13g2_nor2_1 _4782_ (.A(_1364_),
    .B(_1362_),
    .Y(_1586_));
 sg13g2_nor2_1 _4783_ (.A(_1382_),
    .B(net36),
    .Y(_1587_));
 sg13g2_nor2_1 _4784_ (.A(_1367_),
    .B(_1368_),
    .Y(_1588_));
 sg13g2_nor4_1 _4785_ (.A(_1364_),
    .B(net36),
    .C(_1588_),
    .D(_1371_),
    .Y(_1589_));
 sg13g2_a221oi_1 _4786_ (.B2(\g.g_y[2].g_x[3].t.out_sc ),
    .C1(_1589_),
    .B1(_1587_),
    .A1(_1585_),
    .Y(_1590_),
    .A2(_1586_));
 sg13g2_nand3_1 _4787_ (.B(_1583_),
    .C(_1590_),
    .A(_1298_),
    .Y(_1591_));
 sg13g2_mux2_1 _4788_ (.A0(_0937_),
    .A1(_1206_),
    .S(_1204_),
    .X(_1592_));
 sg13g2_nand2_1 _4789_ (.Y(_1593_),
    .A(_1291_),
    .B(_1592_));
 sg13g2_nor2_1 _4790_ (.A(_1290_),
    .B(_1539_),
    .Y(_1594_));
 sg13g2_o21ai_1 _4791_ (.B1(_1594_),
    .Y(_1595_),
    .A1(_1288_),
    .A2(_1593_));
 sg13g2_o21ai_1 _4792_ (.B1(_1290_),
    .Y(_1596_),
    .A1(_1291_),
    .A2(_1592_));
 sg13g2_or2_1 _4793_ (.X(_1597_),
    .B(_1596_),
    .A(_1349_));
 sg13g2_buf_1 _4794_ (.A(_1597_),
    .X(_1598_));
 sg13g2_nand3_1 _4795_ (.B(_1595_),
    .C(_1598_),
    .A(_1295_),
    .Y(_1599_));
 sg13g2_nand3_1 _4796_ (.B(_1591_),
    .C(_1599_),
    .A(_1554_),
    .Y(_1600_));
 sg13g2_a21oi_1 _4797_ (.A1(_1581_),
    .A2(_1600_),
    .Y(_0048_),
    .B1(net135));
 sg13g2_a21oi_1 _4798_ (.A1(_1583_),
    .A2(_1590_),
    .Y(_1601_),
    .B1(_1298_));
 sg13g2_a21oi_1 _4799_ (.A1(_1595_),
    .A2(_1598_),
    .Y(_1602_),
    .B1(_1295_));
 sg13g2_or2_1 _4800_ (.X(_1603_),
    .B(_1602_),
    .A(_1601_));
 sg13g2_a22oi_1 _4801_ (.Y(_1604_),
    .B1(_1555_),
    .B2(_1056_),
    .A2(_1405_),
    .A1(net46));
 sg13g2_a221oi_1 _4802_ (.B2(_1579_),
    .C1(_1326_),
    .B1(_1576_),
    .A1(_1558_),
    .Y(_1605_),
    .A2(_1571_));
 sg13g2_a21oi_1 _4803_ (.A1(_1326_),
    .A2(_1604_),
    .Y(_1606_),
    .B1(_1605_));
 sg13g2_buf_1 _4804_ (.A(net154),
    .X(_1607_));
 sg13g2_a21oi_1 _4805_ (.A1(_1603_),
    .A2(_1606_),
    .Y(_0049_),
    .B1(net134));
 sg13g2_and2_1 _4806_ (.A(\g.g_y[2].g_x[4].t.out_sc ),
    .B(net149),
    .X(_0047_));
 sg13g2_and2_1 _4807_ (.A(\g.g_y[2].g_x[3].t.out_sc ),
    .B(net165),
    .X(_0046_));
 sg13g2_nand2_1 _4808_ (.Y(_1608_),
    .A(_1097_),
    .B(_1078_));
 sg13g2_a21oi_1 _4809_ (.A1(_1063_),
    .A2(_1090_),
    .Y(_1609_),
    .B1(net44));
 sg13g2_o21ai_1 _4810_ (.B1(_1609_),
    .Y(_1610_),
    .A1(_1074_),
    .A2(_1608_));
 sg13g2_o21ai_1 _4811_ (.B1(net44),
    .Y(_1611_),
    .A1(_1097_),
    .A2(_1078_));
 sg13g2_or2_1 _4812_ (.X(_1612_),
    .B(_1611_),
    .A(_1095_));
 sg13g2_nand3_1 _4813_ (.B(_1610_),
    .C(_1612_),
    .A(_1079_),
    .Y(_1613_));
 sg13g2_buf_2 _4814_ (.A(\g.g_y[1].g_x[2].t.r_v ),
    .X(_1614_));
 sg13g2_mux2_1 _4815_ (.A0(_1085_),
    .A1(_1082_),
    .S(_1080_),
    .X(_1615_));
 sg13g2_buf_1 _4816_ (.A(_1615_),
    .X(_1616_));
 sg13g2_or2_1 _4817_ (.X(_1617_),
    .B(_2789_),
    .A(_0204_));
 sg13g2_nor2_1 _4818_ (.A(_2695_),
    .B(_2787_),
    .Y(_1618_));
 sg13g2_nor2_1 _4819_ (.A(_1614_),
    .B(_1618_),
    .Y(_1619_));
 sg13g2_buf_2 _4820_ (.A(\g.g_y[1].g_x[2].t.r_d ),
    .X(_1620_));
 sg13g2_inv_2 _4821_ (.Y(_1621_),
    .A(_1620_));
 sg13g2_a221oi_1 _4822_ (.B2(_1619_),
    .C1(_1621_),
    .B1(_1617_),
    .A1(_1614_),
    .Y(_1622_),
    .A2(_1616_));
 sg13g2_buf_2 _4823_ (.A(\g.g_y[1].g_x[2].t.r_h ),
    .X(_1623_));
 sg13g2_inv_1 _4824_ (.Y(_1624_),
    .A(_1564_));
 sg13g2_mux2_1 _4825_ (.A0(_2706_),
    .A1(_1563_),
    .S(_1624_),
    .X(_1625_));
 sg13g2_buf_2 _4826_ (.A(_1625_),
    .X(_1626_));
 sg13g2_buf_1 _4827_ (.A(\g.g_y[1].g_x[1].t.r_h ),
    .X(_1627_));
 sg13g2_inv_1 _4828_ (.Y(_1628_),
    .A(net33));
 sg13g2_mux2_1 _4829_ (.A0(\g.g_y[1].g_x[1].t.out_sc ),
    .A1(\g.g_y[1].g_x[1].t.r_gnl ),
    .S(_0230_),
    .X(_1629_));
 sg13g2_buf_1 _4830_ (.A(_1629_),
    .X(_1630_));
 sg13g2_or2_1 _4831_ (.X(_1631_),
    .B(_1630_),
    .A(_1628_));
 sg13g2_buf_1 _4832_ (.A(_1631_),
    .X(_1632_));
 sg13g2_nor2_1 _4833_ (.A(_0233_),
    .B(net33),
    .Y(_1633_));
 sg13g2_nor2_1 _4834_ (.A(_1623_),
    .B(_1633_),
    .Y(_1634_));
 sg13g2_a221oi_1 _4835_ (.B2(_1634_),
    .C1(_1620_),
    .B1(_1632_),
    .A1(_1623_),
    .Y(_1635_),
    .A2(_1626_));
 sg13g2_or3_1 _4836_ (.A(_1614_),
    .B(_1622_),
    .C(_1635_),
    .X(_1636_));
 sg13g2_inv_1 _4837_ (.Y(_1637_),
    .A(_1623_));
 sg13g2_nor2_1 _4838_ (.A(_1637_),
    .B(_1633_),
    .Y(_1638_));
 sg13g2_a22oi_1 _4839_ (.Y(_1639_),
    .B1(_1632_),
    .B2(_1638_),
    .A2(_1626_),
    .A1(_1637_));
 sg13g2_buf_1 _4840_ (.A(_1639_),
    .X(_1640_));
 sg13g2_mux2_1 _4841_ (.A0(_2695_),
    .A1(_2789_),
    .S(_2787_),
    .X(_1641_));
 sg13g2_nand2_1 _4842_ (.Y(_1642_),
    .A(_1621_),
    .B(_1641_));
 sg13g2_buf_2 _4843_ (.A(\g.g_y[1].g_x[2].t.out_sc ),
    .X(_1643_));
 sg13g2_inv_1 _4844_ (.Y(_1644_),
    .A(_1643_));
 sg13g2_inv_2 _4845_ (.Y(_1645_),
    .A(_1614_));
 sg13g2_a21oi_1 _4846_ (.A1(_1620_),
    .A2(_1644_),
    .Y(_1646_),
    .B1(_1645_));
 sg13g2_o21ai_1 _4847_ (.B1(_1646_),
    .Y(_1647_),
    .A1(_1640_),
    .A2(_1642_));
 sg13g2_nand3_1 _4848_ (.B(_1636_),
    .C(_1647_),
    .A(_1080_),
    .Y(_1648_));
 sg13g2_nand3_1 _4849_ (.B(_1613_),
    .C(_1648_),
    .A(_1081_),
    .Y(_1649_));
 sg13g2_nand2b_1 _4850_ (.Y(_1650_),
    .B(_0858_),
    .A_N(_0862_));
 sg13g2_o21ai_1 _4851_ (.B1(_1650_),
    .Y(_1651_),
    .A1(_0858_),
    .A2(_0861_));
 sg13g2_mux2_1 _4852_ (.A0(_1651_),
    .A1(_1453_),
    .S(_1446_),
    .X(_1652_));
 sg13g2_nor2_1 _4853_ (.A(_1438_),
    .B(_1442_),
    .Y(_1653_));
 sg13g2_o21ai_1 _4854_ (.B1(_1653_),
    .Y(_1654_),
    .A1(_1440_),
    .A2(_1652_));
 sg13g2_mux2_1 _4855_ (.A0(_0861_),
    .A1(_0862_),
    .S(net50),
    .X(_1655_));
 sg13g2_mux2_1 _4856_ (.A0(_1443_),
    .A1(_1655_),
    .S(_1446_),
    .X(_1656_));
 sg13g2_nor2_1 _4857_ (.A(_1432_),
    .B(_1442_),
    .Y(_1657_));
 sg13g2_nor2_1 _4858_ (.A(_1438_),
    .B(_1441_),
    .Y(_1658_));
 sg13g2_and4_1 _4859_ (.A(_1438_),
    .B(_1442_),
    .C(_1431_),
    .D(_1434_),
    .X(_1659_));
 sg13g2_a221oi_1 _4860_ (.B2(\g.g_y[2].g_x[1].t.out_sc ),
    .C1(_1659_),
    .B1(_1658_),
    .A1(_1656_),
    .Y(_1660_),
    .A2(_1657_));
 sg13g2_nand3_1 _4861_ (.B(_1654_),
    .C(_1660_),
    .A(_1367_),
    .Y(_1661_));
 sg13g2_o21ai_1 _4862_ (.B1(_1586_),
    .Y(_1662_),
    .A1(_1381_),
    .A2(_1385_));
 sg13g2_nand2_1 _4863_ (.Y(_1663_),
    .A(_1585_),
    .B(_1582_));
 sg13g2_nor2_1 _4864_ (.A(_1364_),
    .B(_1361_),
    .Y(_1664_));
 sg13g2_a22oi_1 _4865_ (.Y(_1665_),
    .B1(_1587_),
    .B2(_1366_),
    .A2(_1664_),
    .A1(\g.g_y[2].g_x[3].t.out_sc ));
 sg13g2_nand4_1 _4866_ (.B(_1662_),
    .C(_1663_),
    .A(\g.g_y[2].g_x[2].t.r_h ),
    .Y(_1666_),
    .D(_1665_));
 sg13g2_nand3b_1 _4867_ (.B(_1661_),
    .C(_1666_),
    .Y(_1667_),
    .A_N(_1081_));
 sg13g2_a21oi_1 _4868_ (.A1(_1649_),
    .A2(_1667_),
    .Y(_0044_),
    .B1(net134));
 sg13g2_nand3_1 _4869_ (.B(_1654_),
    .C(_1660_),
    .A(\g.g_y[2].g_x[2].t.r_h ),
    .Y(_1668_));
 sg13g2_nand4_1 _4870_ (.B(_1662_),
    .C(_1663_),
    .A(_1367_),
    .Y(_1669_),
    .D(_1665_));
 sg13g2_and2_1 _4871_ (.A(_1668_),
    .B(_1669_),
    .X(_1670_));
 sg13g2_nand3_1 _4872_ (.B(_1636_),
    .C(_1647_),
    .A(_1079_),
    .Y(_1671_));
 sg13g2_nand3_1 _4873_ (.B(_1610_),
    .C(_1612_),
    .A(_1080_),
    .Y(_1672_));
 sg13g2_and2_1 _4874_ (.A(_1671_),
    .B(_1672_),
    .X(_1673_));
 sg13g2_a21oi_1 _4875_ (.A1(_1670_),
    .A2(_1673_),
    .Y(_0045_),
    .B1(net134));
 sg13g2_and2_1 _4876_ (.A(\g.g_y[2].g_x[2].t.out_sc ),
    .B(net149),
    .X(_0043_));
 sg13g2_inv_1 _4877_ (.Y(_1674_),
    .A(\g.g_y[2].g_x[1].t.out_sc ));
 sg13g2_nor2_1 _4878_ (.A(_1674_),
    .B(net138),
    .Y(_0042_));
 sg13g2_o21ai_1 _4879_ (.B1(_1238_),
    .Y(_1675_),
    .A1(_0567_),
    .A2(_0571_));
 sg13g2_nor2b_1 _4880_ (.A(net42),
    .B_N(_1174_),
    .Y(_1676_));
 sg13g2_o21ai_1 _4881_ (.B1(_1676_),
    .Y(_1677_),
    .A1(_1173_),
    .A2(_1675_));
 sg13g2_nand2_1 _4882_ (.Y(_1678_),
    .A(net43),
    .B(_1675_));
 sg13g2_nand3_1 _4883_ (.B(_1156_),
    .C(_1678_),
    .A(net42),
    .Y(_1679_));
 sg13g2_nand3_1 _4884_ (.B(_1677_),
    .C(_1679_),
    .A(_1157_),
    .Y(_1680_));
 sg13g2_buf_1 _4885_ (.A(\g.g_y[1].g_x[0].t.r_v ),
    .X(_1681_));
 sg13g2_inv_1 _4886_ (.Y(_1682_),
    .A(_1681_));
 sg13g2_inv_1 _4887_ (.Y(_1683_),
    .A(\g.g_y[1].g_x[0].t.r_d ));
 sg13g2_buf_1 _4888_ (.A(\g.g_y[1].g_x[0].t.r_h ),
    .X(_1684_));
 sg13g2_inv_1 _4889_ (.Y(_1685_),
    .A(_1684_));
 sg13g2_nor2b_1 _4890_ (.A(net33),
    .B_N(_1684_),
    .Y(_1686_));
 sg13g2_and3_1 _4891_ (.X(_1687_),
    .A(_0233_),
    .B(net33),
    .C(_1684_));
 sg13g2_a221oi_1 _4892_ (.B2(_1686_),
    .C1(_1687_),
    .B1(_1630_),
    .A1(net2),
    .Y(_1688_),
    .A2(_1685_));
 sg13g2_and2_1 _4893_ (.A(_1683_),
    .B(_1688_),
    .X(_1689_));
 sg13g2_nand2b_1 _4894_ (.Y(_1690_),
    .B(net33),
    .A_N(_0233_));
 sg13g2_o21ai_1 _4895_ (.B1(_1690_),
    .Y(_1691_),
    .A1(net33),
    .A2(_1630_));
 sg13g2_nand2_1 _4896_ (.Y(_1692_),
    .A(net2),
    .B(_1684_));
 sg13g2_o21ai_1 _4897_ (.B1(_1692_),
    .Y(_1693_),
    .A1(_1684_),
    .A2(_1691_));
 sg13g2_buf_1 _4898_ (.A(\g.g_y[1].g_x[0].t.r_d ),
    .X(_1694_));
 sg13g2_or2_1 _4899_ (.X(_1695_),
    .B(_2394_),
    .A(_2400_));
 sg13g2_buf_1 _4900_ (.A(_1695_),
    .X(_1696_));
 sg13g2_o21ai_1 _4901_ (.B1(_1696_),
    .Y(_1697_),
    .A1(_2395_),
    .A2(_2393_));
 sg13g2_nor3_1 _4902_ (.A(_1682_),
    .B(net32),
    .C(_1697_),
    .Y(_1698_));
 sg13g2_nor2_1 _4903_ (.A(_1681_),
    .B(_1683_),
    .Y(_1699_));
 sg13g2_nor3_1 _4904_ (.A(_1682_),
    .B(_1683_),
    .C(\g.g_y[1].g_x[0].t.out_sc ),
    .Y(_1700_));
 sg13g2_a21o_1 _4905_ (.A2(_1699_),
    .A1(_1697_),
    .B1(_1700_),
    .X(_1701_));
 sg13g2_a221oi_1 _4906_ (.B2(_1698_),
    .C1(_1701_),
    .B1(_1693_),
    .A1(_1682_),
    .Y(_1702_),
    .A2(_1689_));
 sg13g2_nand2b_1 _4907_ (.Y(_1703_),
    .B(_1158_),
    .A_N(_1702_));
 sg13g2_nand3_1 _4908_ (.B(_1680_),
    .C(_1703_),
    .A(_1159_),
    .Y(_1704_));
 sg13g2_o21ai_1 _4909_ (.B1(_1657_),
    .Y(_1705_),
    .A1(_1440_),
    .A2(_1652_));
 sg13g2_nor3_1 _4910_ (.A(_1432_),
    .B(_1441_),
    .C(_1674_),
    .Y(_1706_));
 sg13g2_a221oi_1 _4911_ (.B2(_1437_),
    .C1(_1706_),
    .B1(_1658_),
    .A1(_1656_),
    .Y(_1707_),
    .A2(_1653_));
 sg13g2_a21oi_1 _4912_ (.A1(_1705_),
    .A2(_1707_),
    .Y(_1708_),
    .B1(_1213_));
 sg13g2_nor2b_1 _4913_ (.A(_1199_),
    .B_N(net3),
    .Y(_1709_));
 sg13g2_inv_1 _4914_ (.Y(_1710_),
    .A(_1159_));
 sg13g2_o21ai_1 _4915_ (.B1(_1710_),
    .Y(_1711_),
    .A1(_1708_),
    .A2(_1709_));
 sg13g2_a21oi_1 _4916_ (.A1(_1704_),
    .A2(_1711_),
    .Y(_0040_),
    .B1(net134));
 sg13g2_a21oi_1 _4917_ (.A1(_1705_),
    .A2(_1707_),
    .Y(_1712_),
    .B1(_1199_));
 sg13g2_a21o_1 _4918_ (.A2(net3),
    .A1(_1199_),
    .B1(_1712_),
    .X(_1713_));
 sg13g2_a21oi_1 _4919_ (.A1(_1677_),
    .A2(_1679_),
    .Y(_1714_),
    .B1(_1157_));
 sg13g2_a21o_1 _4920_ (.A2(_1702_),
    .A1(_1157_),
    .B1(_1714_),
    .X(_1715_));
 sg13g2_a21oi_1 _4921_ (.A1(_1713_),
    .A2(_1715_),
    .Y(_0041_),
    .B1(net134));
 sg13g2_and2_1 _4922_ (.A(\g.g_y[2].g_x[0].t.out_sc ),
    .B(net149),
    .X(_0039_));
 sg13g2_mux2_1 _4923_ (.A0(_1194_),
    .A1(_1519_),
    .S(_1522_),
    .X(_1716_));
 sg13g2_mux2_1 _4924_ (.A0(net41),
    .A1(_1195_),
    .S(_1522_),
    .X(_1717_));
 sg13g2_o21ai_1 _4925_ (.B1(_1717_),
    .Y(_1718_),
    .A1(_1221_),
    .A2(_1716_));
 sg13g2_nor2_1 _4926_ (.A(_1195_),
    .B(net41),
    .Y(_1719_));
 sg13g2_nor2_1 _4927_ (.A(_1216_),
    .B(_1196_),
    .Y(_1720_));
 sg13g2_a21oi_1 _4928_ (.A1(_1194_),
    .A2(_1209_),
    .Y(_1721_),
    .B1(_1215_));
 sg13g2_nand2_1 _4929_ (.Y(_1722_),
    .A(net40),
    .B(_1519_));
 sg13g2_a221oi_1 _4930_ (.B2(_1208_),
    .C1(_1722_),
    .B1(_1527_),
    .A1(_1194_),
    .Y(_1723_),
    .A2(_1202_));
 sg13g2_a221oi_1 _4931_ (.B2(_1721_),
    .C1(_1723_),
    .B1(_1720_),
    .A1(_1217_),
    .Y(_1724_),
    .A2(_1719_));
 sg13g2_a21oi_1 _4932_ (.A1(_1718_),
    .A2(_1724_),
    .Y(_1725_),
    .B1(_2503_));
 sg13g2_nor3_1 _4933_ (.A(net81),
    .B(_2510_),
    .C(_2512_),
    .Y(_1726_));
 sg13g2_nor2_1 _4934_ (.A(_2491_),
    .B(_2519_),
    .Y(_1727_));
 sg13g2_or3_1 _4935_ (.A(_2471_),
    .B(_2483_),
    .C(_1727_),
    .X(_1728_));
 sg13g2_a221oi_1 _4936_ (.B2(_2517_),
    .C1(_2486_),
    .B1(_2516_),
    .A1(_2511_),
    .Y(_1729_),
    .A2(_2514_));
 sg13g2_a21oi_1 _4937_ (.A1(_2508_),
    .A2(_2485_),
    .Y(_1730_),
    .B1(_2482_));
 sg13g2_a221oi_1 _4938_ (.B2(_1730_),
    .C1(_2519_),
    .B1(_2507_),
    .A1(_2482_),
    .Y(_1731_),
    .A2(_2504_));
 sg13g2_or4_1 _4939_ (.A(_2471_),
    .B(_2482_),
    .C(_1729_),
    .D(_1731_),
    .X(_1732_));
 sg13g2_o21ai_1 _4940_ (.B1(_1732_),
    .Y(_1733_),
    .A1(_1726_),
    .A2(_1728_));
 sg13g2_o21ai_1 _4941_ (.B1(_2472_),
    .Y(_1734_),
    .A1(_1725_),
    .A2(_1733_));
 sg13g2_and2_1 _4942_ (.A(_1503_),
    .B(net35),
    .X(_1735_));
 sg13g2_o21ai_1 _4943_ (.B1(_1735_),
    .Y(_1736_),
    .A1(_1491_),
    .A2(_1504_));
 sg13g2_mux2_1 _4944_ (.A0(_0937_),
    .A1(_0936_),
    .S(_0933_),
    .X(_1737_));
 sg13g2_buf_1 _4945_ (.A(_1737_),
    .X(_1738_));
 sg13g2_mux2_1 _4946_ (.A0(_1487_),
    .A1(_1738_),
    .S(_1486_),
    .X(_1739_));
 sg13g2_nor2b_1 _4947_ (.A(_1503_),
    .B_N(\g.g_y[1].g_x[6].t.r_d ),
    .Y(_1740_));
 sg13g2_nor2_1 _4948_ (.A(_1503_),
    .B(_1505_),
    .Y(_1741_));
 sg13g2_inv_1 _4949_ (.Y(_1742_),
    .A(_1514_));
 sg13g2_nand2b_1 _4950_ (.Y(_1743_),
    .B(_1503_),
    .A_N(\g.g_y[1].g_x[6].t.r_d ));
 sg13g2_nor2_1 _4951_ (.A(_1742_),
    .B(_1743_),
    .Y(_1744_));
 sg13g2_a221oi_1 _4952_ (.B2(_1509_),
    .C1(_1744_),
    .B1(_1741_),
    .A1(_1739_),
    .Y(_1745_),
    .A2(_1740_));
 sg13g2_nand3b_1 _4953_ (.B(_1736_),
    .C(_1745_),
    .Y(_1746_),
    .A_N(_1492_));
 sg13g2_nand2b_1 _4954_ (.Y(_1747_),
    .B(_1158_),
    .A_N(_1161_));
 sg13g2_nand2b_1 _4955_ (.Y(_1748_),
    .B(_1157_),
    .A_N(_1162_));
 sg13g2_and3_1 _4956_ (.X(_1749_),
    .A(_1682_),
    .B(_1694_),
    .C(_1748_));
 sg13g2_and3_1 _4957_ (.X(_1750_),
    .A(_1681_),
    .B(net32),
    .C(_1696_));
 sg13g2_or2_1 _4958_ (.X(_1751_),
    .B(_2393_),
    .A(_2395_));
 sg13g2_buf_1 _4959_ (.A(_1751_),
    .X(_1752_));
 sg13g2_a22oi_1 _4960_ (.Y(_1753_),
    .B1(_1750_),
    .B2(_1752_),
    .A2(_1749_),
    .A1(_1747_));
 sg13g2_nor2_1 _4961_ (.A(net32),
    .B(\g.g_y[1].g_x[0].t.out_sc ),
    .Y(_1754_));
 sg13g2_nor2_1 _4962_ (.A(_1684_),
    .B(_1754_),
    .Y(_1755_));
 sg13g2_o21ai_1 _4963_ (.B1(_1755_),
    .Y(_1756_),
    .A1(_1691_),
    .A2(_1753_));
 sg13g2_mux2_1 _4964_ (.A0(_1162_),
    .A1(_1161_),
    .S(_1158_),
    .X(_1757_));
 sg13g2_and2_1 _4965_ (.A(_1682_),
    .B(_1696_),
    .X(_1758_));
 sg13g2_a221oi_1 _4966_ (.B2(_1752_),
    .C1(_1683_),
    .B1(_1758_),
    .A1(_1681_),
    .Y(_1759_),
    .A2(_1757_));
 sg13g2_or3_1 _4967_ (.A(_1685_),
    .B(_1689_),
    .C(_1759_),
    .X(_1760_));
 sg13g2_nand3_1 _4968_ (.B(_1756_),
    .C(_1760_),
    .A(_1492_),
    .Y(_1761_));
 sg13g2_nand3b_1 _4969_ (.B(_1746_),
    .C(_1761_),
    .Y(_1762_),
    .A_N(_2472_));
 sg13g2_a21oi_1 _4970_ (.A1(_1734_),
    .A2(_1762_),
    .Y(_0037_),
    .B1(_1607_));
 sg13g2_nor3_1 _4971_ (.A(_2483_),
    .B(_1727_),
    .C(_1726_),
    .Y(_1763_));
 sg13g2_or2_1 _4972_ (.X(_1764_),
    .B(_1731_),
    .A(_1729_));
 sg13g2_buf_1 _4973_ (.A(_1764_),
    .X(_1765_));
 sg13g2_nor2_1 _4974_ (.A(_2482_),
    .B(_1765_),
    .Y(_1766_));
 sg13g2_or3_1 _4975_ (.A(_2503_),
    .B(_1763_),
    .C(_1766_),
    .X(_1767_));
 sg13g2_nand3b_1 _4976_ (.B(_1756_),
    .C(_1760_),
    .Y(_1768_),
    .A_N(_1492_));
 sg13g2_nand3_1 _4977_ (.B(_1736_),
    .C(_1745_),
    .A(_1492_),
    .Y(_1769_));
 sg13g2_nand3_1 _4978_ (.B(_1718_),
    .C(_1724_),
    .A(_2503_),
    .Y(_1770_));
 sg13g2_and3_1 _4979_ (.X(_1771_),
    .A(_1768_),
    .B(_1769_),
    .C(_1770_));
 sg13g2_a21oi_1 _4980_ (.A1(_1767_),
    .A2(_1771_),
    .Y(_0038_),
    .B1(_1607_));
 sg13g2_and2_1 _4981_ (.A(\g.g_y[1].g_x[7].t.out_sc ),
    .B(_1479_),
    .X(_0036_));
 sg13g2_nor2_1 _4982_ (.A(_1742_),
    .B(_2546_),
    .Y(_0035_));
 sg13g2_nor3_1 _4983_ (.A(_1279_),
    .B(_1288_),
    .C(_1301_),
    .Y(_1772_));
 sg13g2_mux2_1 _4984_ (.A0(_1314_),
    .A1(_1592_),
    .S(_1290_),
    .X(_1773_));
 sg13g2_nand2_1 _4985_ (.Y(_1774_),
    .A(net39),
    .B(_1310_));
 sg13g2_nand3b_1 _4986_ (.B(net38),
    .C(net39),
    .Y(_1775_),
    .A_N(_1282_));
 sg13g2_o21ai_1 _4987_ (.B1(_1775_),
    .Y(_1776_),
    .A1(_1773_),
    .A2(_1774_));
 sg13g2_o21ai_1 _4988_ (.B1(_2551_),
    .Y(_1777_),
    .A1(_1279_),
    .A2(_1302_));
 sg13g2_nor3_1 _4989_ (.A(_1772_),
    .B(_1776_),
    .C(_1777_),
    .Y(_1778_));
 sg13g2_inv_1 _4990_ (.Y(_1779_),
    .A(_2547_));
 sg13g2_nor3_1 _4991_ (.A(_2551_),
    .B(_1779_),
    .C(_2559_),
    .Y(_1780_));
 sg13g2_nand3_1 _4992_ (.B(_2580_),
    .C(_1780_),
    .A(_2576_),
    .Y(_1781_));
 sg13g2_o21ai_1 _4993_ (.B1(_1779_),
    .Y(_1782_),
    .A1(_2561_),
    .A2(_2572_));
 sg13g2_a21oi_1 _4994_ (.A1(_2547_),
    .A2(_2582_),
    .Y(_1783_),
    .B1(_2551_));
 sg13g2_and3_1 _4995_ (.X(_1784_),
    .A(_1781_),
    .B(_1782_),
    .C(_1783_));
 sg13g2_o21ai_1 _4996_ (.B1(_2549_),
    .Y(_1785_),
    .A1(_1778_),
    .A2(_1784_));
 sg13g2_nand3_1 _4997_ (.B(_1574_),
    .C(_1575_),
    .A(net34),
    .Y(_1786_));
 sg13g2_o21ai_1 _4998_ (.B1(_1566_),
    .Y(_1787_),
    .A1(net34),
    .A2(_1577_));
 sg13g2_inv_1 _4999_ (.Y(_1788_),
    .A(_1787_));
 sg13g2_nand2b_1 _5000_ (.Y(_1789_),
    .B(_1326_),
    .A_N(_0995_));
 sg13g2_nand2b_1 _5001_ (.Y(_1790_),
    .B(_0996_),
    .A_N(_0992_));
 sg13g2_and2_1 _5002_ (.A(_1557_),
    .B(_1790_),
    .X(_1791_));
 sg13g2_a221oi_1 _5003_ (.B2(_1791_),
    .C1(_1570_),
    .B1(_1789_),
    .A1(_1558_),
    .Y(_1792_),
    .A2(_1560_));
 sg13g2_o21ai_1 _5004_ (.B1(_1567_),
    .Y(_1793_),
    .A1(net34),
    .A2(_1565_));
 sg13g2_o21ai_1 _5005_ (.B1(_1498_),
    .Y(_1794_),
    .A1(_1792_),
    .A2(_1793_));
 sg13g2_a21o_1 _5006_ (.A2(_1788_),
    .A1(_1786_),
    .B1(_1794_),
    .X(_1795_));
 sg13g2_o21ai_1 _5007_ (.B1(_1740_),
    .Y(_1796_),
    .A1(_1491_),
    .A2(_1504_));
 sg13g2_nor2_1 _5008_ (.A(_1496_),
    .B(_1743_),
    .Y(_1797_));
 sg13g2_a221oi_1 _5009_ (.B2(_1514_),
    .C1(_1797_),
    .B1(_1741_),
    .A1(_1739_),
    .Y(_1798_),
    .A2(_1735_));
 sg13g2_nand3_1 _5010_ (.B(_1796_),
    .C(_1798_),
    .A(_1497_),
    .Y(_1799_));
 sg13g2_nand3b_1 _5011_ (.B(_1795_),
    .C(_1799_),
    .Y(_1800_),
    .A_N(_2549_));
 sg13g2_a21oi_1 _5012_ (.A1(_1785_),
    .A2(_1800_),
    .Y(_0033_),
    .B1(net134));
 sg13g2_mux2_1 _5013_ (.A0(_1303_),
    .A1(_1350_),
    .S(net39),
    .X(_1801_));
 sg13g2_nor2_1 _5014_ (.A(_1779_),
    .B(_2582_),
    .Y(_1802_));
 sg13g2_a221oi_1 _5015_ (.B2(_1802_),
    .C1(_2552_),
    .B1(_2581_),
    .A1(_1779_),
    .Y(_1803_),
    .A2(_2573_));
 sg13g2_a21oi_1 _5016_ (.A1(_2552_),
    .A2(_1801_),
    .Y(_1804_),
    .B1(_1803_));
 sg13g2_nor2_1 _5017_ (.A(_1792_),
    .B(_1793_),
    .Y(_1805_));
 sg13g2_a21o_1 _5018_ (.A2(_1788_),
    .A1(_1786_),
    .B1(_1805_),
    .X(_1806_));
 sg13g2_a21oi_1 _5019_ (.A1(_1796_),
    .A2(_1798_),
    .Y(_1807_),
    .B1(_1497_));
 sg13g2_a21o_1 _5020_ (.A2(_1806_),
    .A1(_1497_),
    .B1(_1807_),
    .X(_1808_));
 sg13g2_a21oi_1 _5021_ (.A1(_1804_),
    .A2(_1808_),
    .Y(_0034_),
    .B1(net134));
 sg13g2_and2_1 _5022_ (.A(\g.g_y[1].g_x[5].t.out_sc ),
    .B(net149),
    .X(_0032_));
 sg13g2_nor2_1 _5023_ (.A(_1578_),
    .B(net138),
    .Y(_0031_));
 sg13g2_and2_1 _5024_ (.A(_2714_),
    .B(_2727_),
    .X(_1809_));
 sg13g2_a22oi_1 _5025_ (.Y(_1810_),
    .B1(_0216_),
    .B2(_1809_),
    .A2(_0215_),
    .A1(_2724_));
 sg13g2_nor2_1 _5026_ (.A(_1363_),
    .B(_1373_),
    .Y(_1811_));
 sg13g2_and2_1 _5027_ (.A(_1378_),
    .B(_1387_),
    .X(_1812_));
 sg13g2_a221oi_1 _5028_ (.B2(_1812_),
    .C1(_2710_),
    .B1(_1416_),
    .A1(net37),
    .Y(_1813_),
    .A2(_1811_));
 sg13g2_a21o_1 _5029_ (.A2(_1810_),
    .A1(_2710_),
    .B1(_1813_),
    .X(_1814_));
 sg13g2_nand2_1 _5030_ (.Y(_1815_),
    .A(_2707_),
    .B(net166));
 sg13g2_inv_1 _5031_ (.Y(_1816_),
    .A(_2707_));
 sg13g2_nand2b_1 _5032_ (.Y(_1817_),
    .B(_1497_),
    .A_N(_2548_));
 sg13g2_o21ai_1 _5033_ (.B1(_1817_),
    .Y(_1818_),
    .A1(_1497_),
    .A2(_1500_));
 sg13g2_and2_1 _5034_ (.A(_1558_),
    .B(_1790_),
    .X(_1819_));
 sg13g2_a22oi_1 _5035_ (.Y(_1820_),
    .B1(_1789_),
    .B2(_1819_),
    .A2(_1560_),
    .A1(_1557_));
 sg13g2_nor4_1 _5036_ (.A(_1566_),
    .B(_1570_),
    .C(_1818_),
    .D(_1820_),
    .Y(_1821_));
 sg13g2_mux2_1 _5037_ (.A0(_1560_),
    .A1(_1573_),
    .S(_1557_),
    .X(_1822_));
 sg13g2_nand2_1 _5038_ (.Y(_1823_),
    .A(_1566_),
    .B(_1569_));
 sg13g2_nor2_1 _5039_ (.A(net34),
    .B(_1577_),
    .Y(_1824_));
 sg13g2_nor2_1 _5040_ (.A(_1567_),
    .B(net34),
    .Y(_1825_));
 sg13g2_a22oi_1 _5041_ (.Y(_1826_),
    .B1(_1825_),
    .B2(_1818_),
    .A2(_1824_),
    .A1(_1567_));
 sg13g2_o21ai_1 _5042_ (.B1(_1826_),
    .Y(_1827_),
    .A1(_1822_),
    .A2(_1823_));
 sg13g2_o21ai_1 _5043_ (.B1(_1564_),
    .Y(_1828_),
    .A1(_1821_),
    .A2(_1827_));
 sg13g2_nor2_1 _5044_ (.A(_1645_),
    .B(_1618_),
    .Y(_1829_));
 sg13g2_a22oi_1 _5045_ (.Y(_1830_),
    .B1(_1617_),
    .B2(_1829_),
    .A2(_1616_),
    .A1(_1645_));
 sg13g2_nor2_1 _5046_ (.A(_1637_),
    .B(_1621_),
    .Y(_1831_));
 sg13g2_o21ai_1 _5047_ (.B1(_1831_),
    .Y(_1832_),
    .A1(_1640_),
    .A2(_1830_));
 sg13g2_mux2_1 _5048_ (.A0(_1616_),
    .A1(_1641_),
    .S(_1645_),
    .X(_1833_));
 sg13g2_buf_1 _5049_ (.A(_1833_),
    .X(_1834_));
 sg13g2_nor2_1 _5050_ (.A(_1623_),
    .B(_1621_),
    .Y(_1835_));
 sg13g2_nor2_1 _5051_ (.A(_1637_),
    .B(_1620_),
    .Y(_1836_));
 sg13g2_mux2_1 _5052_ (.A0(_0233_),
    .A1(_1630_),
    .S(net33),
    .X(_1837_));
 sg13g2_nor2_1 _5053_ (.A(_1623_),
    .B(_1620_),
    .Y(_1838_));
 sg13g2_and2_1 _5054_ (.A(_1837_),
    .B(_1838_),
    .X(_1839_));
 sg13g2_a221oi_1 _5055_ (.B2(_1643_),
    .C1(_1839_),
    .B1(_1836_),
    .A1(_1834_),
    .Y(_1840_),
    .A2(_1835_));
 sg13g2_nand3_1 _5056_ (.B(_1832_),
    .C(_1840_),
    .A(_1624_),
    .Y(_1841_));
 sg13g2_nand4_1 _5057_ (.B(net166),
    .C(_1828_),
    .A(_1816_),
    .Y(_1842_),
    .D(_1841_));
 sg13g2_o21ai_1 _5058_ (.B1(_1842_),
    .Y(_0028_),
    .A1(_1814_),
    .A2(_1815_));
 sg13g2_a21oi_1 _5059_ (.A1(_1832_),
    .A2(_1840_),
    .Y(_1843_),
    .B1(_1624_));
 sg13g2_nor3_1 _5060_ (.A(_1564_),
    .B(_1821_),
    .C(_1827_),
    .Y(_1844_));
 sg13g2_or2_1 _5061_ (.X(_1845_),
    .B(_1844_),
    .A(_1843_));
 sg13g2_a221oi_1 _5062_ (.B2(_1812_),
    .C1(_2709_),
    .B1(_1416_),
    .A1(net37),
    .Y(_1846_),
    .A2(_1811_));
 sg13g2_a21oi_1 _5063_ (.A1(_2709_),
    .A2(_1810_),
    .Y(_1847_),
    .B1(_1846_));
 sg13g2_a21oi_1 _5064_ (.A1(_1845_),
    .A2(_1847_),
    .Y(_0029_),
    .B1(net134));
 sg13g2_and2_1 _5065_ (.A(\g.g_y[1].g_x[3].t.out_sc ),
    .B(net149),
    .X(_0027_));
 sg13g2_inv_1 _5066_ (.Y(_1848_),
    .A(net13));
 sg13g2_nand2_1 _5067_ (.Y(_1849_),
    .A(net166),
    .B(net11));
 sg13g2_a21oi_1 _5068_ (.A1(net12),
    .A2(_1848_),
    .Y(_0030_),
    .B1(_1849_));
 sg13g2_nor2_1 _5069_ (.A(_1644_),
    .B(net138),
    .Y(_0026_));
 sg13g2_mux2_1 _5070_ (.A0(_1453_),
    .A1(_1651_),
    .S(_1446_),
    .X(_1850_));
 sg13g2_a21oi_1 _5071_ (.A1(_1441_),
    .A2(_1850_),
    .Y(_1851_),
    .B1(_1450_));
 sg13g2_or3_1 _5072_ (.A(_1441_),
    .B(_1440_),
    .C(_1652_),
    .X(_1852_));
 sg13g2_nor2_1 _5073_ (.A(_1446_),
    .B(_1445_),
    .Y(_1853_));
 sg13g2_a221oi_1 _5074_ (.B2(_1853_),
    .C1(_1451_),
    .B1(_1852_),
    .A1(_1446_),
    .Y(_1854_),
    .A2(_1851_));
 sg13g2_nor2b_1 _5075_ (.A(\g.g_y[7].g_x[1].t.r_v ),
    .B_N(_2388_),
    .Y(_1855_));
 sg13g2_a21oi_1 _5076_ (.A1(_0228_),
    .A2(_0518_),
    .Y(_1856_),
    .B1(_1855_));
 sg13g2_a21oi_1 _5077_ (.A1(net70),
    .A2(_1856_),
    .Y(_1857_),
    .B1(\g.g_y[0].g_x[1].t.r_v ));
 sg13g2_nand2b_1 _5078_ (.Y(_1858_),
    .B(_1857_),
    .A_N(_0254_));
 sg13g2_a21oi_1 _5079_ (.A1(_0249_),
    .A2(net70),
    .Y(_1859_),
    .B1(_0255_));
 sg13g2_o21ai_1 _5080_ (.B1(_1859_),
    .Y(_1860_),
    .A1(_0248_),
    .A2(_1856_));
 sg13g2_nand3_1 _5081_ (.B(_1858_),
    .C(_1860_),
    .A(_1451_),
    .Y(_1861_));
 sg13g2_nand3b_1 _5082_ (.B(_1861_),
    .C(_0230_),
    .Y(_1862_),
    .A_N(_1854_));
 sg13g2_o21ai_1 _5083_ (.B1(_1835_),
    .Y(_1863_),
    .A1(_1640_),
    .A2(_1830_));
 sg13g2_nand2_1 _5084_ (.Y(_1864_),
    .A(_1834_),
    .B(_1831_));
 sg13g2_a22oi_1 _5085_ (.Y(_1865_),
    .B1(_1836_),
    .B2(_1626_),
    .A2(_1838_),
    .A1(_1643_));
 sg13g2_nand4_1 _5086_ (.B(_1863_),
    .C(_1864_),
    .A(net33),
    .Y(_1866_),
    .D(_1865_));
 sg13g2_o21ai_1 _5087_ (.B1(_1685_),
    .Y(_1867_),
    .A1(net2),
    .A2(net32));
 sg13g2_or2_1 _5088_ (.X(_1868_),
    .B(_1867_),
    .A(_1759_));
 sg13g2_inv_1 _5089_ (.Y(_1869_),
    .A(net2));
 sg13g2_nor2_1 _5090_ (.A(_1685_),
    .B(_1754_),
    .Y(_1870_));
 sg13g2_o21ai_1 _5091_ (.B1(_1870_),
    .Y(_1871_),
    .A1(_1869_),
    .A2(_1753_));
 sg13g2_nand3_1 _5092_ (.B(_1868_),
    .C(_1871_),
    .A(_1628_),
    .Y(_1872_));
 sg13g2_nand3b_1 _5093_ (.B(_1866_),
    .C(_1872_),
    .Y(_1873_),
    .A_N(_0230_));
 sg13g2_buf_1 _5094_ (.A(net156),
    .X(_1874_));
 sg13g2_a21oi_1 _5095_ (.A1(_1862_),
    .A2(_1873_),
    .Y(_0023_),
    .B1(net131));
 sg13g2_nand4_1 _5096_ (.B(_1863_),
    .C(_1864_),
    .A(_1628_),
    .Y(_1875_),
    .D(_1865_));
 sg13g2_a22oi_1 _5097_ (.Y(_1876_),
    .B1(_1852_),
    .B2(_1853_),
    .A2(_1851_),
    .A1(_1446_));
 sg13g2_and2_1 _5098_ (.A(_1868_),
    .B(_1871_),
    .X(_1877_));
 sg13g2_and3_1 _5099_ (.X(_1878_),
    .A(_0229_),
    .B(_1858_),
    .C(_1860_));
 sg13g2_a221oi_1 _5100_ (.B2(_1627_),
    .C1(_1878_),
    .B1(_1877_),
    .A1(_1451_),
    .Y(_1879_),
    .A2(_1876_));
 sg13g2_a21oi_1 _5101_ (.A1(_1875_),
    .A2(_1879_),
    .Y(_0024_),
    .B1(net131));
 sg13g2_and2_1 _5102_ (.A(\g.g_y[1].g_x[1].t.out_sc ),
    .B(_1479_),
    .X(_0022_));
 sg13g2_inv_1 _5103_ (.Y(_1880_),
    .A(net12));
 sg13g2_a21oi_1 _5104_ (.A1(_1880_),
    .A2(net13),
    .Y(_0025_),
    .B1(_1849_));
 sg13g2_inv_1 _5105_ (.Y(_1881_),
    .A(\g.g_y[1].g_x[0].t.out_sc ));
 sg13g2_nor2_1 _5106_ (.A(_1881_),
    .B(net138),
    .Y(_0021_));
 sg13g2_nor2_1 _5107_ (.A(_2502_),
    .B(_2546_),
    .Y(_0020_));
 sg13g2_a21oi_1 _5108_ (.A1(net89),
    .A2(_2544_),
    .Y(_1882_),
    .B1(_2363_));
 sg13g2_a221oi_1 _5109_ (.B2(_1882_),
    .C1(_2359_),
    .B1(_0362_),
    .A1(_2363_),
    .Y(_1883_),
    .A2(_0360_));
 sg13g2_nand2_1 _5110_ (.Y(_1884_),
    .A(_1506_),
    .B(_1502_));
 sg13g2_nand3b_1 _5111_ (.B(_1510_),
    .C(_1738_),
    .Y(_1885_),
    .A_N(_1506_));
 sg13g2_nand3_1 _5112_ (.B(_1884_),
    .C(_1885_),
    .A(_1741_),
    .Y(_1886_));
 sg13g2_a221oi_1 _5113_ (.B2(_1738_),
    .C1(_1743_),
    .B1(_1509_),
    .A1(net24),
    .Y(_1887_),
    .A2(_1496_));
 sg13g2_nand2_1 _5114_ (.Y(_1888_),
    .A(_1503_),
    .B(_1486_));
 sg13g2_nor3_1 _5115_ (.A(net35),
    .B(_1496_),
    .C(_1888_),
    .Y(_1889_));
 sg13g2_and3_1 _5116_ (.X(_1890_),
    .A(net24),
    .B(net35),
    .C(_1738_));
 sg13g2_nand2_1 _5117_ (.Y(_1891_),
    .A(net35),
    .B(_1514_));
 sg13g2_o21ai_1 _5118_ (.B1(_2359_),
    .Y(_1892_),
    .A1(net24),
    .A2(_1891_));
 sg13g2_nor4_1 _5119_ (.A(_1887_),
    .B(_1889_),
    .C(_1890_),
    .D(_1892_),
    .Y(_1893_));
 sg13g2_nand2_1 _5120_ (.Y(_1894_),
    .A(_1886_),
    .B(_1893_));
 sg13g2_nand3b_1 _5121_ (.B(_1894_),
    .C(_2357_),
    .Y(_1895_),
    .A_N(_1883_));
 sg13g2_nor2_1 _5122_ (.A(_2461_),
    .B(_2511_),
    .Y(_1896_));
 sg13g2_nor3_1 _5123_ (.A(_2460_),
    .B(_2578_),
    .C(_2560_),
    .Y(_1897_));
 sg13g2_and2_1 _5124_ (.A(_2576_),
    .B(_2580_),
    .X(_1898_));
 sg13g2_a22oi_1 _5125_ (.Y(_1899_),
    .B1(_1897_),
    .B2(_1898_),
    .A2(_1896_),
    .A1(_1765_));
 sg13g2_nor3_1 _5126_ (.A(_2461_),
    .B(_2481_),
    .C(_2519_),
    .Y(_1900_));
 sg13g2_nor3_1 _5127_ (.A(_2460_),
    .B(_2569_),
    .C(_2560_),
    .Y(_1901_));
 sg13g2_mux2_1 _5128_ (.A0(_2553_),
    .A1(_2574_),
    .S(_1779_),
    .X(_1902_));
 sg13g2_inv_1 _5129_ (.Y(_1903_),
    .A(_1902_));
 sg13g2_nor4_1 _5130_ (.A(_2461_),
    .B(_2481_),
    .C(_2491_),
    .D(net81),
    .Y(_1904_));
 sg13g2_nand2_1 _5131_ (.Y(_1905_),
    .A(_2461_),
    .B(_2560_));
 sg13g2_a221oi_1 _5132_ (.B2(_2570_),
    .C1(_1905_),
    .B1(_2566_),
    .A1(net80),
    .Y(_1906_),
    .A2(\g.g_y[0].g_x[5].t.out_sc ));
 sg13g2_or2_1 _5133_ (.X(_1907_),
    .B(_1906_),
    .A(_1904_));
 sg13g2_a221oi_1 _5134_ (.B2(_1903_),
    .C1(_1907_),
    .B1(_1901_),
    .A1(_2513_),
    .Y(_1908_),
    .A2(_1900_));
 sg13g2_nand3b_1 _5135_ (.B(_1899_),
    .C(_1908_),
    .Y(_1909_),
    .A_N(_2357_));
 sg13g2_a21oi_1 _5136_ (.A1(_1895_),
    .A2(_1909_),
    .Y(_0018_),
    .B1(_1874_));
 sg13g2_a22oi_1 _5137_ (.Y(_1910_),
    .B1(_2507_),
    .B2(_1730_),
    .A2(_2504_),
    .A1(_2482_));
 sg13g2_mux4_1 _5138_ (.S0(_2481_),
    .A0(_2502_),
    .A1(_2470_),
    .A2(_2513_),
    .A3(_1910_),
    .S1(net81),
    .X(_1911_));
 sg13g2_nand3_1 _5139_ (.B(_2576_),
    .C(_2580_),
    .A(_2559_),
    .Y(_1912_));
 sg13g2_nor2_1 _5140_ (.A(\g.g_y[0].g_x[5].t.out_sc ),
    .B(_2559_),
    .Y(_1913_));
 sg13g2_nor2_1 _5141_ (.A(_2578_),
    .B(_1913_),
    .Y(_1914_));
 sg13g2_a221oi_1 _5142_ (.B2(_1914_),
    .C1(_2461_),
    .B1(_1912_),
    .A1(_2578_),
    .Y(_1915_),
    .A2(_2573_));
 sg13g2_a21oi_1 _5143_ (.A1(_2461_),
    .A2(_1911_),
    .Y(_1916_),
    .B1(_1915_));
 sg13g2_a22oi_1 _5144_ (.Y(_1917_),
    .B1(_0362_),
    .B2(_1882_),
    .A2(_0360_),
    .A1(_2363_));
 sg13g2_o21ai_1 _5145_ (.B1(_2360_),
    .Y(_1918_),
    .A1(net24),
    .A2(_1891_));
 sg13g2_nor4_1 _5146_ (.A(_1887_),
    .B(_1889_),
    .C(_1890_),
    .D(_1918_),
    .Y(_1919_));
 sg13g2_a22oi_1 _5147_ (.Y(_1920_),
    .B1(_1886_),
    .B2(_1919_),
    .A2(_1917_),
    .A1(_2359_));
 sg13g2_a21oi_1 _5148_ (.A1(_1916_),
    .A2(_1920_),
    .Y(_0019_),
    .B1(_1874_));
 sg13g2_buf_1 _5149_ (.A(net165),
    .X(_1921_));
 sg13g2_and2_1 _5150_ (.A(\g.g_y[0].g_x[6].t.out_sc ),
    .B(_1921_),
    .X(_0017_));
 sg13g2_and2_1 _5151_ (.A(\g.g_y[0].g_x[5].t.out_sc ),
    .B(net168),
    .X(_0016_));
 sg13g2_inv_1 _5152_ (.Y(_1922_),
    .A(_2564_));
 sg13g2_nand3_1 _5153_ (.B(_1561_),
    .C(_1573_),
    .A(_1558_),
    .Y(_1923_));
 sg13g2_or2_1 _5154_ (.X(_1924_),
    .B(_1564_),
    .A(_2706_));
 sg13g2_o21ai_1 _5155_ (.B1(_1924_),
    .Y(_1925_),
    .A1(_1624_),
    .A2(_1563_));
 sg13g2_a21oi_1 _5156_ (.A1(_1557_),
    .A2(_1925_),
    .Y(_1926_),
    .B1(_1566_));
 sg13g2_nand3_1 _5157_ (.B(_1923_),
    .C(_1926_),
    .A(_1570_),
    .Y(_1927_));
 sg13g2_mux2_1 _5158_ (.A0(_1577_),
    .A1(_1573_),
    .S(_1557_),
    .X(_1928_));
 sg13g2_nand2_1 _5159_ (.Y(_1929_),
    .A(_1566_),
    .B(_1570_));
 sg13g2_a21oi_1 _5160_ (.A1(_1557_),
    .A2(_1818_),
    .Y(_1930_),
    .B1(_1929_));
 sg13g2_or2_1 _5161_ (.X(_1931_),
    .B(_1563_),
    .A(_1624_));
 sg13g2_and2_1 _5162_ (.A(_1924_),
    .B(_1790_),
    .X(_1932_));
 sg13g2_nand4_1 _5163_ (.B(_1931_),
    .C(_1789_),
    .A(_1558_),
    .Y(_1933_),
    .D(_1932_));
 sg13g2_a22oi_1 _5164_ (.Y(_1934_),
    .B1(_1930_),
    .B2(_1933_),
    .A2(_1928_),
    .A1(net34));
 sg13g2_and3_1 _5165_ (.X(_1935_),
    .A(_2646_),
    .B(_1927_),
    .C(_1934_));
 sg13g2_and2_1 _5166_ (.A(net78),
    .B(_0430_),
    .X(_1936_));
 sg13g2_a221oi_1 _5167_ (.B2(_1936_),
    .C1(_2646_),
    .B1(_0463_),
    .A1(_2644_),
    .Y(_1937_),
    .A2(_0461_));
 sg13g2_or3_1 _5168_ (.A(_1922_),
    .B(_1935_),
    .C(_1937_),
    .X(_1938_));
 sg13g2_nor2_1 _5169_ (.A(net80),
    .B(_1913_),
    .Y(_1939_));
 sg13g2_a221oi_1 _5170_ (.B2(_1939_),
    .C1(_2563_),
    .B1(_1912_),
    .A1(net80),
    .Y(_1940_),
    .A2(_2573_));
 sg13g2_nand4_1 _5171_ (.B(net31),
    .C(_2701_),
    .A(net77),
    .Y(_1941_),
    .D(_2722_));
 sg13g2_nor2_1 _5172_ (.A(\g.g_y[0].g_x[3].t.out_sc ),
    .B(_2693_),
    .Y(_1942_));
 sg13g2_nor2b_1 _5173_ (.A(net77),
    .B_N(_2693_),
    .Y(_1943_));
 sg13g2_or2_1 _5174_ (.X(_1944_),
    .B(_2719_),
    .A(_2728_));
 sg13g2_inv_1 _5175_ (.Y(_1945_),
    .A(_2631_));
 sg13g2_a21oi_1 _5176_ (.A1(_1945_),
    .A2(_2728_),
    .Y(_1946_),
    .B1(_2714_));
 sg13g2_a22oi_1 _5177_ (.Y(_1947_),
    .B1(_1944_),
    .B2(_1946_),
    .A2(_2712_),
    .A1(_2714_));
 sg13g2_nor3_1 _5178_ (.A(net77),
    .B(_2693_),
    .C(_2701_),
    .Y(_1948_));
 sg13g2_a221oi_1 _5179_ (.B2(_1947_),
    .C1(_1948_),
    .B1(_1943_),
    .A1(net77),
    .Y(_1949_),
    .A2(_1942_));
 sg13g2_a21oi_1 _5180_ (.A1(_1941_),
    .A2(_1949_),
    .Y(_1950_),
    .B1(_2562_));
 sg13g2_or3_1 _5181_ (.A(_2564_),
    .B(_1940_),
    .C(_1950_),
    .X(_1951_));
 sg13g2_a21oi_1 _5182_ (.A1(_1938_),
    .A2(_1951_),
    .Y(_0014_),
    .B1(net131));
 sg13g2_a22oi_1 _5183_ (.Y(_1952_),
    .B1(_0463_),
    .B2(_1936_),
    .A2(_0461_),
    .A1(_2644_));
 sg13g2_a22oi_1 _5184_ (.Y(_1953_),
    .B1(_1912_),
    .B2(_1939_),
    .A2(_2573_),
    .A1(net80));
 sg13g2_a22oi_1 _5185_ (.Y(_1954_),
    .B1(_1953_),
    .B2(_2563_),
    .A2(_1952_),
    .A1(_2646_));
 sg13g2_and2_1 _5186_ (.A(_1927_),
    .B(_1934_),
    .X(_1955_));
 sg13g2_nand2_1 _5187_ (.Y(_1956_),
    .A(_1941_),
    .B(_1949_));
 sg13g2_a22oi_1 _5188_ (.Y(_1957_),
    .B1(_1956_),
    .B2(_2562_),
    .A2(_1955_),
    .A1(_2647_));
 sg13g2_a21oi_1 _5189_ (.A1(_1954_),
    .A2(_1957_),
    .Y(_0015_),
    .B1(net131));
 sg13g2_and2_1 _5190_ (.A(\g.g_y[0].g_x[4].t.out_sc ),
    .B(net148),
    .X(_0013_));
 sg13g2_and2_1 _5191_ (.A(\g.g_y[0].g_x[3].t.out_sc ),
    .B(net148),
    .X(_0012_));
 sg13g2_nand2_1 _5192_ (.Y(_1958_),
    .A(_1614_),
    .B(_1616_));
 sg13g2_a21oi_1 _5193_ (.A1(_1645_),
    .A2(_1643_),
    .Y(_1959_),
    .B1(_1621_));
 sg13g2_mux2_1 _5194_ (.A0(_1626_),
    .A1(_1837_),
    .S(_1623_),
    .X(_1960_));
 sg13g2_and2_1 _5195_ (.A(_1645_),
    .B(_1616_),
    .X(_1961_));
 sg13g2_a221oi_1 _5196_ (.B2(_1634_),
    .C1(_1645_),
    .B1(_1632_),
    .A1(_1623_),
    .Y(_1962_),
    .A2(_1626_));
 sg13g2_a21o_1 _5197_ (.A2(_1961_),
    .A1(_1960_),
    .B1(_1962_),
    .X(_1963_));
 sg13g2_a221oi_1 _5198_ (.B2(_1621_),
    .C1(_0204_),
    .B1(_1963_),
    .A1(_1958_),
    .Y(_1964_),
    .A2(_1959_));
 sg13g2_nor3_1 _5199_ (.A(_2792_),
    .B(net73),
    .C(_0472_),
    .Y(_1965_));
 sg13g2_nor3_1 _5200_ (.A(_2792_),
    .B(_2773_),
    .C(_0295_),
    .Y(_1966_));
 sg13g2_nor4_1 _5201_ (.A(_2793_),
    .B(_2772_),
    .C(_2780_),
    .D(_2786_),
    .Y(_1967_));
 sg13g2_nand2_1 _5202_ (.Y(_1968_),
    .A(_2772_),
    .B(_0227_));
 sg13g2_o21ai_1 _5203_ (.B1(_0204_),
    .Y(_1969_),
    .A1(_2793_),
    .A2(_1968_));
 sg13g2_nor4_1 _5204_ (.A(_1965_),
    .B(_1966_),
    .C(_1967_),
    .D(_1969_),
    .Y(_1970_));
 sg13g2_nor2_1 _5205_ (.A(_1964_),
    .B(_1970_),
    .Y(_1971_));
 sg13g2_nand2_1 _5206_ (.Y(_1972_),
    .A(_2696_),
    .B(net168));
 sg13g2_nand3_1 _5207_ (.B(_2717_),
    .C(_2722_),
    .A(net31),
    .Y(_1973_));
 sg13g2_nor2_1 _5208_ (.A(net77),
    .B(_1942_),
    .Y(_1974_));
 sg13g2_nor2_1 _5209_ (.A(net31),
    .B(_2702_),
    .Y(_1975_));
 sg13g2_a21oi_1 _5210_ (.A1(net31),
    .A2(_1947_),
    .Y(_1976_),
    .B1(_1975_));
 sg13g2_a221oi_1 _5211_ (.B2(net77),
    .C1(_0236_),
    .B1(_1976_),
    .A1(_1973_),
    .Y(_1977_),
    .A2(_1974_));
 sg13g2_or2_1 _5212_ (.X(_1978_),
    .B(net82),
    .A(_2400_));
 sg13g2_o21ai_1 _5213_ (.B1(_1978_),
    .Y(_1979_),
    .A1(_2515_),
    .A2(_2467_));
 sg13g2_a21o_1 _5214_ (.A2(_0518_),
    .A1(net71),
    .B1(_1855_),
    .X(_1980_));
 sg13g2_nor2_1 _5215_ (.A(_0255_),
    .B(_0241_),
    .Y(_1981_));
 sg13g2_nor2_1 _5216_ (.A(\g.g_y[0].g_x[1].t.r_v ),
    .B(_0241_),
    .Y(_1982_));
 sg13g2_mux2_1 _5217_ (.A0(_0233_),
    .A1(_0232_),
    .S(_1451_),
    .X(_1983_));
 sg13g2_a22oi_1 _5218_ (.Y(_1984_),
    .B1(_1982_),
    .B2(_1983_),
    .A2(_1981_),
    .A1(_1980_));
 sg13g2_or2_1 _5219_ (.X(_1985_),
    .B(_0240_),
    .A(\g.g_y[0].g_x[1].t.out_sc ));
 sg13g2_nand2_1 _5220_ (.Y(_1986_),
    .A(_0238_),
    .B(_1985_));
 sg13g2_inv_1 _5221_ (.Y(_1987_),
    .A(_1986_));
 sg13g2_o21ai_1 _5222_ (.B1(_1987_),
    .Y(_1988_),
    .A1(_1979_),
    .A2(_1984_));
 sg13g2_mux2_1 _5223_ (.A0(_1983_),
    .A1(_1980_),
    .S(_0255_),
    .X(_1989_));
 sg13g2_a21oi_1 _5224_ (.A1(_0241_),
    .A2(_1979_),
    .Y(_1990_),
    .B1(_0238_));
 sg13g2_o21ai_1 _5225_ (.B1(_1990_),
    .Y(_1991_),
    .A1(_0241_),
    .A2(_1989_));
 sg13g2_nand3_1 _5226_ (.B(_1988_),
    .C(_1991_),
    .A(_0236_),
    .Y(_1992_));
 sg13g2_nor2_1 _5227_ (.A(_2696_),
    .B(_2500_),
    .Y(_1993_));
 sg13g2_nand3b_1 _5228_ (.B(_1992_),
    .C(_1993_),
    .Y(_1994_),
    .A_N(_1977_));
 sg13g2_o21ai_1 _5229_ (.B1(_1994_),
    .Y(_0009_),
    .A1(_1971_),
    .A2(_1972_));
 sg13g2_or2_1 _5230_ (.X(_1995_),
    .B(_1830_),
    .A(_1640_));
 sg13g2_mux2_1 _5231_ (.A0(_1626_),
    .A1(_1837_),
    .S(_1637_),
    .X(_1996_));
 sg13g2_mux4_1 _5232_ (.S0(_1614_),
    .A0(_1643_),
    .A1(_1834_),
    .A2(_1995_),
    .A3(_1996_),
    .S1(_1621_),
    .X(_1997_));
 sg13g2_or2_1 _5233_ (.X(_1998_),
    .B(_2795_),
    .A(_2780_));
 sg13g2_mux4_1 _5234_ (.S0(_2773_),
    .A0(_0200_),
    .A1(_1998_),
    .A2(_0296_),
    .A3(_0472_),
    .S1(_2793_),
    .X(_1999_));
 sg13g2_mux2_1 _5235_ (.A0(_1997_),
    .A1(_1999_),
    .S(_2787_),
    .X(_2000_));
 sg13g2_a221oi_1 _5236_ (.B2(_2703_),
    .C1(_2699_),
    .B1(_1976_),
    .A1(_1973_),
    .Y(_2001_),
    .A2(_1974_));
 sg13g2_nand3_1 _5237_ (.B(_1988_),
    .C(_1991_),
    .A(_2699_),
    .Y(_2002_));
 sg13g2_nor2b_1 _5238_ (.A(_2001_),
    .B_N(_2002_),
    .Y(_2003_));
 sg13g2_a21oi_1 _5239_ (.A1(_2000_),
    .A2(_2003_),
    .Y(_0010_),
    .B1(net131));
 sg13g2_and2_1 _5240_ (.A(\g.g_y[0].g_x[2].t.out_sc ),
    .B(net148),
    .X(_0008_));
 sg13g2_a21oi_1 _5241_ (.A1(net12),
    .A2(net13),
    .Y(_0011_),
    .B1(_1849_));
 sg13g2_nor2_1 _5242_ (.A(_0249_),
    .B(_2499_),
    .Y(_0007_));
 sg13g2_inv_1 _5243_ (.Y(_2004_),
    .A(net9));
 sg13g2_a21oi_1 _5244_ (.A1(net10),
    .A2(_2004_),
    .Y(_0005_),
    .B1(net131));
 sg13g2_or2_1 _5245_ (.X(_2005_),
    .B(_2404_),
    .A(_2403_));
 sg13g2_o21ai_1 _5246_ (.B1(_2005_),
    .Y(_2006_),
    .A1(_2408_),
    .A2(_2411_));
 sg13g2_a21oi_1 _5247_ (.A1(net86),
    .A2(_2006_),
    .Y(_2007_),
    .B1(_2428_));
 sg13g2_nor2_1 _5248_ (.A(net86),
    .B(_2006_),
    .Y(_2008_));
 sg13g2_a21oi_1 _5249_ (.A1(_0553_),
    .A2(_2008_),
    .Y(_2009_),
    .B1(_0556_));
 sg13g2_mux2_1 _5250_ (.A0(_2007_),
    .A1(_2009_),
    .S(_2397_),
    .X(_2010_));
 sg13g2_o21ai_1 _5251_ (.B1(_1748_),
    .Y(_2011_),
    .A1(_1157_),
    .A2(_1161_));
 sg13g2_nor2_1 _5252_ (.A(net32),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_a221oi_1 _5253_ (.B2(_2012_),
    .C1(_1681_),
    .B1(_1693_),
    .A1(net32),
    .Y(_2013_),
    .A2(_1881_));
 sg13g2_nand2_1 _5254_ (.Y(_2014_),
    .A(_1694_),
    .B(_2011_));
 sg13g2_nand3b_1 _5255_ (.B(_2014_),
    .C(_1681_),
    .Y(_2015_),
    .A_N(_1689_));
 sg13g2_nand3b_1 _5256_ (.B(_2015_),
    .C(_2394_),
    .Y(_2016_),
    .A_N(_2013_));
 sg13g2_o21ai_1 _5257_ (.B1(_2016_),
    .Y(_2017_),
    .A1(_2394_),
    .A2(_2010_));
 sg13g2_nand2_1 _5258_ (.Y(_2018_),
    .A(_2391_),
    .B(net166));
 sg13g2_o21ai_1 _5259_ (.B1(_0242_),
    .Y(_2019_),
    .A1(_2699_),
    .A2(_2698_));
 sg13g2_o21ai_1 _5260_ (.B1(_1985_),
    .Y(_2020_),
    .A1(_2019_),
    .A2(_1984_));
 sg13g2_nand2_1 _5261_ (.Y(_2021_),
    .A(_0241_),
    .B(_2019_));
 sg13g2_o21ai_1 _5262_ (.B1(_2021_),
    .Y(_2022_),
    .A1(_0241_),
    .A2(_1989_));
 sg13g2_mux2_1 _5263_ (.A0(_2020_),
    .A1(_2022_),
    .S(_0238_),
    .X(_2023_));
 sg13g2_nor2_1 _5264_ (.A(_2465_),
    .B(net1),
    .Y(_2024_));
 sg13g2_or3_1 _5265_ (.A(_2391_),
    .B(_2499_),
    .C(_2024_),
    .X(_2025_));
 sg13g2_a21o_1 _5266_ (.A2(_2023_),
    .A1(net82),
    .B1(_2025_),
    .X(_2026_));
 sg13g2_o21ai_1 _5267_ (.B1(_2026_),
    .Y(_0001_),
    .A1(_2017_),
    .A2(_2018_));
 sg13g2_nand2b_1 _5268_ (.Y(_2027_),
    .B(_2015_),
    .A_N(_2013_));
 sg13g2_mux2_1 _5269_ (.A0(_2027_),
    .A1(_2010_),
    .S(_2394_),
    .X(_2028_));
 sg13g2_nand2_1 _5270_ (.Y(_2029_),
    .A(_2465_),
    .B(net1));
 sg13g2_o21ai_1 _5271_ (.B1(_2029_),
    .Y(_2030_),
    .A1(net82),
    .A2(_2023_));
 sg13g2_a21oi_1 _5272_ (.A1(_2028_),
    .A2(_2030_),
    .Y(_0002_),
    .B1(net131));
 sg13g2_inv_1 _5273_ (.Y(_2031_),
    .A(net10));
 sg13g2_a21oi_1 _5274_ (.A1(_2031_),
    .A2(net9),
    .Y(_0006_),
    .B1(net131));
 sg13g2_buf_1 _5275_ (.A(net156),
    .X(_2032_));
 sg13g2_a21oi_1 _5276_ (.A1(net10),
    .A2(net9),
    .Y(_0004_),
    .B1(net126));
 sg13g2_and2_1 _5277_ (.A(\g.g_y[0].g_x[0].t.out_sc ),
    .B(net148),
    .X(_0000_));
 sg13g2_o21ai_1 _5278_ (.B1(_1921_),
    .Y(_2033_),
    .A1(net12),
    .A2(net13));
 sg13g2_inv_1 _5279_ (.Y(_0003_),
    .A(_2033_));
 sg13g2_buf_1 _5280_ (.A(uio_in[0]),
    .X(_2034_));
 sg13g2_buf_1 _5281_ (.A(net167),
    .X(_2035_));
 sg13g2_nor2_1 _5282_ (.A(_2391_),
    .B(net163),
    .Y(_2036_));
 sg13g2_inv_1 _5283_ (.Y(_2037_),
    .A(net167));
 sg13g2_buf_1 _5284_ (.A(_2037_),
    .X(_2038_));
 sg13g2_and3_1 _5285_ (.X(_2039_),
    .A(_2391_),
    .B(net82),
    .C(net147));
 sg13g2_buf_1 _5286_ (.A(_2037_),
    .X(_2040_));
 sg13g2_o21ai_1 _5287_ (.B1(_0515_),
    .Y(_2041_),
    .A1(net8),
    .A2(_2040_));
 sg13g2_nand3_1 _5288_ (.B(net146),
    .C(_2024_),
    .A(_2391_),
    .Y(_2042_));
 sg13g2_nand2b_1 _5289_ (.Y(_2043_),
    .B(_2042_),
    .A_N(_2041_));
 sg13g2_a221oi_1 _5290_ (.B2(_2023_),
    .C1(_2043_),
    .B1(_2039_),
    .A1(_2017_),
    .Y(_0135_),
    .A2(_2036_));
 sg13g2_a221oi_1 _5291_ (.B2(_0247_),
    .C1(_0241_),
    .B1(_0253_),
    .A1(_0238_),
    .Y(_2044_),
    .A2(_0252_));
 sg13g2_nor2_1 _5292_ (.A(net70),
    .B(_1989_),
    .Y(_2045_));
 sg13g2_or2_1 _5293_ (.X(_2046_),
    .B(_2045_),
    .A(_2044_));
 sg13g2_buf_1 _5294_ (.A(net167),
    .X(_2047_));
 sg13g2_nand2_1 _5295_ (.Y(_2048_),
    .A(\g.g_y[0].g_x[0].t.out_sc ),
    .B(net162));
 sg13g2_o21ai_1 _5296_ (.B1(_2048_),
    .Y(_2049_),
    .A1(net163),
    .A2(_2046_));
 sg13g2_and2_1 _5297_ (.A(net155),
    .B(_2049_),
    .X(_0136_));
 sg13g2_nor2_1 _5298_ (.A(net162),
    .B(_1972_),
    .Y(_2050_));
 sg13g2_nand3b_1 _5299_ (.B(_1992_),
    .C(_2050_),
    .Y(_2051_),
    .A_N(_1977_));
 sg13g2_buf_1 _5300_ (.A(net167),
    .X(_2052_));
 sg13g2_nor3_1 _5301_ (.A(_2696_),
    .B(_2500_),
    .C(net161),
    .Y(_2053_));
 sg13g2_o21ai_1 _5302_ (.B1(_2053_),
    .Y(_2054_),
    .A1(_1964_),
    .A2(_1970_));
 sg13g2_buf_1 _5303_ (.A(net161),
    .X(_2055_));
 sg13g2_nand2_1 _5304_ (.Y(_2056_),
    .A(net145),
    .B(_0007_));
 sg13g2_nand3_1 _5305_ (.B(_2054_),
    .C(_2056_),
    .A(_2051_),
    .Y(_0137_));
 sg13g2_nor2_1 _5306_ (.A(_2694_),
    .B(_1947_),
    .Y(_2057_));
 sg13g2_a21oi_1 _5307_ (.A1(_2694_),
    .A2(_2704_),
    .Y(_2058_),
    .B1(_2057_));
 sg13g2_nand2_1 _5308_ (.Y(_2059_),
    .A(\g.g_y[0].g_x[2].t.out_sc ),
    .B(net162));
 sg13g2_o21ai_1 _5309_ (.B1(_2059_),
    .Y(_2060_),
    .A1(_2035_),
    .A2(_2058_));
 sg13g2_and2_1 _5310_ (.A(_2543_),
    .B(_2060_),
    .X(_0138_));
 sg13g2_buf_1 _5311_ (.A(net167),
    .X(_2061_));
 sg13g2_nor2_1 _5312_ (.A(_1922_),
    .B(net160),
    .Y(_2062_));
 sg13g2_o21ai_1 _5313_ (.B1(_2062_),
    .Y(_2063_),
    .A1(_1940_),
    .A2(_1950_));
 sg13g2_nor2_1 _5314_ (.A(_2564_),
    .B(net160),
    .Y(_2064_));
 sg13g2_o21ai_1 _5315_ (.B1(_2064_),
    .Y(_2065_),
    .A1(_1935_),
    .A2(_1937_));
 sg13g2_buf_8 _5316_ (.A(net167),
    .X(_2066_));
 sg13g2_nand2b_1 _5317_ (.Y(_2067_),
    .B(net159),
    .A_N(\g.g_y[0].g_x[3].t.out_sc ));
 sg13g2_and4_1 _5318_ (.A(net148),
    .B(_2063_),
    .C(_2065_),
    .D(_2067_),
    .X(_0139_));
 sg13g2_nand2_1 _5319_ (.Y(_2068_),
    .A(\g.g_y[0].g_x[4].t.out_sc ),
    .B(net145));
 sg13g2_buf_1 _5320_ (.A(net146),
    .X(_2069_));
 sg13g2_mux2_1 _5321_ (.A0(_2577_),
    .A1(_2571_),
    .S(net80),
    .X(_2070_));
 sg13g2_nand2_1 _5322_ (.Y(_2071_),
    .A(_2559_),
    .B(_2070_));
 sg13g2_o21ai_1 _5323_ (.B1(_2071_),
    .Y(_2072_),
    .A1(_2559_),
    .A2(_1903_));
 sg13g2_nand2_1 _5324_ (.Y(_2073_),
    .A(net125),
    .B(_2072_));
 sg13g2_a21oi_1 _5325_ (.A1(_2068_),
    .A2(_2073_),
    .Y(_0140_),
    .B1(net126));
 sg13g2_a21oi_1 _5326_ (.A1(_1886_),
    .A2(_1893_),
    .Y(_2074_),
    .B1(_2357_));
 sg13g2_nor2_1 _5327_ (.A(_2499_),
    .B(net160),
    .Y(_2075_));
 sg13g2_nand3b_1 _5328_ (.B(_2074_),
    .C(_2075_),
    .Y(_2076_),
    .A_N(_1883_));
 sg13g2_buf_1 _5329_ (.A(_2037_),
    .X(_2077_));
 sg13g2_and2_1 _5330_ (.A(_2357_),
    .B(_2498_),
    .X(_2078_));
 sg13g2_nand4_1 _5331_ (.B(_1899_),
    .C(_1908_),
    .A(net144),
    .Y(_2079_),
    .D(_2078_));
 sg13g2_nand2_1 _5332_ (.Y(_2080_),
    .A(net145),
    .B(_0016_));
 sg13g2_nand3_1 _5333_ (.B(_2079_),
    .C(_2080_),
    .A(_2076_),
    .Y(_0141_));
 sg13g2_buf_1 _5334_ (.A(net160),
    .X(_2081_));
 sg13g2_buf_1 _5335_ (.A(net167),
    .X(_2082_));
 sg13g2_mux2_1 _5336_ (.A0(_2518_),
    .A1(_1910_),
    .S(_2519_),
    .X(_2083_));
 sg13g2_nor2_1 _5337_ (.A(_2082_),
    .B(_2083_),
    .Y(_2084_));
 sg13g2_a21oi_1 _5338_ (.A1(\g.g_y[0].g_x[6].t.out_sc ),
    .A2(net143),
    .Y(_2085_),
    .B1(_2084_));
 sg13g2_nor2_1 _5339_ (.A(net139),
    .B(_2085_),
    .Y(_0142_));
 sg13g2_and2_1 _5340_ (.A(net32),
    .B(_1688_),
    .X(_2086_));
 sg13g2_a221oi_1 _5341_ (.B2(_1752_),
    .C1(net32),
    .B1(_1758_),
    .A1(_1681_),
    .Y(_2087_),
    .A2(_1757_));
 sg13g2_nor3_1 _5342_ (.A(net162),
    .B(_2086_),
    .C(_2087_),
    .Y(_2088_));
 sg13g2_a21oi_1 _5343_ (.A1(_2491_),
    .A2(net143),
    .Y(_2089_),
    .B1(_2088_));
 sg13g2_nor2_1 _5344_ (.A(net139),
    .B(_2089_),
    .Y(_0143_));
 sg13g2_nand2b_1 _5345_ (.Y(_2090_),
    .B(_1861_),
    .A_N(_1854_));
 sg13g2_nor2_1 _5346_ (.A(_0230_),
    .B(net163),
    .Y(_2091_));
 sg13g2_buf_1 _5347_ (.A(_2034_),
    .X(_2092_));
 sg13g2_nor2b_1 _5348_ (.A(net157),
    .B_N(_0230_),
    .Y(_2093_));
 sg13g2_nand2_1 _5349_ (.Y(_2094_),
    .A(_1866_),
    .B(_1872_));
 sg13g2_buf_1 _5350_ (.A(_2037_),
    .X(_2095_));
 sg13g2_buf_1 _5351_ (.A(net165),
    .X(_2096_));
 sg13g2_o21ai_1 _5352_ (.B1(net141),
    .Y(_2097_),
    .A1(\g.g_y[1].g_x[0].t.out_sc ),
    .A2(_2095_));
 sg13g2_a221oi_1 _5353_ (.B2(_2094_),
    .C1(_2097_),
    .B1(_2093_),
    .A1(_2090_),
    .Y(_0144_),
    .A2(_2091_));
 sg13g2_nand2_1 _5354_ (.Y(_2098_),
    .A(\g.g_y[1].g_x[1].t.out_sc ),
    .B(_2055_));
 sg13g2_mux2_1 _5355_ (.A0(_1834_),
    .A1(_1996_),
    .S(_1620_),
    .X(_2099_));
 sg13g2_nand2_1 _5356_ (.Y(_2100_),
    .A(net125),
    .B(_2099_));
 sg13g2_a21oi_1 _5357_ (.A1(_2098_),
    .A2(_2100_),
    .Y(_0145_),
    .B1(net126));
 sg13g2_nor2_1 _5358_ (.A(_2707_),
    .B(net163),
    .Y(_2101_));
 sg13g2_nor2_1 _5359_ (.A(_1816_),
    .B(net157),
    .Y(_2102_));
 sg13g2_nand2_1 _5360_ (.Y(_2103_),
    .A(_1828_),
    .B(_1841_));
 sg13g2_o21ai_1 _5361_ (.B1(net141),
    .Y(_2104_),
    .A1(_1643_),
    .A2(net142));
 sg13g2_a221oi_1 _5362_ (.B2(_2103_),
    .C1(_2104_),
    .B1(_2102_),
    .A1(_1814_),
    .Y(_0146_),
    .A2(_2101_));
 sg13g2_nand2_1 _5363_ (.Y(_2105_),
    .A(\g.g_y[1].g_x[3].t.out_sc ),
    .B(net145));
 sg13g2_mux2_1 _5364_ (.A0(_1568_),
    .A1(_1822_),
    .S(_1570_),
    .X(_2106_));
 sg13g2_nand2_1 _5365_ (.Y(_2107_),
    .A(net125),
    .B(_2106_));
 sg13g2_a21oi_1 _5366_ (.A1(_2105_),
    .A2(_2107_),
    .Y(_0147_),
    .B1(net126));
 sg13g2_nor4_1 _5367_ (.A(_2549_),
    .B(net159),
    .C(_1778_),
    .D(_1784_),
    .Y(_2108_));
 sg13g2_nand2_1 _5368_ (.Y(_2109_),
    .A(_2549_),
    .B(net147));
 sg13g2_a21oi_1 _5369_ (.A1(_1795_),
    .A2(_1799_),
    .Y(_2110_),
    .B1(_2109_));
 sg13g2_buf_1 _5370_ (.A(net146),
    .X(_2111_));
 sg13g2_o21ai_1 _5371_ (.B1(net152),
    .Y(_2112_),
    .A1(_1577_),
    .A2(net124));
 sg13g2_nor3_1 _5372_ (.A(_2108_),
    .B(_2110_),
    .C(_2112_),
    .Y(_0148_));
 sg13g2_buf_1 _5373_ (.A(net161),
    .X(_2113_));
 sg13g2_nand2_1 _5374_ (.Y(_2114_),
    .A(\g.g_y[1].g_x[5].t.out_sc ),
    .B(net140));
 sg13g2_mux2_1 _5375_ (.A0(_1739_),
    .A1(_1511_),
    .S(_1505_),
    .X(_2115_));
 sg13g2_nand2_1 _5376_ (.Y(_2116_),
    .A(net125),
    .B(_2115_));
 sg13g2_a21oi_1 _5377_ (.A1(_2114_),
    .A2(_2116_),
    .Y(_0149_),
    .B1(net126));
 sg13g2_nand2_1 _5378_ (.Y(_2117_),
    .A(_2472_),
    .B(net147));
 sg13g2_a21oi_1 _5379_ (.A1(_1746_),
    .A2(_1761_),
    .Y(_2118_),
    .B1(_2117_));
 sg13g2_nor4_1 _5380_ (.A(_2472_),
    .B(net159),
    .C(_1725_),
    .D(_1733_),
    .Y(_2119_));
 sg13g2_o21ai_1 _5381_ (.B1(_0516_),
    .Y(_2120_),
    .A1(_1514_),
    .A2(_2111_));
 sg13g2_nor3_1 _5382_ (.A(_2118_),
    .B(_2119_),
    .C(_2120_),
    .Y(_0150_));
 sg13g2_nor4_1 _5383_ (.A(_1710_),
    .B(net159),
    .C(_1708_),
    .D(_1709_),
    .Y(_2121_));
 sg13g2_nand2_1 _5384_ (.Y(_2122_),
    .A(_1710_),
    .B(net147));
 sg13g2_a21oi_1 _5385_ (.A1(_1680_),
    .A2(_1703_),
    .Y(_2123_),
    .B1(_2122_));
 sg13g2_o21ai_1 _5386_ (.B1(_0516_),
    .Y(_2124_),
    .A1(\g.g_y[1].g_x[7].t.out_sc ),
    .A2(net124));
 sg13g2_nor3_1 _5387_ (.A(_2121_),
    .B(_2123_),
    .C(_2124_),
    .Y(_0151_));
 sg13g2_a221oi_1 _5388_ (.B2(_1431_),
    .C1(_1442_),
    .B1(_1449_),
    .A1(_1432_),
    .Y(_2125_),
    .A2(_1437_));
 sg13g2_a21o_1 _5389_ (.A2(_1850_),
    .A1(_1442_),
    .B1(_2125_),
    .X(_2126_));
 sg13g2_nand2_1 _5390_ (.Y(_2127_),
    .A(\g.g_y[2].g_x[0].t.out_sc ),
    .B(net162));
 sg13g2_o21ai_1 _5391_ (.B1(_2127_),
    .Y(_2128_),
    .A1(net163),
    .A2(_2126_));
 sg13g2_and2_1 _5392_ (.A(net155),
    .B(_2128_),
    .X(_0152_));
 sg13g2_nand2_1 _5393_ (.Y(_2129_),
    .A(_1081_),
    .B(net147));
 sg13g2_a21oi_1 _5394_ (.A1(_1661_),
    .A2(_1666_),
    .Y(_2130_),
    .B1(_2129_));
 sg13g2_or2_1 _5395_ (.X(_2131_),
    .B(_2061_),
    .A(_1081_));
 sg13g2_a21oi_1 _5396_ (.A1(_1613_),
    .A2(_1648_),
    .Y(_2132_),
    .B1(_2131_));
 sg13g2_o21ai_1 _5397_ (.B1(net152),
    .Y(_2133_),
    .A1(\g.g_y[2].g_x[1].t.out_sc ),
    .A2(net124));
 sg13g2_nor3_1 _5398_ (.A(_2130_),
    .B(_2132_),
    .C(_2133_),
    .Y(_0153_));
 sg13g2_nand2_1 _5399_ (.Y(_2134_),
    .A(\g.g_y[2].g_x[2].t.out_sc ),
    .B(net140));
 sg13g2_nor2_1 _5400_ (.A(net36),
    .B(_1585_),
    .Y(_2135_));
 sg13g2_a221oi_1 _5401_ (.B2(_1372_),
    .C1(_1362_),
    .B1(_1370_),
    .A1(_1364_),
    .Y(_2136_),
    .A2(_1366_));
 sg13g2_or3_1 _5402_ (.A(net158),
    .B(_2135_),
    .C(_2136_),
    .X(_2137_));
 sg13g2_a21oi_1 _5403_ (.A1(_2134_),
    .A2(_2137_),
    .Y(_0154_),
    .B1(net126));
 sg13g2_nand2_1 _5404_ (.Y(_2138_),
    .A(_1554_),
    .B(_0996_));
 sg13g2_a221oi_1 _5405_ (.B2(_1056_),
    .C1(_2138_),
    .B1(_1555_),
    .A1(_1013_),
    .Y(_2139_),
    .A2(_1405_));
 sg13g2_nand4_1 _5406_ (.B(_1295_),
    .C(_1595_),
    .A(_0993_),
    .Y(_2140_),
    .D(_1598_));
 sg13g2_nand3b_1 _5407_ (.B(_2140_),
    .C(_2075_),
    .Y(_2141_),
    .A_N(_2139_));
 sg13g2_and4_1 _5408_ (.A(_0993_),
    .B(_1298_),
    .C(_1583_),
    .D(_1590_),
    .X(_2142_));
 sg13g2_a21o_1 _5409_ (.A2(_1580_),
    .A1(_1554_),
    .B1(_2142_),
    .X(_2143_));
 sg13g2_nand2_1 _5410_ (.Y(_2144_),
    .A(net145),
    .B(_0046_));
 sg13g2_o21ai_1 _5411_ (.B1(_2144_),
    .Y(_0155_),
    .A1(_2141_),
    .A2(_2143_));
 sg13g2_nand2_1 _5412_ (.Y(_2145_),
    .A(\g.g_y[2].g_x[4].t.out_sc ),
    .B(net140));
 sg13g2_nor2_1 _5413_ (.A(_1310_),
    .B(_1773_),
    .Y(_2146_));
 sg13g2_a221oi_1 _5414_ (.B2(_1348_),
    .C1(net38),
    .B1(_1284_),
    .A1(net39),
    .Y(_2147_),
    .A2(_1282_));
 sg13g2_or3_1 _5415_ (.A(net158),
    .B(_2146_),
    .C(_2147_),
    .X(_2148_));
 sg13g2_a21oi_1 _5416_ (.A1(_2145_),
    .A2(_2148_),
    .Y(_0156_),
    .B1(net126));
 sg13g2_nor4_1 _5417_ (.A(_1543_),
    .B(net159),
    .C(_1535_),
    .D(_1542_),
    .Y(_2149_));
 sg13g2_nand2_1 _5418_ (.Y(_2150_),
    .A(_1543_),
    .B(net147));
 sg13g2_a21oi_1 _5419_ (.A1(_1485_),
    .A2(_1517_),
    .Y(_2151_),
    .B1(_2150_));
 sg13g2_o21ai_1 _5420_ (.B1(net152),
    .Y(_2152_),
    .A1(\g.g_y[2].g_x[5].t.out_sc ),
    .A2(net124));
 sg13g2_nor3_1 _5421_ (.A(_2149_),
    .B(_2151_),
    .C(_2152_),
    .Y(_0157_));
 sg13g2_nand2_1 _5422_ (.Y(_2153_),
    .A(\g.g_y[2].g_x[6].t.out_sc ),
    .B(net140));
 sg13g2_mux2_1 _5423_ (.A0(_1217_),
    .A1(_1547_),
    .S(_1519_),
    .X(_2154_));
 sg13g2_nand2_1 _5424_ (.Y(_2155_),
    .A(net125),
    .B(_2154_));
 sg13g2_a21oi_1 _5425_ (.A1(_2153_),
    .A2(_2155_),
    .Y(_0158_),
    .B1(_2032_));
 sg13g2_nand2_1 _5426_ (.Y(_2156_),
    .A(_1221_),
    .B(_2113_));
 sg13g2_o21ai_1 _5427_ (.B1(net43),
    .Y(_2157_),
    .A1(_1150_),
    .A2(_1153_));
 sg13g2_a22oi_1 _5428_ (.Y(_2158_),
    .B1(_1249_),
    .B2(_1243_),
    .A2(_1248_),
    .A1(net42));
 sg13g2_nand2_1 _5429_ (.Y(_2159_),
    .A(_1155_),
    .B(_2158_));
 sg13g2_nand3_1 _5430_ (.B(_2157_),
    .C(_2159_),
    .A(net144),
    .Y(_2160_));
 sg13g2_a21oi_1 _5431_ (.A1(_2156_),
    .A2(_2160_),
    .Y(_0159_),
    .B1(_2032_));
 sg13g2_nand2_1 _5432_ (.Y(_2161_),
    .A(_0859_),
    .B(net147));
 sg13g2_a21oi_1 _5433_ (.A1(_1467_),
    .A2(_1472_),
    .Y(_2162_),
    .B1(_2161_));
 sg13g2_or2_1 _5434_ (.X(_2163_),
    .B(_2061_),
    .A(_0859_));
 sg13g2_a21oi_1 _5435_ (.A1(_1429_),
    .A2(_1456_),
    .Y(_2164_),
    .B1(_2163_));
 sg13g2_o21ai_1 _5436_ (.B1(net152),
    .Y(_2165_),
    .A1(\g.g_y[3].g_x[0].t.out_sc ),
    .A2(net124));
 sg13g2_nor3_1 _5437_ (.A(_2162_),
    .B(_2164_),
    .C(_2165_),
    .Y(_0160_));
 sg13g2_nand2_1 _5438_ (.Y(_2166_),
    .A(\g.g_y[3].g_x[1].t.out_sc ),
    .B(net140));
 sg13g2_a221oi_1 _5439_ (.B2(_1093_),
    .C1(_1097_),
    .B1(_1071_),
    .A1(_1064_),
    .Y(_2167_),
    .A2(_1066_));
 sg13g2_nor2_1 _5440_ (.A(net45),
    .B(_1462_),
    .Y(_2168_));
 sg13g2_or3_1 _5441_ (.A(_2082_),
    .B(_2167_),
    .C(_2168_),
    .X(_2169_));
 sg13g2_a21oi_1 _5442_ (.A1(_2166_),
    .A2(_2169_),
    .Y(_0161_),
    .B1(net126));
 sg13g2_a22oi_1 _5443_ (.Y(_2170_),
    .B1(_1403_),
    .B2(_1407_),
    .A2(_1401_),
    .A1(_1397_));
 sg13g2_nor2_1 _5444_ (.A(_1395_),
    .B(net163),
    .Y(_2171_));
 sg13g2_nor2_1 _5445_ (.A(_0796_),
    .B(net157),
    .Y(_2172_));
 sg13g2_nand2_1 _5446_ (.Y(_2173_),
    .A(_1389_),
    .B(_1394_));
 sg13g2_o21ai_1 _5447_ (.B1(net141),
    .Y(_2174_),
    .A1(\g.g_y[3].g_x[2].t.out_sc ),
    .A2(net142));
 sg13g2_a221oi_1 _5448_ (.B2(_2173_),
    .C1(_2174_),
    .B1(_2172_),
    .A1(_2170_),
    .Y(_0162_),
    .A2(_2171_));
 sg13g2_nand2_1 _5449_ (.Y(_2175_),
    .A(\g.g_y[3].g_x[3].t.out_sc ),
    .B(net140));
 sg13g2_a221oi_1 _5450_ (.B2(_1010_),
    .C1(_0991_),
    .B1(_1005_),
    .A1(net47),
    .Y(_2176_),
    .A2(_1002_));
 sg13g2_a21oi_1 _5451_ (.A1(net25),
    .A2(_1404_),
    .Y(_2177_),
    .B1(_2176_));
 sg13g2_nand2_1 _5452_ (.Y(_2178_),
    .A(net125),
    .B(_2177_));
 sg13g2_buf_1 _5453_ (.A(net156),
    .X(_2179_));
 sg13g2_a21oi_1 _5454_ (.A1(_2175_),
    .A2(_2178_),
    .Y(_0163_),
    .B1(net123));
 sg13g2_o21ai_1 _5455_ (.B1(_0703_),
    .Y(_2180_),
    .A1(_1335_),
    .A2(_1340_));
 sg13g2_a21oi_1 _5456_ (.A1(_1303_),
    .A2(_1304_),
    .Y(_2181_),
    .B1(_0703_));
 sg13g2_a21oi_1 _5457_ (.A1(_1319_),
    .A2(_2181_),
    .Y(_2182_),
    .B1(net157));
 sg13g2_o21ai_1 _5458_ (.B1(net148),
    .Y(_2183_),
    .A1(\g.g_y[3].g_x[4].t.out_sc ),
    .A2(net144));
 sg13g2_a21oi_1 _5459_ (.A1(_2180_),
    .A2(_2182_),
    .Y(_0164_),
    .B1(_2183_));
 sg13g2_nand2_1 _5460_ (.Y(_2184_),
    .A(\g.g_y[3].g_x[5].t.out_sc ),
    .B(net140));
 sg13g2_a221oi_1 _5461_ (.B2(_0918_),
    .C1(_1258_),
    .B1(_0946_),
    .A1(_0919_),
    .Y(_2185_),
    .A2(_0927_));
 sg13g2_a221oi_1 _5462_ (.B2(_1257_),
    .C1(_0931_),
    .B1(_1255_),
    .A1(_0942_),
    .Y(_2186_),
    .A2(_1254_));
 sg13g2_or3_1 _5463_ (.A(net158),
    .B(_2185_),
    .C(_2186_),
    .X(_2187_));
 sg13g2_a21oi_1 _5464_ (.A1(_2184_),
    .A2(_2187_),
    .Y(_0165_),
    .B1(net123));
 sg13g2_nand2_1 _5465_ (.Y(_2188_),
    .A(_0616_),
    .B(net147));
 sg13g2_a21oi_1 _5466_ (.A1(_1252_),
    .A2(_1271_),
    .Y(_2189_),
    .B1(_2188_));
 sg13g2_nor4_1 _5467_ (.A(_0616_),
    .B(_2066_),
    .C(_1224_),
    .D(_1234_),
    .Y(_2190_));
 sg13g2_o21ai_1 _5468_ (.B1(net152),
    .Y(_2191_),
    .A1(\g.g_y[3].g_x[6].t.out_sc ),
    .A2(_2111_));
 sg13g2_nor3_1 _5469_ (.A(_2189_),
    .B(_2190_),
    .C(_2191_),
    .Y(_0166_));
 sg13g2_nand3_1 _5470_ (.B(_0515_),
    .C(net146),
    .A(_0569_),
    .Y(_2192_));
 sg13g2_a221oi_1 _5471_ (.B2(_1184_),
    .C1(_2192_),
    .B1(_1182_),
    .A1(_0867_),
    .Y(_2193_),
    .A2(_1185_));
 sg13g2_nor3_1 _5472_ (.A(_0569_),
    .B(_2499_),
    .C(net161),
    .Y(_2194_));
 sg13g2_nand3_1 _5473_ (.B(_1177_),
    .C(_2194_),
    .A(_1148_),
    .Y(_2195_));
 sg13g2_nand2_1 _5474_ (.Y(_2196_),
    .A(_2055_),
    .B(_0068_));
 sg13g2_nand3b_1 _5475_ (.B(_2195_),
    .C(_2196_),
    .Y(_0167_),
    .A_N(_2193_));
 sg13g2_nor2_1 _5476_ (.A(_0857_),
    .B(_1113_),
    .Y(_2197_));
 sg13g2_a21oi_1 _5477_ (.A1(_0857_),
    .A2(_0878_),
    .Y(_2198_),
    .B1(_2197_));
 sg13g2_nand2_1 _5478_ (.Y(_2199_),
    .A(\g.g_y[4].g_x[0].t.out_sc ),
    .B(_2052_));
 sg13g2_o21ai_1 _5479_ (.B1(_2199_),
    .Y(_2200_),
    .A1(_2035_),
    .A2(_2198_));
 sg13g2_and2_1 _5480_ (.A(_2543_),
    .B(_2200_),
    .X(_0168_));
 sg13g2_nand2_1 _5481_ (.Y(_2201_),
    .A(_0478_),
    .B(net146));
 sg13g2_a21oi_1 _5482_ (.A1(_1127_),
    .A2(_1131_),
    .Y(_2202_),
    .B1(_2201_));
 sg13g2_nor4_1 _5483_ (.A(_0478_),
    .B(net159),
    .C(_1100_),
    .D(_1108_),
    .Y(_2203_));
 sg13g2_o21ai_1 _5484_ (.B1(net152),
    .Y(_2204_),
    .A1(_0882_),
    .A2(net124));
 sg13g2_nor3_1 _5485_ (.A(_2202_),
    .B(_2203_),
    .C(_2204_),
    .Y(_0169_));
 sg13g2_mux2_1 _5486_ (.A0(_0838_),
    .A1(_0844_),
    .S(net54),
    .X(_2205_));
 sg13g2_and2_1 _5487_ (.A(\g.g_y[4].g_x[2].t.out_sc ),
    .B(_2052_),
    .X(_2206_));
 sg13g2_a21oi_1 _5488_ (.A1(net125),
    .A2(_2205_),
    .Y(_2207_),
    .B1(_2206_));
 sg13g2_nor2_1 _5489_ (.A(net139),
    .B(_2207_),
    .Y(_0170_));
 sg13g2_nor4_1 _5490_ (.A(_1045_),
    .B(net159),
    .C(_1037_),
    .D(_1044_),
    .Y(_2208_));
 sg13g2_nor4_1 _5491_ (.A(_0398_),
    .B(net159),
    .C(_1022_),
    .D(_1032_),
    .Y(_2209_));
 sg13g2_o21ai_1 _5492_ (.B1(net141),
    .Y(_2210_),
    .A1(net164),
    .A2(net124));
 sg13g2_nor3_1 _5493_ (.A(_2208_),
    .B(_2209_),
    .C(_2210_),
    .Y(_0171_));
 sg13g2_nand2_1 _5494_ (.Y(_2211_),
    .A(\g.g_y[4].g_x[4].t.out_sc ),
    .B(net140));
 sg13g2_a221oi_1 _5495_ (.B2(_0706_),
    .C1(_0707_),
    .B1(_0702_),
    .A1(net57),
    .Y(_2212_),
    .A2(_0697_));
 sg13g2_a221oi_1 _5496_ (.B2(_0720_),
    .C1(_0708_),
    .B1(_0718_),
    .A1(net28),
    .Y(_2213_),
    .A2(_0716_));
 sg13g2_or3_1 _5497_ (.A(net158),
    .B(_2212_),
    .C(_2213_),
    .X(_2214_));
 sg13g2_a21oi_1 _5498_ (.A1(_2211_),
    .A2(_2214_),
    .Y(_0172_),
    .B1(net123));
 sg13g2_nand2_1 _5499_ (.Y(_2215_),
    .A(_0328_),
    .B(net165));
 sg13g2_or3_1 _5500_ (.A(net158),
    .B(_0974_),
    .C(_2215_),
    .X(_2216_));
 sg13g2_nor3_1 _5501_ (.A(_0328_),
    .B(net156),
    .C(net161),
    .Y(_2217_));
 sg13g2_nand3_1 _5502_ (.B(_0950_),
    .C(_2217_),
    .A(_0914_),
    .Y(_2218_));
 sg13g2_nand2_1 _5503_ (.Y(_2219_),
    .A(net145),
    .B(_0082_));
 sg13g2_nand3_1 _5504_ (.B(_2218_),
    .C(_2219_),
    .A(_2216_),
    .Y(_0173_));
 sg13g2_mux2_1 _5505_ (.A0(_0638_),
    .A1(net23),
    .S(net58),
    .X(_2220_));
 sg13g2_nand2_1 _5506_ (.Y(_2221_),
    .A(net59),
    .B(_2220_));
 sg13g2_o21ai_1 _5507_ (.B1(_2221_),
    .Y(_2222_),
    .A1(net59),
    .A2(_0980_));
 sg13g2_nand2_1 _5508_ (.Y(_2223_),
    .A(\g.g_y[4].g_x[6].t.out_sc ),
    .B(net161));
 sg13g2_o21ai_1 _5509_ (.B1(_2223_),
    .Y(_2224_),
    .A1(net163),
    .A2(_2222_));
 sg13g2_and2_1 _5510_ (.A(net155),
    .B(_2224_),
    .X(_0174_));
 sg13g2_nor2_1 _5511_ (.A(_0579_),
    .B(_0566_),
    .Y(_2225_));
 sg13g2_a221oi_1 _5512_ (.B2(_0653_),
    .C1(net61),
    .B1(_0651_),
    .A1(_0576_),
    .Y(_2226_),
    .A2(_0649_));
 sg13g2_nor2_1 _5513_ (.A(_2225_),
    .B(_2226_),
    .Y(_2227_));
 sg13g2_nor2_1 _5514_ (.A(_0623_),
    .B(_2095_),
    .Y(_2228_));
 sg13g2_a21oi_1 _5515_ (.A1(_2069_),
    .A2(_2227_),
    .Y(_2229_),
    .B1(_2228_));
 sg13g2_nor2_1 _5516_ (.A(net139),
    .B(_2229_),
    .Y(_0175_));
 sg13g2_nand2_1 _5517_ (.Y(_2230_),
    .A(_0271_),
    .B(net146));
 sg13g2_a21oi_1 _5518_ (.A1(_0895_),
    .A2(_0900_),
    .Y(_2231_),
    .B1(_2230_));
 sg13g2_or2_1 _5519_ (.X(_2232_),
    .B(net160),
    .A(_0271_));
 sg13g2_a21oi_1 _5520_ (.A1(_0853_),
    .A2(_0887_),
    .Y(_2233_),
    .B1(_2232_));
 sg13g2_o21ai_1 _5521_ (.B1(net141),
    .Y(_2234_),
    .A1(\g.g_y[5].g_x[0].t.out_sc ),
    .A2(net124));
 sg13g2_nor3_1 _5522_ (.A(_2231_),
    .B(_2233_),
    .C(_2234_),
    .Y(_0176_));
 sg13g2_nand2_1 _5523_ (.Y(_2235_),
    .A(\g.g_y[5].g_x[1].t.out_sc ),
    .B(_2113_));
 sg13g2_a221oi_1 _5524_ (.B2(_0503_),
    .C1(_0509_),
    .B1(_0501_),
    .A1(_0484_),
    .Y(_2236_),
    .A2(_0483_));
 sg13g2_a21oi_1 _5525_ (.A1(net29),
    .A2(_1102_),
    .Y(_2237_),
    .B1(_2236_));
 sg13g2_nand2_1 _5526_ (.Y(_2238_),
    .A(net125),
    .B(_2237_));
 sg13g2_a21oi_1 _5527_ (.A1(_2235_),
    .A2(_2238_),
    .Y(_0177_),
    .B1(net123));
 sg13g2_nand2_1 _5528_ (.Y(_2239_),
    .A(_2741_),
    .B(net165));
 sg13g2_or3_1 _5529_ (.A(net158),
    .B(_0827_),
    .C(_2239_),
    .X(_2240_));
 sg13g2_nor3_1 _5530_ (.A(_2741_),
    .B(net156),
    .C(net161),
    .Y(_2241_));
 sg13g2_nand3_1 _5531_ (.B(_0812_),
    .C(_2241_),
    .A(_0775_),
    .Y(_2242_));
 sg13g2_nand2_1 _5532_ (.Y(_2243_),
    .A(net145),
    .B(_0091_));
 sg13g2_nand3_1 _5533_ (.B(_2242_),
    .C(_2243_),
    .A(_2240_),
    .Y(_0178_));
 sg13g2_nand2_1 _5534_ (.Y(_2244_),
    .A(\g.g_y[5].g_x[3].t.out_sc ),
    .B(net143));
 sg13g2_nand2_1 _5535_ (.Y(_2245_),
    .A(net63),
    .B(_1026_));
 sg13g2_o21ai_1 _5536_ (.B1(_2245_),
    .Y(_2246_),
    .A1(net63),
    .A2(_0814_));
 sg13g2_nand2_1 _5537_ (.Y(_2247_),
    .A(net144),
    .B(_2246_));
 sg13g2_a21oi_1 _5538_ (.A1(_2244_),
    .A2(_2247_),
    .Y(_0179_),
    .B1(net123));
 sg13g2_nand3b_1 _5539_ (.B(_0694_),
    .C(_0737_),
    .Y(_2248_),
    .A_N(_2599_));
 sg13g2_a21oi_1 _5540_ (.A1(_2599_),
    .A2(_0755_),
    .Y(_2249_),
    .B1(net157));
 sg13g2_o21ai_1 _5541_ (.B1(net148),
    .Y(_2250_),
    .A1(_0390_),
    .A2(net144));
 sg13g2_a21oi_1 _5542_ (.A1(_2248_),
    .A2(_2249_),
    .Y(_0180_),
    .B1(_2250_));
 sg13g2_nand2_1 _5543_ (.Y(_2251_),
    .A(\g.g_y[5].g_x[5].t.out_sc ),
    .B(net143));
 sg13g2_a221oi_1 _5544_ (.B2(_0344_),
    .C1(_0349_),
    .B1(_0342_),
    .A1(net66),
    .Y(_2252_),
    .A2(_0337_));
 sg13g2_a221oi_1 _5545_ (.B2(_0331_),
    .C1(net67),
    .B1(_0679_),
    .A1(_0356_),
    .Y(_2253_),
    .A2(_0678_));
 sg13g2_or3_1 _5546_ (.A(net158),
    .B(_2252_),
    .C(_2253_),
    .X(_2254_));
 sg13g2_a21oi_1 _5547_ (.A1(_2251_),
    .A2(_2254_),
    .Y(_0181_),
    .B1(net123));
 sg13g2_nand2_1 _5548_ (.Y(_2255_),
    .A(_2446_),
    .B(_2040_));
 sg13g2_a21oi_1 _5549_ (.A1(_0665_),
    .A2(_0683_),
    .Y(_2256_),
    .B1(_2255_));
 sg13g2_or2_1 _5550_ (.X(_2257_),
    .B(net160),
    .A(_2446_));
 sg13g2_a21oi_1 _5551_ (.A1(_0613_),
    .A2(_0647_),
    .Y(_2258_),
    .B1(_2257_));
 sg13g2_o21ai_1 _5552_ (.B1(net141),
    .Y(_2259_),
    .A1(\g.g_y[5].g_x[6].t.out_sc ),
    .A2(net142));
 sg13g2_nor3_1 _5553_ (.A(_2256_),
    .B(_2258_),
    .C(_2259_),
    .Y(_0182_));
 sg13g2_nor4_1 _5554_ (.A(_0597_),
    .B(_2066_),
    .C(_0592_),
    .D(_0596_),
    .Y(_2260_));
 sg13g2_nand2_1 _5555_ (.Y(_2261_),
    .A(_0597_),
    .B(_2038_));
 sg13g2_a21oi_1 _5556_ (.A1(_0560_),
    .A2(_0588_),
    .Y(_2262_),
    .B1(_2261_));
 sg13g2_o21ai_1 _5557_ (.B1(net141),
    .Y(_2263_),
    .A1(\g.g_y[5].g_x[7].t.out_sc ),
    .A2(net142));
 sg13g2_nor3_1 _5558_ (.A(_2260_),
    .B(_2262_),
    .C(_2263_),
    .Y(_0183_));
 sg13g2_a221oi_1 _5559_ (.B2(_0286_),
    .C1(net30),
    .B1(_0285_),
    .A1(_0265_),
    .Y(_2264_),
    .A2(_0284_));
 sg13g2_and2_1 _5560_ (.A(net30),
    .B(_0527_),
    .X(_2265_));
 sg13g2_nor3_1 _5561_ (.A(_2047_),
    .B(_2264_),
    .C(_2265_),
    .Y(_2266_));
 sg13g2_a21oi_1 _5562_ (.A1(\g.g_y[6].g_x[0].t.out_sc ),
    .A2(net157),
    .Y(_2267_),
    .B1(_2266_));
 sg13g2_nor2_1 _5563_ (.A(_2501_),
    .B(_2267_),
    .Y(_0184_));
 sg13g2_nand3b_1 _5564_ (.B(net166),
    .C(net142),
    .Y(_2268_),
    .A_N(_2753_));
 sg13g2_nor2_1 _5565_ (.A(net162),
    .B(_0514_),
    .Y(_2269_));
 sg13g2_a22oi_1 _5566_ (.Y(_2270_),
    .B1(_2269_),
    .B2(_0539_),
    .A2(_0106_),
    .A1(net157));
 sg13g2_o21ai_1 _5567_ (.B1(_2270_),
    .Y(_0185_),
    .A1(_0513_),
    .A2(_2268_));
 sg13g2_nand2_1 _5568_ (.Y(_2271_),
    .A(\g.g_y[6].g_x[2].t.out_sc ),
    .B(net143));
 sg13g2_nand2_1 _5569_ (.Y(_2272_),
    .A(_2757_),
    .B(_2756_));
 sg13g2_nand3_1 _5570_ (.B(_0534_),
    .C(_2272_),
    .A(_2730_),
    .Y(_2273_));
 sg13g2_nand2_1 _5571_ (.Y(_2274_),
    .A(_2731_),
    .B(_0446_));
 sg13g2_nand3_1 _5572_ (.B(_2273_),
    .C(_2274_),
    .A(net144),
    .Y(_2275_));
 sg13g2_a21oi_1 _5573_ (.A1(_2271_),
    .A2(_2275_),
    .Y(_0186_),
    .B1(net123));
 sg13g2_nand2_1 _5574_ (.Y(_2276_),
    .A(_2588_),
    .B(net146));
 sg13g2_a21oi_1 _5575_ (.A1(_0449_),
    .A2(_0456_),
    .Y(_2277_),
    .B1(_2276_));
 sg13g2_or2_1 _5576_ (.X(_2278_),
    .B(net160),
    .A(_2588_));
 sg13g2_a21oi_1 _5577_ (.A1(_0421_),
    .A2(_0436_),
    .Y(_2279_),
    .B1(_2278_));
 sg13g2_o21ai_1 _5578_ (.B1(net141),
    .Y(_2280_),
    .A1(_2732_),
    .A2(net142));
 sg13g2_nor3_1 _5579_ (.A(_2277_),
    .B(_2279_),
    .C(_2280_),
    .Y(_0187_));
 sg13g2_nand2_1 _5580_ (.Y(_2281_),
    .A(\g.g_y[6].g_x[4].t.out_sc ),
    .B(net143));
 sg13g2_and2_1 _5581_ (.A(_2586_),
    .B(_0380_),
    .X(_2282_));
 sg13g2_a221oi_1 _5582_ (.B2(_2619_),
    .C1(_2586_),
    .B1(_2618_),
    .A1(_2595_),
    .Y(_2283_),
    .A2(_2594_));
 sg13g2_or3_1 _5583_ (.A(net158),
    .B(_2282_),
    .C(_2283_),
    .X(_2284_));
 sg13g2_a21oi_1 _5584_ (.A1(_2281_),
    .A2(_2284_),
    .Y(_0188_),
    .B1(_2179_));
 sg13g2_nor2_1 _5585_ (.A(_2352_),
    .B(net163),
    .Y(_2285_));
 sg13g2_nand2_1 _5586_ (.Y(_2286_),
    .A(_2352_),
    .B(net146));
 sg13g2_a221oi_1 _5587_ (.B2(_0381_),
    .C1(_2286_),
    .B1(_0379_),
    .A1(_0375_),
    .Y(_2287_),
    .A2(_0377_));
 sg13g2_o21ai_1 _5588_ (.B1(_2096_),
    .Y(_2288_),
    .A1(\g.g_y[6].g_x[5].t.out_sc ),
    .A2(net142));
 sg13g2_a221oi_1 _5589_ (.B2(_0374_),
    .C1(_2288_),
    .B1(_2287_),
    .A1(_0365_),
    .Y(_0189_),
    .A2(_2285_));
 sg13g2_nand2_1 _5590_ (.Y(_2289_),
    .A(\g.g_y[6].g_x[6].t.out_sc ),
    .B(net143));
 sg13g2_a22oi_1 _5591_ (.Y(_2290_),
    .B1(_2530_),
    .B2(net84),
    .A2(_0369_),
    .A1(_0368_));
 sg13g2_nand2_1 _5592_ (.Y(_2291_),
    .A(net83),
    .B(_2526_));
 sg13g2_o21ai_1 _5593_ (.B1(_2291_),
    .Y(_2292_),
    .A1(net83),
    .A2(_2290_));
 sg13g2_nand2_1 _5594_ (.Y(_2293_),
    .A(_2077_),
    .B(_2292_));
 sg13g2_a21oi_1 _5595_ (.A1(_2289_),
    .A2(_2293_),
    .Y(_0190_),
    .B1(_2179_));
 sg13g2_and2_1 _5596_ (.A(net86),
    .B(_2427_),
    .X(_2294_));
 sg13g2_a221oi_1 _5597_ (.B2(_2413_),
    .C1(net86),
    .B1(_2422_),
    .A1(net87),
    .Y(_2295_),
    .A2(_2421_));
 sg13g2_nor3_1 _5598_ (.A(_2047_),
    .B(_2294_),
    .C(_2295_),
    .Y(_2296_));
 sg13g2_a21oi_1 _5599_ (.A1(_2489_),
    .A2(_2092_),
    .Y(_2297_),
    .B1(_2296_));
 sg13g2_nor2_1 _5600_ (.A(_2501_),
    .B(_2297_),
    .Y(_0191_));
 sg13g2_inv_1 _5601_ (.Y(_2298_),
    .A(_2386_));
 sg13g2_nor3_1 _5602_ (.A(_2298_),
    .B(_0307_),
    .C(_0310_),
    .Y(_2299_));
 sg13g2_nor2_1 _5603_ (.A(_2386_),
    .B(net71),
    .Y(_2300_));
 sg13g2_nand2_1 _5604_ (.Y(_2301_),
    .A(_0282_),
    .B(_0290_));
 sg13g2_nand2_1 _5605_ (.Y(_2302_),
    .A(_2298_),
    .B(net71));
 sg13g2_a21oi_1 _5606_ (.A1(_0251_),
    .A2(_0257_),
    .Y(_2303_),
    .B1(_2302_));
 sg13g2_a221oi_1 _5607_ (.B2(_2301_),
    .C1(_2303_),
    .B1(_2300_),
    .A1(_0302_),
    .Y(_2304_),
    .A2(_2299_));
 sg13g2_o21ai_1 _5608_ (.B1(net152),
    .Y(_2305_),
    .A1(\g.g_y[7].g_x[0].t.out_sc ),
    .A2(net144));
 sg13g2_a21oi_1 _5609_ (.A1(_2069_),
    .A2(_2304_),
    .Y(_0192_),
    .B1(_2305_));
 sg13g2_nand2_1 _5610_ (.Y(_2306_),
    .A(\g.g_y[7].g_x[1].t.out_sc ),
    .B(_2081_));
 sg13g2_nand2_1 _5611_ (.Y(_2307_),
    .A(_2773_),
    .B(_0296_));
 sg13g2_o21ai_1 _5612_ (.B1(_2307_),
    .Y(_2308_),
    .A1(_2773_),
    .A2(_0473_));
 sg13g2_nand2_1 _5613_ (.Y(_2309_),
    .A(net144),
    .B(_2308_));
 sg13g2_a21oi_1 _5614_ (.A1(_2306_),
    .A2(_2309_),
    .Y(_0193_),
    .B1(net123));
 sg13g2_nor3_1 _5615_ (.A(_2766_),
    .B(net156),
    .C(net162),
    .Y(_2310_));
 sg13g2_o21ai_1 _5616_ (.B1(_2310_),
    .Y(_2311_),
    .A1(_2771_),
    .A2(_0210_));
 sg13g2_nor3_1 _5617_ (.A(_2632_),
    .B(net156),
    .C(net161),
    .Y(_2312_));
 sg13g2_nand3_1 _5618_ (.B(_2765_),
    .C(_2312_),
    .A(_2736_),
    .Y(_2313_));
 sg13g2_nand2_1 _5619_ (.Y(_2314_),
    .A(net145),
    .B(_0123_));
 sg13g2_nand3_1 _5620_ (.B(_2313_),
    .C(_2314_),
    .A(_2311_),
    .Y(_0194_));
 sg13g2_nand2_1 _5621_ (.Y(_2315_),
    .A(\g.g_y[7].g_x[3].t.out_sc ),
    .B(net143));
 sg13g2_a221oi_1 _5622_ (.B2(_2665_),
    .C1(_2629_),
    .B1(_2654_),
    .A1(net78),
    .Y(_2316_),
    .A2(_2649_));
 sg13g2_a221oi_1 _5623_ (.B2(_2627_),
    .C1(_2630_),
    .B1(_2637_),
    .A1(_2641_),
    .Y(_2317_),
    .A2(_2662_));
 sg13g2_or3_1 _5624_ (.A(net162),
    .B(_2316_),
    .C(_2317_),
    .X(_2318_));
 sg13g2_a21oi_1 _5625_ (.A1(_2315_),
    .A2(_2318_),
    .Y(_0195_),
    .B1(_2545_));
 sg13g2_nand2b_1 _5626_ (.Y(_2319_),
    .B(net157),
    .A_N(_2676_));
 sg13g2_nand2_1 _5627_ (.Y(_2320_),
    .A(_2367_),
    .B(_2037_));
 sg13g2_a21o_1 _5628_ (.A2(_2681_),
    .A1(_2660_),
    .B1(_2320_),
    .X(_2321_));
 sg13g2_nor3_1 _5629_ (.A(_2367_),
    .B(_2554_),
    .C(net167),
    .Y(_2322_));
 sg13g2_nor3_1 _5630_ (.A(_2367_),
    .B(\g.g_y[7].g_x[5].t.r_v ),
    .C(net160),
    .Y(_2323_));
 sg13g2_a22oi_1 _5631_ (.Y(_2324_),
    .B1(_2323_),
    .B2(_2622_),
    .A2(_2322_),
    .A1(_2584_));
 sg13g2_and4_1 _5632_ (.A(net148),
    .B(_2319_),
    .C(_2321_),
    .D(_2324_),
    .X(_0196_));
 sg13g2_nand2_1 _5633_ (.Y(_2325_),
    .A(\g.g_y[7].g_x[5].t.out_sc ),
    .B(_2081_));
 sg13g2_nand2_1 _5634_ (.Y(_2326_),
    .A(net89),
    .B(_0358_));
 sg13g2_o21ai_1 _5635_ (.B1(_2326_),
    .Y(_2327_),
    .A1(net89),
    .A2(_2378_));
 sg13g2_nand2_1 _5636_ (.Y(_2328_),
    .A(_2077_),
    .B(_2327_));
 sg13g2_a21oi_1 _5637_ (.A1(_2325_),
    .A2(_2328_),
    .Y(_0197_),
    .B1(_2545_));
 sg13g2_nor3_1 _5638_ (.A(_2348_),
    .B(_2092_),
    .C(_2496_),
    .Y(_2329_));
 sg13g2_nand2_1 _5639_ (.Y(_2330_),
    .A(_2348_),
    .B(_2038_));
 sg13g2_a21oi_1 _5640_ (.A1(_2384_),
    .A2(_2430_),
    .Y(_2331_),
    .B1(_2330_));
 sg13g2_o21ai_1 _5641_ (.B1(_2096_),
    .Y(_2332_),
    .A1(_2373_),
    .A2(net142));
 sg13g2_nor3_1 _5642_ (.A(_2329_),
    .B(_2331_),
    .C(_2332_),
    .Y(_0198_));
 sg13g2_nor2_1 _5643_ (.A(_2491_),
    .B(net81),
    .Y(_2333_));
 sg13g2_a21oi_1 _5644_ (.A1(net81),
    .A2(_2513_),
    .Y(_2334_),
    .B1(_2333_));
 sg13g2_nor2_1 _5645_ (.A(_2481_),
    .B(_1765_),
    .Y(_2335_));
 sg13g2_a21oi_1 _5646_ (.A1(_2481_),
    .A2(_2334_),
    .Y(_2336_),
    .B1(_2335_));
 sg13g2_inv_1 _5647_ (.Y(\g.g_y[0].g_x[7].t.out_r ),
    .A(_2336_));
 sg13g2_mux2_1 _5648_ (.A0(_2475_),
    .A1(_1493_),
    .S(_1492_),
    .X(\g.g_y[1].g_x[7].t.out_r ));
 sg13g2_nor2_1 _5649_ (.A(_1524_),
    .B(_1525_),
    .Y(_2337_));
 sg13g2_nor3_1 _5650_ (.A(net40),
    .B(_1529_),
    .C(_1532_),
    .Y(_2338_));
 sg13g2_a21o_1 _5651_ (.A2(_2337_),
    .A1(_1216_),
    .B1(_2338_),
    .X(\g.g_y[2].g_x[7].t.out_r ));
 sg13g2_nand2_1 _5652_ (.Y(_2339_),
    .A(_0924_),
    .B(_0923_));
 sg13g2_o21ai_1 _5653_ (.B1(_2339_),
    .Y(\g.g_y[3].g_x[7].t.out_r ),
    .A1(_0954_),
    .A2(_0924_));
 sg13g2_a21o_1 _5654_ (.A2(_0638_),
    .A1(_0958_),
    .B1(_0959_),
    .X(_2340_));
 sg13g2_mux2_1 _5655_ (.A0(\g.g_y[4].g_x[7].t.out_sc ),
    .A1(_0979_),
    .S(net59),
    .X(_2341_));
 sg13g2_nand2_1 _5656_ (.Y(_2342_),
    .A(net58),
    .B(_2341_));
 sg13g2_o21ai_1 _5657_ (.B1(_2342_),
    .Y(\g.g_y[4].g_x[7].t.out_r ),
    .A1(_0642_),
    .A2(_2340_));
 sg13g2_inv_1 _5658_ (.Y(_2343_),
    .A(_2449_));
 sg13g2_nand2_1 _5659_ (.Y(_2344_),
    .A(net65),
    .B(_0334_));
 sg13g2_o21ai_1 _5660_ (.B1(_2344_),
    .Y(\g.g_y[5].g_x[7].t.out_r ),
    .A1(_2343_),
    .A2(_0335_));
 sg13g2_a21oi_1 _5661_ (.A1(_2527_),
    .A2(_2438_),
    .Y(_2345_),
    .B1(_0370_));
 sg13g2_mux2_1 _5662_ (.A0(_2489_),
    .A1(_2533_),
    .S(_2458_),
    .X(_2346_));
 sg13g2_mux2_1 _5663_ (.A0(_2345_),
    .A1(_2346_),
    .S(_2454_),
    .X(\g.g_y[6].g_x[7].t.out_r ));
 sg13g2_nand2_1 _5664_ (.Y(_2347_),
    .A(_2383_),
    .B(_2670_));
 sg13g2_o21ai_1 _5665_ (.B1(_2347_),
    .Y(\g.g_y[7].g_x[7].t.out_r ),
    .A1(_2508_),
    .A2(_2383_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _5675__183 (.L_HI(net183));
 sg13g2_buf_1 _5668_ (.A(net169),
    .X(uio_oe[0]));
 sg13g2_buf_1 _5669_ (.A(net170),
    .X(uio_oe[1]));
 sg13g2_buf_1 _5670_ (.A(net171),
    .X(uio_oe[2]));
 sg13g2_buf_1 _5671_ (.A(net172),
    .X(uio_oe[3]));
 sg13g2_buf_1 _5672_ (.A(net173),
    .X(uio_oe[4]));
 sg13g2_buf_1 _5673_ (.A(net174),
    .X(uio_oe[5]));
 sg13g2_buf_1 _5674_ (.A(net175),
    .X(uio_oe[6]));
 sg13g2_buf_1 _5675_ (.A(net183),
    .X(uio_oe[7]));
 sg13g2_buf_1 _5676_ (.A(net176),
    .X(uio_out[0]));
 sg13g2_buf_1 _5677_ (.A(net177),
    .X(uio_out[1]));
 sg13g2_buf_1 _5678_ (.A(net178),
    .X(uio_out[2]));
 sg13g2_buf_1 _5679_ (.A(net179),
    .X(uio_out[3]));
 sg13g2_buf_1 _5680_ (.A(net180),
    .X(uio_out[4]));
 sg13g2_buf_1 _5681_ (.A(net181),
    .X(uio_out[5]));
 sg13g2_buf_1 _5682_ (.A(net182),
    .X(uio_out[6]));
 sg13g2_buf_1 _5683_ (.A(\g.g_y[7].g_x[7].t.out_sc ),
    .X(net14));
 sg13g2_buf_1 _5684_ (.A(\g.g_y[0].g_x[7].t.out_r ),
    .X(net15));
 sg13g2_buf_1 _5685_ (.A(\g.g_y[1].g_x[7].t.out_r ),
    .X(net16));
 sg13g2_buf_1 _5686_ (.A(\g.g_y[2].g_x[7].t.out_r ),
    .X(net17));
 sg13g2_buf_1 _5687_ (.A(\g.g_y[3].g_x[7].t.out_r ),
    .X(net18));
 sg13g2_buf_1 _5688_ (.A(\g.g_y[4].g_x[7].t.out_r ),
    .X(net19));
 sg13g2_buf_1 _5689_ (.A(\g.g_y[5].g_x[7].t.out_r ),
    .X(net20));
 sg13g2_buf_1 _5690_ (.A(\g.g_y[6].g_x[7].t.out_r ),
    .X(net21));
 sg13g2_buf_1 _5691_ (.A(\g.g_y[7].g_x[7].t.out_r ),
    .X(net22));
 sg13g2_dllrq_1 \g.g_y[0].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0000_),
    .GATE_N(net100),
    .RESET_B(net184),
    .Q(\g.g_y[0].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0001_),
    .GATE_N(net92),
    .RESET_B(net185),
    .Q(\g.g_y[0].g_x[0].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0002_),
    .GATE_N(net92),
    .RESET_B(net186),
    .Q(\g.g_y[0].g_x[0].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0000_),
    .GATE_N(net121),
    .RESET_B(net187),
    .Q(\g.g_y[0].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[0].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net188),
    .D(_0135_),
    .Q_N(_2859_),
    .Q(\g.g_y[0].g_x[0].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0000_),
    .GATE_N(net110),
    .RESET_B(net189),
    .Q(\g.g_y[0].g_x[0].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0007_),
    .GATE_N(net100),
    .RESET_B(net190),
    .Q(\g.g_y[0].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0007_),
    .GATE_N(net121),
    .RESET_B(net191),
    .Q(\g.g_y[0].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[1].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net192),
    .D(_0136_),
    .Q_N(_2858_),
    .Q(\g.g_y[0].g_x[1].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0007_),
    .GATE_N(net110),
    .RESET_B(net193),
    .Q(\g.g_y[0].g_x[1].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0008_),
    .GATE_N(net101),
    .RESET_B(net194),
    .Q(\g.g_y[0].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0009_),
    .GATE_N(net128),
    .RESET_B(net195),
    .Q(\g.g_y[0].g_x[2].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0010_),
    .GATE_N(net128),
    .RESET_B(net196),
    .Q(\g.g_y[0].g_x[2].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0008_),
    .GATE_N(net120),
    .RESET_B(net197),
    .Q(\g.g_y[0].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[2].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net198),
    .D(_0137_),
    .Q_N(_2857_),
    .Q(\g.g_y[0].g_x[2].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0008_),
    .GATE_N(net111),
    .RESET_B(net199),
    .Q(\g.g_y[0].g_x[2].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0012_),
    .GATE_N(net101),
    .RESET_B(net200),
    .Q(\g.g_y[0].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0012_),
    .GATE_N(net120),
    .RESET_B(net201),
    .Q(\g.g_y[0].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[3].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net202),
    .D(_0138_),
    .Q_N(_2856_),
    .Q(\g.g_y[0].g_x[3].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0012_),
    .GATE_N(net111),
    .RESET_B(net203),
    .Q(\g.g_y[0].g_x[3].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0013_),
    .GATE_N(net93),
    .RESET_B(net204),
    .Q(\g.g_y[0].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0014_),
    .GATE_N(net91),
    .RESET_B(net205),
    .Q(\g.g_y[0].g_x[4].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0015_),
    .GATE_N(net91),
    .RESET_B(net206),
    .Q(\g.g_y[0].g_x[4].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0013_),
    .GATE_N(net113),
    .RESET_B(net207),
    .Q(\g.g_y[0].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[4].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net208),
    .D(_0139_),
    .Q_N(_2855_),
    .Q(\g.g_y[0].g_x[4].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0013_),
    .GATE_N(net103),
    .RESET_B(net209),
    .Q(\g.g_y[0].g_x[4].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0016_),
    .GATE_N(net99),
    .RESET_B(net210),
    .Q(\g.g_y[0].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0016_),
    .GATE_N(net122),
    .RESET_B(net211),
    .Q(\g.g_y[0].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[5].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net212),
    .D(_0140_),
    .Q_N(_2854_),
    .Q(\g.g_y[0].g_x[5].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0016_),
    .GATE_N(net109),
    .RESET_B(net213),
    .Q(\g.g_y[0].g_x[5].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0017_),
    .GATE_N(net98),
    .RESET_B(net214),
    .Q(\g.g_y[0].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0018_),
    .GATE_N(net128),
    .RESET_B(net215),
    .Q(\g.g_y[0].g_x[6].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0019_),
    .GATE_N(net128),
    .RESET_B(net216),
    .Q(\g.g_y[0].g_x[6].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0017_),
    .GATE_N(net118),
    .RESET_B(net217),
    .Q(\g.g_y[0].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[6].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net218),
    .D(_0141_),
    .Q_N(_2853_),
    .Q(\g.g_y[0].g_x[6].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0017_),
    .GATE_N(net108),
    .RESET_B(net219),
    .Q(\g.g_y[0].g_x[6].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0020_),
    .GATE_N(net102),
    .RESET_B(net220),
    .Q(\g.g_y[0].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0020_),
    .GATE_N(net122),
    .RESET_B(net221),
    .Q(\g.g_y[0].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[7].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net222),
    .D(_0142_),
    .Q_N(_2852_),
    .Q(\g.g_y[0].g_x[7].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0020_),
    .GATE_N(net108),
    .RESET_B(net223),
    .Q(\g.g_y[0].g_x[7].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0021_),
    .GATE_N(net100),
    .RESET_B(net224),
    .Q(\g.g_y[1].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0021_),
    .GATE_N(net121),
    .RESET_B(net225),
    .Q(\g.g_y[1].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[0].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net226),
    .D(_0143_),
    .Q_N(_2851_),
    .Q(\g.g_y[1].g_x[0].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0021_),
    .GATE_N(net110),
    .RESET_B(net227),
    .Q(\g.g_y[1].g_x[0].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0022_),
    .GATE_N(net102),
    .RESET_B(net228),
    .Q(\g.g_y[1].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0023_),
    .GATE_N(net130),
    .RESET_B(net229),
    .Q(\g.g_y[1].g_x[1].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0024_),
    .GATE_N(net130),
    .RESET_B(net230),
    .Q(\g.g_y[1].g_x[1].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0022_),
    .GATE_N(net122),
    .RESET_B(net231),
    .Q(\g.g_y[1].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[1].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net232),
    .D(_0144_),
    .Q_N(_2850_),
    .Q(\g.g_y[1].g_x[1].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0022_),
    .GATE_N(net110),
    .RESET_B(net233),
    .Q(\g.g_y[1].g_x[1].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0026_),
    .GATE_N(net101),
    .RESET_B(net234),
    .Q(\g.g_y[1].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0026_),
    .GATE_N(net121),
    .RESET_B(net235),
    .Q(\g.g_y[1].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[2].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net236),
    .D(_0145_),
    .Q_N(_2849_),
    .Q(\g.g_y[1].g_x[2].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0026_),
    .GATE_N(net111),
    .RESET_B(net237),
    .Q(\g.g_y[1].g_x[2].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0027_),
    .GATE_N(net95),
    .RESET_B(net238),
    .Q(\g.g_y[1].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0028_),
    .GATE_N(net132),
    .RESET_B(net239),
    .Q(\g.g_y[1].g_x[3].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0029_),
    .GATE_N(net132),
    .RESET_B(net240),
    .Q(\g.g_y[1].g_x[3].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0027_),
    .GATE_N(net115),
    .RESET_B(net241),
    .Q(\g.g_y[1].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[3].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net242),
    .D(_0146_),
    .Q_N(_2848_),
    .Q(\g.g_y[1].g_x[3].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0027_),
    .GATE_N(net105),
    .RESET_B(net243),
    .Q(\g.g_y[1].g_x[3].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0031_),
    .GATE_N(net95),
    .RESET_B(net244),
    .Q(\g.g_y[1].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0031_),
    .GATE_N(net115),
    .RESET_B(net245),
    .Q(\g.g_y[1].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[4].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net246),
    .D(_0147_),
    .Q_N(_2847_),
    .Q(\g.g_y[1].g_x[4].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0031_),
    .GATE_N(net105),
    .RESET_B(net247),
    .Q(\g.g_y[1].g_x[4].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0032_),
    .GATE_N(net93),
    .RESET_B(net248),
    .Q(\g.g_y[1].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0033_),
    .GATE_N(net129),
    .RESET_B(net249),
    .Q(\g.g_y[1].g_x[5].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0034_),
    .GATE_N(net129),
    .RESET_B(net250),
    .Q(\g.g_y[1].g_x[5].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0032_),
    .GATE_N(net114),
    .RESET_B(net251),
    .Q(\g.g_y[1].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[5].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net252),
    .D(_0148_),
    .Q_N(_2846_),
    .Q(\g.g_y[1].g_x[5].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0032_),
    .GATE_N(net103),
    .RESET_B(net253),
    .Q(\g.g_y[1].g_x[5].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0035_),
    .GATE_N(net98),
    .RESET_B(net254),
    .Q(\g.g_y[1].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0035_),
    .GATE_N(net122),
    .RESET_B(net255),
    .Q(\g.g_y[1].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[6].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net256),
    .D(_0149_),
    .Q_N(_2845_),
    .Q(\g.g_y[1].g_x[6].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0035_),
    .GATE_N(net112),
    .RESET_B(net257),
    .Q(\g.g_y[1].g_x[6].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0036_),
    .GATE_N(net98),
    .RESET_B(net258),
    .Q(\g.g_y[1].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0037_),
    .GATE_N(net133),
    .RESET_B(net259),
    .Q(\g.g_y[1].g_x[7].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0038_),
    .GATE_N(net133),
    .RESET_B(net260),
    .Q(\g.g_y[1].g_x[7].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0036_),
    .GATE_N(net118),
    .RESET_B(net261),
    .Q(\g.g_y[1].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[7].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net262),
    .D(_0150_),
    .Q_N(_2844_),
    .Q(\g.g_y[1].g_x[7].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0036_),
    .GATE_N(net108),
    .RESET_B(net263),
    .Q(\g.g_y[1].g_x[7].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0039_),
    .GATE_N(net100),
    .RESET_B(net264),
    .Q(\g.g_y[2].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0040_),
    .GATE_N(net128),
    .RESET_B(net265),
    .Q(\g.g_y[2].g_x[0].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0041_),
    .GATE_N(net128),
    .RESET_B(net266),
    .Q(\g.g_y[2].g_x[0].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0039_),
    .GATE_N(net121),
    .RESET_B(net267),
    .Q(\g.g_y[2].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[0].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net268),
    .D(_0151_),
    .Q_N(_2843_),
    .Q(\g.g_y[2].g_x[0].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0039_),
    .GATE_N(net112),
    .RESET_B(net269),
    .Q(\g.g_y[2].g_x[0].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0042_),
    .GATE_N(net101),
    .RESET_B(net270),
    .Q(\g.g_y[2].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0042_),
    .GATE_N(net120),
    .RESET_B(net271),
    .Q(\g.g_y[2].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[1].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net272),
    .D(_0152_),
    .Q_N(_2842_),
    .Q(\g.g_y[2].g_x[1].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0042_),
    .GATE_N(net111),
    .RESET_B(net273),
    .Q(\g.g_y[2].g_x[1].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0043_),
    .GATE_N(net95),
    .RESET_B(net274),
    .Q(\g.g_y[2].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0044_),
    .GATE_N(net91),
    .RESET_B(net275),
    .Q(\g.g_y[2].g_x[2].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0045_),
    .GATE_N(net91),
    .RESET_B(net276),
    .Q(\g.g_y[2].g_x[2].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0043_),
    .GATE_N(net115),
    .RESET_B(net277),
    .Q(\g.g_y[2].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[2].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net278),
    .D(_0153_),
    .Q_N(_2841_),
    .Q(\g.g_y[2].g_x[2].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0043_),
    .GATE_N(net105),
    .RESET_B(net279),
    .Q(\g.g_y[2].g_x[2].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0046_),
    .GATE_N(net95),
    .RESET_B(net280),
    .Q(\g.g_y[2].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0046_),
    .GATE_N(net115),
    .RESET_B(net281),
    .Q(\g.g_y[2].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[3].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net282),
    .D(_0154_),
    .Q_N(_2840_),
    .Q(\g.g_y[2].g_x[3].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0046_),
    .GATE_N(net105),
    .RESET_B(net283),
    .Q(\g.g_y[2].g_x[3].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0047_),
    .GATE_N(net95),
    .RESET_B(net284),
    .Q(\g.g_y[2].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0048_),
    .GATE_N(net127),
    .RESET_B(net285),
    .Q(\g.g_y[2].g_x[4].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0049_),
    .GATE_N(net127),
    .RESET_B(net286),
    .Q(\g.g_y[2].g_x[4].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0047_),
    .GATE_N(net115),
    .RESET_B(net287),
    .Q(\g.g_y[2].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[4].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net288),
    .D(_0155_),
    .Q_N(_2839_),
    .Q(\g.g_y[2].g_x[4].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0047_),
    .GATE_N(net105),
    .RESET_B(net289),
    .Q(\g.g_y[2].g_x[4].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0050_),
    .GATE_N(net94),
    .RESET_B(net290),
    .Q(\g.g_y[2].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0050_),
    .GATE_N(net113),
    .RESET_B(net291),
    .Q(\g.g_y[2].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[5].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net292),
    .D(_0156_),
    .Q_N(_2838_),
    .Q(\g.g_y[2].g_x[5].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0050_),
    .GATE_N(net104),
    .RESET_B(net293),
    .Q(\g.g_y[2].g_x[5].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0051_),
    .GATE_N(net97),
    .RESET_B(net294),
    .Q(\g.g_y[2].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0052_),
    .GATE_N(net91),
    .RESET_B(net295),
    .Q(\g.g_y[2].g_x[6].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0053_),
    .GATE_N(net91),
    .RESET_B(net296),
    .Q(\g.g_y[2].g_x[6].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0051_),
    .GATE_N(net114),
    .RESET_B(net297),
    .Q(\g.g_y[2].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[6].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net298),
    .D(_0157_),
    .Q_N(_2837_),
    .Q(\g.g_y[2].g_x[6].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0051_),
    .GATE_N(net107),
    .RESET_B(net299),
    .Q(\g.g_y[2].g_x[6].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0054_),
    .GATE_N(net98),
    .RESET_B(net300),
    .Q(\g.g_y[2].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0054_),
    .GATE_N(net118),
    .RESET_B(net301),
    .Q(\g.g_y[2].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[7].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net302),
    .D(_0158_),
    .Q_N(_2836_),
    .Q(\g.g_y[2].g_x[7].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0054_),
    .GATE_N(net108),
    .RESET_B(net303),
    .Q(\g.g_y[2].g_x[7].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0055_),
    .GATE_N(net101),
    .RESET_B(net304),
    .Q(\g.g_y[3].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0055_),
    .GATE_N(net120),
    .RESET_B(net305),
    .Q(\g.g_y[3].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[0].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net306),
    .D(_0159_),
    .Q_N(_2835_),
    .Q(\g.g_y[3].g_x[0].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0055_),
    .GATE_N(net111),
    .RESET_B(net307),
    .Q(\g.g_y[3].g_x[0].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0056_),
    .GATE_N(net96),
    .RESET_B(net308),
    .Q(\g.g_y[3].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0057_),
    .GATE_N(net132),
    .RESET_B(net309),
    .Q(\g.g_y[3].g_x[1].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0058_),
    .GATE_N(net133),
    .RESET_B(net310),
    .Q(\g.g_y[3].g_x[1].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0056_),
    .GATE_N(net116),
    .RESET_B(net311),
    .Q(\g.g_y[3].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[1].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net312),
    .D(_0160_),
    .Q_N(_2834_),
    .Q(\g.g_y[3].g_x[1].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0056_),
    .GATE_N(net106),
    .RESET_B(net313),
    .Q(\g.g_y[3].g_x[1].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0059_),
    .GATE_N(net95),
    .RESET_B(net314),
    .Q(\g.g_y[3].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0059_),
    .GATE_N(net115),
    .RESET_B(net315),
    .Q(\g.g_y[3].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[2].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net316),
    .D(_0161_),
    .Q_N(_2833_),
    .Q(\g.g_y[3].g_x[2].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0059_),
    .GATE_N(net105),
    .RESET_B(net317),
    .Q(\g.g_y[3].g_x[2].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0060_),
    .GATE_N(net95),
    .RESET_B(net318),
    .Q(\g.g_y[3].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0061_),
    .GATE_N(net129),
    .RESET_B(net319),
    .Q(\g.g_y[3].g_x[3].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0062_),
    .GATE_N(net129),
    .RESET_B(net320),
    .Q(\g.g_y[3].g_x[3].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0060_),
    .GATE_N(net115),
    .RESET_B(net321),
    .Q(\g.g_y[3].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[3].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net322),
    .D(_0162_),
    .Q_N(_2832_),
    .Q(\g.g_y[3].g_x[3].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0060_),
    .GATE_N(net105),
    .RESET_B(net323),
    .Q(\g.g_y[3].g_x[3].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0063_),
    .GATE_N(net94),
    .RESET_B(net324),
    .Q(\g.g_y[3].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0063_),
    .GATE_N(net113),
    .RESET_B(net325),
    .Q(\g.g_y[3].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[4].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net326),
    .D(_0163_),
    .Q_N(_2831_),
    .Q(\g.g_y[3].g_x[4].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0063_),
    .GATE_N(net104),
    .RESET_B(net327),
    .Q(\g.g_y[3].g_x[4].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0064_),
    .GATE_N(net94),
    .RESET_B(net328),
    .Q(\g.g_y[3].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0065_),
    .GATE_N(net132),
    .RESET_B(net329),
    .Q(\g.g_y[3].g_x[5].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0066_),
    .GATE_N(net132),
    .RESET_B(net330),
    .Q(\g.g_y[3].g_x[5].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0064_),
    .GATE_N(net113),
    .RESET_B(net331),
    .Q(\g.g_y[3].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[5].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net332),
    .D(_0164_),
    .Q_N(_2830_),
    .Q(\g.g_y[3].g_x[5].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0064_),
    .GATE_N(net104),
    .RESET_B(net333),
    .Q(\g.g_y[3].g_x[5].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0067_),
    .GATE_N(net93),
    .RESET_B(net334),
    .Q(\g.g_y[3].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0067_),
    .GATE_N(net114),
    .RESET_B(net335),
    .Q(\g.g_y[3].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[6].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net336),
    .D(_0165_),
    .Q_N(_2829_),
    .Q(\g.g_y[3].g_x[6].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0067_),
    .GATE_N(net103),
    .RESET_B(net337),
    .Q(\g.g_y[3].g_x[6].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0068_),
    .GATE_N(net99),
    .RESET_B(net338),
    .Q(\g.g_y[3].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0069_),
    .GATE_N(net130),
    .RESET_B(net339),
    .Q(\g.g_y[3].g_x[7].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0070_),
    .GATE_N(net130),
    .RESET_B(net340),
    .Q(\g.g_y[3].g_x[7].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0068_),
    .GATE_N(net119),
    .RESET_B(net341),
    .Q(\g.g_y[3].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[7].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net342),
    .D(_0166_),
    .Q_N(_2828_),
    .Q(\g.g_y[3].g_x[7].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0068_),
    .GATE_N(net109),
    .RESET_B(net343),
    .Q(\g.g_y[3].g_x[7].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0071_),
    .GATE_N(net101),
    .RESET_B(net344),
    .Q(\g.g_y[4].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0072_),
    .GATE_N(net92),
    .RESET_B(net345),
    .Q(\g.g_y[4].g_x[0].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0073_),
    .GATE_N(net92),
    .RESET_B(net346),
    .Q(\g.g_y[4].g_x[0].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0071_),
    .GATE_N(net120),
    .RESET_B(net347),
    .Q(\g.g_y[4].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[0].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net348),
    .D(_0167_),
    .Q_N(_2827_),
    .Q(\g.g_y[4].g_x[0].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0071_),
    .GATE_N(net111),
    .RESET_B(net349),
    .Q(\g.g_y[4].g_x[0].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0074_),
    .GATE_N(net96),
    .RESET_B(net350),
    .Q(\g.g_y[4].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0074_),
    .GATE_N(net116),
    .RESET_B(net351),
    .Q(\g.g_y[4].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[1].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net352),
    .D(_0168_),
    .Q_N(_2826_),
    .Q(\g.g_y[4].g_x[1].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0074_),
    .GATE_N(net106),
    .RESET_B(net353),
    .Q(\g.g_y[4].g_x[1].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0075_),
    .GATE_N(net96),
    .RESET_B(net354),
    .Q(\g.g_y[4].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0076_),
    .GATE_N(net127),
    .RESET_B(net355),
    .Q(\g.g_y[4].g_x[2].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0077_),
    .GATE_N(net127),
    .RESET_B(net356),
    .Q(\g.g_y[4].g_x[2].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0075_),
    .GATE_N(net116),
    .RESET_B(net357),
    .Q(\g.g_y[4].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[2].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net358),
    .D(_0169_),
    .Q_N(_2825_),
    .Q(\g.g_y[4].g_x[2].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0075_),
    .GATE_N(net106),
    .RESET_B(net359),
    .Q(\g.g_y[4].g_x[2].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0078_),
    .GATE_N(net95),
    .RESET_B(net360),
    .Q(\g.g_y[4].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0078_),
    .GATE_N(net115),
    .RESET_B(net361),
    .Q(\g.g_y[4].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[3].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net362),
    .D(_0170_),
    .Q_N(_2824_),
    .Q(\g.g_y[4].g_x[3].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0078_),
    .GATE_N(net105),
    .RESET_B(net363),
    .Q(\g.g_y[4].g_x[3].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0079_),
    .GATE_N(net94),
    .RESET_B(net364),
    .Q(\g.g_y[4].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0080_),
    .GATE_N(net91),
    .RESET_B(net365),
    .Q(\g.g_y[4].g_x[4].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0081_),
    .GATE_N(net91),
    .RESET_B(net366),
    .Q(\g.g_y[4].g_x[4].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0079_),
    .GATE_N(net113),
    .RESET_B(net367),
    .Q(\g.g_y[4].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[4].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net368),
    .D(_0171_),
    .Q_N(_2823_),
    .Q(\g.g_y[4].g_x[4].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0079_),
    .GATE_N(net104),
    .RESET_B(net369),
    .Q(\g.g_y[4].g_x[4].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0082_),
    .GATE_N(net94),
    .RESET_B(net370),
    .Q(\g.g_y[4].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0082_),
    .GATE_N(net113),
    .RESET_B(net371),
    .Q(\g.g_y[4].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[5].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net372),
    .D(_0172_),
    .Q_N(_2822_),
    .Q(\g.g_y[4].g_x[5].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0082_),
    .GATE_N(net104),
    .RESET_B(net373),
    .Q(\g.g_y[4].g_x[5].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0083_),
    .GATE_N(net93),
    .RESET_B(net374),
    .Q(\g.g_y[4].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0084_),
    .GATE_N(net127),
    .RESET_B(net375),
    .Q(\g.g_y[4].g_x[6].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0085_),
    .GATE_N(net127),
    .RESET_B(net376),
    .Q(\g.g_y[4].g_x[6].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0083_),
    .GATE_N(net114),
    .RESET_B(net377),
    .Q(\g.g_y[4].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[6].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net378),
    .D(_0173_),
    .Q_N(_2821_),
    .Q(\g.g_y[4].g_x[6].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0083_),
    .GATE_N(net103),
    .RESET_B(net379),
    .Q(\g.g_y[4].g_x[6].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0086_),
    .GATE_N(net99),
    .RESET_B(net380),
    .Q(\g.g_y[4].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0086_),
    .GATE_N(net119),
    .RESET_B(net381),
    .Q(\g.g_y[4].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[7].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net382),
    .D(_0174_),
    .Q_N(_2820_),
    .Q(\g.g_y[4].g_x[7].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0086_),
    .GATE_N(net109),
    .RESET_B(net383),
    .Q(\g.g_y[4].g_x[7].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0087_),
    .GATE_N(net100),
    .RESET_B(net384),
    .Q(\g.g_y[5].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0087_),
    .GATE_N(net120),
    .RESET_B(net385),
    .Q(\g.g_y[5].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[0].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net386),
    .D(_0175_),
    .Q_N(_2819_),
    .Q(\g.g_y[5].g_x[0].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0087_),
    .GATE_N(net110),
    .RESET_B(net387),
    .Q(\g.g_y[5].g_x[0].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0088_),
    .GATE_N(net96),
    .RESET_B(net388),
    .Q(\g.g_y[5].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0089_),
    .GATE_N(net129),
    .RESET_B(net389),
    .Q(\g.g_y[5].g_x[1].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0090_),
    .GATE_N(net129),
    .RESET_B(net390),
    .Q(\g.g_y[5].g_x[1].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0088_),
    .GATE_N(net116),
    .RESET_B(net391),
    .Q(\g.g_y[5].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[1].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net392),
    .D(_0176_),
    .Q_N(_2818_),
    .Q(\g.g_y[5].g_x[1].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0088_),
    .GATE_N(net106),
    .RESET_B(net393),
    .Q(\g.g_y[5].g_x[1].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0091_),
    .GATE_N(net96),
    .RESET_B(net394),
    .Q(\g.g_y[5].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0091_),
    .GATE_N(net116),
    .RESET_B(net395),
    .Q(\g.g_y[5].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[2].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net396),
    .D(_0177_),
    .Q_N(_2817_),
    .Q(\g.g_y[5].g_x[2].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0091_),
    .GATE_N(net106),
    .RESET_B(net397),
    .Q(\g.g_y[5].g_x[2].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0092_),
    .GATE_N(net96),
    .RESET_B(net398),
    .Q(\g.g_y[5].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0093_),
    .GATE_N(net132),
    .RESET_B(net399),
    .Q(\g.g_y[5].g_x[3].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0094_),
    .GATE_N(net132),
    .RESET_B(net400),
    .Q(\g.g_y[5].g_x[3].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0092_),
    .GATE_N(net116),
    .RESET_B(net401),
    .Q(\g.g_y[5].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[3].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net402),
    .D(_0178_),
    .Q_N(_2816_),
    .Q(\g.g_y[5].g_x[3].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0092_),
    .GATE_N(net106),
    .RESET_B(net403),
    .Q(\g.g_y[5].g_x[3].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0095_),
    .GATE_N(net94),
    .RESET_B(net404),
    .Q(\g.g_y[5].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0095_),
    .GATE_N(net113),
    .RESET_B(net405),
    .Q(\g.g_y[5].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[4].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net406),
    .D(_0179_),
    .Q_N(_2815_),
    .Q(\g.g_y[5].g_x[4].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0095_),
    .GATE_N(net104),
    .RESET_B(net407),
    .Q(\g.g_y[5].g_x[4].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0096_),
    .GATE_N(net94),
    .RESET_B(net408),
    .Q(\g.g_y[5].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0097_),
    .GATE_N(net129),
    .RESET_B(net409),
    .Q(\g.g_y[5].g_x[5].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0098_),
    .GATE_N(net129),
    .RESET_B(net410),
    .Q(\g.g_y[5].g_x[5].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0096_),
    .GATE_N(net113),
    .RESET_B(net411),
    .Q(\g.g_y[5].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[5].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net412),
    .D(_0180_),
    .Q_N(_2814_),
    .Q(\g.g_y[5].g_x[5].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0096_),
    .GATE_N(net104),
    .RESET_B(net413),
    .Q(\g.g_y[5].g_x[5].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0099_),
    .GATE_N(net93),
    .RESET_B(net414),
    .Q(\g.g_y[5].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0099_),
    .GATE_N(net114),
    .RESET_B(net415),
    .Q(\g.g_y[5].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[6].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net416),
    .D(_0181_),
    .Q_N(_2813_),
    .Q(\g.g_y[5].g_x[6].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0099_),
    .GATE_N(net103),
    .RESET_B(net417),
    .Q(\g.g_y[5].g_x[6].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0100_),
    .GATE_N(net98),
    .RESET_B(net418),
    .Q(\g.g_y[5].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0101_),
    .GATE_N(net133),
    .RESET_B(net419),
    .Q(\g.g_y[5].g_x[7].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0102_),
    .GATE_N(net133),
    .RESET_B(net420),
    .Q(\g.g_y[5].g_x[7].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0100_),
    .GATE_N(net118),
    .RESET_B(net421),
    .Q(\g.g_y[5].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[7].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net422),
    .D(_0182_),
    .Q_N(_2812_),
    .Q(\g.g_y[5].g_x[7].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0100_),
    .GATE_N(net108),
    .RESET_B(net423),
    .Q(\g.g_y[5].g_x[7].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0103_),
    .GATE_N(net100),
    .RESET_B(net424),
    .Q(\g.g_y[6].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0104_),
    .GATE_N(net128),
    .RESET_B(net425),
    .Q(\g.g_y[6].g_x[0].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0105_),
    .GATE_N(net128),
    .RESET_B(net426),
    .Q(\g.g_y[6].g_x[0].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0103_),
    .GATE_N(net118),
    .RESET_B(net427),
    .Q(\g.g_y[6].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[0].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net428),
    .D(_0183_),
    .Q_N(_2811_),
    .Q(\g.g_y[6].g_x[0].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0103_),
    .GATE_N(net110),
    .RESET_B(net429),
    .Q(\g.g_y[6].g_x[0].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0106_),
    .GATE_N(net101),
    .RESET_B(net430),
    .Q(\g.g_y[6].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0106_),
    .GATE_N(net120),
    .RESET_B(net431),
    .Q(\g.g_y[6].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[1].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net432),
    .D(_0184_),
    .Q_N(_2810_),
    .Q(\g.g_y[6].g_x[1].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0106_),
    .GATE_N(net111),
    .RESET_B(net433),
    .Q(\g.g_y[6].g_x[1].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0107_),
    .GATE_N(net96),
    .RESET_B(net434),
    .Q(\g.g_y[6].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0108_),
    .GATE_N(net92),
    .RESET_B(net435),
    .Q(\g.g_y[6].g_x[2].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0109_),
    .GATE_N(net92),
    .RESET_B(net436),
    .Q(\g.g_y[6].g_x[2].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0107_),
    .GATE_N(net116),
    .RESET_B(net437),
    .Q(\g.g_y[6].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[2].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net438),
    .D(_0185_),
    .Q_N(_2809_),
    .Q(\g.g_y[6].g_x[2].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0107_),
    .GATE_N(net106),
    .RESET_B(net439),
    .Q(\g.g_y[6].g_x[2].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0110_),
    .GATE_N(net93),
    .RESET_B(net440),
    .Q(\g.g_y[6].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0110_),
    .GATE_N(net114),
    .RESET_B(net441),
    .Q(\g.g_y[6].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[3].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net442),
    .D(_0186_),
    .Q_N(_2808_),
    .Q(\g.g_y[6].g_x[3].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0110_),
    .GATE_N(net103),
    .RESET_B(net443),
    .Q(\g.g_y[6].g_x[3].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0111_),
    .GATE_N(net93),
    .RESET_B(net444),
    .Q(\g.g_y[6].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0112_),
    .GATE_N(net127),
    .RESET_B(net445),
    .Q(\g.g_y[6].g_x[4].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0113_),
    .GATE_N(net127),
    .RESET_B(net446),
    .Q(\g.g_y[6].g_x[4].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0111_),
    .GATE_N(net114),
    .RESET_B(net447),
    .Q(\g.g_y[6].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[4].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net448),
    .D(_0187_),
    .Q_N(_2807_),
    .Q(\g.g_y[6].g_x[4].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0111_),
    .GATE_N(net103),
    .RESET_B(net449),
    .Q(\g.g_y[6].g_x[4].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0114_),
    .GATE_N(net99),
    .RESET_B(net450),
    .Q(\g.g_y[6].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0114_),
    .GATE_N(net119),
    .RESET_B(net451),
    .Q(\g.g_y[6].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[5].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net452),
    .D(_0188_),
    .Q_N(_2806_),
    .Q(\g.g_y[6].g_x[5].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0114_),
    .GATE_N(net109),
    .RESET_B(net453),
    .Q(\g.g_y[6].g_x[5].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0115_),
    .GATE_N(net99),
    .RESET_B(net454),
    .Q(\g.g_y[6].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0116_),
    .GATE_N(net92),
    .RESET_B(net455),
    .Q(\g.g_y[6].g_x[6].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0117_),
    .GATE_N(_0003_),
    .RESET_B(net456),
    .Q(\g.g_y[6].g_x[6].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0115_),
    .GATE_N(net119),
    .RESET_B(net457),
    .Q(\g.g_y[6].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[6].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net458),
    .D(_0189_),
    .Q_N(_2805_),
    .Q(\g.g_y[6].g_x[6].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0115_),
    .GATE_N(net109),
    .RESET_B(net459),
    .Q(\g.g_y[6].g_x[6].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0118_),
    .GATE_N(net98),
    .RESET_B(net460),
    .Q(\g.g_y[6].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0118_),
    .GATE_N(net118),
    .RESET_B(net461),
    .Q(\g.g_y[6].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[7].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net462),
    .D(_0190_),
    .Q_N(_2804_),
    .Q(\g.g_y[6].g_x[7].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0118_),
    .GATE_N(net108),
    .RESET_B(net463),
    .Q(\g.g_y[6].g_x[7].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0119_),
    .GATE_N(net100),
    .RESET_B(net464),
    .Q(\g.g_y[7].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0119_),
    .GATE_N(net121),
    .RESET_B(net465),
    .Q(\g.g_y[7].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[0].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net466),
    .D(_0191_),
    .Q_N(_2803_),
    .Q(\g.g_y[7].g_x[0].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0119_),
    .GATE_N(net110),
    .RESET_B(net467),
    .Q(\g.g_y[7].g_x[0].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0120_),
    .GATE_N(net100),
    .RESET_B(net468),
    .Q(\g.g_y[7].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0121_),
    .GATE_N(net133),
    .RESET_B(net469),
    .Q(\g.g_y[7].g_x[1].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0122_),
    .GATE_N(net133),
    .RESET_B(net470),
    .Q(\g.g_y[7].g_x[1].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0120_),
    .GATE_N(net121),
    .RESET_B(net471),
    .Q(\g.g_y[7].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[1].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net472),
    .D(_0192_),
    .Q_N(_2802_),
    .Q(\g.g_y[7].g_x[1].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0120_),
    .GATE_N(net110),
    .RESET_B(net473),
    .Q(\g.g_y[7].g_x[1].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0123_),
    .GATE_N(net101),
    .RESET_B(net474),
    .Q(\g.g_y[7].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0123_),
    .GATE_N(net120),
    .RESET_B(net475),
    .Q(\g.g_y[7].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[2].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net476),
    .D(_0193_),
    .Q_N(_2801_),
    .Q(\g.g_y[7].g_x[2].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0123_),
    .GATE_N(net111),
    .RESET_B(net477),
    .Q(\g.g_y[7].g_x[2].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0124_),
    .GATE_N(net99),
    .RESET_B(net478),
    .Q(\g.g_y[7].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0125_),
    .GATE_N(net130),
    .RESET_B(net479),
    .Q(\g.g_y[7].g_x[3].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0126_),
    .GATE_N(net130),
    .RESET_B(net480),
    .Q(\g.g_y[7].g_x[3].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0124_),
    .GATE_N(net119),
    .RESET_B(net481),
    .Q(\g.g_y[7].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[3].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net482),
    .D(_0194_),
    .Q_N(_2800_),
    .Q(\g.g_y[7].g_x[3].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0124_),
    .GATE_N(net109),
    .RESET_B(net483),
    .Q(\g.g_y[7].g_x[3].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0127_),
    .GATE_N(net93),
    .RESET_B(net484),
    .Q(\g.g_y[7].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0127_),
    .GATE_N(net119),
    .RESET_B(net485),
    .Q(\g.g_y[7].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[4].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net486),
    .D(_0195_),
    .Q_N(_2799_),
    .Q(\g.g_y[7].g_x[4].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0127_),
    .GATE_N(net103),
    .RESET_B(net487),
    .Q(\g.g_y[7].g_x[4].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0128_),
    .GATE_N(net99),
    .RESET_B(net488),
    .Q(\g.g_y[7].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0129_),
    .GATE_N(_0030_),
    .RESET_B(net489),
    .Q(\g.g_y[7].g_x[5].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0130_),
    .GATE_N(net132),
    .RESET_B(net490),
    .Q(\g.g_y[7].g_x[5].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0128_),
    .GATE_N(net119),
    .RESET_B(net491),
    .Q(\g.g_y[7].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[5].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net492),
    .D(_0196_),
    .Q_N(_2798_),
    .Q(\g.g_y[7].g_x[5].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0128_),
    .GATE_N(net109),
    .RESET_B(net493),
    .Q(\g.g_y[7].g_x[5].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0131_),
    .GATE_N(net98),
    .RESET_B(net494),
    .Q(\g.g_y[7].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0131_),
    .GATE_N(net118),
    .RESET_B(net495),
    .Q(\g.g_y[7].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[6].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net496),
    .D(_0197_),
    .Q_N(_2797_),
    .Q(\g.g_y[7].g_x[6].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0131_),
    .GATE_N(net108),
    .RESET_B(net497),
    .Q(\g.g_y[7].g_x[6].t.r_v ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0132_),
    .GATE_N(net98),
    .RESET_B(net498),
    .Q(\g.g_y[7].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0133_),
    .GATE_N(net130),
    .RESET_B(net499),
    .Q(\g.g_y[7].g_x[7].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0134_),
    .GATE_N(_0025_),
    .RESET_B(net500),
    .Q(\g.g_y[7].g_x[7].t.r_gnl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0132_),
    .GATE_N(net118),
    .RESET_B(net501),
    .Q(\g.g_y[7].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[7].t.r_sc$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net502),
    .D(_0198_),
    .Q_N(_2796_),
    .Q(\g.g_y[7].g_x[7].t.out_sc ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0132_),
    .GATE_N(net108),
    .RESET_B(net503),
    .Q(\g.g_y[7].g_x[7].t.r_v ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[6]),
    .X(net13));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[7]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[0]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[1]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[2]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[3]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[4]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[5]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[6]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout23 (.A(_0632_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1506_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0991_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0877_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0857_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0712_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0509_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0269_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_2694_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1694_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1627_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1569_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1505_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1361_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1356_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1291_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1279_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1216_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1196_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1166_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1154_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1075_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1063_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1013_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1000_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0942_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0931_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0858_),
    .X(net50));
 sg13g2_buf_1 fanout51 (.A(_0856_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0854_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0778_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0776_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0714_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0707_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0695_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0642_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0625_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0614_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0561_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0392_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0388_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0356_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0335_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0333_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0323_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0268_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0261_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0240_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0228_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_2778_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2772_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2749_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_2740_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_2713_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_2703_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_2643_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_2635_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_2569_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_2486_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_2465_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_2458_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_2455_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_2439_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_2398_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_2397_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_2369_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_2350_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_2349_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(net92),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0003_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net97),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(net97),
    .X(net95));
 sg13g2_buf_1 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_1 fanout97 (.A(_0004_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(net99),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net102),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(net102),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_1 fanout102 (.A(_0004_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(net107),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(net107),
    .X(net105));
 sg13g2_buf_1 fanout106 (.A(net107),
    .X(net106));
 sg13g2_buf_1 fanout107 (.A(_0006_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(net112),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(net112),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_1 fanout112 (.A(_0006_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net117),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(net117),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(net117),
    .X(net115));
 sg13g2_buf_1 fanout116 (.A(net117),
    .X(net116));
 sg13g2_buf_1 fanout117 (.A(_0005_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(net119),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(net122),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(net121),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_1 fanout122 (.A(_0005_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_2179_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_2111_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_2069_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_2032_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_0011_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_0011_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0025_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_1874_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(net133),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_0030_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_1607_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_1193_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_0829_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_0313_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_2546_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_2501_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_2113_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_2096_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_2095_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_2081_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_2077_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_2055_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_2040_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_2038_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_1921_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_1479_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_1062_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_0551_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0516_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_2692_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_2545_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_2543_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_2500_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_2092_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_2082_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_2066_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_2061_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_2052_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_2047_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_2035_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_0810_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_0515_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_2542_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_2034_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_2498_),
    .X(net168));
 sg13g2_tielo _5668__169 (.L_LO(net169));
 sg13g2_tielo _5669__170 (.L_LO(net170));
 sg13g2_tielo _5670__171 (.L_LO(net171));
 sg13g2_tielo _5671__172 (.L_LO(net172));
 sg13g2_tielo _5672__173 (.L_LO(net173));
 sg13g2_tielo _5673__174 (.L_LO(net174));
 sg13g2_tielo _5674__175 (.L_LO(net175));
 sg13g2_tielo _5676__176 (.L_LO(net176));
 sg13g2_tielo _5677__177 (.L_LO(net177));
 sg13g2_tielo _5678__178 (.L_LO(net178));
 sg13g2_tielo _5679__179 (.L_LO(net179));
 sg13g2_tielo _5680__180 (.L_LO(net180));
 sg13g2_tielo _5681__181 (.L_LO(net181));
 sg13g2_tielo _5682__182 (.L_LO(net182));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_184  (.L_HI(net184));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_185  (.L_HI(net185));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_186  (.L_HI(net186));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_187  (.L_HI(net187));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_sc$_SDFF_PN0__188  (.L_HI(net188));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_189  (.L_HI(net189));
 sg13g2_tiehi \g.g_y[0].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_190  (.L_HI(net190));
 sg13g2_tiehi \g.g_y[0].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_191  (.L_HI(net191));
 sg13g2_tiehi \g.g_y[0].g_x[1].t.r_sc$_SDFF_PN0__192  (.L_HI(net192));
 sg13g2_tiehi \g.g_y[0].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_193  (.L_HI(net193));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_194  (.L_HI(net194));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_195  (.L_HI(net195));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_196  (.L_HI(net196));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_197  (.L_HI(net197));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_sc$_SDFF_PN0__198  (.L_HI(net198));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_199  (.L_HI(net199));
 sg13g2_tiehi \g.g_y[0].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_200  (.L_HI(net200));
 sg13g2_tiehi \g.g_y[0].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_201  (.L_HI(net201));
 sg13g2_tiehi \g.g_y[0].g_x[3].t.r_sc$_SDFF_PN0__202  (.L_HI(net202));
 sg13g2_tiehi \g.g_y[0].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_203  (.L_HI(net203));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_204  (.L_HI(net204));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_205  (.L_HI(net205));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_206  (.L_HI(net206));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_207  (.L_HI(net207));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_sc$_SDFF_PN0__208  (.L_HI(net208));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_209  (.L_HI(net209));
 sg13g2_tiehi \g.g_y[0].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_210  (.L_HI(net210));
 sg13g2_tiehi \g.g_y[0].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_211  (.L_HI(net211));
 sg13g2_tiehi \g.g_y[0].g_x[5].t.r_sc$_SDFF_PN0__212  (.L_HI(net212));
 sg13g2_tiehi \g.g_y[0].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_213  (.L_HI(net213));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_214  (.L_HI(net214));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_215  (.L_HI(net215));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_216  (.L_HI(net216));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_217  (.L_HI(net217));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_sc$_SDFF_PN0__218  (.L_HI(net218));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_219  (.L_HI(net219));
 sg13g2_tiehi \g.g_y[0].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_220  (.L_HI(net220));
 sg13g2_tiehi \g.g_y[0].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_221  (.L_HI(net221));
 sg13g2_tiehi \g.g_y[0].g_x[7].t.r_sc$_SDFF_PN0__222  (.L_HI(net222));
 sg13g2_tiehi \g.g_y[0].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_223  (.L_HI(net223));
 sg13g2_tiehi \g.g_y[1].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_224  (.L_HI(net224));
 sg13g2_tiehi \g.g_y[1].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_225  (.L_HI(net225));
 sg13g2_tiehi \g.g_y[1].g_x[0].t.r_sc$_SDFF_PN0__226  (.L_HI(net226));
 sg13g2_tiehi \g.g_y[1].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_227  (.L_HI(net227));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_228  (.L_HI(net228));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_229  (.L_HI(net229));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_230  (.L_HI(net230));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_231  (.L_HI(net231));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_sc$_SDFF_PN0__232  (.L_HI(net232));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_233  (.L_HI(net233));
 sg13g2_tiehi \g.g_y[1].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_234  (.L_HI(net234));
 sg13g2_tiehi \g.g_y[1].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_235  (.L_HI(net235));
 sg13g2_tiehi \g.g_y[1].g_x[2].t.r_sc$_SDFF_PN0__236  (.L_HI(net236));
 sg13g2_tiehi \g.g_y[1].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_237  (.L_HI(net237));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_238  (.L_HI(net238));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_239  (.L_HI(net239));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_240  (.L_HI(net240));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_241  (.L_HI(net241));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_sc$_SDFF_PN0__242  (.L_HI(net242));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_243  (.L_HI(net243));
 sg13g2_tiehi \g.g_y[1].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_244  (.L_HI(net244));
 sg13g2_tiehi \g.g_y[1].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_245  (.L_HI(net245));
 sg13g2_tiehi \g.g_y[1].g_x[4].t.r_sc$_SDFF_PN0__246  (.L_HI(net246));
 sg13g2_tiehi \g.g_y[1].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_247  (.L_HI(net247));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_248  (.L_HI(net248));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_249  (.L_HI(net249));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_250  (.L_HI(net250));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_251  (.L_HI(net251));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_sc$_SDFF_PN0__252  (.L_HI(net252));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_253  (.L_HI(net253));
 sg13g2_tiehi \g.g_y[1].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_254  (.L_HI(net254));
 sg13g2_tiehi \g.g_y[1].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_255  (.L_HI(net255));
 sg13g2_tiehi \g.g_y[1].g_x[6].t.r_sc$_SDFF_PN0__256  (.L_HI(net256));
 sg13g2_tiehi \g.g_y[1].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_257  (.L_HI(net257));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_258  (.L_HI(net258));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_259  (.L_HI(net259));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_260  (.L_HI(net260));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_261  (.L_HI(net261));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_sc$_SDFF_PN0__262  (.L_HI(net262));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_263  (.L_HI(net263));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_264  (.L_HI(net264));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_265  (.L_HI(net265));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_266  (.L_HI(net266));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_267  (.L_HI(net267));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_sc$_SDFF_PN0__268  (.L_HI(net268));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_269  (.L_HI(net269));
 sg13g2_tiehi \g.g_y[2].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_270  (.L_HI(net270));
 sg13g2_tiehi \g.g_y[2].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_271  (.L_HI(net271));
 sg13g2_tiehi \g.g_y[2].g_x[1].t.r_sc$_SDFF_PN0__272  (.L_HI(net272));
 sg13g2_tiehi \g.g_y[2].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_273  (.L_HI(net273));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_274  (.L_HI(net274));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_275  (.L_HI(net275));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_276  (.L_HI(net276));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_277  (.L_HI(net277));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_sc$_SDFF_PN0__278  (.L_HI(net278));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_279  (.L_HI(net279));
 sg13g2_tiehi \g.g_y[2].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_280  (.L_HI(net280));
 sg13g2_tiehi \g.g_y[2].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_281  (.L_HI(net281));
 sg13g2_tiehi \g.g_y[2].g_x[3].t.r_sc$_SDFF_PN0__282  (.L_HI(net282));
 sg13g2_tiehi \g.g_y[2].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_283  (.L_HI(net283));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_284  (.L_HI(net284));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_285  (.L_HI(net285));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_286  (.L_HI(net286));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_287  (.L_HI(net287));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_sc$_SDFF_PN0__288  (.L_HI(net288));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_289  (.L_HI(net289));
 sg13g2_tiehi \g.g_y[2].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_290  (.L_HI(net290));
 sg13g2_tiehi \g.g_y[2].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_291  (.L_HI(net291));
 sg13g2_tiehi \g.g_y[2].g_x[5].t.r_sc$_SDFF_PN0__292  (.L_HI(net292));
 sg13g2_tiehi \g.g_y[2].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_293  (.L_HI(net293));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_294  (.L_HI(net294));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_295  (.L_HI(net295));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_296  (.L_HI(net296));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_297  (.L_HI(net297));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_sc$_SDFF_PN0__298  (.L_HI(net298));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_299  (.L_HI(net299));
 sg13g2_tiehi \g.g_y[2].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_300  (.L_HI(net300));
 sg13g2_tiehi \g.g_y[2].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_301  (.L_HI(net301));
 sg13g2_tiehi \g.g_y[2].g_x[7].t.r_sc$_SDFF_PN0__302  (.L_HI(net302));
 sg13g2_tiehi \g.g_y[2].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_303  (.L_HI(net303));
 sg13g2_tiehi \g.g_y[3].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_304  (.L_HI(net304));
 sg13g2_tiehi \g.g_y[3].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_305  (.L_HI(net305));
 sg13g2_tiehi \g.g_y[3].g_x[0].t.r_sc$_SDFF_PN0__306  (.L_HI(net306));
 sg13g2_tiehi \g.g_y[3].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_307  (.L_HI(net307));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_308  (.L_HI(net308));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_309  (.L_HI(net309));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_310  (.L_HI(net310));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_311  (.L_HI(net311));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_sc$_SDFF_PN0__312  (.L_HI(net312));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_313  (.L_HI(net313));
 sg13g2_tiehi \g.g_y[3].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_314  (.L_HI(net314));
 sg13g2_tiehi \g.g_y[3].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_315  (.L_HI(net315));
 sg13g2_tiehi \g.g_y[3].g_x[2].t.r_sc$_SDFF_PN0__316  (.L_HI(net316));
 sg13g2_tiehi \g.g_y[3].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_317  (.L_HI(net317));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_318  (.L_HI(net318));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_319  (.L_HI(net319));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_320  (.L_HI(net320));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_321  (.L_HI(net321));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_sc$_SDFF_PN0__322  (.L_HI(net322));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_323  (.L_HI(net323));
 sg13g2_tiehi \g.g_y[3].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_324  (.L_HI(net324));
 sg13g2_tiehi \g.g_y[3].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_325  (.L_HI(net325));
 sg13g2_tiehi \g.g_y[3].g_x[4].t.r_sc$_SDFF_PN0__326  (.L_HI(net326));
 sg13g2_tiehi \g.g_y[3].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_327  (.L_HI(net327));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_328  (.L_HI(net328));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_329  (.L_HI(net329));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_330  (.L_HI(net330));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_331  (.L_HI(net331));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_sc$_SDFF_PN0__332  (.L_HI(net332));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_333  (.L_HI(net333));
 sg13g2_tiehi \g.g_y[3].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_334  (.L_HI(net334));
 sg13g2_tiehi \g.g_y[3].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_335  (.L_HI(net335));
 sg13g2_tiehi \g.g_y[3].g_x[6].t.r_sc$_SDFF_PN0__336  (.L_HI(net336));
 sg13g2_tiehi \g.g_y[3].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_337  (.L_HI(net337));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_338  (.L_HI(net338));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_339  (.L_HI(net339));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_340  (.L_HI(net340));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_341  (.L_HI(net341));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_sc$_SDFF_PN0__342  (.L_HI(net342));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_343  (.L_HI(net343));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_344  (.L_HI(net344));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_345  (.L_HI(net345));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_346  (.L_HI(net346));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_347  (.L_HI(net347));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_sc$_SDFF_PN0__348  (.L_HI(net348));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_349  (.L_HI(net349));
 sg13g2_tiehi \g.g_y[4].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_350  (.L_HI(net350));
 sg13g2_tiehi \g.g_y[4].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_351  (.L_HI(net351));
 sg13g2_tiehi \g.g_y[4].g_x[1].t.r_sc$_SDFF_PN0__352  (.L_HI(net352));
 sg13g2_tiehi \g.g_y[4].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_353  (.L_HI(net353));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_354  (.L_HI(net354));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_355  (.L_HI(net355));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_356  (.L_HI(net356));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_357  (.L_HI(net357));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_sc$_SDFF_PN0__358  (.L_HI(net358));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_359  (.L_HI(net359));
 sg13g2_tiehi \g.g_y[4].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_360  (.L_HI(net360));
 sg13g2_tiehi \g.g_y[4].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_361  (.L_HI(net361));
 sg13g2_tiehi \g.g_y[4].g_x[3].t.r_sc$_SDFF_PN0__362  (.L_HI(net362));
 sg13g2_tiehi \g.g_y[4].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_363  (.L_HI(net363));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_364  (.L_HI(net364));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_365  (.L_HI(net365));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_366  (.L_HI(net366));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_367  (.L_HI(net367));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_sc$_SDFF_PN0__368  (.L_HI(net368));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_369  (.L_HI(net369));
 sg13g2_tiehi \g.g_y[4].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_370  (.L_HI(net370));
 sg13g2_tiehi \g.g_y[4].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_371  (.L_HI(net371));
 sg13g2_tiehi \g.g_y[4].g_x[5].t.r_sc$_SDFF_PN0__372  (.L_HI(net372));
 sg13g2_tiehi \g.g_y[4].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_373  (.L_HI(net373));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_374  (.L_HI(net374));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_375  (.L_HI(net375));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_376  (.L_HI(net376));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_377  (.L_HI(net377));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_sc$_SDFF_PN0__378  (.L_HI(net378));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_379  (.L_HI(net379));
 sg13g2_tiehi \g.g_y[4].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_380  (.L_HI(net380));
 sg13g2_tiehi \g.g_y[4].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_381  (.L_HI(net381));
 sg13g2_tiehi \g.g_y[4].g_x[7].t.r_sc$_SDFF_PN0__382  (.L_HI(net382));
 sg13g2_tiehi \g.g_y[4].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_383  (.L_HI(net383));
 sg13g2_tiehi \g.g_y[5].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_384  (.L_HI(net384));
 sg13g2_tiehi \g.g_y[5].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_385  (.L_HI(net385));
 sg13g2_tiehi \g.g_y[5].g_x[0].t.r_sc$_SDFF_PN0__386  (.L_HI(net386));
 sg13g2_tiehi \g.g_y[5].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_387  (.L_HI(net387));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_388  (.L_HI(net388));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_389  (.L_HI(net389));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_390  (.L_HI(net390));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_391  (.L_HI(net391));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_sc$_SDFF_PN0__392  (.L_HI(net392));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_393  (.L_HI(net393));
 sg13g2_tiehi \g.g_y[5].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_394  (.L_HI(net394));
 sg13g2_tiehi \g.g_y[5].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_395  (.L_HI(net395));
 sg13g2_tiehi \g.g_y[5].g_x[2].t.r_sc$_SDFF_PN0__396  (.L_HI(net396));
 sg13g2_tiehi \g.g_y[5].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_397  (.L_HI(net397));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_398  (.L_HI(net398));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_399  (.L_HI(net399));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_400  (.L_HI(net400));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_401  (.L_HI(net401));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_sc$_SDFF_PN0__402  (.L_HI(net402));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_403  (.L_HI(net403));
 sg13g2_tiehi \g.g_y[5].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_404  (.L_HI(net404));
 sg13g2_tiehi \g.g_y[5].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_405  (.L_HI(net405));
 sg13g2_tiehi \g.g_y[5].g_x[4].t.r_sc$_SDFF_PN0__406  (.L_HI(net406));
 sg13g2_tiehi \g.g_y[5].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_407  (.L_HI(net407));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_408  (.L_HI(net408));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_409  (.L_HI(net409));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_410  (.L_HI(net410));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_411  (.L_HI(net411));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_sc$_SDFF_PN0__412  (.L_HI(net412));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_413  (.L_HI(net413));
 sg13g2_tiehi \g.g_y[5].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_414  (.L_HI(net414));
 sg13g2_tiehi \g.g_y[5].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_415  (.L_HI(net415));
 sg13g2_tiehi \g.g_y[5].g_x[6].t.r_sc$_SDFF_PN0__416  (.L_HI(net416));
 sg13g2_tiehi \g.g_y[5].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_417  (.L_HI(net417));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_418  (.L_HI(net418));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_419  (.L_HI(net419));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_420  (.L_HI(net420));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_421  (.L_HI(net421));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_sc$_SDFF_PN0__422  (.L_HI(net422));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_423  (.L_HI(net423));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_424  (.L_HI(net424));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_425  (.L_HI(net425));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_426  (.L_HI(net426));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_427  (.L_HI(net427));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_sc$_SDFF_PN0__428  (.L_HI(net428));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_429  (.L_HI(net429));
 sg13g2_tiehi \g.g_y[6].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_430  (.L_HI(net430));
 sg13g2_tiehi \g.g_y[6].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_431  (.L_HI(net431));
 sg13g2_tiehi \g.g_y[6].g_x[1].t.r_sc$_SDFF_PN0__432  (.L_HI(net432));
 sg13g2_tiehi \g.g_y[6].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_433  (.L_HI(net433));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_434  (.L_HI(net434));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_435  (.L_HI(net435));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_436  (.L_HI(net436));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_437  (.L_HI(net437));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_sc$_SDFF_PN0__438  (.L_HI(net438));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_439  (.L_HI(net439));
 sg13g2_tiehi \g.g_y[6].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_440  (.L_HI(net440));
 sg13g2_tiehi \g.g_y[6].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_441  (.L_HI(net441));
 sg13g2_tiehi \g.g_y[6].g_x[3].t.r_sc$_SDFF_PN0__442  (.L_HI(net442));
 sg13g2_tiehi \g.g_y[6].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_443  (.L_HI(net443));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_444  (.L_HI(net444));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_445  (.L_HI(net445));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_446  (.L_HI(net446));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_447  (.L_HI(net447));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_sc$_SDFF_PN0__448  (.L_HI(net448));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_449  (.L_HI(net449));
 sg13g2_tiehi \g.g_y[6].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_450  (.L_HI(net450));
 sg13g2_tiehi \g.g_y[6].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_451  (.L_HI(net451));
 sg13g2_tiehi \g.g_y[6].g_x[5].t.r_sc$_SDFF_PN0__452  (.L_HI(net452));
 sg13g2_tiehi \g.g_y[6].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_453  (.L_HI(net453));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_454  (.L_HI(net454));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_455  (.L_HI(net455));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_456  (.L_HI(net456));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_457  (.L_HI(net457));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_sc$_SDFF_PN0__458  (.L_HI(net458));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_459  (.L_HI(net459));
 sg13g2_tiehi \g.g_y[6].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_460  (.L_HI(net460));
 sg13g2_tiehi \g.g_y[6].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_461  (.L_HI(net461));
 sg13g2_tiehi \g.g_y[6].g_x[7].t.r_sc$_SDFF_PN0__462  (.L_HI(net462));
 sg13g2_tiehi \g.g_y[6].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_463  (.L_HI(net463));
 sg13g2_tiehi \g.g_y[7].g_x[0].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_464  (.L_HI(net464));
 sg13g2_tiehi \g.g_y[7].g_x[0].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_465  (.L_HI(net465));
 sg13g2_tiehi \g.g_y[7].g_x[0].t.r_sc$_SDFF_PN0__466  (.L_HI(net466));
 sg13g2_tiehi \g.g_y[7].g_x[0].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_467  (.L_HI(net467));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_468  (.L_HI(net468));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_469  (.L_HI(net469));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_470  (.L_HI(net470));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_471  (.L_HI(net471));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_sc$_SDFF_PN0__472  (.L_HI(net472));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_473  (.L_HI(net473));
 sg13g2_tiehi \g.g_y[7].g_x[2].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_474  (.L_HI(net474));
 sg13g2_tiehi \g.g_y[7].g_x[2].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_475  (.L_HI(net475));
 sg13g2_tiehi \g.g_y[7].g_x[2].t.r_sc$_SDFF_PN0__476  (.L_HI(net476));
 sg13g2_tiehi \g.g_y[7].g_x[2].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_477  (.L_HI(net477));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_478  (.L_HI(net478));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_479  (.L_HI(net479));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_480  (.L_HI(net480));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_481  (.L_HI(net481));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_sc$_SDFF_PN0__482  (.L_HI(net482));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_483  (.L_HI(net483));
 sg13g2_tiehi \g.g_y[7].g_x[4].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_484  (.L_HI(net484));
 sg13g2_tiehi \g.g_y[7].g_x[4].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_485  (.L_HI(net485));
 sg13g2_tiehi \g.g_y[7].g_x[4].t.r_sc$_SDFF_PN0__486  (.L_HI(net486));
 sg13g2_tiehi \g.g_y[7].g_x[4].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_487  (.L_HI(net487));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_488  (.L_HI(net488));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_489  (.L_HI(net489));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_490  (.L_HI(net490));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_491  (.L_HI(net491));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_sc$_SDFF_PN0__492  (.L_HI(net492));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_493  (.L_HI(net493));
 sg13g2_tiehi \g.g_y[7].g_x[6].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_494  (.L_HI(net494));
 sg13g2_tiehi \g.g_y[7].g_x[6].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_495  (.L_HI(net495));
 sg13g2_tiehi \g.g_y[7].g_x[6].t.r_sc$_SDFF_PN0__496  (.L_HI(net496));
 sg13g2_tiehi \g.g_y[7].g_x[6].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_497  (.L_HI(net497));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_d$_DLATCH_N_._TECHMAP_DLATCH_N_498  (.L_HI(net498));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_499  (.L_HI(net499));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_500  (.L_HI(net500));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_h$_DLATCH_N_._TECHMAP_DLATCH_N_501  (.L_HI(net501));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_sc$_SDFF_PN0__502  (.L_HI(net502));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_v$_DLATCH_N_._TECHMAP_DLATCH_N_503  (.L_HI(net503));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_fill_1 FILLER_0_147 ();
 sg13g2_fill_1 FILLER_0_153 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_fill_2 FILLER_0_179 ();
 sg13g2_fill_1 FILLER_0_181 ();
 sg13g2_decap_4 FILLER_0_210 ();
 sg13g2_fill_1 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_decap_8 FILLER_0_237 ();
 sg13g2_decap_8 FILLER_0_244 ();
 sg13g2_decap_8 FILLER_0_251 ();
 sg13g2_decap_8 FILLER_0_258 ();
 sg13g2_decap_8 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_272 ();
 sg13g2_decap_8 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_311 ();
 sg13g2_decap_8 FILLER_0_318 ();
 sg13g2_decap_8 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_0_409 ();
 sg13g2_decap_8 FILLER_0_416 ();
 sg13g2_decap_8 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_fill_2 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_125 ();
 sg13g2_decap_8 FILLER_1_132 ();
 sg13g2_fill_2 FILLER_1_139 ();
 sg13g2_fill_1 FILLER_1_170 ();
 sg13g2_fill_1 FILLER_1_181 ();
 sg13g2_fill_2 FILLER_1_186 ();
 sg13g2_fill_1 FILLER_1_204 ();
 sg13g2_fill_2 FILLER_1_210 ();
 sg13g2_fill_1 FILLER_1_228 ();
 sg13g2_decap_4 FILLER_1_239 ();
 sg13g2_decap_8 FILLER_1_251 ();
 sg13g2_decap_8 FILLER_1_258 ();
 sg13g2_decap_8 FILLER_1_265 ();
 sg13g2_decap_8 FILLER_1_272 ();
 sg13g2_decap_4 FILLER_1_279 ();
 sg13g2_decap_8 FILLER_1_303 ();
 sg13g2_fill_1 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_4 FILLER_2_128 ();
 sg13g2_fill_1 FILLER_2_152 ();
 sg13g2_decap_4 FILLER_2_212 ();
 sg13g2_fill_1 FILLER_2_216 ();
 sg13g2_fill_2 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_decap_8 FILLER_2_272 ();
 sg13g2_decap_4 FILLER_2_279 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_8 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_2_412 ();
 sg13g2_decap_8 FILLER_2_419 ();
 sg13g2_decap_4 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_4 FILLER_3_140 ();
 sg13g2_fill_2 FILLER_3_144 ();
 sg13g2_fill_2 FILLER_3_150 ();
 sg13g2_fill_1 FILLER_3_152 ();
 sg13g2_fill_1 FILLER_3_213 ();
 sg13g2_fill_1 FILLER_3_229 ();
 sg13g2_decap_8 FILLER_3_246 ();
 sg13g2_decap_4 FILLER_3_253 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_fill_2 FILLER_3_268 ();
 sg13g2_decap_4 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_278 ();
 sg13g2_fill_2 FILLER_3_305 ();
 sg13g2_fill_1 FILLER_3_307 ();
 sg13g2_decap_4 FILLER_3_313 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_fill_1 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_4 FILLER_4_133 ();
 sg13g2_fill_1 FILLER_4_137 ();
 sg13g2_fill_1 FILLER_4_166 ();
 sg13g2_fill_2 FILLER_4_177 ();
 sg13g2_fill_1 FILLER_4_199 ();
 sg13g2_fill_1 FILLER_4_230 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_fill_2 FILLER_4_252 ();
 sg13g2_fill_2 FILLER_4_279 ();
 sg13g2_decap_4 FILLER_4_316 ();
 sg13g2_fill_2 FILLER_4_320 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_130 ();
 sg13g2_fill_2 FILLER_5_151 ();
 sg13g2_fill_1 FILLER_5_153 ();
 sg13g2_fill_1 FILLER_5_174 ();
 sg13g2_fill_2 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_184 ();
 sg13g2_fill_2 FILLER_5_206 ();
 sg13g2_fill_1 FILLER_5_233 ();
 sg13g2_fill_1 FILLER_5_258 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_fill_1 FILLER_5_296 ();
 sg13g2_fill_1 FILLER_5_312 ();
 sg13g2_decap_4 FILLER_5_339 ();
 sg13g2_fill_2 FILLER_5_363 ();
 sg13g2_fill_1 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_8 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_5_412 ();
 sg13g2_decap_8 FILLER_5_419 ();
 sg13g2_decap_4 FILLER_5_426 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_4 FILLER_6_105 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_fill_1 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_142 ();
 sg13g2_fill_1 FILLER_6_144 ();
 sg13g2_fill_1 FILLER_6_165 ();
 sg13g2_fill_1 FILLER_6_188 ();
 sg13g2_fill_1 FILLER_6_205 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_fill_1 FILLER_6_216 ();
 sg13g2_fill_1 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_249 ();
 sg13g2_fill_2 FILLER_6_269 ();
 sg13g2_fill_2 FILLER_6_299 ();
 sg13g2_fill_1 FILLER_6_301 ();
 sg13g2_fill_1 FILLER_6_313 ();
 sg13g2_fill_1 FILLER_6_319 ();
 sg13g2_fill_2 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_8 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_411 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_decap_4 FILLER_6_425 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_4 FILLER_7_98 ();
 sg13g2_fill_2 FILLER_7_122 ();
 sg13g2_fill_1 FILLER_7_136 ();
 sg13g2_fill_2 FILLER_7_149 ();
 sg13g2_fill_2 FILLER_7_155 ();
 sg13g2_fill_1 FILLER_7_157 ();
 sg13g2_fill_2 FILLER_7_163 ();
 sg13g2_fill_2 FILLER_7_170 ();
 sg13g2_fill_1 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_210 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_fill_2 FILLER_7_250 ();
 sg13g2_fill_1 FILLER_7_252 ();
 sg13g2_fill_2 FILLER_7_256 ();
 sg13g2_fill_1 FILLER_7_258 ();
 sg13g2_decap_8 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_271 ();
 sg13g2_fill_1 FILLER_7_311 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_fill_1 FILLER_7_323 ();
 sg13g2_fill_1 FILLER_7_329 ();
 sg13g2_fill_1 FILLER_7_334 ();
 sg13g2_fill_1 FILLER_7_340 ();
 sg13g2_fill_2 FILLER_7_346 ();
 sg13g2_fill_2 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_fill_1 FILLER_8_105 ();
 sg13g2_fill_2 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_160 ();
 sg13g2_fill_1 FILLER_8_162 ();
 sg13g2_fill_1 FILLER_8_183 ();
 sg13g2_decap_8 FILLER_8_188 ();
 sg13g2_fill_2 FILLER_8_195 ();
 sg13g2_fill_1 FILLER_8_197 ();
 sg13g2_decap_8 FILLER_8_202 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_decap_4 FILLER_8_216 ();
 sg13g2_fill_2 FILLER_8_229 ();
 sg13g2_fill_2 FILLER_8_268 ();
 sg13g2_decap_4 FILLER_8_278 ();
 sg13g2_fill_1 FILLER_8_290 ();
 sg13g2_fill_1 FILLER_8_296 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_338 ();
 sg13g2_fill_1 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_8 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_8_412 ();
 sg13g2_decap_8 FILLER_8_419 ();
 sg13g2_decap_4 FILLER_8_426 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_4 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_109 ();
 sg13g2_fill_2 FILLER_9_175 ();
 sg13g2_fill_1 FILLER_9_177 ();
 sg13g2_fill_2 FILLER_9_182 ();
 sg13g2_decap_4 FILLER_9_188 ();
 sg13g2_decap_4 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_fill_1 FILLER_9_234 ();
 sg13g2_fill_1 FILLER_9_240 ();
 sg13g2_fill_1 FILLER_9_263 ();
 sg13g2_decap_4 FILLER_9_280 ();
 sg13g2_fill_1 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_decap_8 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_9_414 ();
 sg13g2_decap_8 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_fill_1 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_132 ();
 sg13g2_fill_1 FILLER_10_141 ();
 sg13g2_fill_1 FILLER_10_151 ();
 sg13g2_fill_2 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_200 ();
 sg13g2_fill_2 FILLER_10_228 ();
 sg13g2_fill_2 FILLER_10_246 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_301 ();
 sg13g2_fill_2 FILLER_10_331 ();
 sg13g2_fill_2 FILLER_10_339 ();
 sg13g2_fill_1 FILLER_10_366 ();
 sg13g2_fill_2 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_4 FILLER_11_112 ();
 sg13g2_fill_1 FILLER_11_152 ();
 sg13g2_fill_1 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_fill_1 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_185 ();
 sg13g2_fill_2 FILLER_11_203 ();
 sg13g2_fill_1 FILLER_11_205 ();
 sg13g2_fill_2 FILLER_11_226 ();
 sg13g2_fill_1 FILLER_11_266 ();
 sg13g2_decap_4 FILLER_11_272 ();
 sg13g2_fill_1 FILLER_11_319 ();
 sg13g2_fill_2 FILLER_11_331 ();
 sg13g2_fill_1 FILLER_11_361 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_decap_8 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_421 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_fill_1 FILLER_12_119 ();
 sg13g2_fill_1 FILLER_12_159 ();
 sg13g2_fill_1 FILLER_12_170 ();
 sg13g2_fill_2 FILLER_12_202 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_fill_2 FILLER_12_225 ();
 sg13g2_fill_1 FILLER_12_227 ();
 sg13g2_fill_1 FILLER_12_254 ();
 sg13g2_fill_1 FILLER_12_260 ();
 sg13g2_decap_4 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_fill_2 FILLER_12_328 ();
 sg13g2_fill_2 FILLER_12_355 ();
 sg13g2_fill_1 FILLER_12_357 ();
 sg13g2_decap_4 FILLER_12_384 ();
 sg13g2_fill_2 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_decap_8 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_fill_1 FILLER_13_81 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_1 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_127 ();
 sg13g2_fill_2 FILLER_13_174 ();
 sg13g2_decap_4 FILLER_13_190 ();
 sg13g2_fill_2 FILLER_13_194 ();
 sg13g2_fill_2 FILLER_13_214 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_2 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_fill_1 FILLER_13_238 ();
 sg13g2_fill_1 FILLER_13_249 ();
 sg13g2_decap_4 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_fill_2 FILLER_13_301 ();
 sg13g2_fill_1 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_fill_2 FILLER_13_315 ();
 sg13g2_fill_1 FILLER_13_322 ();
 sg13g2_fill_1 FILLER_13_328 ();
 sg13g2_fill_2 FILLER_13_336 ();
 sg13g2_fill_2 FILLER_13_347 ();
 sg13g2_fill_2 FILLER_13_358 ();
 sg13g2_fill_1 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_4 FILLER_13_377 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_decap_4 FILLER_13_402 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_8 FILLER_13_419 ();
 sg13g2_decap_4 FILLER_13_426 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_fill_2 FILLER_14_70 ();
 sg13g2_fill_2 FILLER_14_88 ();
 sg13g2_fill_1 FILLER_14_90 ();
 sg13g2_fill_2 FILLER_14_107 ();
 sg13g2_fill_1 FILLER_14_109 ();
 sg13g2_fill_1 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_161 ();
 sg13g2_fill_1 FILLER_14_166 ();
 sg13g2_fill_1 FILLER_14_229 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_240 ();
 sg13g2_fill_2 FILLER_14_259 ();
 sg13g2_fill_1 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_fill_1 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_fill_2 FILLER_14_365 ();
 sg13g2_fill_1 FILLER_14_367 ();
 sg13g2_decap_4 FILLER_14_372 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_418 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_4 FILLER_15_63 ();
 sg13g2_fill_1 FILLER_15_108 ();
 sg13g2_fill_2 FILLER_15_115 ();
 sg13g2_fill_1 FILLER_15_129 ();
 sg13g2_fill_1 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_2 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_fill_2 FILLER_15_188 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_fill_1 FILLER_15_234 ();
 sg13g2_fill_2 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_fill_1 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_4 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_fill_1 FILLER_16_88 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_101 ();
 sg13g2_fill_2 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_134 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_2 FILLER_16_172 ();
 sg13g2_fill_1 FILLER_16_179 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_fill_2 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_262 ();
 sg13g2_fill_1 FILLER_16_286 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_fill_2 FILLER_16_298 ();
 sg13g2_fill_1 FILLER_16_316 ();
 sg13g2_fill_1 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_fill_1 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_384 ();
 sg13g2_fill_1 FILLER_16_389 ();
 sg13g2_fill_2 FILLER_16_411 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_4 FILLER_16_424 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_fill_2 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_77 ();
 sg13g2_fill_1 FILLER_17_79 ();
 sg13g2_fill_2 FILLER_17_85 ();
 sg13g2_fill_2 FILLER_17_108 ();
 sg13g2_decap_8 FILLER_17_138 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_decap_4 FILLER_17_152 ();
 sg13g2_fill_2 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_200 ();
 sg13g2_fill_2 FILLER_17_217 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_decap_4 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_2 FILLER_17_245 ();
 sg13g2_fill_1 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_304 ();
 sg13g2_decap_4 FILLER_17_314 ();
 sg13g2_fill_2 FILLER_17_334 ();
 sg13g2_fill_1 FILLER_17_394 ();
 sg13g2_fill_2 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_418 ();
 sg13g2_decap_4 FILLER_17_425 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_4 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_78 ();
 sg13g2_decap_4 FILLER_18_85 ();
 sg13g2_fill_1 FILLER_18_89 ();
 sg13g2_fill_1 FILLER_18_100 ();
 sg13g2_fill_2 FILLER_18_106 ();
 sg13g2_fill_1 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_118 ();
 sg13g2_fill_2 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_181 ();
 sg13g2_decap_8 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_218 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_232 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_fill_1 FILLER_18_314 ();
 sg13g2_fill_1 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_fill_2 FILLER_18_360 ();
 sg13g2_fill_1 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_405 ();
 sg13g2_decap_4 FILLER_18_425 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_96 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_153 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_decap_4 FILLER_19_163 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_decap_4 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_decap_4 FILLER_19_186 ();
 sg13g2_fill_2 FILLER_19_190 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_decap_8 FILLER_19_199 ();
 sg13g2_fill_2 FILLER_19_206 ();
 sg13g2_fill_1 FILLER_19_208 ();
 sg13g2_fill_1 FILLER_19_219 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_fill_1 FILLER_19_325 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_decap_4 FILLER_19_363 ();
 sg13g2_fill_1 FILLER_19_392 ();
 sg13g2_decap_4 FILLER_19_397 ();
 sg13g2_decap_8 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_19_412 ();
 sg13g2_decap_8 FILLER_19_419 ();
 sg13g2_decap_4 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_fill_2 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_127 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_decap_4 FILLER_20_161 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_262 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_fill_1 FILLER_20_294 ();
 sg13g2_fill_1 FILLER_20_300 ();
 sg13g2_fill_2 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_331 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_fill_2 FILLER_20_363 ();
 sg13g2_fill_1 FILLER_20_365 ();
 sg13g2_fill_2 FILLER_20_400 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_4 FILLER_21_104 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_fill_2 FILLER_21_117 ();
 sg13g2_fill_1 FILLER_21_119 ();
 sg13g2_fill_2 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_171 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_decap_4 FILLER_21_207 ();
 sg13g2_decap_4 FILLER_21_225 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_fill_1 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_291 ();
 sg13g2_fill_1 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_decap_4 FILLER_21_329 ();
 sg13g2_decap_4 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_342 ();
 sg13g2_decap_4 FILLER_21_353 ();
 sg13g2_fill_1 FILLER_21_357 ();
 sg13g2_fill_1 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_414 ();
 sg13g2_decap_8 FILLER_21_421 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_fill_1 FILLER_22_95 ();
 sg13g2_fill_1 FILLER_22_103 ();
 sg13g2_decap_4 FILLER_22_113 ();
 sg13g2_fill_2 FILLER_22_122 ();
 sg13g2_decap_4 FILLER_22_153 ();
 sg13g2_fill_2 FILLER_22_165 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_fill_1 FILLER_22_216 ();
 sg13g2_decap_4 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_fill_2 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_4 FILLER_22_424 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_87 ();
 sg13g2_fill_1 FILLER_23_92 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_fill_2 FILLER_23_114 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_122 ();
 sg13g2_fill_2 FILLER_23_129 ();
 sg13g2_decap_4 FILLER_23_145 ();
 sg13g2_fill_2 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_fill_2 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_370 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_23_418 ();
 sg13g2_decap_4 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_4 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_90 ();
 sg13g2_fill_1 FILLER_24_141 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_187 ();
 sg13g2_fill_1 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_248 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_fill_2 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_342 ();
 sg13g2_decap_4 FILLER_24_348 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_24_392 ();
 sg13g2_fill_2 FILLER_24_409 ();
 sg13g2_fill_1 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_416 ();
 sg13g2_decap_8 FILLER_24_423 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_4 FILLER_25_63 ();
 sg13g2_fill_2 FILLER_25_72 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_136 ();
 sg13g2_decap_4 FILLER_25_141 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_206 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_314 ();
 sg13g2_fill_1 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_333 ();
 sg13g2_fill_2 FILLER_25_351 ();
 sg13g2_fill_2 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_decap_4 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_416 ();
 sg13g2_decap_8 FILLER_25_423 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_106 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_194 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_205 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_228 ();
 sg13g2_fill_1 FILLER_26_230 ();
 sg13g2_fill_2 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_decap_4 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_300 ();
 sg13g2_decap_4 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_67 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_83 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_fill_2 FILLER_27_99 ();
 sg13g2_decap_8 FILLER_27_107 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_fill_2 FILLER_27_153 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_fill_2 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_247 ();
 sg13g2_decap_8 FILLER_27_254 ();
 sg13g2_decap_4 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_345 ();
 sg13g2_fill_2 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_27_411 ();
 sg13g2_decap_8 FILLER_27_418 ();
 sg13g2_decap_4 FILLER_27_425 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_fill_2 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_58 ();
 sg13g2_fill_1 FILLER_28_82 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_decap_4 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_116 ();
 sg13g2_fill_1 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_164 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_190 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_259 ();
 sg13g2_decap_4 FILLER_28_264 ();
 sg13g2_fill_1 FILLER_28_268 ();
 sg13g2_decap_4 FILLER_28_281 ();
 sg13g2_decap_4 FILLER_28_289 ();
 sg13g2_fill_1 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_2 FILLER_28_374 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_404 ();
 sg13g2_decap_8 FILLER_28_411 ();
 sg13g2_decap_8 FILLER_28_418 ();
 sg13g2_decap_4 FILLER_28_425 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_75 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_2 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_2 FILLER_29_196 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_350 ();
 sg13g2_fill_2 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_409 ();
 sg13g2_decap_8 FILLER_29_416 ();
 sg13g2_decap_8 FILLER_29_423 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_58 ();
 sg13g2_fill_2 FILLER_30_79 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_decap_8 FILLER_30_103 ();
 sg13g2_decap_4 FILLER_30_110 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_2 FILLER_30_120 ();
 sg13g2_fill_1 FILLER_30_127 ();
 sg13g2_fill_1 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_314 ();
 sg13g2_fill_2 FILLER_30_319 ();
 sg13g2_decap_4 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_342 ();
 sg13g2_fill_1 FILLER_30_375 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_8 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_30_412 ();
 sg13g2_decap_8 FILLER_30_419 ();
 sg13g2_decap_4 FILLER_30_426 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_fill_1 FILLER_31_78 ();
 sg13g2_fill_2 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_366 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_fill_2 FILLER_32_78 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_fill_2 FILLER_32_101 ();
 sg13g2_fill_2 FILLER_32_108 ();
 sg13g2_fill_1 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_145 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_decap_4 FILLER_32_251 ();
 sg13g2_decap_4 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_318 ();
 sg13g2_fill_2 FILLER_32_332 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_388 ();
 sg13g2_fill_2 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_decap_4 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_decap_8 FILLER_33_144 ();
 sg13g2_decap_4 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_187 ();
 sg13g2_decap_4 FILLER_33_194 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_fill_2 FILLER_33_209 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_decap_4 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_286 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_364 ();
 sg13g2_fill_2 FILLER_33_369 ();
 sg13g2_fill_1 FILLER_33_380 ();
 sg13g2_fill_2 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_33_400 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_60 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_decap_4 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_146 ();
 sg13g2_decap_4 FILLER_34_153 ();
 sg13g2_decap_8 FILLER_34_181 ();
 sg13g2_decap_8 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_211 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_312 ();
 sg13g2_decap_4 FILLER_34_412 ();
 sg13g2_decap_4 FILLER_34_425 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_81 ();
 sg13g2_fill_1 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_103 ();
 sg13g2_fill_1 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_115 ();
 sg13g2_fill_2 FILLER_35_122 ();
 sg13g2_fill_2 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_162 ();
 sg13g2_fill_2 FILLER_35_169 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_212 ();
 sg13g2_fill_1 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_223 ();
 sg13g2_fill_1 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_2 FILLER_35_269 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_fill_2 FILLER_35_315 ();
 sg13g2_fill_1 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_fill_1 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_406 ();
 sg13g2_fill_2 FILLER_35_427 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_92 ();
 sg13g2_fill_1 FILLER_36_94 ();
 sg13g2_fill_2 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_163 ();
 sg13g2_fill_1 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_decap_4 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_decap_8 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_407 ();
 sg13g2_fill_1 FILLER_36_424 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_78 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_133 ();
 sg13g2_fill_2 FILLER_37_203 ();
 sg13g2_fill_2 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_281 ();
 sg13g2_decap_4 FILLER_37_286 ();
 sg13g2_fill_1 FILLER_37_307 ();
 sg13g2_fill_2 FILLER_37_314 ();
 sg13g2_fill_1 FILLER_37_321 ();
 sg13g2_fill_1 FILLER_37_353 ();
 sg13g2_fill_2 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_372 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_4 FILLER_38_63 ();
 sg13g2_fill_1 FILLER_38_67 ();
 sg13g2_decap_8 FILLER_38_72 ();
 sg13g2_decap_4 FILLER_38_79 ();
 sg13g2_fill_1 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_89 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_101 ();
 sg13g2_fill_1 FILLER_38_118 ();
 sg13g2_fill_1 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_128 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_163 ();
 sg13g2_fill_1 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_413 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_4 FILLER_39_63 ();
 sg13g2_fill_2 FILLER_39_67 ();
 sg13g2_fill_1 FILLER_39_81 ();
 sg13g2_fill_1 FILLER_39_90 ();
 sg13g2_fill_2 FILLER_39_105 ();
 sg13g2_fill_1 FILLER_39_123 ();
 sg13g2_fill_2 FILLER_39_128 ();
 sg13g2_fill_2 FILLER_39_153 ();
 sg13g2_fill_1 FILLER_39_155 ();
 sg13g2_decap_4 FILLER_39_160 ();
 sg13g2_fill_2 FILLER_39_164 ();
 sg13g2_fill_1 FILLER_39_239 ();
 sg13g2_fill_1 FILLER_39_257 ();
 sg13g2_fill_1 FILLER_39_264 ();
 sg13g2_fill_1 FILLER_39_275 ();
 sg13g2_fill_2 FILLER_39_291 ();
 sg13g2_fill_1 FILLER_39_366 ();
 sg13g2_decap_8 FILLER_39_381 ();
 sg13g2_fill_2 FILLER_39_388 ();
 sg13g2_fill_1 FILLER_39_390 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_fill_1 FILLER_40_56 ();
 sg13g2_fill_1 FILLER_40_83 ();
 sg13g2_fill_1 FILLER_40_92 ();
 sg13g2_fill_1 FILLER_40_100 ();
 sg13g2_fill_1 FILLER_40_117 ();
 sg13g2_fill_1 FILLER_40_123 ();
 sg13g2_fill_2 FILLER_40_137 ();
 sg13g2_decap_4 FILLER_40_146 ();
 sg13g2_decap_4 FILLER_40_176 ();
 sg13g2_fill_2 FILLER_40_180 ();
 sg13g2_fill_2 FILLER_40_189 ();
 sg13g2_fill_1 FILLER_40_191 ();
 sg13g2_decap_4 FILLER_40_226 ();
 sg13g2_fill_1 FILLER_40_230 ();
 sg13g2_decap_8 FILLER_40_241 ();
 sg13g2_fill_1 FILLER_40_248 ();
 sg13g2_fill_1 FILLER_40_254 ();
 sg13g2_fill_2 FILLER_40_260 ();
 sg13g2_fill_1 FILLER_40_262 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_4 FILLER_40_273 ();
 sg13g2_fill_2 FILLER_40_277 ();
 sg13g2_fill_1 FILLER_40_282 ();
 sg13g2_fill_1 FILLER_40_316 ();
 sg13g2_decap_4 FILLER_40_359 ();
 sg13g2_fill_1 FILLER_40_363 ();
 sg13g2_decap_8 FILLER_40_380 ();
 sg13g2_decap_4 FILLER_40_407 ();
 sg13g2_fill_1 FILLER_40_411 ();
 sg13g2_decap_4 FILLER_40_426 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_fill_1 FILLER_41_63 ();
 sg13g2_fill_1 FILLER_41_68 ();
 sg13g2_decap_8 FILLER_41_73 ();
 sg13g2_decap_4 FILLER_41_102 ();
 sg13g2_fill_1 FILLER_41_106 ();
 sg13g2_fill_1 FILLER_41_112 ();
 sg13g2_fill_2 FILLER_41_117 ();
 sg13g2_fill_1 FILLER_41_132 ();
 sg13g2_fill_1 FILLER_41_159 ();
 sg13g2_decap_8 FILLER_41_164 ();
 sg13g2_fill_1 FILLER_41_171 ();
 sg13g2_decap_4 FILLER_41_185 ();
 sg13g2_decap_8 FILLER_41_205 ();
 sg13g2_decap_8 FILLER_41_212 ();
 sg13g2_fill_2 FILLER_41_219 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_fill_2 FILLER_41_238 ();
 sg13g2_fill_1 FILLER_41_240 ();
 sg13g2_decap_8 FILLER_41_264 ();
 sg13g2_decap_8 FILLER_41_271 ();
 sg13g2_fill_2 FILLER_41_278 ();
 sg13g2_fill_1 FILLER_41_280 ();
 sg13g2_decap_4 FILLER_41_290 ();
 sg13g2_fill_1 FILLER_41_294 ();
 sg13g2_fill_1 FILLER_41_300 ();
 sg13g2_fill_2 FILLER_41_305 ();
 sg13g2_fill_2 FILLER_41_311 ();
 sg13g2_fill_2 FILLER_41_318 ();
 sg13g2_fill_2 FILLER_41_325 ();
 sg13g2_fill_1 FILLER_41_327 ();
 sg13g2_decap_4 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_347 ();
 sg13g2_decap_8 FILLER_41_352 ();
 sg13g2_decap_4 FILLER_41_359 ();
 sg13g2_fill_1 FILLER_41_363 ();
 sg13g2_fill_1 FILLER_41_373 ();
 sg13g2_fill_1 FILLER_41_384 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_fill_2 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_106 ();
 sg13g2_decap_8 FILLER_42_113 ();
 sg13g2_fill_1 FILLER_42_120 ();
 sg13g2_fill_1 FILLER_42_125 ();
 sg13g2_decap_8 FILLER_42_145 ();
 sg13g2_decap_8 FILLER_42_152 ();
 sg13g2_decap_8 FILLER_42_159 ();
 sg13g2_fill_2 FILLER_42_166 ();
 sg13g2_fill_2 FILLER_42_173 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_fill_2 FILLER_42_189 ();
 sg13g2_fill_2 FILLER_42_215 ();
 sg13g2_fill_1 FILLER_42_217 ();
 sg13g2_fill_2 FILLER_42_238 ();
 sg13g2_decap_4 FILLER_42_266 ();
 sg13g2_fill_1 FILLER_42_270 ();
 sg13g2_fill_1 FILLER_42_319 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_355 ();
 sg13g2_fill_1 FILLER_42_362 ();
 sg13g2_fill_1 FILLER_42_373 ();
 sg13g2_fill_2 FILLER_42_384 ();
 sg13g2_fill_1 FILLER_42_391 ();
 sg13g2_fill_2 FILLER_42_397 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_fill_2 FILLER_43_56 ();
 sg13g2_fill_1 FILLER_43_58 ();
 sg13g2_fill_1 FILLER_43_80 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_4 FILLER_43_112 ();
 sg13g2_fill_1 FILLER_43_116 ();
 sg13g2_fill_1 FILLER_43_121 ();
 sg13g2_fill_2 FILLER_43_132 ();
 sg13g2_fill_1 FILLER_43_134 ();
 sg13g2_fill_1 FILLER_43_145 ();
 sg13g2_decap_4 FILLER_43_186 ();
 sg13g2_fill_1 FILLER_43_190 ();
 sg13g2_fill_1 FILLER_43_209 ();
 sg13g2_fill_2 FILLER_43_214 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_fill_2 FILLER_43_250 ();
 sg13g2_fill_1 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_257 ();
 sg13g2_fill_2 FILLER_43_268 ();
 sg13g2_decap_4 FILLER_43_344 ();
 sg13g2_fill_1 FILLER_43_369 ();
 sg13g2_decap_8 FILLER_43_373 ();
 sg13g2_fill_1 FILLER_43_380 ();
 sg13g2_fill_1 FILLER_43_386 ();
 sg13g2_fill_1 FILLER_43_391 ();
 sg13g2_fill_1 FILLER_43_397 ();
 sg13g2_fill_2 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_fill_2 FILLER_44_56 ();
 sg13g2_fill_2 FILLER_44_78 ();
 sg13g2_fill_1 FILLER_44_90 ();
 sg13g2_fill_1 FILLER_44_102 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_fill_1 FILLER_44_140 ();
 sg13g2_fill_2 FILLER_44_172 ();
 sg13g2_fill_1 FILLER_44_179 ();
 sg13g2_decap_4 FILLER_44_197 ();
 sg13g2_fill_1 FILLER_44_201 ();
 sg13g2_fill_1 FILLER_44_218 ();
 sg13g2_fill_2 FILLER_44_223 ();
 sg13g2_fill_2 FILLER_44_304 ();
 sg13g2_fill_1 FILLER_44_319 ();
 sg13g2_fill_2 FILLER_44_345 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_44_364 ();
 sg13g2_fill_2 FILLER_44_380 ();
 sg13g2_fill_1 FILLER_44_382 ();
 sg13g2_fill_2 FILLER_44_388 ();
 sg13g2_fill_1 FILLER_44_390 ();
 sg13g2_fill_1 FILLER_44_398 ();
 sg13g2_fill_2 FILLER_44_414 ();
 sg13g2_fill_1 FILLER_44_416 ();
 sg13g2_fill_2 FILLER_44_420 ();
 sg13g2_decap_4 FILLER_44_426 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_4 FILLER_45_63 ();
 sg13g2_fill_1 FILLER_45_67 ();
 sg13g2_decap_4 FILLER_45_72 ();
 sg13g2_fill_2 FILLER_45_100 ();
 sg13g2_fill_1 FILLER_45_102 ();
 sg13g2_fill_1 FILLER_45_123 ();
 sg13g2_fill_1 FILLER_45_129 ();
 sg13g2_fill_1 FILLER_45_144 ();
 sg13g2_fill_2 FILLER_45_150 ();
 sg13g2_fill_1 FILLER_45_152 ();
 sg13g2_fill_1 FILLER_45_167 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_188 ();
 sg13g2_fill_1 FILLER_45_194 ();
 sg13g2_fill_2 FILLER_45_205 ();
 sg13g2_fill_2 FILLER_45_212 ();
 sg13g2_fill_2 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_245 ();
 sg13g2_fill_2 FILLER_45_252 ();
 sg13g2_fill_2 FILLER_45_267 ();
 sg13g2_fill_1 FILLER_45_269 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_4 FILLER_45_287 ();
 sg13g2_fill_1 FILLER_45_291 ();
 sg13g2_decap_4 FILLER_45_297 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_fill_1 FILLER_45_320 ();
 sg13g2_decap_4 FILLER_45_325 ();
 sg13g2_decap_4 FILLER_45_362 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_fill_1 FILLER_45_389 ();
 sg13g2_fill_2 FILLER_45_395 ();
 sg13g2_fill_2 FILLER_45_412 ();
 sg13g2_decap_8 FILLER_45_419 ();
 sg13g2_decap_4 FILLER_45_426 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_4 FILLER_46_70 ();
 sg13g2_fill_2 FILLER_46_74 ();
 sg13g2_fill_1 FILLER_46_113 ();
 sg13g2_fill_2 FILLER_46_162 ();
 sg13g2_fill_1 FILLER_46_277 ();
 sg13g2_decap_4 FILLER_46_288 ();
 sg13g2_fill_2 FILLER_46_292 ();
 sg13g2_fill_2 FILLER_46_309 ();
 sg13g2_decap_4 FILLER_46_327 ();
 sg13g2_fill_1 FILLER_46_335 ();
 sg13g2_fill_1 FILLER_46_357 ();
 sg13g2_fill_1 FILLER_46_362 ();
 sg13g2_fill_1 FILLER_46_373 ();
 sg13g2_fill_2 FILLER_46_409 ();
 sg13g2_fill_1 FILLER_46_411 ();
 sg13g2_fill_1 FILLER_46_417 ();
 sg13g2_decap_8 FILLER_46_423 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_fill_2 FILLER_47_70 ();
 sg13g2_fill_1 FILLER_47_72 ();
 sg13g2_decap_4 FILLER_47_87 ();
 sg13g2_fill_1 FILLER_47_122 ();
 sg13g2_fill_2 FILLER_47_133 ();
 sg13g2_fill_1 FILLER_47_139 ();
 sg13g2_fill_1 FILLER_47_145 ();
 sg13g2_fill_1 FILLER_47_181 ();
 sg13g2_fill_1 FILLER_47_191 ();
 sg13g2_fill_1 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_202 ();
 sg13g2_decap_8 FILLER_47_213 ();
 sg13g2_fill_1 FILLER_47_228 ();
 sg13g2_fill_1 FILLER_47_233 ();
 sg13g2_fill_2 FILLER_47_261 ();
 sg13g2_fill_1 FILLER_47_268 ();
 sg13g2_fill_1 FILLER_47_275 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_286 ();
 sg13g2_fill_2 FILLER_47_293 ();
 sg13g2_decap_4 FILLER_47_300 ();
 sg13g2_fill_1 FILLER_47_304 ();
 sg13g2_fill_2 FILLER_47_350 ();
 sg13g2_fill_1 FILLER_47_352 ();
 sg13g2_fill_1 FILLER_47_358 ();
 sg13g2_fill_2 FILLER_47_427 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_4 FILLER_48_70 ();
 sg13g2_fill_2 FILLER_48_74 ();
 sg13g2_decap_4 FILLER_48_104 ();
 sg13g2_fill_1 FILLER_48_108 ();
 sg13g2_fill_1 FILLER_48_117 ();
 sg13g2_fill_1 FILLER_48_123 ();
 sg13g2_fill_1 FILLER_48_129 ();
 sg13g2_fill_1 FILLER_48_135 ();
 sg13g2_fill_1 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_4 FILLER_48_196 ();
 sg13g2_fill_1 FILLER_48_200 ();
 sg13g2_fill_2 FILLER_48_204 ();
 sg13g2_fill_1 FILLER_48_206 ();
 sg13g2_fill_1 FILLER_48_286 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_fill_1 FILLER_48_301 ();
 sg13g2_fill_2 FILLER_48_341 ();
 sg13g2_fill_2 FILLER_48_411 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_4 FILLER_49_77 ();
 sg13g2_fill_1 FILLER_49_81 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_96 ();
 sg13g2_fill_1 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_104 ();
 sg13g2_fill_2 FILLER_49_149 ();
 sg13g2_fill_2 FILLER_49_156 ();
 sg13g2_fill_2 FILLER_49_162 ();
 sg13g2_fill_2 FILLER_49_168 ();
 sg13g2_fill_1 FILLER_49_170 ();
 sg13g2_decap_8 FILLER_49_176 ();
 sg13g2_fill_2 FILLER_49_183 ();
 sg13g2_fill_1 FILLER_49_321 ();
 sg13g2_fill_1 FILLER_49_326 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_fill_1 FILLER_49_348 ();
 sg13g2_fill_2 FILLER_49_359 ();
 sg13g2_fill_2 FILLER_49_365 ();
 sg13g2_fill_1 FILLER_49_367 ();
 sg13g2_fill_1 FILLER_49_372 ();
 sg13g2_fill_1 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_402 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_fill_1 FILLER_50_70 ();
 sg13g2_fill_1 FILLER_50_75 ();
 sg13g2_fill_1 FILLER_50_80 ();
 sg13g2_fill_1 FILLER_50_86 ();
 sg13g2_fill_1 FILLER_50_124 ();
 sg13g2_fill_1 FILLER_50_129 ();
 sg13g2_decap_4 FILLER_50_146 ();
 sg13g2_fill_2 FILLER_50_178 ();
 sg13g2_fill_2 FILLER_50_195 ();
 sg13g2_fill_2 FILLER_50_232 ();
 sg13g2_fill_2 FILLER_50_238 ();
 sg13g2_fill_1 FILLER_50_240 ();
 sg13g2_fill_2 FILLER_50_314 ();
 sg13g2_fill_2 FILLER_50_326 ();
 sg13g2_fill_1 FILLER_50_340 ();
 sg13g2_decap_4 FILLER_50_346 ();
 sg13g2_fill_1 FILLER_50_350 ();
 sg13g2_decap_4 FILLER_50_356 ();
 sg13g2_fill_1 FILLER_50_360 ();
 sg13g2_decap_4 FILLER_50_366 ();
 sg13g2_decap_8 FILLER_50_379 ();
 sg13g2_fill_2 FILLER_50_386 ();
 sg13g2_decap_4 FILLER_50_393 ();
 sg13g2_decap_4 FILLER_50_411 ();
 sg13g2_fill_1 FILLER_50_425 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_4 FILLER_51_63 ();
 sg13g2_fill_1 FILLER_51_96 ();
 sg13g2_fill_2 FILLER_51_137 ();
 sg13g2_fill_2 FILLER_51_143 ();
 sg13g2_fill_1 FILLER_51_150 ();
 sg13g2_fill_2 FILLER_51_216 ();
 sg13g2_fill_1 FILLER_51_218 ();
 sg13g2_decap_4 FILLER_51_232 ();
 sg13g2_fill_1 FILLER_51_236 ();
 sg13g2_fill_2 FILLER_51_245 ();
 sg13g2_fill_1 FILLER_51_247 ();
 sg13g2_fill_2 FILLER_51_253 ();
 sg13g2_fill_1 FILLER_51_255 ();
 sg13g2_fill_2 FILLER_51_260 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_fill_2 FILLER_51_310 ();
 sg13g2_fill_1 FILLER_51_352 ();
 sg13g2_fill_1 FILLER_51_358 ();
 sg13g2_fill_2 FILLER_51_366 ();
 sg13g2_fill_2 FILLER_51_394 ();
 sg13g2_fill_2 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_56 ();
 sg13g2_fill_1 FILLER_52_83 ();
 sg13g2_fill_2 FILLER_52_128 ();
 sg13g2_fill_1 FILLER_52_181 ();
 sg13g2_fill_2 FILLER_52_229 ();
 sg13g2_fill_1 FILLER_52_240 ();
 sg13g2_fill_2 FILLER_52_301 ();
 sg13g2_decap_4 FILLER_52_307 ();
 sg13g2_fill_1 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_372 ();
 sg13g2_fill_2 FILLER_52_378 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_fill_1 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_68 ();
 sg13g2_fill_2 FILLER_53_79 ();
 sg13g2_decap_8 FILLER_53_86 ();
 sg13g2_fill_1 FILLER_53_93 ();
 sg13g2_decap_4 FILLER_53_104 ();
 sg13g2_fill_1 FILLER_53_108 ();
 sg13g2_fill_1 FILLER_53_113 ();
 sg13g2_fill_2 FILLER_53_118 ();
 sg13g2_fill_1 FILLER_53_120 ();
 sg13g2_fill_1 FILLER_53_125 ();
 sg13g2_fill_2 FILLER_53_130 ();
 sg13g2_fill_2 FILLER_53_143 ();
 sg13g2_fill_1 FILLER_53_178 ();
 sg13g2_fill_1 FILLER_53_206 ();
 sg13g2_decap_4 FILLER_53_211 ();
 sg13g2_fill_1 FILLER_53_247 ();
 sg13g2_decap_4 FILLER_53_252 ();
 sg13g2_fill_2 FILLER_53_264 ();
 sg13g2_fill_1 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_271 ();
 sg13g2_fill_2 FILLER_53_276 ();
 sg13g2_fill_1 FILLER_53_278 ();
 sg13g2_fill_2 FILLER_53_295 ();
 sg13g2_fill_2 FILLER_53_301 ();
 sg13g2_fill_1 FILLER_53_303 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_fill_2 FILLER_53_315 ();
 sg13g2_fill_1 FILLER_53_317 ();
 sg13g2_decap_4 FILLER_53_328 ();
 sg13g2_decap_4 FILLER_53_336 ();
 sg13g2_fill_2 FILLER_53_376 ();
 sg13g2_fill_1 FILLER_53_378 ();
 sg13g2_fill_2 FILLER_53_386 ();
 sg13g2_fill_2 FILLER_53_410 ();
 sg13g2_fill_1 FILLER_53_412 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_4 FILLER_54_63 ();
 sg13g2_fill_1 FILLER_54_67 ();
 sg13g2_fill_2 FILLER_54_94 ();
 sg13g2_fill_1 FILLER_54_101 ();
 sg13g2_fill_2 FILLER_54_111 ();
 sg13g2_decap_8 FILLER_54_118 ();
 sg13g2_fill_2 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_fill_1 FILLER_54_136 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_fill_1 FILLER_54_165 ();
 sg13g2_fill_1 FILLER_54_173 ();
 sg13g2_fill_2 FILLER_54_179 ();
 sg13g2_fill_2 FILLER_54_185 ();
 sg13g2_fill_1 FILLER_54_187 ();
 sg13g2_fill_2 FILLER_54_205 ();
 sg13g2_fill_1 FILLER_54_207 ();
 sg13g2_fill_2 FILLER_54_241 ();
 sg13g2_fill_1 FILLER_54_243 ();
 sg13g2_decap_8 FILLER_54_249 ();
 sg13g2_decap_8 FILLER_54_256 ();
 sg13g2_decap_4 FILLER_54_263 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_fill_1 FILLER_54_297 ();
 sg13g2_fill_1 FILLER_54_324 ();
 sg13g2_fill_1 FILLER_54_329 ();
 sg13g2_fill_1 FILLER_54_340 ();
 sg13g2_fill_1 FILLER_54_345 ();
 sg13g2_decap_8 FILLER_54_376 ();
 sg13g2_decap_4 FILLER_54_383 ();
 sg13g2_fill_2 FILLER_54_387 ();
 sg13g2_fill_1 FILLER_54_394 ();
 sg13g2_fill_2 FILLER_54_410 ();
 sg13g2_fill_1 FILLER_54_422 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_4 FILLER_55_63 ();
 sg13g2_fill_2 FILLER_55_67 ();
 sg13g2_fill_2 FILLER_55_148 ();
 sg13g2_fill_2 FILLER_55_159 ();
 sg13g2_decap_4 FILLER_55_189 ();
 sg13g2_fill_1 FILLER_55_193 ();
 sg13g2_fill_1 FILLER_55_197 ();
 sg13g2_fill_1 FILLER_55_207 ();
 sg13g2_fill_1 FILLER_55_216 ();
 sg13g2_fill_2 FILLER_55_278 ();
 sg13g2_fill_1 FILLER_55_280 ();
 sg13g2_fill_1 FILLER_55_306 ();
 sg13g2_fill_2 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_55_383 ();
 sg13g2_decap_8 FILLER_55_390 ();
 sg13g2_decap_4 FILLER_55_397 ();
 sg13g2_fill_1 FILLER_55_401 ();
 sg13g2_fill_1 FILLER_55_421 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_4 FILLER_56_63 ();
 sg13g2_fill_2 FILLER_56_77 ();
 sg13g2_fill_1 FILLER_56_79 ();
 sg13g2_fill_1 FILLER_56_84 ();
 sg13g2_fill_1 FILLER_56_89 ();
 sg13g2_fill_1 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_174 ();
 sg13g2_fill_2 FILLER_56_181 ();
 sg13g2_fill_2 FILLER_56_187 ();
 sg13g2_fill_1 FILLER_56_194 ();
 sg13g2_fill_1 FILLER_56_201 ();
 sg13g2_fill_1 FILLER_56_212 ();
 sg13g2_fill_1 FILLER_56_223 ();
 sg13g2_decap_4 FILLER_56_248 ();
 sg13g2_fill_2 FILLER_56_252 ();
 sg13g2_fill_1 FILLER_56_258 ();
 sg13g2_fill_1 FILLER_56_294 ();
 sg13g2_fill_1 FILLER_56_300 ();
 sg13g2_fill_2 FILLER_56_305 ();
 sg13g2_fill_1 FILLER_56_307 ();
 sg13g2_fill_1 FILLER_56_338 ();
 sg13g2_fill_2 FILLER_56_374 ();
 sg13g2_fill_1 FILLER_56_383 ();
 sg13g2_fill_2 FILLER_56_388 ();
 sg13g2_fill_2 FILLER_56_395 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_2 FILLER_56_419 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_fill_2 FILLER_57_83 ();
 sg13g2_fill_2 FILLER_57_150 ();
 sg13g2_fill_1 FILLER_57_172 ();
 sg13g2_fill_1 FILLER_57_191 ();
 sg13g2_fill_1 FILLER_57_207 ();
 sg13g2_fill_2 FILLER_57_241 ();
 sg13g2_decap_4 FILLER_57_248 ();
 sg13g2_fill_1 FILLER_57_252 ();
 sg13g2_fill_1 FILLER_57_259 ();
 sg13g2_fill_2 FILLER_57_305 ();
 sg13g2_fill_1 FILLER_57_307 ();
 sg13g2_fill_1 FILLER_57_312 ();
 sg13g2_fill_1 FILLER_57_318 ();
 sg13g2_fill_1 FILLER_57_324 ();
 sg13g2_fill_1 FILLER_57_375 ();
 sg13g2_fill_2 FILLER_57_423 ();
 sg13g2_fill_1 FILLER_57_425 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_4 FILLER_58_56 ();
 sg13g2_fill_2 FILLER_58_60 ();
 sg13g2_decap_8 FILLER_58_87 ();
 sg13g2_fill_2 FILLER_58_94 ();
 sg13g2_fill_1 FILLER_58_123 ();
 sg13g2_fill_2 FILLER_58_133 ();
 sg13g2_fill_1 FILLER_58_135 ();
 sg13g2_fill_1 FILLER_58_143 ();
 sg13g2_fill_1 FILLER_58_187 ();
 sg13g2_fill_1 FILLER_58_228 ();
 sg13g2_decap_4 FILLER_58_245 ();
 sg13g2_fill_2 FILLER_58_346 ();
 sg13g2_fill_2 FILLER_58_381 ();
 sg13g2_fill_1 FILLER_58_383 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_4 FILLER_59_56 ();
 sg13g2_fill_2 FILLER_59_60 ();
 sg13g2_fill_1 FILLER_59_91 ();
 sg13g2_fill_2 FILLER_59_102 ();
 sg13g2_fill_1 FILLER_59_104 ();
 sg13g2_fill_1 FILLER_59_115 ();
 sg13g2_fill_2 FILLER_59_121 ();
 sg13g2_fill_1 FILLER_59_123 ();
 sg13g2_fill_1 FILLER_59_150 ();
 sg13g2_fill_2 FILLER_59_168 ();
 sg13g2_decap_4 FILLER_59_175 ();
 sg13g2_fill_2 FILLER_59_179 ();
 sg13g2_decap_8 FILLER_59_185 ();
 sg13g2_fill_1 FILLER_59_192 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_decap_8 FILLER_59_245 ();
 sg13g2_fill_2 FILLER_59_272 ();
 sg13g2_fill_1 FILLER_59_274 ();
 sg13g2_fill_1 FILLER_59_286 ();
 sg13g2_fill_2 FILLER_59_350 ();
 sg13g2_fill_1 FILLER_59_352 ();
 sg13g2_fill_1 FILLER_59_368 ();
 sg13g2_fill_1 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_409 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_fill_2 FILLER_60_63 ();
 sg13g2_decap_4 FILLER_60_119 ();
 sg13g2_fill_1 FILLER_60_123 ();
 sg13g2_fill_2 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_172 ();
 sg13g2_decap_4 FILLER_60_179 ();
 sg13g2_decap_8 FILLER_60_187 ();
 sg13g2_fill_2 FILLER_60_194 ();
 sg13g2_fill_1 FILLER_60_196 ();
 sg13g2_fill_1 FILLER_60_252 ();
 sg13g2_decap_4 FILLER_60_257 ();
 sg13g2_fill_1 FILLER_60_261 ();
 sg13g2_fill_2 FILLER_60_267 ();
 sg13g2_fill_2 FILLER_60_274 ();
 sg13g2_fill_1 FILLER_60_297 ();
 sg13g2_fill_1 FILLER_60_301 ();
 sg13g2_fill_1 FILLER_60_306 ();
 sg13g2_fill_1 FILLER_60_316 ();
 sg13g2_fill_1 FILLER_60_321 ();
 sg13g2_fill_2 FILLER_60_359 ();
 sg13g2_fill_1 FILLER_60_361 ();
 sg13g2_fill_2 FILLER_60_386 ();
 sg13g2_fill_1 FILLER_60_393 ();
 sg13g2_fill_1 FILLER_60_398 ();
 sg13g2_fill_2 FILLER_60_404 ();
 sg13g2_fill_2 FILLER_60_411 ();
 sg13g2_fill_2 FILLER_60_418 ();
 sg13g2_fill_2 FILLER_60_428 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_fill_2 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_65 ();
 sg13g2_fill_2 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_124 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_fill_2 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_190 ();
 sg13g2_decap_4 FILLER_61_197 ();
 sg13g2_fill_1 FILLER_61_201 ();
 sg13g2_fill_1 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_214 ();
 sg13g2_fill_1 FILLER_61_231 ();
 sg13g2_fill_1 FILLER_61_237 ();
 sg13g2_fill_2 FILLER_61_241 ();
 sg13g2_fill_2 FILLER_61_248 ();
 sg13g2_fill_2 FILLER_61_254 ();
 sg13g2_fill_1 FILLER_61_256 ();
 sg13g2_decap_8 FILLER_61_272 ();
 sg13g2_fill_1 FILLER_61_287 ();
 sg13g2_fill_2 FILLER_61_293 ();
 sg13g2_fill_1 FILLER_61_295 ();
 sg13g2_decap_4 FILLER_61_316 ();
 sg13g2_fill_2 FILLER_61_351 ();
 sg13g2_fill_2 FILLER_61_362 ();
 sg13g2_decap_4 FILLER_61_370 ();
 sg13g2_fill_2 FILLER_61_390 ();
 sg13g2_fill_1 FILLER_61_397 ();
 sg13g2_fill_1 FILLER_61_403 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_fill_1 FILLER_61_419 ();
 sg13g2_fill_2 FILLER_61_427 ();
 sg13g2_fill_1 FILLER_61_429 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_fill_1 FILLER_62_63 ();
 sg13g2_fill_2 FILLER_62_124 ();
 sg13g2_fill_1 FILLER_62_142 ();
 sg13g2_fill_1 FILLER_62_153 ();
 sg13g2_fill_1 FILLER_62_158 ();
 sg13g2_decap_4 FILLER_62_197 ();
 sg13g2_fill_1 FILLER_62_205 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_decap_4 FILLER_62_217 ();
 sg13g2_fill_1 FILLER_62_272 ();
 sg13g2_fill_1 FILLER_62_283 ();
 sg13g2_fill_2 FILLER_62_302 ();
 sg13g2_fill_1 FILLER_62_314 ();
 sg13g2_fill_2 FILLER_62_319 ();
 sg13g2_fill_2 FILLER_62_326 ();
 sg13g2_fill_2 FILLER_62_333 ();
 sg13g2_fill_2 FILLER_62_382 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_fill_2 FILLER_62_394 ();
 sg13g2_fill_1 FILLER_62_396 ();
 sg13g2_fill_1 FILLER_62_407 ();
 sg13g2_fill_1 FILLER_62_413 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_4 FILLER_63_63 ();
 sg13g2_fill_1 FILLER_63_96 ();
 sg13g2_decap_4 FILLER_63_107 ();
 sg13g2_fill_2 FILLER_63_114 ();
 sg13g2_fill_2 FILLER_63_119 ();
 sg13g2_fill_1 FILLER_63_125 ();
 sg13g2_decap_4 FILLER_63_155 ();
 sg13g2_fill_1 FILLER_63_159 ();
 sg13g2_fill_2 FILLER_63_173 ();
 sg13g2_fill_2 FILLER_63_190 ();
 sg13g2_fill_2 FILLER_63_197 ();
 sg13g2_fill_1 FILLER_63_204 ();
 sg13g2_fill_1 FILLER_63_209 ();
 sg13g2_fill_2 FILLER_63_220 ();
 sg13g2_decap_8 FILLER_63_227 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_fill_1 FILLER_63_236 ();
 sg13g2_decap_4 FILLER_63_241 ();
 sg13g2_fill_2 FILLER_63_249 ();
 sg13g2_fill_1 FILLER_63_251 ();
 sg13g2_fill_1 FILLER_63_285 ();
 sg13g2_fill_1 FILLER_63_318 ();
 sg13g2_fill_2 FILLER_63_334 ();
 sg13g2_decap_4 FILLER_63_340 ();
 sg13g2_fill_2 FILLER_63_344 ();
 sg13g2_decap_4 FILLER_63_351 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_4 FILLER_64_70 ();
 sg13g2_fill_1 FILLER_64_74 ();
 sg13g2_decap_4 FILLER_64_80 ();
 sg13g2_fill_2 FILLER_64_105 ();
 sg13g2_fill_1 FILLER_64_156 ();
 sg13g2_fill_1 FILLER_64_160 ();
 sg13g2_fill_1 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_185 ();
 sg13g2_decap_4 FILLER_64_231 ();
 sg13g2_fill_1 FILLER_64_235 ();
 sg13g2_fill_2 FILLER_64_259 ();
 sg13g2_fill_1 FILLER_64_301 ();
 sg13g2_fill_1 FILLER_64_311 ();
 sg13g2_fill_2 FILLER_64_330 ();
 sg13g2_fill_2 FILLER_64_342 ();
 sg13g2_fill_1 FILLER_64_411 ();
 sg13g2_fill_2 FILLER_64_420 ();
 sg13g2_fill_1 FILLER_64_426 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_fill_2 FILLER_65_77 ();
 sg13g2_fill_1 FILLER_65_79 ();
 sg13g2_fill_2 FILLER_65_152 ();
 sg13g2_fill_1 FILLER_65_154 ();
 sg13g2_fill_1 FILLER_65_183 ();
 sg13g2_decap_4 FILLER_65_230 ();
 sg13g2_fill_1 FILLER_65_234 ();
 sg13g2_fill_2 FILLER_65_265 ();
 sg13g2_fill_2 FILLER_65_283 ();
 sg13g2_fill_2 FILLER_65_290 ();
 sg13g2_fill_2 FILLER_65_297 ();
 sg13g2_fill_2 FILLER_65_304 ();
 sg13g2_decap_4 FILLER_65_316 ();
 sg13g2_fill_1 FILLER_65_320 ();
 sg13g2_fill_2 FILLER_65_326 ();
 sg13g2_fill_1 FILLER_65_333 ();
 sg13g2_fill_2 FILLER_65_339 ();
 sg13g2_fill_1 FILLER_65_341 ();
 sg13g2_fill_2 FILLER_65_354 ();
 sg13g2_fill_1 FILLER_65_356 ();
 sg13g2_fill_1 FILLER_65_384 ();
 sg13g2_fill_2 FILLER_65_410 ();
 sg13g2_fill_2 FILLER_65_420 ();
 sg13g2_fill_1 FILLER_65_422 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_fill_1 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_87 ();
 sg13g2_fill_2 FILLER_66_94 ();
 sg13g2_fill_1 FILLER_66_96 ();
 sg13g2_fill_1 FILLER_66_101 ();
 sg13g2_fill_1 FILLER_66_107 ();
 sg13g2_fill_2 FILLER_66_113 ();
 sg13g2_fill_1 FILLER_66_234 ();
 sg13g2_fill_2 FILLER_66_240 ();
 sg13g2_fill_1 FILLER_66_246 ();
 sg13g2_fill_2 FILLER_66_251 ();
 sg13g2_fill_2 FILLER_66_263 ();
 sg13g2_fill_1 FILLER_66_270 ();
 sg13g2_fill_2 FILLER_66_275 ();
 sg13g2_fill_1 FILLER_66_277 ();
 sg13g2_fill_2 FILLER_66_282 ();
 sg13g2_fill_1 FILLER_66_284 ();
 sg13g2_fill_2 FILLER_66_289 ();
 sg13g2_decap_8 FILLER_66_302 ();
 sg13g2_decap_8 FILLER_66_309 ();
 sg13g2_fill_2 FILLER_66_316 ();
 sg13g2_fill_1 FILLER_66_318 ();
 sg13g2_decap_4 FILLER_66_324 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_fill_2 FILLER_66_343 ();
 sg13g2_fill_2 FILLER_66_350 ();
 sg13g2_fill_1 FILLER_66_352 ();
 sg13g2_fill_2 FILLER_66_377 ();
 sg13g2_fill_2 FILLER_66_402 ();
 sg13g2_fill_1 FILLER_66_404 ();
 sg13g2_fill_2 FILLER_66_428 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_4 FILLER_67_77 ();
 sg13g2_fill_1 FILLER_67_81 ();
 sg13g2_fill_1 FILLER_67_87 ();
 sg13g2_fill_1 FILLER_67_96 ();
 sg13g2_fill_1 FILLER_67_102 ();
 sg13g2_fill_1 FILLER_67_107 ();
 sg13g2_fill_2 FILLER_67_114 ();
 sg13g2_fill_1 FILLER_67_116 ();
 sg13g2_fill_2 FILLER_67_129 ();
 sg13g2_fill_2 FILLER_67_135 ();
 sg13g2_fill_2 FILLER_67_153 ();
 sg13g2_fill_2 FILLER_67_160 ();
 sg13g2_decap_4 FILLER_67_193 ();
 sg13g2_fill_2 FILLER_67_197 ();
 sg13g2_fill_1 FILLER_67_213 ();
 sg13g2_fill_1 FILLER_67_218 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_fill_2 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_266 ();
 sg13g2_fill_1 FILLER_67_282 ();
 sg13g2_fill_2 FILLER_67_288 ();
 sg13g2_fill_2 FILLER_67_304 ();
 sg13g2_fill_1 FILLER_67_339 ();
 sg13g2_fill_1 FILLER_67_361 ();
 sg13g2_fill_1 FILLER_67_369 ();
 sg13g2_decap_4 FILLER_67_424 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_4 FILLER_68_77 ();
 sg13g2_fill_1 FILLER_68_81 ();
 sg13g2_fill_1 FILLER_68_119 ();
 sg13g2_fill_2 FILLER_68_128 ();
 sg13g2_fill_1 FILLER_68_134 ();
 sg13g2_fill_1 FILLER_68_164 ();
 sg13g2_decap_4 FILLER_68_190 ();
 sg13g2_fill_1 FILLER_68_194 ();
 sg13g2_fill_1 FILLER_68_220 ();
 sg13g2_fill_2 FILLER_68_230 ();
 sg13g2_fill_1 FILLER_68_232 ();
 sg13g2_fill_1 FILLER_68_237 ();
 sg13g2_fill_1 FILLER_68_259 ();
 sg13g2_fill_1 FILLER_68_270 ();
 sg13g2_fill_1 FILLER_68_276 ();
 sg13g2_fill_1 FILLER_68_282 ();
 sg13g2_fill_1 FILLER_68_312 ();
 sg13g2_fill_1 FILLER_68_318 ();
 sg13g2_fill_2 FILLER_68_401 ();
 sg13g2_fill_1 FILLER_68_403 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_fill_1 FILLER_69_104 ();
 sg13g2_decap_4 FILLER_69_126 ();
 sg13g2_fill_1 FILLER_69_130 ();
 sg13g2_fill_2 FILLER_69_160 ();
 sg13g2_fill_2 FILLER_69_192 ();
 sg13g2_fill_1 FILLER_69_194 ();
 sg13g2_fill_1 FILLER_69_315 ();
 sg13g2_fill_2 FILLER_69_355 ();
 sg13g2_fill_2 FILLER_69_361 ();
 sg13g2_fill_1 FILLER_69_363 ();
 sg13g2_fill_1 FILLER_69_368 ();
 sg13g2_fill_1 FILLER_69_374 ();
 sg13g2_fill_1 FILLER_69_388 ();
 sg13g2_fill_2 FILLER_69_416 ();
 sg13g2_fill_2 FILLER_69_428 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_115 ();
 sg13g2_decap_4 FILLER_70_122 ();
 sg13g2_fill_1 FILLER_70_126 ();
 sg13g2_fill_1 FILLER_70_134 ();
 sg13g2_fill_1 FILLER_70_140 ();
 sg13g2_fill_1 FILLER_70_183 ();
 sg13g2_fill_2 FILLER_70_189 ();
 sg13g2_fill_1 FILLER_70_191 ();
 sg13g2_fill_2 FILLER_70_216 ();
 sg13g2_fill_1 FILLER_70_218 ();
 sg13g2_fill_1 FILLER_70_223 ();
 sg13g2_fill_1 FILLER_70_249 ();
 sg13g2_fill_1 FILLER_70_254 ();
 sg13g2_fill_1 FILLER_70_275 ();
 sg13g2_fill_1 FILLER_70_284 ();
 sg13g2_fill_1 FILLER_70_318 ();
 sg13g2_fill_1 FILLER_70_344 ();
 sg13g2_fill_1 FILLER_70_362 ();
 sg13g2_fill_1 FILLER_70_373 ();
 sg13g2_decap_4 FILLER_70_379 ();
 sg13g2_fill_1 FILLER_70_383 ();
 sg13g2_fill_1 FILLER_70_388 ();
 sg13g2_fill_1 FILLER_70_397 ();
 sg13g2_fill_1 FILLER_70_416 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_fill_2 FILLER_71_84 ();
 sg13g2_fill_1 FILLER_71_86 ();
 sg13g2_fill_1 FILLER_71_98 ();
 sg13g2_fill_2 FILLER_71_124 ();
 sg13g2_decap_4 FILLER_71_135 ();
 sg13g2_fill_2 FILLER_71_139 ();
 sg13g2_fill_1 FILLER_71_171 ();
 sg13g2_fill_1 FILLER_71_178 ();
 sg13g2_fill_1 FILLER_71_184 ();
 sg13g2_fill_1 FILLER_71_189 ();
 sg13g2_fill_2 FILLER_71_193 ();
 sg13g2_fill_2 FILLER_71_199 ();
 sg13g2_fill_1 FILLER_71_201 ();
 sg13g2_fill_1 FILLER_71_206 ();
 sg13g2_decap_8 FILLER_71_211 ();
 sg13g2_decap_8 FILLER_71_218 ();
 sg13g2_fill_2 FILLER_71_225 ();
 sg13g2_decap_8 FILLER_71_232 ();
 sg13g2_decap_8 FILLER_71_239 ();
 sg13g2_fill_1 FILLER_71_292 ();
 sg13g2_fill_2 FILLER_71_297 ();
 sg13g2_fill_1 FILLER_71_304 ();
 sg13g2_decap_8 FILLER_71_309 ();
 sg13g2_fill_2 FILLER_71_316 ();
 sg13g2_fill_1 FILLER_71_318 ();
 sg13g2_fill_2 FILLER_71_355 ();
 sg13g2_fill_1 FILLER_71_357 ();
 sg13g2_fill_2 FILLER_71_373 ();
 sg13g2_fill_1 FILLER_71_394 ();
 sg13g2_fill_1 FILLER_71_425 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_84 ();
 sg13g2_fill_1 FILLER_72_86 ();
 sg13g2_fill_1 FILLER_72_112 ();
 sg13g2_fill_1 FILLER_72_118 ();
 sg13g2_fill_1 FILLER_72_124 ();
 sg13g2_decap_4 FILLER_72_141 ();
 sg13g2_fill_2 FILLER_72_145 ();
 sg13g2_decap_8 FILLER_72_151 ();
 sg13g2_decap_8 FILLER_72_158 ();
 sg13g2_decap_8 FILLER_72_165 ();
 sg13g2_decap_8 FILLER_72_172 ();
 sg13g2_fill_2 FILLER_72_179 ();
 sg13g2_fill_2 FILLER_72_185 ();
 sg13g2_decap_4 FILLER_72_191 ();
 sg13g2_fill_2 FILLER_72_195 ();
 sg13g2_fill_1 FILLER_72_245 ();
 sg13g2_fill_1 FILLER_72_251 ();
 sg13g2_decap_8 FILLER_72_261 ();
 sg13g2_fill_1 FILLER_72_277 ();
 sg13g2_fill_1 FILLER_72_295 ();
 sg13g2_decap_8 FILLER_72_305 ();
 sg13g2_decap_8 FILLER_72_312 ();
 sg13g2_fill_2 FILLER_72_319 ();
 sg13g2_fill_2 FILLER_72_325 ();
 sg13g2_decap_4 FILLER_72_332 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_4 FILLER_73_63 ();
 sg13g2_fill_2 FILLER_73_67 ();
 sg13g2_fill_1 FILLER_73_90 ();
 sg13g2_fill_2 FILLER_73_95 ();
 sg13g2_fill_1 FILLER_73_137 ();
 sg13g2_decap_4 FILLER_73_166 ();
 sg13g2_fill_2 FILLER_73_195 ();
 sg13g2_decap_4 FILLER_73_212 ();
 sg13g2_fill_2 FILLER_73_244 ();
 sg13g2_fill_2 FILLER_73_347 ();
 sg13g2_fill_2 FILLER_73_377 ();
 sg13g2_fill_1 FILLER_73_403 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_fill_1 FILLER_74_111 ();
 sg13g2_fill_2 FILLER_74_150 ();
 sg13g2_fill_2 FILLER_74_259 ();
 sg13g2_fill_2 FILLER_74_303 ();
 sg13g2_fill_1 FILLER_74_305 ();
 sg13g2_fill_1 FILLER_74_311 ();
 sg13g2_fill_2 FILLER_74_371 ();
 sg13g2_fill_1 FILLER_74_419 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_fill_2 FILLER_75_70 ();
 sg13g2_fill_1 FILLER_75_72 ();
 sg13g2_fill_2 FILLER_75_97 ();
 sg13g2_decap_8 FILLER_75_103 ();
 sg13g2_fill_1 FILLER_75_110 ();
 sg13g2_fill_1 FILLER_75_116 ();
 sg13g2_fill_1 FILLER_75_122 ();
 sg13g2_fill_1 FILLER_75_128 ();
 sg13g2_fill_1 FILLER_75_134 ();
 sg13g2_fill_2 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_192 ();
 sg13g2_fill_2 FILLER_75_210 ();
 sg13g2_fill_1 FILLER_75_212 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_fill_2 FILLER_75_259 ();
 sg13g2_fill_2 FILLER_75_323 ();
 sg13g2_fill_2 FILLER_75_418 ();
 sg13g2_fill_1 FILLER_75_425 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_4 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_109 ();
 sg13g2_fill_1 FILLER_76_114 ();
 sg13g2_fill_1 FILLER_76_125 ();
 sg13g2_fill_1 FILLER_76_130 ();
 sg13g2_fill_1 FILLER_76_141 ();
 sg13g2_fill_1 FILLER_76_146 ();
 sg13g2_fill_2 FILLER_76_161 ();
 sg13g2_fill_2 FILLER_76_182 ();
 sg13g2_fill_2 FILLER_76_197 ();
 sg13g2_fill_2 FILLER_76_216 ();
 sg13g2_fill_1 FILLER_76_227 ();
 sg13g2_fill_1 FILLER_76_233 ();
 sg13g2_fill_1 FILLER_76_238 ();
 sg13g2_fill_1 FILLER_76_253 ();
 sg13g2_fill_1 FILLER_76_259 ();
 sg13g2_decap_4 FILLER_76_264 ();
 sg13g2_fill_1 FILLER_76_304 ();
 sg13g2_fill_1 FILLER_76_309 ();
 sg13g2_fill_1 FILLER_76_315 ();
 sg13g2_fill_1 FILLER_76_320 ();
 sg13g2_fill_1 FILLER_76_360 ();
 sg13g2_fill_2 FILLER_76_366 ();
 sg13g2_fill_1 FILLER_76_388 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_fill_2 FILLER_77_98 ();
 sg13g2_fill_1 FILLER_77_100 ();
 sg13g2_fill_1 FILLER_77_117 ();
 sg13g2_fill_2 FILLER_77_143 ();
 sg13g2_fill_1 FILLER_77_195 ();
 sg13g2_fill_1 FILLER_77_203 ();
 sg13g2_fill_1 FILLER_77_209 ();
 sg13g2_fill_1 FILLER_77_219 ();
 sg13g2_fill_1 FILLER_77_241 ();
 sg13g2_fill_1 FILLER_77_303 ();
 sg13g2_fill_2 FILLER_77_356 ();
 sg13g2_fill_2 FILLER_77_428 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_4 FILLER_78_84 ();
 sg13g2_fill_1 FILLER_78_88 ();
 sg13g2_fill_1 FILLER_78_175 ();
 sg13g2_fill_1 FILLER_78_185 ();
 sg13g2_fill_1 FILLER_78_213 ();
 sg13g2_fill_1 FILLER_78_218 ();
 sg13g2_fill_1 FILLER_78_222 ();
 sg13g2_fill_1 FILLER_78_228 ();
 sg13g2_fill_1 FILLER_78_322 ();
 sg13g2_fill_1 FILLER_78_405 ();
 sg13g2_fill_2 FILLER_78_427 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_fill_2 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_83 ();
 sg13g2_fill_1 FILLER_79_90 ();
 sg13g2_fill_2 FILLER_79_197 ();
 sg13g2_fill_1 FILLER_79_245 ();
 sg13g2_fill_2 FILLER_79_323 ();
 sg13g2_fill_1 FILLER_79_325 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_78 ();
 sg13g2_fill_1 FILLER_80_80 ();
 sg13g2_fill_1 FILLER_80_139 ();
 sg13g2_fill_1 FILLER_80_222 ();
 sg13g2_fill_2 FILLER_80_232 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_fill_1 FILLER_80_264 ();
 sg13g2_fill_1 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_275 ();
 sg13g2_fill_1 FILLER_80_280 ();
 sg13g2_fill_1 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_423 ();
endmodule
