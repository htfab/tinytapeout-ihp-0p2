module tt_um_calonso88_rsa (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire clknet_leaf_0_clk;
 wire net156;
 wire eoc_rsa;
 wire \gpio_wrapper_i.gpio_start_cmd_i.data ;
 wire \gpio_wrapper_i.gpio_start_cmd_i.data_dly ;
 wire \gpio_wrapper_i.gpio_stop_cmd_i.data ;
 wire \gpio_wrapper_i.gpio_stop_cmd_i.data_dly ;
 wire \gpio_wrapper_i.sync_gpio_start.data_sync[1] ;
 wire \gpio_wrapper_i.sync_gpio_stop.data_sync[1] ;
 wire irq;
 wire \rsa_c[0] ;
 wire \rsa_c[1] ;
 wire \rsa_c[2] ;
 wire \rsa_c[3] ;
 wire \rsa_c[4] ;
 wire \rsa_c[5] ;
 wire \rsa_c[6] ;
 wire \rsa_c[7] ;
 wire \rsa_const[0] ;
 wire \rsa_const[1] ;
 wire \rsa_const[2] ;
 wire \rsa_const[3] ;
 wire \rsa_const[4] ;
 wire \rsa_const[5] ;
 wire \rsa_const[6] ;
 wire \rsa_const[7] ;
 wire \rsa_e[0] ;
 wire \rsa_e[1] ;
 wire \rsa_e[2] ;
 wire \rsa_e[3] ;
 wire \rsa_e[4] ;
 wire \rsa_e[5] ;
 wire \rsa_e[6] ;
 wire \rsa_e[7] ;
 wire \rsa_en_logic_i.state[0] ;
 wire \rsa_en_logic_i.state[1] ;
 wire \rsa_en_logic_i.state[2] ;
 wire \rsa_en_logic_i.state[3] ;
 wire \rsa_en_logic_i.state[4] ;
 wire \rsa_en_logic_i.state[5] ;
 wire \rsa_p[0] ;
 wire \rsa_p[1] ;
 wire \rsa_p[2] ;
 wire \rsa_p[3] ;
 wire \rsa_p[4] ;
 wire \rsa_p[5] ;
 wire \rsa_p[6] ;
 wire \rsa_p[7] ;
 wire \rsa_spi_wrapper_i.config_regs[0] ;
 wire \rsa_spi_wrapper_i.config_regs[10] ;
 wire \rsa_spi_wrapper_i.config_regs[11] ;
 wire \rsa_spi_wrapper_i.config_regs[12] ;
 wire \rsa_spi_wrapper_i.config_regs[13] ;
 wire \rsa_spi_wrapper_i.config_regs[14] ;
 wire \rsa_spi_wrapper_i.config_regs[15] ;
 wire \rsa_spi_wrapper_i.config_regs[1] ;
 wire \rsa_spi_wrapper_i.config_regs[2] ;
 wire \rsa_spi_wrapper_i.config_regs[32] ;
 wire \rsa_spi_wrapper_i.config_regs[33] ;
 wire \rsa_spi_wrapper_i.config_regs[34] ;
 wire \rsa_spi_wrapper_i.config_regs[35] ;
 wire \rsa_spi_wrapper_i.config_regs[36] ;
 wire \rsa_spi_wrapper_i.config_regs[37] ;
 wire \rsa_spi_wrapper_i.config_regs[38] ;
 wire \rsa_spi_wrapper_i.config_regs[39] ;
 wire \rsa_spi_wrapper_i.config_regs[3] ;
 wire \rsa_spi_wrapper_i.config_regs[48] ;
 wire \rsa_spi_wrapper_i.config_regs[49] ;
 wire \rsa_spi_wrapper_i.config_regs[4] ;
 wire \rsa_spi_wrapper_i.config_regs[50] ;
 wire \rsa_spi_wrapper_i.config_regs[51] ;
 wire \rsa_spi_wrapper_i.config_regs[52] ;
 wire \rsa_spi_wrapper_i.config_regs[53] ;
 wire \rsa_spi_wrapper_i.config_regs[54] ;
 wire \rsa_spi_wrapper_i.config_regs[55] ;
 wire \rsa_spi_wrapper_i.config_regs[56] ;
 wire \rsa_spi_wrapper_i.config_regs[57] ;
 wire \rsa_spi_wrapper_i.config_regs[58] ;
 wire \rsa_spi_wrapper_i.config_regs[59] ;
 wire \rsa_spi_wrapper_i.config_regs[5] ;
 wire \rsa_spi_wrapper_i.config_regs[60] ;
 wire \rsa_spi_wrapper_i.config_regs[61] ;
 wire \rsa_spi_wrapper_i.config_regs[62] ;
 wire \rsa_spi_wrapper_i.config_regs[63] ;
 wire \rsa_spi_wrapper_i.config_regs[6] ;
 wire \rsa_spi_wrapper_i.config_regs[7] ;
 wire \rsa_spi_wrapper_i.config_regs[8] ;
 wire \rsa_spi_wrapper_i.config_regs[9] ;
 wire \rsa_spi_wrapper_i.spi_clk ;
 wire \rsa_spi_wrapper_i.spi_cs_n ;
 wire \rsa_spi_wrapper_i.spi_miso ;
 wire \rsa_spi_wrapper_i.spi_mosi ;
 wire \rsa_spi_wrapper_i.spi_start_cmd_i.data_dly ;
 wire \rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[4] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[5] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[6] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[7] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o_vld ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[4] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[5] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[6] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ;
 wire \rsa_unit_i.P_i[0] ;
 wire \rsa_unit_i.P_i[1] ;
 wire \rsa_unit_i.P_i[2] ;
 wire \rsa_unit_i.P_i[3] ;
 wire \rsa_unit_i.P_i[4] ;
 wire \rsa_unit_i.P_i[5] ;
 wire \rsa_unit_i.P_i[6] ;
 wire \rsa_unit_i.P_i[7] ;
 wire \rsa_unit_i.P_i[8] ;
 wire \rsa_unit_i.P_i[9] ;
 wire \rsa_unit_i.R_i[0] ;
 wire \rsa_unit_i.R_i[1] ;
 wire \rsa_unit_i.R_i[2] ;
 wire \rsa_unit_i.R_i[3] ;
 wire \rsa_unit_i.R_i[4] ;
 wire \rsa_unit_i.R_i[5] ;
 wire \rsa_unit_i.R_i[6] ;
 wire \rsa_unit_i.R_i[7] ;
 wire \rsa_unit_i.R_i[8] ;
 wire \rsa_unit_i.R_i[9] ;
 wire \rsa_unit_i.mmm_multiply.A_bit ;
 wire \rsa_unit_i.mmm_multiply.adder2.fa_bit0.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[1].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[2].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[3].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[4].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[5].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[6].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[7].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[8].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[1] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[2] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[3] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[4] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[5] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[6] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[7] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[8] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[9] ;
 wire \rsa_unit_i.mmm_square.A_bit ;
 wire \rsa_unit_i.mmm_square.adder2.fa_bit0.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[1].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[2].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[3].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[4].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[5].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[6].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[7].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[8].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[1] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[2] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[3] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[4] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[5] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[6] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[7] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[8] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[9] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_rounds[0] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_rounds[1] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_rounds[2] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_rounds[3] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_steps[0] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_steps[1] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_steps[2] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_steps[3] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[0] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[1] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[2] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[3] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[4] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[5] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[6] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[7] ;
 wire \rsa_unit_i.rsa_control_fsm.increment_rounds ;
 wire \rsa_unit_i.rsa_control_fsm.load_exp ;
 wire \rsa_unit_i.rsa_control_fsm.state[0] ;
 wire \rsa_unit_i.rsa_control_fsm.state[10] ;
 wire \rsa_unit_i.rsa_control_fsm.state[11] ;
 wire \rsa_unit_i.rsa_control_fsm.state[1] ;
 wire \rsa_unit_i.rsa_control_fsm.state[2] ;
 wire \rsa_unit_i.rsa_control_fsm.state[3] ;
 wire \rsa_unit_i.rsa_control_fsm.state[6] ;
 wire \rsa_unit_i.rsa_control_fsm.state[7] ;
 wire \rsa_unit_i.rsa_control_fsm.state[8] ;
 wire \synchronizer_spi_clk_inst.data_sync[1] ;
 wire \synchronizer_spi_cs_n_inst.data_sync[1] ;
 wire \synchronizer_spi_mosi_inst.data_sync[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_1 _1756_ (.A(ena),
    .X(_1307_));
 sg13g2_inv_2 _1757_ (.Y(_1308_),
    .A(net111));
 sg13g2_inv_1 _1758_ (.Y(_1309_),
    .A(\gpio_wrapper_i.gpio_start_cmd_i.data_dly ));
 sg13g2_inv_1 _1759_ (.Y(_1310_),
    .A(\rsa_spi_wrapper_i.spi_start_cmd_i.data_dly ));
 sg13g2_a22oi_1 _1760_ (.Y(_1311_),
    .B1(\rsa_spi_wrapper_i.config_regs[8] ),
    .B2(_1310_),
    .A2(_1309_),
    .A1(\gpio_wrapper_i.gpio_start_cmd_i.data ));
 sg13g2_nor2_1 _1761_ (.A(_1308_),
    .B(_1311_),
    .Y(_1312_));
 sg13g2_a22oi_1 _1762_ (.Y(_1313_),
    .B1(\rsa_en_logic_i.state[3] ),
    .B2(_1312_),
    .A2(_1308_),
    .A1(\rsa_en_logic_i.state[2] ));
 sg13g2_inv_1 _1763_ (.Y(_0001_),
    .A(_1313_));
 sg13g2_buf_1 _1764_ (.A(net111),
    .X(_1314_));
 sg13g2_buf_1 _1765_ (.A(net110),
    .X(_1315_));
 sg13g2_nand2_1 _1766_ (.Y(_1316_),
    .A(net87),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_buf_1 _1767_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .X(_1317_));
 sg13g2_buf_2 _1768_ (.A(\rsa_spi_wrapper_i.spi_cs_n ),
    .X(_1318_));
 sg13g2_nor2b_1 _1769_ (.A(_1317_),
    .B_N(_1318_),
    .Y(_1319_));
 sg13g2_buf_1 _1770_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .X(_1320_));
 sg13g2_buf_2 _1771_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .X(_1321_));
 sg13g2_buf_2 _1772_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ),
    .X(_1322_));
 sg13g2_buf_2 _1773_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .X(_1323_));
 sg13g2_nor3_2 _1774_ (.A(_1321_),
    .B(_1322_),
    .C(_1323_),
    .Y(_1324_));
 sg13g2_mux2_1 _1775_ (.A0(_1319_),
    .A1(_1320_),
    .S(_1324_),
    .X(_1325_));
 sg13g2_nand2_1 _1776_ (.Y(_1326_),
    .A(net87),
    .B(_1325_));
 sg13g2_nand2_1 _1777_ (.Y(_1327_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ),
    .B(_1326_));
 sg13g2_o21ai_1 _1778_ (.B1(_1327_),
    .Y(_0005_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ),
    .A2(_1316_));
 sg13g2_buf_2 _1779_ (.A(\rsa_unit_i.rsa_control_fsm.state[1] ),
    .X(_1328_));
 sg13g2_buf_2 _1780_ (.A(\rsa_en_logic_i.state[4] ),
    .X(_1329_));
 sg13g2_buf_1 _1781_ (.A(\rsa_en_logic_i.state[1] ),
    .X(_1330_));
 sg13g2_nand2b_1 _1782_ (.Y(_1331_),
    .B(_0053_),
    .A_N(_1330_));
 sg13g2_nor2_2 _1783_ (.A(_1329_),
    .B(_1331_),
    .Y(_1332_));
 sg13g2_buf_1 _1784_ (.A(\rsa_unit_i.rsa_control_fsm.counter_steps[1] ),
    .X(_1333_));
 sg13g2_buf_2 _1785_ (.A(\rsa_unit_i.rsa_control_fsm.counter_steps[0] ),
    .X(_1334_));
 sg13g2_nand2b_1 _1786_ (.Y(_1335_),
    .B(_1334_),
    .A_N(_1333_));
 sg13g2_nor2b_1 _1787_ (.A(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ),
    .B_N(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ),
    .Y(_1336_));
 sg13g2_nand2b_1 _1788_ (.Y(_1337_),
    .B(_1336_),
    .A_N(_1335_));
 sg13g2_inv_1 _1789_ (.Y(_1338_),
    .A(_1337_));
 sg13g2_or2_1 _1790_ (.X(_1339_),
    .B(\rsa_en_logic_i.state[5] ),
    .A(\rsa_en_logic_i.state[2] ));
 sg13g2_buf_1 _1791_ (.A(_1339_),
    .X(_1340_));
 sg13g2_or3_1 _1792_ (.A(_1330_),
    .B(_1329_),
    .C(_1340_),
    .X(_1341_));
 sg13g2_buf_1 _1793_ (.A(_1341_),
    .X(_1342_));
 sg13g2_o21ai_1 _1794_ (.B1(net58),
    .Y(_1343_),
    .A1(_1332_),
    .A2(_1338_));
 sg13g2_nor3_2 _1795_ (.A(_1330_),
    .B(_1329_),
    .C(_1340_),
    .Y(_1344_));
 sg13g2_or2_1 _1796_ (.X(_1345_),
    .B(_1332_),
    .A(_1344_));
 sg13g2_buf_1 _1797_ (.A(_1345_),
    .X(_1346_));
 sg13g2_nor2_1 _1798_ (.A(_0052_),
    .B(_1346_),
    .Y(_1347_));
 sg13g2_a21o_1 _1799_ (.A2(_1343_),
    .A1(_1328_),
    .B1(_1347_),
    .X(_0011_));
 sg13g2_inv_1 _1800_ (.Y(_1348_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_inv_1 _1801_ (.Y(_1349_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_buf_1 _1802_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ),
    .X(_1350_));
 sg13g2_buf_1 _1803_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .X(_1351_));
 sg13g2_nor2_1 _1804_ (.A(_1351_),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .Y(_1352_));
 sg13g2_nand2b_1 _1805_ (.Y(_1353_),
    .B(_1352_),
    .A_N(_1350_));
 sg13g2_nor2_1 _1806_ (.A(_1349_),
    .B(_1353_),
    .Y(_1354_));
 sg13g2_buf_2 _1807_ (.A(_1354_),
    .X(_1355_));
 sg13g2_o21ai_1 _1808_ (.B1(net87),
    .Y(_1356_),
    .A1(_1319_),
    .A2(_1355_));
 sg13g2_nand2_1 _1809_ (.Y(_1357_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ),
    .B(_1356_));
 sg13g2_o21ai_1 _1810_ (.B1(_1357_),
    .Y(_0008_),
    .A1(_1348_),
    .A2(_1316_));
 sg13g2_o21ai_1 _1811_ (.B1(net110),
    .Y(_1358_),
    .A1(_1318_),
    .A2(_1355_));
 sg13g2_inv_1 _1812_ (.Y(_1359_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0] ));
 sg13g2_nand2b_1 _1813_ (.Y(_1360_),
    .B(net111),
    .A_N(_1318_));
 sg13g2_o21ai_1 _1814_ (.B1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ),
    .Y(_1361_),
    .A1(_1349_),
    .A2(_1353_));
 sg13g2_o21ai_1 _1815_ (.B1(_1361_),
    .Y(_1362_),
    .A1(_1359_),
    .A2(_1360_));
 sg13g2_a22oi_1 _1816_ (.Y(_1363_),
    .B1(_1362_),
    .B2(_1317_),
    .A2(_1358_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_inv_1 _1817_ (.Y(_0007_),
    .A(_1363_));
 sg13g2_buf_1 _1818_ (.A(net110),
    .X(_1364_));
 sg13g2_inv_1 _1819_ (.Y(_1365_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_nand3_1 _1820_ (.B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ),
    .C(_1355_),
    .A(net111),
    .Y(_1366_));
 sg13g2_buf_2 _1821_ (.A(_1366_),
    .X(_1367_));
 sg13g2_o21ai_1 _1822_ (.B1(_1367_),
    .Y(_0006_),
    .A1(net86),
    .A2(_1365_));
 sg13g2_nor2_1 _1823_ (.A(_1346_),
    .B(_1337_),
    .Y(_1368_));
 sg13g2_nand2_1 _1824_ (.Y(_1369_),
    .A(\rsa_unit_i.rsa_control_fsm.state[3] ),
    .B(_1368_));
 sg13g2_o21ai_1 _1825_ (.B1(_1369_),
    .Y(_0019_),
    .A1(_0051_),
    .A2(net58));
 sg13g2_buf_1 _1826_ (.A(eoc_rsa),
    .X(_1370_));
 sg13g2_nand2_1 _1827_ (.Y(_1371_),
    .A(net109),
    .B(net58));
 sg13g2_buf_1 _1828_ (.A(_1371_),
    .X(_1372_));
 sg13g2_inv_1 _1829_ (.Y(_1373_),
    .A(\rsa_unit_i.rsa_control_fsm.state[10] ));
 sg13g2_a22oi_1 _1830_ (.Y(_0009_),
    .B1(net40),
    .B2(_1373_),
    .A2(_1332_),
    .A1(_1340_));
 sg13g2_buf_8 _1831_ (.A(\rsa_unit_i.rsa_control_fsm.increment_rounds ),
    .X(_1374_));
 sg13g2_buf_1 _1832_ (.A(_1344_),
    .X(_1375_));
 sg13g2_nor2_2 _1833_ (.A(net57),
    .B(_1332_),
    .Y(_1376_));
 sg13g2_inv_1 _1834_ (.Y(_1377_),
    .A(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ));
 sg13g2_buf_1 _1835_ (.A(\rsa_unit_i.rsa_control_fsm.counter_rounds[1] ),
    .X(_1378_));
 sg13g2_buf_2 _1836_ (.A(\rsa_unit_i.rsa_control_fsm.counter_rounds[0] ),
    .X(_1379_));
 sg13g2_nand2b_1 _1837_ (.Y(_1380_),
    .B(_1379_),
    .A_N(_1378_));
 sg13g2_nor3_1 _1838_ (.A(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ),
    .B(_1377_),
    .C(_1380_),
    .Y(_1381_));
 sg13g2_nand3_1 _1839_ (.B(_1376_),
    .C(_1381_),
    .A(net108),
    .Y(_1382_));
 sg13g2_o21ai_1 _1840_ (.B1(_1382_),
    .Y(_0010_),
    .A1(_0052_),
    .A2(net58));
 sg13g2_inv_1 _1841_ (.Y(_1383_),
    .A(\gpio_wrapper_i.gpio_stop_cmd_i.data ));
 sg13g2_nand2b_1 _1842_ (.Y(_1384_),
    .B(\rsa_spi_wrapper_i.config_regs[9] ),
    .A_N(\rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly ));
 sg13g2_o21ai_1 _1843_ (.B1(_1384_),
    .Y(_1385_),
    .A1(_1383_),
    .A2(\gpio_wrapper_i.gpio_stop_cmd_i.data_dly ));
 sg13g2_buf_1 _1844_ (.A(_1385_),
    .X(_1386_));
 sg13g2_nand2_1 _1845_ (.Y(_1387_),
    .A(\rsa_en_logic_i.state[5] ),
    .B(_1315_));
 sg13g2_o21ai_1 _1846_ (.B1(net110),
    .Y(_1388_),
    .A1(_1370_),
    .A2(_1386_));
 sg13g2_nand2_1 _1847_ (.Y(_1389_),
    .A(_1330_),
    .B(_1388_));
 sg13g2_o21ai_1 _1848_ (.B1(_1389_),
    .Y(_0000_),
    .A1(_1386_),
    .A2(_1387_));
 sg13g2_buf_1 _1849_ (.A(_1375_),
    .X(_1390_));
 sg13g2_buf_2 _1850_ (.A(\rsa_unit_i.rsa_control_fsm.state[8] ),
    .X(_1391_));
 sg13g2_a22oi_1 _1851_ (.Y(_1392_),
    .B1(_1368_),
    .B2(_1391_),
    .A2(net49),
    .A1(net108));
 sg13g2_inv_1 _1852_ (.Y(_0015_),
    .A(_1392_));
 sg13g2_a22oi_1 _1853_ (.Y(_1393_),
    .B1(_1376_),
    .B2(\rsa_unit_i.rsa_control_fsm.state[0] ),
    .A2(net49),
    .A1(\rsa_unit_i.rsa_control_fsm.state[6] ));
 sg13g2_inv_1 _1854_ (.Y(_0016_),
    .A(_1393_));
 sg13g2_buf_2 _1855_ (.A(\rsa_unit_i.rsa_control_fsm.state[7] ),
    .X(_1394_));
 sg13g2_a22oi_1 _1856_ (.Y(_1395_),
    .B1(_1368_),
    .B2(_1328_),
    .A2(_1390_),
    .A1(_1394_));
 sg13g2_inv_1 _1857_ (.Y(_0017_),
    .A(_1395_));
 sg13g2_buf_2 _1858_ (.A(\rsa_unit_i.rsa_control_fsm.state[2] ),
    .X(_1396_));
 sg13g2_a21oi_1 _1859_ (.A1(_1391_),
    .A2(_1337_),
    .Y(_1397_),
    .B1(_1396_));
 sg13g2_buf_2 _1860_ (.A(_0054_),
    .X(_1398_));
 sg13g2_inv_1 _1861_ (.Y(_1399_),
    .A(_1398_));
 sg13g2_buf_1 _1862_ (.A(_1399_),
    .X(_1400_));
 sg13g2_buf_1 _1863_ (.A(net57),
    .X(_1401_));
 sg13g2_nand2_1 _1864_ (.Y(_1402_),
    .A(_1400_),
    .B(_1401_));
 sg13g2_o21ai_1 _1865_ (.B1(_1402_),
    .Y(_0018_),
    .A1(_1346_),
    .A2(_1397_));
 sg13g2_inv_1 _1866_ (.Y(_1403_),
    .A(net108));
 sg13g2_o21ai_1 _1867_ (.B1(_0051_),
    .Y(_1404_),
    .A1(_1403_),
    .A2(_1381_));
 sg13g2_a22oi_1 _1868_ (.Y(_1405_),
    .B1(_1376_),
    .B2(_1404_),
    .A2(_1390_),
    .A1(_1396_));
 sg13g2_inv_1 _1869_ (.Y(_0012_),
    .A(_1405_));
 sg13g2_a22oi_1 _1870_ (.Y(_1406_),
    .B1(_1343_),
    .B2(\rsa_unit_i.rsa_control_fsm.state[3] ),
    .A2(_1376_),
    .A1(\rsa_unit_i.rsa_control_fsm.state[6] ));
 sg13g2_inv_1 _1871_ (.Y(_0013_),
    .A(_1406_));
 sg13g2_nand2_1 _1872_ (.Y(_1407_),
    .A(_1394_),
    .B(_1376_));
 sg13g2_o21ai_1 _1873_ (.B1(_1407_),
    .Y(_0014_),
    .A1(_0055_),
    .A2(net58));
 sg13g2_nand2_1 _1874_ (.Y(_1408_),
    .A(\rsa_en_logic_i.state[2] ),
    .B(net87));
 sg13g2_nand2_1 _1875_ (.Y(_1409_),
    .A(\rsa_en_logic_i.state[5] ),
    .B(_1308_));
 sg13g2_o21ai_1 _1876_ (.B1(_1409_),
    .Y(_0004_),
    .A1(_1386_),
    .A2(_1408_));
 sg13g2_nand3_1 _1877_ (.B(net87),
    .C(net109),
    .A(_1330_),
    .Y(_1410_));
 sg13g2_nand2_1 _1878_ (.Y(_1411_),
    .A(_1329_),
    .B(_1308_));
 sg13g2_o21ai_1 _1879_ (.B1(_1411_),
    .Y(_0003_),
    .A1(_1386_),
    .A2(_1410_));
 sg13g2_inv_1 _1880_ (.Y(_1412_),
    .A(_1312_));
 sg13g2_nor2_1 _1881_ (.A(_1329_),
    .B(\rsa_en_logic_i.state[0] ),
    .Y(_1413_));
 sg13g2_o21ai_1 _1882_ (.B1(_1386_),
    .Y(_1414_),
    .A1(\rsa_en_logic_i.state[2] ),
    .A2(_1331_));
 sg13g2_nand2_1 _1883_ (.Y(_1415_),
    .A(_1413_),
    .B(_1414_));
 sg13g2_a22oi_1 _1884_ (.Y(_1416_),
    .B1(_1415_),
    .B2(net86),
    .A2(_1412_),
    .A1(\rsa_en_logic_i.state[3] ));
 sg13g2_inv_1 _1885_ (.Y(_0002_),
    .A(_1416_));
 sg13g2_buf_1 _1886_ (.A(net110),
    .X(_1417_));
 sg13g2_nand2_1 _1887_ (.Y(_1418_),
    .A(net85),
    .B(\gpio_wrapper_i.gpio_start_cmd_i.data ));
 sg13g2_o21ai_1 _1888_ (.B1(_1418_),
    .Y(_0121_),
    .A1(net86),
    .A2(_1309_));
 sg13g2_mux2_1 _1889_ (.A0(\gpio_wrapper_i.gpio_stop_cmd_i.data_dly ),
    .A1(\gpio_wrapper_i.gpio_stop_cmd_i.data ),
    .S(net86),
    .X(_0122_));
 sg13g2_mux2_1 _1890_ (.A0(\gpio_wrapper_i.sync_gpio_start.data_sync[1] ),
    .A1(net5),
    .S(net86),
    .X(_0123_));
 sg13g2_mux2_1 _1891_ (.A0(\gpio_wrapper_i.gpio_start_cmd_i.data ),
    .A1(\gpio_wrapper_i.sync_gpio_start.data_sync[1] ),
    .S(_1364_),
    .X(_0124_));
 sg13g2_mux2_1 _1892_ (.A0(\gpio_wrapper_i.sync_gpio_stop.data_sync[1] ),
    .A1(net6),
    .S(net85),
    .X(_0125_));
 sg13g2_nand2_1 _1893_ (.Y(_1419_),
    .A(net87),
    .B(\gpio_wrapper_i.sync_gpio_stop.data_sync[1] ));
 sg13g2_o21ai_1 _1894_ (.B1(_1419_),
    .Y(_0126_),
    .A1(net86),
    .A2(_1383_));
 sg13g2_a21oi_1 _1895_ (.A1(_1329_),
    .A2(net110),
    .Y(_1420_),
    .B1(irq));
 sg13g2_a21oi_1 _1896_ (.A1(net87),
    .A2(_1386_),
    .Y(_1421_),
    .B1(_1420_));
 sg13g2_nor2b_1 _1897_ (.A(_1312_),
    .B_N(_1421_),
    .Y(_0127_));
 sg13g2_nand2_1 _1898_ (.Y(_1422_),
    .A(net87),
    .B(\rsa_spi_wrapper_i.config_regs[8] ));
 sg13g2_o21ai_1 _1899_ (.B1(_1422_),
    .Y(_0128_),
    .A1(_1364_),
    .A2(_1310_));
 sg13g2_mux2_1 _1900_ (.A0(\rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly ),
    .A1(\rsa_spi_wrapper_i.config_regs[9] ),
    .S(net85),
    .X(_0129_));
 sg13g2_buf_1 _1901_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[0] ),
    .X(_1423_));
 sg13g2_buf_1 _1902_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[2] ),
    .X(_1424_));
 sg13g2_buf_1 _1903_ (.A(_1424_),
    .X(_1425_));
 sg13g2_buf_1 _1904_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[0] ),
    .X(_1426_));
 sg13g2_buf_1 _1905_ (.A(_1426_),
    .X(_1427_));
 sg13g2_nor2_1 _1906_ (.A(_1308_),
    .B(_1427_),
    .Y(_1428_));
 sg13g2_buf_1 _1907_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[1] ),
    .X(_1429_));
 sg13g2_buf_1 _1908_ (.A(_1429_),
    .X(_1430_));
 sg13g2_buf_1 _1909_ (.A(net82),
    .X(_1431_));
 sg13g2_buf_1 _1910_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o_vld ),
    .X(_1432_));
 sg13g2_nor2b_1 _1911_ (.A(net68),
    .B_N(_1432_),
    .Y(_1433_));
 sg13g2_nand2_1 _1912_ (.Y(_1434_),
    .A(_1428_),
    .B(_1433_));
 sg13g2_nor2_1 _1913_ (.A(net84),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_buf_4 _1914_ (.X(_1436_),
    .A(_1435_));
 sg13g2_mux2_1 _1915_ (.A0(\rsa_spi_wrapper_i.config_regs[0] ),
    .A1(net107),
    .S(_1436_),
    .X(_0130_));
 sg13g2_buf_1 _1916_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[1] ),
    .X(_1437_));
 sg13g2_mux2_1 _1917_ (.A0(\rsa_spi_wrapper_i.config_regs[1] ),
    .A1(net106),
    .S(_1436_),
    .X(_0131_));
 sg13g2_buf_1 _1918_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[2] ),
    .X(_1438_));
 sg13g2_mux2_1 _1919_ (.A0(\rsa_spi_wrapper_i.config_regs[2] ),
    .A1(net105),
    .S(_1436_),
    .X(_0132_));
 sg13g2_buf_1 _1920_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[3] ),
    .X(_1439_));
 sg13g2_mux2_1 _1921_ (.A0(\rsa_spi_wrapper_i.config_regs[3] ),
    .A1(net104),
    .S(_1436_),
    .X(_0133_));
 sg13g2_buf_1 _1922_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[4] ),
    .X(_1440_));
 sg13g2_mux2_1 _1923_ (.A0(\rsa_spi_wrapper_i.config_regs[4] ),
    .A1(net103),
    .S(_1436_),
    .X(_0134_));
 sg13g2_buf_1 _1924_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[5] ),
    .X(_1441_));
 sg13g2_mux2_1 _1925_ (.A0(\rsa_spi_wrapper_i.config_regs[5] ),
    .A1(_1441_),
    .S(_1436_),
    .X(_0135_));
 sg13g2_buf_1 _1926_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[6] ),
    .X(_1442_));
 sg13g2_mux2_1 _1927_ (.A0(\rsa_spi_wrapper_i.config_regs[6] ),
    .A1(_1442_),
    .S(_1436_),
    .X(_0136_));
 sg13g2_buf_1 _1928_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[7] ),
    .X(_1443_));
 sg13g2_mux2_1 _1929_ (.A0(\rsa_spi_wrapper_i.config_regs[7] ),
    .A1(net100),
    .S(_1436_),
    .X(_0137_));
 sg13g2_buf_1 _1930_ (.A(net83),
    .X(_1444_));
 sg13g2_buf_1 _1931_ (.A(net67),
    .X(_1445_));
 sg13g2_buf_2 _1932_ (.A(_0050_),
    .X(_1446_));
 sg13g2_buf_1 _1933_ (.A(_1446_),
    .X(_1447_));
 sg13g2_nand4_1 _1934_ (.B(net56),
    .C(net81),
    .A(net111),
    .Y(_1448_),
    .D(_1433_));
 sg13g2_buf_4 _1935_ (.X(_1449_),
    .A(_1448_));
 sg13g2_mux2_1 _1936_ (.A0(net107),
    .A1(\rsa_spi_wrapper_i.config_regs[8] ),
    .S(_1449_),
    .X(_0138_));
 sg13g2_mux2_1 _1937_ (.A0(net106),
    .A1(\rsa_spi_wrapper_i.config_regs[9] ),
    .S(_1449_),
    .X(_0139_));
 sg13g2_mux2_1 _1938_ (.A0(net105),
    .A1(\rsa_spi_wrapper_i.config_regs[10] ),
    .S(_1449_),
    .X(_0140_));
 sg13g2_mux2_1 _1939_ (.A0(net104),
    .A1(\rsa_spi_wrapper_i.config_regs[11] ),
    .S(_1449_),
    .X(_0141_));
 sg13g2_mux2_1 _1940_ (.A0(net103),
    .A1(\rsa_spi_wrapper_i.config_regs[12] ),
    .S(_1449_),
    .X(_0142_));
 sg13g2_mux2_1 _1941_ (.A0(net102),
    .A1(\rsa_spi_wrapper_i.config_regs[13] ),
    .S(_1449_),
    .X(_0143_));
 sg13g2_mux2_1 _1942_ (.A0(net101),
    .A1(\rsa_spi_wrapper_i.config_regs[14] ),
    .S(_1449_),
    .X(_0144_));
 sg13g2_mux2_1 _1943_ (.A0(net100),
    .A1(\rsa_spi_wrapper_i.config_regs[15] ),
    .S(_1449_),
    .X(_0145_));
 sg13g2_inv_1 _1944_ (.Y(_1450_),
    .A(_1429_));
 sg13g2_nor2_2 _1945_ (.A(_1450_),
    .B(net84),
    .Y(_1451_));
 sg13g2_and3_1 _1946_ (.X(_1452_),
    .A(_1432_),
    .B(_1428_),
    .C(_1451_));
 sg13g2_buf_1 _1947_ (.A(_1452_),
    .X(_1453_));
 sg13g2_mux2_1 _1948_ (.A0(\rsa_p[0] ),
    .A1(net107),
    .S(net47),
    .X(_0146_));
 sg13g2_buf_1 _1949_ (.A(\rsa_p[1] ),
    .X(_1454_));
 sg13g2_inv_1 _1950_ (.Y(_1455_),
    .A(net99));
 sg13g2_nand2_1 _1951_ (.Y(_1456_),
    .A(net106),
    .B(net47));
 sg13g2_o21ai_1 _1952_ (.B1(_1456_),
    .Y(_0147_),
    .A1(_1455_),
    .A2(net47));
 sg13g2_mux2_1 _1953_ (.A0(\rsa_p[2] ),
    .A1(net105),
    .S(net47),
    .X(_0148_));
 sg13g2_mux2_1 _1954_ (.A0(\rsa_p[3] ),
    .A1(net104),
    .S(net47),
    .X(_0149_));
 sg13g2_mux2_1 _1955_ (.A0(\rsa_p[4] ),
    .A1(net103),
    .S(_1453_),
    .X(_0150_));
 sg13g2_mux2_1 _1956_ (.A0(\rsa_p[5] ),
    .A1(net102),
    .S(net47),
    .X(_0151_));
 sg13g2_mux2_1 _1957_ (.A0(\rsa_p[6] ),
    .A1(net101),
    .S(net47),
    .X(_0152_));
 sg13g2_mux2_1 _1958_ (.A0(\rsa_p[7] ),
    .A1(net100),
    .S(net47),
    .X(_0153_));
 sg13g2_and4_1 _1959_ (.A(net111),
    .B(net56),
    .C(_1432_),
    .D(_1451_),
    .X(_1457_));
 sg13g2_buf_4 _1960_ (.X(_1458_),
    .A(_1457_));
 sg13g2_mux2_1 _1961_ (.A0(\rsa_e[0] ),
    .A1(net107),
    .S(_1458_),
    .X(_0154_));
 sg13g2_mux2_1 _1962_ (.A0(\rsa_e[1] ),
    .A1(net106),
    .S(_1458_),
    .X(_0155_));
 sg13g2_mux2_1 _1963_ (.A0(\rsa_e[2] ),
    .A1(net105),
    .S(_1458_),
    .X(_0156_));
 sg13g2_mux2_1 _1964_ (.A0(\rsa_e[3] ),
    .A1(net104),
    .S(_1458_),
    .X(_0157_));
 sg13g2_mux2_1 _1965_ (.A0(\rsa_e[4] ),
    .A1(net103),
    .S(_1458_),
    .X(_0158_));
 sg13g2_mux2_1 _1966_ (.A0(\rsa_e[5] ),
    .A1(net102),
    .S(_1458_),
    .X(_0159_));
 sg13g2_mux2_1 _1967_ (.A0(\rsa_e[6] ),
    .A1(net101),
    .S(_1458_),
    .X(_0160_));
 sg13g2_mux2_1 _1968_ (.A0(\rsa_e[7] ),
    .A1(net100),
    .S(_1458_),
    .X(_0161_));
 sg13g2_buf_2 _1969_ (.A(\rsa_spi_wrapper_i.config_regs[32] ),
    .X(_1459_));
 sg13g2_inv_2 _1970_ (.Y(_1460_),
    .A(_1459_));
 sg13g2_inv_1 _1971_ (.Y(_1461_),
    .A(_1424_));
 sg13g2_buf_1 _1972_ (.A(_1461_),
    .X(_1462_));
 sg13g2_nor2_1 _1973_ (.A(_1462_),
    .B(_1434_),
    .Y(_1463_));
 sg13g2_buf_1 _1974_ (.A(_1463_),
    .X(_1464_));
 sg13g2_nand2_1 _1975_ (.Y(_1465_),
    .A(net107),
    .B(net34));
 sg13g2_o21ai_1 _1976_ (.B1(_1465_),
    .Y(_0162_),
    .A1(_1460_),
    .A2(net34));
 sg13g2_buf_1 _1977_ (.A(\rsa_spi_wrapper_i.config_regs[33] ),
    .X(_1466_));
 sg13g2_inv_1 _1978_ (.Y(_1467_),
    .A(_1466_));
 sg13g2_nand2_1 _1979_ (.Y(_1468_),
    .A(net106),
    .B(_1464_));
 sg13g2_o21ai_1 _1980_ (.B1(_1468_),
    .Y(_0163_),
    .A1(_1467_),
    .A2(_1464_));
 sg13g2_mux2_1 _1981_ (.A0(\rsa_spi_wrapper_i.config_regs[34] ),
    .A1(net105),
    .S(net34),
    .X(_0164_));
 sg13g2_mux2_1 _1982_ (.A0(\rsa_spi_wrapper_i.config_regs[35] ),
    .A1(net104),
    .S(net34),
    .X(_0165_));
 sg13g2_mux2_1 _1983_ (.A0(\rsa_spi_wrapper_i.config_regs[36] ),
    .A1(net103),
    .S(net34),
    .X(_0166_));
 sg13g2_mux2_1 _1984_ (.A0(\rsa_spi_wrapper_i.config_regs[37] ),
    .A1(net102),
    .S(net34),
    .X(_0167_));
 sg13g2_mux2_1 _1985_ (.A0(\rsa_spi_wrapper_i.config_regs[38] ),
    .A1(net101),
    .S(net34),
    .X(_0168_));
 sg13g2_mux2_1 _1986_ (.A0(\rsa_spi_wrapper_i.config_regs[39] ),
    .A1(net100),
    .S(net34),
    .X(_0169_));
 sg13g2_inv_2 _1987_ (.Y(_1469_),
    .A(_1446_));
 sg13g2_buf_1 _1988_ (.A(_1469_),
    .X(_1470_));
 sg13g2_and4_1 _1989_ (.A(net111),
    .B(net56),
    .C(_1470_),
    .D(_1433_),
    .X(_1471_));
 sg13g2_buf_4 _1990_ (.X(_1472_),
    .A(_1471_));
 sg13g2_mux2_1 _1991_ (.A0(\rsa_const[0] ),
    .A1(_1423_),
    .S(_1472_),
    .X(_0170_));
 sg13g2_mux2_1 _1992_ (.A0(\rsa_const[1] ),
    .A1(net106),
    .S(_1472_),
    .X(_0171_));
 sg13g2_mux2_1 _1993_ (.A0(\rsa_const[2] ),
    .A1(net105),
    .S(_1472_),
    .X(_0172_));
 sg13g2_mux2_1 _1994_ (.A0(\rsa_const[3] ),
    .A1(net104),
    .S(_1472_),
    .X(_0173_));
 sg13g2_mux2_1 _1995_ (.A0(\rsa_const[4] ),
    .A1(_1440_),
    .S(_1472_),
    .X(_0174_));
 sg13g2_mux2_1 _1996_ (.A0(\rsa_const[5] ),
    .A1(net102),
    .S(_1472_),
    .X(_0175_));
 sg13g2_mux2_1 _1997_ (.A0(\rsa_const[6] ),
    .A1(net101),
    .S(_1472_),
    .X(_0176_));
 sg13g2_mux2_1 _1998_ (.A0(\rsa_const[7] ),
    .A1(_1443_),
    .S(_1472_),
    .X(_0177_));
 sg13g2_nor2_1 _1999_ (.A(_1450_),
    .B(_1446_),
    .Y(_1473_));
 sg13g2_buf_2 _2000_ (.A(_1473_),
    .X(_1474_));
 sg13g2_and3_1 _2001_ (.X(_1475_),
    .A(_1432_),
    .B(_1428_),
    .C(_1474_));
 sg13g2_buf_4 _2002_ (.X(_1476_),
    .A(_1475_));
 sg13g2_mux2_1 _2003_ (.A0(\rsa_spi_wrapper_i.config_regs[48] ),
    .A1(net107),
    .S(_1476_),
    .X(_0178_));
 sg13g2_mux2_1 _2004_ (.A0(\rsa_spi_wrapper_i.config_regs[49] ),
    .A1(_1437_),
    .S(_1476_),
    .X(_0179_));
 sg13g2_mux2_1 _2005_ (.A0(\rsa_spi_wrapper_i.config_regs[50] ),
    .A1(_1438_),
    .S(_1476_),
    .X(_0180_));
 sg13g2_mux2_1 _2006_ (.A0(\rsa_spi_wrapper_i.config_regs[51] ),
    .A1(net104),
    .S(_1476_),
    .X(_0181_));
 sg13g2_mux2_1 _2007_ (.A0(\rsa_spi_wrapper_i.config_regs[52] ),
    .A1(net103),
    .S(_1476_),
    .X(_0182_));
 sg13g2_mux2_1 _2008_ (.A0(\rsa_spi_wrapper_i.config_regs[53] ),
    .A1(net102),
    .S(_1476_),
    .X(_0183_));
 sg13g2_mux2_1 _2009_ (.A0(\rsa_spi_wrapper_i.config_regs[54] ),
    .A1(net101),
    .S(_1476_),
    .X(_0184_));
 sg13g2_mux2_1 _2010_ (.A0(\rsa_spi_wrapper_i.config_regs[55] ),
    .A1(net100),
    .S(_1476_),
    .X(_0185_));
 sg13g2_and4_1 _2011_ (.A(net111),
    .B(_1445_),
    .C(_1432_),
    .D(_1474_),
    .X(_1477_));
 sg13g2_buf_4 _2012_ (.X(_1478_),
    .A(_1477_));
 sg13g2_mux2_1 _2013_ (.A0(\rsa_spi_wrapper_i.config_regs[56] ),
    .A1(net107),
    .S(_1478_),
    .X(_0186_));
 sg13g2_mux2_1 _2014_ (.A0(\rsa_spi_wrapper_i.config_regs[57] ),
    .A1(net106),
    .S(_1478_),
    .X(_0187_));
 sg13g2_mux2_1 _2015_ (.A0(\rsa_spi_wrapper_i.config_regs[58] ),
    .A1(net105),
    .S(_1478_),
    .X(_0188_));
 sg13g2_mux2_1 _2016_ (.A0(\rsa_spi_wrapper_i.config_regs[59] ),
    .A1(_1439_),
    .S(_1478_),
    .X(_0189_));
 sg13g2_mux2_1 _2017_ (.A0(\rsa_spi_wrapper_i.config_regs[60] ),
    .A1(net103),
    .S(_1478_),
    .X(_0190_));
 sg13g2_mux2_1 _2018_ (.A0(\rsa_spi_wrapper_i.config_regs[61] ),
    .A1(net102),
    .S(_1478_),
    .X(_0191_));
 sg13g2_mux2_1 _2019_ (.A0(\rsa_spi_wrapper_i.config_regs[62] ),
    .A1(net101),
    .S(_1478_),
    .X(_0192_));
 sg13g2_mux2_1 _2020_ (.A0(\rsa_spi_wrapper_i.config_regs[63] ),
    .A1(net100),
    .S(_1478_),
    .X(_0193_));
 sg13g2_mux2_1 _2021_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .A1(_1445_),
    .S(_1367_),
    .X(_0194_));
 sg13g2_buf_1 _2022_ (.A(net68),
    .X(_1479_));
 sg13g2_mux2_1 _2023_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .A1(net55),
    .S(_1367_),
    .X(_0195_));
 sg13g2_mux2_1 _2024_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .A1(net84),
    .S(_1367_),
    .X(_0196_));
 sg13g2_buf_2 _2025_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[3] ),
    .X(_1480_));
 sg13g2_buf_1 _2026_ (.A(_1480_),
    .X(_1481_));
 sg13g2_mux2_1 _2027_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .A1(net80),
    .S(_1367_),
    .X(_0197_));
 sg13g2_nand3_1 _2028_ (.B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ),
    .C(_1355_),
    .A(_1307_),
    .Y(_1482_));
 sg13g2_buf_1 _2029_ (.A(_1482_),
    .X(_1483_));
 sg13g2_mux2_1 _2030_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .A1(net107),
    .S(net33),
    .X(_0198_));
 sg13g2_mux2_1 _2031_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .A1(net106),
    .S(_1483_),
    .X(_0199_));
 sg13g2_mux2_1 _2032_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .A1(net105),
    .S(net33),
    .X(_0200_));
 sg13g2_mux2_1 _2033_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .A1(net104),
    .S(net33),
    .X(_0201_));
 sg13g2_mux2_1 _2034_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .A1(net103),
    .S(net33),
    .X(_0202_));
 sg13g2_mux2_1 _2035_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .A1(net102),
    .S(net33),
    .X(_0203_));
 sg13g2_mux2_1 _2036_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .A1(net101),
    .S(net33),
    .X(_0204_));
 sg13g2_mux2_1 _2037_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .A1(net100),
    .S(net33),
    .X(_0205_));
 sg13g2_nand2_1 _2038_ (.Y(_1484_),
    .A(_1308_),
    .B(_1432_));
 sg13g2_o21ai_1 _2039_ (.B1(_1484_),
    .Y(_0206_),
    .A1(_1348_),
    .A2(net33));
 sg13g2_mux2_1 _2040_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ),
    .S(_1367_),
    .X(_0207_));
 sg13g2_mux2_1 _2041_ (.A0(_1317_),
    .A1(_1318_),
    .S(net85),
    .X(_0208_));
 sg13g2_mux2_1 _2042_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .A1(\rsa_spi_wrapper_i.spi_clk ),
    .S(net85),
    .X(_0209_));
 sg13g2_inv_1 _2043_ (.Y(_1485_),
    .A(\rsa_spi_wrapper_i.spi_clk ));
 sg13g2_nor3_1 _2044_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .B(_1485_),
    .C(_1360_),
    .Y(_1486_));
 sg13g2_buf_1 _2045_ (.A(_1486_),
    .X(_1487_));
 sg13g2_buf_1 _2046_ (.A(_1487_),
    .X(_1488_));
 sg13g2_mux2_1 _2047_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .A1(\rsa_spi_wrapper_i.spi_mosi ),
    .S(_1488_),
    .X(_0210_));
 sg13g2_mux2_1 _2048_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .S(net46),
    .X(_0211_));
 sg13g2_mux2_1 _2049_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .S(net46),
    .X(_0212_));
 sg13g2_mux2_1 _2050_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .S(net46),
    .X(_0213_));
 sg13g2_mux2_1 _2051_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .S(net46),
    .X(_0214_));
 sg13g2_mux2_1 _2052_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .S(net46),
    .X(_0215_));
 sg13g2_mux2_1 _2053_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .S(net46),
    .X(_0216_));
 sg13g2_mux2_1 _2054_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .S(net46),
    .X(_0217_));
 sg13g2_or3_1 _2055_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .B(_1485_),
    .C(_1360_),
    .X(_1489_));
 sg13g2_nor3_1 _2056_ (.A(_1351_),
    .B(_1355_),
    .C(_1489_),
    .Y(_1490_));
 sg13g2_a21o_1 _2057_ (.A2(_1489_),
    .A1(_1351_),
    .B1(_1490_),
    .X(_0218_));
 sg13g2_and2_1 _2058_ (.A(_1351_),
    .B(_1487_),
    .X(_1491_));
 sg13g2_buf_1 _2059_ (.A(_1491_),
    .X(_1492_));
 sg13g2_xor2_1 _2060_ (.B(_1492_),
    .A(_1350_),
    .X(_0219_));
 sg13g2_nand2_1 _2061_ (.Y(_1493_),
    .A(_1350_),
    .B(_1492_));
 sg13g2_xnor2_1 _2062_ (.Y(_0220_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .B(_1493_));
 sg13g2_a21oi_1 _2063_ (.A1(_1314_),
    .A2(_1352_),
    .Y(_1494_),
    .B1(_1349_));
 sg13g2_nor2_1 _2064_ (.A(_1350_),
    .B(_1494_),
    .Y(_1495_));
 sg13g2_nand4_1 _2065_ (.B(_1351_),
    .C(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .A(_1350_),
    .Y(_1496_),
    .D(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ));
 sg13g2_a21oi_1 _2066_ (.A1(_1353_),
    .A2(_1496_),
    .Y(_1497_),
    .B1(_1489_));
 sg13g2_a21oi_1 _2067_ (.A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .A2(_1492_),
    .Y(_1498_),
    .B1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_nor3_1 _2068_ (.A(_1495_),
    .B(_1497_),
    .C(_1498_),
    .Y(_0221_));
 sg13g2_a21oi_1 _2069_ (.A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .A2(_1485_),
    .Y(_1499_),
    .B1(_1317_));
 sg13g2_inv_1 _2070_ (.Y(_1500_),
    .A(_1320_));
 sg13g2_nand3_1 _2071_ (.B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ),
    .C(_1324_),
    .A(_1500_),
    .Y(_1501_));
 sg13g2_buf_1 _2072_ (.A(_1501_),
    .X(_1502_));
 sg13g2_o21ai_1 _2073_ (.B1(_1502_),
    .Y(_1503_),
    .A1(_1318_),
    .A2(_1499_));
 sg13g2_nand2_1 _2074_ (.Y(_1504_),
    .A(_1307_),
    .B(_1503_));
 sg13g2_buf_2 _2075_ (.A(_1504_),
    .X(_1505_));
 sg13g2_nand2_1 _2076_ (.Y(_1506_),
    .A(_1469_),
    .B(\rsa_spi_wrapper_i.config_regs[48] ));
 sg13g2_nand3_1 _2077_ (.B(net66),
    .C(\rsa_e[0] ),
    .A(net83),
    .Y(_1507_));
 sg13g2_o21ai_1 _2078_ (.B1(_1507_),
    .Y(_1508_),
    .A1(net83),
    .A2(_1506_));
 sg13g2_mux2_1 _2079_ (.A0(\rsa_const[0] ),
    .A1(\rsa_spi_wrapper_i.config_regs[8] ),
    .S(_1446_),
    .X(_1509_));
 sg13g2_a22oi_1 _2080_ (.Y(_1510_),
    .B1(_1509_),
    .B2(_1450_),
    .A2(_1474_),
    .A1(\rsa_spi_wrapper_i.config_regs[56] ));
 sg13g2_nor2_1 _2081_ (.A(_1429_),
    .B(_1461_),
    .Y(_1511_));
 sg13g2_buf_1 _2082_ (.A(_1511_),
    .X(_1512_));
 sg13g2_buf_2 _2083_ (.A(_0057_),
    .X(_1513_));
 sg13g2_inv_1 _2084_ (.Y(_1514_),
    .A(_1513_));
 sg13g2_a221oi_1 _2085_ (.B2(_1514_),
    .C1(_1427_),
    .B1(_1512_),
    .A1(\rsa_p[0] ),
    .Y(_1515_),
    .A2(_1451_));
 sg13g2_a21oi_1 _2086_ (.A1(_1444_),
    .A2(_1510_),
    .Y(_1516_),
    .B1(_1515_));
 sg13g2_a21oi_1 _2087_ (.A1(net55),
    .A2(_1508_),
    .Y(_1517_),
    .B1(_1516_));
 sg13g2_nor2_1 _2088_ (.A(_1426_),
    .B(net84),
    .Y(_1518_));
 sg13g2_inv_1 _2089_ (.Y(_1519_),
    .A(_1518_));
 sg13g2_nand3_1 _2090_ (.B(_1446_),
    .C(_1424_),
    .A(_1429_),
    .Y(_1520_));
 sg13g2_buf_1 _2091_ (.A(_1520_),
    .X(_1521_));
 sg13g2_o21ai_1 _2092_ (.B1(_1521_),
    .Y(_1522_),
    .A1(net82),
    .A2(_1519_));
 sg13g2_buf_2 _2093_ (.A(_1522_),
    .X(_1523_));
 sg13g2_mux2_1 _2094_ (.A0(_1517_),
    .A1(_0056_),
    .S(_1523_),
    .X(_1524_));
 sg13g2_inv_1 _2095_ (.Y(_1525_),
    .A(_1426_));
 sg13g2_nor2_1 _2096_ (.A(net81),
    .B(\rsa_c[0] ),
    .Y(_1526_));
 sg13g2_nand2b_1 _2097_ (.Y(_1527_),
    .B(_1425_),
    .A_N(_0058_));
 sg13g2_a22oi_1 _2098_ (.Y(_1528_),
    .B1(_1527_),
    .B2(net81),
    .A2(_1526_),
    .A1(net79));
 sg13g2_nor2b_1 _2099_ (.A(_1425_),
    .B_N(_0058_),
    .Y(_1529_));
 sg13g2_nor3_1 _2100_ (.A(net56),
    .B(_1479_),
    .C(_1529_),
    .Y(_1530_));
 sg13g2_a21oi_1 _2101_ (.A1(_1479_),
    .A2(_1528_),
    .Y(_1531_),
    .B1(_1530_));
 sg13g2_mux2_1 _2102_ (.A0(_1524_),
    .A1(_1531_),
    .S(net80),
    .X(_1532_));
 sg13g2_buf_1 _2103_ (.A(_1502_),
    .X(_1533_));
 sg13g2_nand2b_1 _2104_ (.Y(_1534_),
    .B(_1317_),
    .A_N(_1318_));
 sg13g2_nand2_1 _2105_ (.Y(_1535_),
    .A(net110),
    .B(_1534_));
 sg13g2_nor3_1 _2106_ (.A(_1532_),
    .B(net45),
    .C(_1535_),
    .Y(_1536_));
 sg13g2_a21o_1 _2107_ (.A2(_1505_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[0] ),
    .B1(_1536_),
    .X(_0222_));
 sg13g2_nand3_1 _2108_ (.B(_1534_),
    .C(_1503_),
    .A(net110),
    .Y(_1537_));
 sg13g2_buf_2 _2109_ (.A(_1537_),
    .X(_1538_));
 sg13g2_mux2_1 _2110_ (.A0(_0060_),
    .A1(_1455_),
    .S(_1430_),
    .X(_1539_));
 sg13g2_inv_1 _2111_ (.Y(_1540_),
    .A(_0061_));
 sg13g2_a22oi_1 _2112_ (.Y(_1541_),
    .B1(_1474_),
    .B2(\rsa_spi_wrapper_i.config_regs[49] ),
    .A2(_1512_),
    .A1(_1540_));
 sg13g2_o21ai_1 _2113_ (.B1(_1541_),
    .Y(_1542_),
    .A1(net84),
    .A2(_1539_));
 sg13g2_a22oi_1 _2114_ (.Y(_1543_),
    .B1(\rsa_e[1] ),
    .B2(net66),
    .A2(\rsa_spi_wrapper_i.config_regs[57] ),
    .A1(_1469_));
 sg13g2_and2_1 _2115_ (.A(net82),
    .B(_1543_),
    .X(_1544_));
 sg13g2_mux2_1 _2116_ (.A0(\rsa_const[1] ),
    .A1(\rsa_spi_wrapper_i.config_regs[9] ),
    .S(_1446_),
    .X(_1545_));
 sg13g2_nor2_1 _2117_ (.A(net68),
    .B(_1545_),
    .Y(_1546_));
 sg13g2_o21ai_1 _2118_ (.B1(_1444_),
    .Y(_1547_),
    .A1(_1544_),
    .A2(_1546_));
 sg13g2_o21ai_1 _2119_ (.B1(_1547_),
    .Y(_1548_),
    .A1(net56),
    .A2(_1542_));
 sg13g2_o21ai_1 _2120_ (.B1(_1548_),
    .Y(_1549_),
    .A1(_0060_),
    .A2(_1521_));
 sg13g2_o21ai_1 _2121_ (.B1(_1521_),
    .Y(_1550_),
    .A1(_1431_),
    .A2(_1447_));
 sg13g2_a21oi_1 _2122_ (.A1(_1470_),
    .A2(\rsa_c[1] ),
    .Y(_1551_),
    .B1(net56));
 sg13g2_o21ai_1 _2123_ (.B1(_1480_),
    .Y(_1552_),
    .A1(_1550_),
    .A2(_1551_));
 sg13g2_o21ai_1 _2124_ (.B1(_1552_),
    .Y(_1553_),
    .A1(net80),
    .A2(_1549_));
 sg13g2_mux2_1 _2125_ (.A0(_1553_),
    .A1(_0059_),
    .S(net45),
    .X(_1554_));
 sg13g2_nand2_1 _2126_ (.Y(_1555_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[1] ),
    .B(_1505_));
 sg13g2_o21ai_1 _2127_ (.B1(_1555_),
    .Y(_0223_),
    .A1(_1538_),
    .A2(_1554_));
 sg13g2_inv_1 _2128_ (.Y(_1556_),
    .A(\rsa_c[2] ));
 sg13g2_o21ai_1 _2129_ (.B1(net83),
    .Y(_1557_),
    .A1(net65),
    .A2(net66));
 sg13g2_o21ai_1 _2130_ (.B1(_1557_),
    .Y(_1558_),
    .A1(net81),
    .A2(_1556_));
 sg13g2_a22oi_1 _2131_ (.Y(_1559_),
    .B1(_1558_),
    .B2(net55),
    .A2(_1512_),
    .A1(net79));
 sg13g2_and2_1 _2132_ (.A(_1446_),
    .B(\rsa_spi_wrapper_i.config_regs[10] ),
    .X(_1560_));
 sg13g2_a21oi_1 _2133_ (.A1(net65),
    .A2(\rsa_const[2] ),
    .Y(_1561_),
    .B1(_1560_));
 sg13g2_a22oi_1 _2134_ (.Y(_1562_),
    .B1(\rsa_e[2] ),
    .B2(net66),
    .A2(\rsa_spi_wrapper_i.config_regs[58] ),
    .A1(net65));
 sg13g2_mux2_1 _2135_ (.A0(_1561_),
    .A1(_1562_),
    .S(net68),
    .X(_1563_));
 sg13g2_inv_2 _2136_ (.Y(_1564_),
    .A(_0064_));
 sg13g2_nor2b_1 _2137_ (.A(net84),
    .B_N(\rsa_p[2] ),
    .Y(_1565_));
 sg13g2_a21o_1 _2138_ (.A2(\rsa_spi_wrapper_i.config_regs[50] ),
    .A1(net65),
    .B1(_1565_),
    .X(_1566_));
 sg13g2_a221oi_1 _2139_ (.B2(_1431_),
    .C1(net67),
    .B1(_1566_),
    .A1(_1564_),
    .Y(_1567_),
    .A2(_1512_));
 sg13g2_a21oi_1 _2140_ (.A1(net56),
    .A2(_1563_),
    .Y(_1568_),
    .B1(_1567_));
 sg13g2_nor2b_1 _2141_ (.A(_0063_),
    .B_N(_1523_),
    .Y(_1569_));
 sg13g2_nor3_1 _2142_ (.A(_1480_),
    .B(_1568_),
    .C(_1569_),
    .Y(_1570_));
 sg13g2_a21oi_1 _2143_ (.A1(_1481_),
    .A2(_1559_),
    .Y(_1571_),
    .B1(_1570_));
 sg13g2_nand2_1 _2144_ (.Y(_1572_),
    .A(_0062_),
    .B(net45));
 sg13g2_o21ai_1 _2145_ (.B1(_1572_),
    .Y(_1573_),
    .A1(net45),
    .A2(_1571_));
 sg13g2_nand2_1 _2146_ (.Y(_1574_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[2] ),
    .B(_1505_));
 sg13g2_o21ai_1 _2147_ (.B1(_1574_),
    .Y(_0224_),
    .A1(_1538_),
    .A2(_1573_));
 sg13g2_inv_1 _2148_ (.Y(_1575_),
    .A(\rsa_c[3] ));
 sg13g2_o21ai_1 _2149_ (.B1(_1557_),
    .Y(_1576_),
    .A1(net81),
    .A2(_1575_));
 sg13g2_nor2_2 _2150_ (.A(net79),
    .B(_1446_),
    .Y(_1577_));
 sg13g2_nor3_1 _2151_ (.A(net55),
    .B(_1518_),
    .C(_1577_),
    .Y(_1578_));
 sg13g2_a21oi_1 _2152_ (.A1(net55),
    .A2(_1576_),
    .Y(_1579_),
    .B1(_1578_));
 sg13g2_nor2_1 _2153_ (.A(_1429_),
    .B(_1469_),
    .Y(_1580_));
 sg13g2_a22oi_1 _2154_ (.Y(_1581_),
    .B1(_1580_),
    .B2(\rsa_spi_wrapper_i.config_regs[11] ),
    .A2(_1451_),
    .A1(\rsa_e[3] ));
 sg13g2_nand3_1 _2155_ (.B(\rsa_spi_wrapper_i.config_regs[51] ),
    .C(_1474_),
    .A(net79),
    .Y(_1582_));
 sg13g2_o21ai_1 _2156_ (.B1(_1582_),
    .Y(_1583_),
    .A1(net79),
    .A2(_1581_));
 sg13g2_a22oi_1 _2157_ (.Y(_1584_),
    .B1(_1577_),
    .B2(\rsa_spi_wrapper_i.config_regs[59] ),
    .A2(_1518_),
    .A1(\rsa_p[3] ));
 sg13g2_buf_1 _2158_ (.A(_0067_),
    .X(_1585_));
 sg13g2_inv_2 _2159_ (.Y(_1586_),
    .A(net97));
 sg13g2_nor2_1 _2160_ (.A(_1426_),
    .B(_1461_),
    .Y(_1587_));
 sg13g2_a221oi_1 _2161_ (.B2(\rsa_const[3] ),
    .C1(net82),
    .B1(_1577_),
    .A1(_1586_),
    .Y(_1588_),
    .A2(_1587_));
 sg13g2_a21oi_1 _2162_ (.A1(net68),
    .A2(_1584_),
    .Y(_1589_),
    .B1(_1588_));
 sg13g2_nor3_1 _2163_ (.A(_1523_),
    .B(_1583_),
    .C(_1589_),
    .Y(_1590_));
 sg13g2_a21oi_1 _2164_ (.A1(_0066_),
    .A2(_1523_),
    .Y(_1591_),
    .B1(_1590_));
 sg13g2_nor2_1 _2165_ (.A(net80),
    .B(_1591_),
    .Y(_1592_));
 sg13g2_a21oi_1 _2166_ (.A1(net80),
    .A2(_1579_),
    .Y(_1593_),
    .B1(_1592_));
 sg13g2_nand2_1 _2167_ (.Y(_1594_),
    .A(_0065_),
    .B(_1533_));
 sg13g2_o21ai_1 _2168_ (.B1(_1594_),
    .Y(_1595_),
    .A1(_1533_),
    .A2(_1593_));
 sg13g2_nand2_1 _2169_ (.Y(_1596_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[3] ),
    .B(_1505_));
 sg13g2_o21ai_1 _2170_ (.B1(_1596_),
    .Y(_0225_),
    .A1(_1538_),
    .A2(_1595_));
 sg13g2_inv_1 _2171_ (.Y(_1597_),
    .A(_0068_));
 sg13g2_o21ai_1 _2172_ (.B1(net65),
    .Y(_1598_),
    .A1(net67),
    .A2(\rsa_c[4] ));
 sg13g2_and3_1 _2173_ (.X(_1599_),
    .A(net84),
    .B(_1480_),
    .C(_1598_));
 sg13g2_nor3_1 _2174_ (.A(net82),
    .B(net84),
    .C(_0069_),
    .Y(_1600_));
 sg13g2_a21oi_1 _2175_ (.A1(\rsa_spi_wrapper_i.config_regs[52] ),
    .A2(_1474_),
    .Y(_1601_),
    .B1(_1600_));
 sg13g2_or2_1 _2176_ (.X(_1602_),
    .B(_1521_),
    .A(_0069_));
 sg13g2_o21ai_1 _2177_ (.B1(_1602_),
    .Y(_1603_),
    .A1(net83),
    .A2(_1601_));
 sg13g2_a22oi_1 _2178_ (.Y(_1604_),
    .B1(\rsa_e[4] ),
    .B2(net66),
    .A2(\rsa_spi_wrapper_i.config_regs[60] ),
    .A1(net65));
 sg13g2_nor2_1 _2179_ (.A(net79),
    .B(_1604_),
    .Y(_1605_));
 sg13g2_and2_1 _2180_ (.A(\rsa_p[4] ),
    .B(_1518_),
    .X(_1606_));
 sg13g2_or4_1 _2181_ (.A(_1480_),
    .B(_1603_),
    .C(_1605_),
    .D(_1606_),
    .X(_1607_));
 sg13g2_buf_2 _2182_ (.A(_0070_),
    .X(_1608_));
 sg13g2_inv_2 _2183_ (.Y(_1609_),
    .A(_1608_));
 sg13g2_mux2_1 _2184_ (.A0(\rsa_const[4] ),
    .A1(\rsa_spi_wrapper_i.config_regs[12] ),
    .S(net81),
    .X(_1610_));
 sg13g2_a221oi_1 _2185_ (.B2(net67),
    .C1(_1603_),
    .B1(_1610_),
    .A1(_1609_),
    .Y(_1611_),
    .A2(_1587_));
 sg13g2_nor3_1 _2186_ (.A(net55),
    .B(_1480_),
    .C(_1611_),
    .Y(_1612_));
 sg13g2_a21oi_1 _2187_ (.A1(net55),
    .A2(_1607_),
    .Y(_1613_),
    .B1(_1612_));
 sg13g2_nor3_1 _2188_ (.A(_1502_),
    .B(_1599_),
    .C(_1613_),
    .Y(_1614_));
 sg13g2_a21oi_1 _2189_ (.A1(_1597_),
    .A2(net45),
    .Y(_1615_),
    .B1(_1614_));
 sg13g2_nand2_1 _2190_ (.Y(_1616_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[4] ),
    .B(_1505_));
 sg13g2_o21ai_1 _2191_ (.B1(_1616_),
    .Y(_0226_),
    .A1(_1538_),
    .A2(_1615_));
 sg13g2_nor2b_1 _2192_ (.A(_1426_),
    .B_N(net82),
    .Y(_1617_));
 sg13g2_nor2_1 _2193_ (.A(_1525_),
    .B(_1430_),
    .Y(_1618_));
 sg13g2_a22oi_1 _2194_ (.Y(_1619_),
    .B1(_1618_),
    .B2(\rsa_const[5] ),
    .A2(_1617_),
    .A1(\rsa_spi_wrapper_i.config_regs[53] ));
 sg13g2_nor2_1 _2195_ (.A(_1447_),
    .B(_1619_),
    .Y(_1620_));
 sg13g2_a22oi_1 _2196_ (.Y(_1621_),
    .B1(\rsa_e[5] ),
    .B2(_1462_),
    .A2(\rsa_spi_wrapper_i.config_regs[61] ),
    .A1(_1469_));
 sg13g2_nor2b_1 _2197_ (.A(_1621_),
    .B_N(net82),
    .Y(_1622_));
 sg13g2_a21oi_1 _2198_ (.A1(\rsa_spi_wrapper_i.config_regs[13] ),
    .A2(_1580_),
    .Y(_1623_),
    .B1(_1622_));
 sg13g2_buf_1 _2199_ (.A(_0073_),
    .X(_1624_));
 sg13g2_inv_1 _2200_ (.Y(_1625_),
    .A(net96));
 sg13g2_a221oi_1 _2201_ (.B2(_1625_),
    .C1(net83),
    .B1(_1512_),
    .A1(\rsa_p[5] ),
    .Y(_1626_),
    .A2(_1451_));
 sg13g2_a21oi_1 _2202_ (.A1(net67),
    .A2(_1623_),
    .Y(_1627_),
    .B1(_1626_));
 sg13g2_nor3_1 _2203_ (.A(_1523_),
    .B(_1620_),
    .C(_1627_),
    .Y(_0322_));
 sg13g2_a21oi_1 _2204_ (.A1(_0072_),
    .A2(_1523_),
    .Y(_0323_),
    .B1(_0322_));
 sg13g2_or2_1 _2205_ (.X(_0324_),
    .B(\rsa_c[5] ),
    .A(net67));
 sg13g2_a22oi_1 _2206_ (.Y(_0325_),
    .B1(_1474_),
    .B2(_0324_),
    .A2(_1512_),
    .A1(net79));
 sg13g2_nand2_1 _2207_ (.Y(_0326_),
    .A(net80),
    .B(_0325_));
 sg13g2_o21ai_1 _2208_ (.B1(_0326_),
    .Y(_0327_),
    .A1(_1481_),
    .A2(_0323_));
 sg13g2_mux2_1 _2209_ (.A0(_0327_),
    .A1(_0071_),
    .S(net45),
    .X(_0328_));
 sg13g2_nand2_1 _2210_ (.Y(_0329_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[5] ),
    .B(_1505_));
 sg13g2_o21ai_1 _2211_ (.B1(_0329_),
    .Y(_0227_),
    .A1(_1538_),
    .A2(_0328_));
 sg13g2_a22oi_1 _2212_ (.Y(_0330_),
    .B1(\rsa_e[6] ),
    .B2(net66),
    .A2(\rsa_spi_wrapper_i.config_regs[62] ),
    .A1(_1469_));
 sg13g2_nor2b_1 _2213_ (.A(_0330_),
    .B_N(net82),
    .Y(_0331_));
 sg13g2_a21oi_1 _2214_ (.A1(\rsa_spi_wrapper_i.config_regs[14] ),
    .A2(_1580_),
    .Y(_0332_),
    .B1(_0331_));
 sg13g2_buf_1 _2215_ (.A(_0076_),
    .X(_0333_));
 sg13g2_inv_1 _2216_ (.Y(_0334_),
    .A(net95));
 sg13g2_a221oi_1 _2217_ (.B2(_0334_),
    .C1(net67),
    .B1(_1512_),
    .A1(\rsa_p[6] ),
    .Y(_0335_),
    .A2(_1451_));
 sg13g2_a21oi_1 _2218_ (.A1(net67),
    .A2(_0332_),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_a22oi_1 _2219_ (.Y(_0337_),
    .B1(_1618_),
    .B2(\rsa_const[6] ),
    .A2(_1617_),
    .A1(\rsa_spi_wrapper_i.config_regs[54] ));
 sg13g2_nand2b_1 _2220_ (.Y(_0338_),
    .B(_1523_),
    .A_N(_0075_));
 sg13g2_o21ai_1 _2221_ (.B1(_0338_),
    .Y(_0339_),
    .A1(net81),
    .A2(_0337_));
 sg13g2_or3_1 _2222_ (.A(_1480_),
    .B(_0336_),
    .C(_0339_),
    .X(_0340_));
 sg13g2_a21oi_1 _2223_ (.A1(net65),
    .A2(\rsa_c[6] ),
    .Y(_0341_),
    .B1(net56));
 sg13g2_o21ai_1 _2224_ (.B1(_1480_),
    .Y(_0342_),
    .A1(_1550_),
    .A2(_0341_));
 sg13g2_a21oi_1 _2225_ (.A1(_0340_),
    .A2(_0342_),
    .Y(_0343_),
    .B1(_1502_));
 sg13g2_a21o_1 _2226_ (.A2(net45),
    .A1(_0074_),
    .B1(_0343_),
    .X(_0344_));
 sg13g2_nand2_1 _2227_ (.Y(_0345_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[6] ),
    .B(_1505_));
 sg13g2_o21ai_1 _2228_ (.B1(_0345_),
    .Y(_0228_),
    .A1(_1538_),
    .A2(_0344_));
 sg13g2_inv_1 _2229_ (.Y(_0346_),
    .A(\rsa_c[7] ));
 sg13g2_o21ai_1 _2230_ (.B1(_1557_),
    .Y(_0347_),
    .A1(net81),
    .A2(_0346_));
 sg13g2_a21oi_1 _2231_ (.A1(net55),
    .A2(_0347_),
    .Y(_0348_),
    .B1(_1578_));
 sg13g2_buf_1 _2232_ (.A(_0079_),
    .X(_0349_));
 sg13g2_inv_2 _2233_ (.Y(_0350_),
    .A(net94));
 sg13g2_nor2_1 _2234_ (.A(net79),
    .B(net65),
    .Y(_0351_));
 sg13g2_a221oi_1 _2235_ (.B2(\rsa_spi_wrapper_i.config_regs[15] ),
    .C1(net68),
    .B1(_0351_),
    .A1(_0350_),
    .Y(_0352_),
    .A2(_1587_));
 sg13g2_nand2_1 _2236_ (.Y(_0353_),
    .A(net66),
    .B(\rsa_e[7] ));
 sg13g2_a221oi_1 _2237_ (.B2(net66),
    .C1(net83),
    .B1(\rsa_p[7] ),
    .A1(_1469_),
    .Y(_0354_),
    .A2(\rsa_spi_wrapper_i.config_regs[55] ));
 sg13g2_a21oi_1 _2238_ (.A1(net83),
    .A2(_0353_),
    .Y(_0355_),
    .B1(_0354_));
 sg13g2_nor2b_1 _2239_ (.A(_0355_),
    .B_N(net68),
    .Y(_0356_));
 sg13g2_inv_1 _2240_ (.Y(_0357_),
    .A(_0078_));
 sg13g2_mux2_1 _2241_ (.A0(\rsa_const[7] ),
    .A1(\rsa_spi_wrapper_i.config_regs[63] ),
    .S(net68),
    .X(_0358_));
 sg13g2_a22oi_1 _2242_ (.Y(_0359_),
    .B1(_1577_),
    .B2(_0358_),
    .A2(_1523_),
    .A1(_0357_));
 sg13g2_o21ai_1 _2243_ (.B1(_0359_),
    .Y(_0360_),
    .A1(_0352_),
    .A2(_0356_));
 sg13g2_nor2_1 _2244_ (.A(net80),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_a21oi_1 _2245_ (.A1(net80),
    .A2(_0348_),
    .Y(_0362_),
    .B1(_0361_));
 sg13g2_nand2_1 _2246_ (.Y(_0363_),
    .A(_0077_),
    .B(_1502_));
 sg13g2_o21ai_1 _2247_ (.B1(_0363_),
    .Y(_0364_),
    .A1(net45),
    .A2(_0362_));
 sg13g2_nand2_1 _2248_ (.Y(_0365_),
    .A(\rsa_spi_wrapper_i.spi_miso ),
    .B(_1505_));
 sg13g2_o21ai_1 _2249_ (.B1(_0365_),
    .Y(_0229_),
    .A1(_1538_),
    .A2(_0364_));
 sg13g2_nor2_1 _2250_ (.A(_1321_),
    .B(_1323_),
    .Y(_0366_));
 sg13g2_a21oi_1 _2251_ (.A1(_1320_),
    .A2(_0366_),
    .Y(_0367_),
    .B1(_1322_));
 sg13g2_mux2_1 _2252_ (.A0(_1322_),
    .A1(_0367_),
    .S(_1488_),
    .X(_0230_));
 sg13g2_nand2_1 _2253_ (.Y(_0368_),
    .A(_1322_),
    .B(_1487_));
 sg13g2_xnor2_1 _2254_ (.Y(_0231_),
    .A(_1321_),
    .B(_0368_));
 sg13g2_nand3_1 _2255_ (.B(_1322_),
    .C(_1487_),
    .A(_1321_),
    .Y(_0369_));
 sg13g2_xnor2_1 _2256_ (.Y(_0232_),
    .A(_1323_),
    .B(_0369_));
 sg13g2_nand4_1 _2257_ (.B(_1322_),
    .C(_1323_),
    .A(_1321_),
    .Y(_0370_),
    .D(_1320_));
 sg13g2_nand2b_1 _2258_ (.Y(_0371_),
    .B(_0370_),
    .A_N(_1324_));
 sg13g2_nand3_1 _2259_ (.B(_1323_),
    .C(_1487_),
    .A(_1322_),
    .Y(_0372_));
 sg13g2_or3_1 _2260_ (.A(_1322_),
    .B(_1323_),
    .C(_1308_),
    .X(_0373_));
 sg13g2_a21oi_1 _2261_ (.A1(_1320_),
    .A2(_0373_),
    .Y(_0374_),
    .B1(_1321_));
 sg13g2_a221oi_1 _2262_ (.B2(_1500_),
    .C1(_0374_),
    .B1(_0372_),
    .A1(net46),
    .Y(_0233_),
    .A2(_0371_));
 sg13g2_buf_1 _2263_ (.A(\rsa_unit_i.rsa_control_fsm.load_exp ),
    .X(_0375_));
 sg13g2_nor4_1 _2264_ (.A(net108),
    .B(net109),
    .C(_1394_),
    .D(net93),
    .Y(_0376_));
 sg13g2_or4_1 _2265_ (.A(net109),
    .B(_1328_),
    .C(_1394_),
    .D(\rsa_unit_i.rsa_control_fsm.state[11] ),
    .X(_0377_));
 sg13g2_buf_1 _2266_ (.A(_0377_),
    .X(_0378_));
 sg13g2_buf_8 _2267_ (.A(_0378_),
    .X(_0379_));
 sg13g2_or3_1 _2268_ (.A(_1374_),
    .B(_1391_),
    .C(_1396_),
    .X(_0380_));
 sg13g2_buf_1 _2269_ (.A(_0380_),
    .X(_0381_));
 sg13g2_nor2_1 _2270_ (.A(net54),
    .B(net64),
    .Y(_0382_));
 sg13g2_buf_1 _2271_ (.A(_0382_),
    .X(_0383_));
 sg13g2_buf_1 _2272_ (.A(net39),
    .X(_0384_));
 sg13g2_nor3_2 _2273_ (.A(\rsa_unit_i.rsa_control_fsm.state[3] ),
    .B(net93),
    .C(\rsa_unit_i.rsa_control_fsm.state[6] ),
    .Y(_0385_));
 sg13g2_nand2_1 _2274_ (.Y(_0386_),
    .A(net32),
    .B(_0385_));
 sg13g2_nand2_1 _2275_ (.Y(_0387_),
    .A(net58),
    .B(_0386_));
 sg13g2_or2_1 _2276_ (.X(_0388_),
    .B(_0387_),
    .A(_0376_));
 sg13g2_buf_1 _2277_ (.A(_0388_),
    .X(_0389_));
 sg13g2_buf_1 _2278_ (.A(_0389_),
    .X(_0390_));
 sg13g2_buf_1 _2279_ (.A(_0042_),
    .X(_0391_));
 sg13g2_inv_1 _2280_ (.Y(_0392_),
    .A(_0391_));
 sg13g2_buf_1 _2281_ (.A(_1398_),
    .X(_0393_));
 sg13g2_nor2_2 _2282_ (.A(net108),
    .B(_1396_),
    .Y(_0394_));
 sg13g2_buf_1 _2283_ (.A(_0394_),
    .X(_0395_));
 sg13g2_nand2_1 _2284_ (.Y(_0396_),
    .A(net78),
    .B(net63));
 sg13g2_nor4_2 _2285_ (.A(net109),
    .B(_1328_),
    .C(_1394_),
    .Y(_0397_),
    .D(\rsa_unit_i.rsa_control_fsm.state[11] ));
 sg13g2_buf_8 _2286_ (.A(_0397_),
    .X(_0398_));
 sg13g2_nand2_1 _2287_ (.Y(_0399_),
    .A(net62),
    .B(_0385_));
 sg13g2_a21oi_1 _2288_ (.A1(\rsa_unit_i.rsa_control_fsm.exp[0] ),
    .A2(_0396_),
    .Y(_0400_),
    .B1(_0399_));
 sg13g2_buf_1 _2289_ (.A(_0400_),
    .X(_0401_));
 sg13g2_buf_1 _2290_ (.A(\rsa_unit_i.R_i[0] ),
    .X(_0402_));
 sg13g2_or2_1 _2291_ (.X(_0403_),
    .B(_1396_),
    .A(net108));
 sg13g2_buf_1 _2292_ (.A(_0403_),
    .X(_0404_));
 sg13g2_buf_1 _2293_ (.A(_0404_),
    .X(_0405_));
 sg13g2_nor2_1 _2294_ (.A(_1399_),
    .B(net53),
    .Y(_0406_));
 sg13g2_buf_1 _2295_ (.A(_0406_),
    .X(_0407_));
 sg13g2_nor3_2 _2296_ (.A(net109),
    .B(_1328_),
    .C(_1394_),
    .Y(_0408_));
 sg13g2_nor2b_1 _2297_ (.A(\rsa_unit_i.rsa_control_fsm.state[10] ),
    .B_N(_0052_),
    .Y(_0409_));
 sg13g2_buf_1 _2298_ (.A(_0409_),
    .X(_0410_));
 sg13g2_nand2_1 _2299_ (.Y(_0411_),
    .A(_0408_),
    .B(_0410_));
 sg13g2_buf_2 _2300_ (.A(_0411_),
    .X(_0412_));
 sg13g2_nor2_1 _2301_ (.A(net37),
    .B(_0412_),
    .Y(_0413_));
 sg13g2_buf_1 _2302_ (.A(_0413_),
    .X(_0414_));
 sg13g2_and2_1 _2303_ (.A(_0408_),
    .B(_0410_),
    .X(_0415_));
 sg13g2_buf_1 _2304_ (.A(_0415_),
    .X(_0416_));
 sg13g2_buf_1 _2305_ (.A(net52),
    .X(_0417_));
 sg13g2_nand2b_1 _2306_ (.Y(_0418_),
    .B(net44),
    .A_N(\rsa_const[0] ));
 sg13g2_buf_1 _2307_ (.A(net37),
    .X(_0419_));
 sg13g2_a22oi_1 _2308_ (.Y(_0420_),
    .B1(_0418_),
    .B2(net31),
    .A2(_0414_),
    .A1(_0402_));
 sg13g2_nand2_1 _2309_ (.Y(_0421_),
    .A(net38),
    .B(_0420_));
 sg13g2_o21ai_1 _2310_ (.B1(_0421_),
    .Y(_0422_),
    .A1(_0392_),
    .A2(net38));
 sg13g2_a21o_1 _2311_ (.A2(_0386_),
    .A1(_0376_),
    .B1(_1344_),
    .X(_0423_));
 sg13g2_buf_1 _2312_ (.A(_0423_),
    .X(_0424_));
 sg13g2_buf_1 _2313_ (.A(_0424_),
    .X(_0425_));
 sg13g2_nand2_1 _2314_ (.Y(_0426_),
    .A(_0402_),
    .B(net22));
 sg13g2_o21ai_1 _2315_ (.B1(_0426_),
    .Y(_0253_),
    .A1(net17),
    .A2(_0422_));
 sg13g2_nand2_1 _2316_ (.Y(_0427_),
    .A(\rsa_const[1] ),
    .B(_0419_));
 sg13g2_o21ai_1 _2317_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0025_),
    .A2(_0419_));
 sg13g2_nand2_1 _2318_ (.Y(_0429_),
    .A(net44),
    .B(_0428_));
 sg13g2_mux2_1 _2319_ (.A0(_0041_),
    .A1(_0429_),
    .S(_0401_),
    .X(_0430_));
 sg13g2_nand2_1 _2320_ (.Y(_0431_),
    .A(\rsa_unit_i.R_i[1] ),
    .B(net22));
 sg13g2_o21ai_1 _2321_ (.B1(_0431_),
    .Y(_0254_),
    .A1(net17),
    .A2(_0430_));
 sg13g2_nand2_1 _2322_ (.Y(_0432_),
    .A(\rsa_const[2] ),
    .B(net31));
 sg13g2_o21ai_1 _2323_ (.B1(_0432_),
    .Y(_0433_),
    .A1(_0027_),
    .A2(net31));
 sg13g2_nand2_1 _2324_ (.Y(_0434_),
    .A(net44),
    .B(_0433_));
 sg13g2_mux2_1 _2325_ (.A0(_0043_),
    .A1(_0434_),
    .S(net38),
    .X(_0435_));
 sg13g2_nand2_1 _2326_ (.Y(_0436_),
    .A(\rsa_unit_i.R_i[2] ),
    .B(net22));
 sg13g2_o21ai_1 _2327_ (.B1(_0436_),
    .Y(_0255_),
    .A1(net17),
    .A2(_0435_));
 sg13g2_buf_1 _2328_ (.A(_0044_),
    .X(_0437_));
 sg13g2_nand2_1 _2329_ (.Y(_0438_),
    .A(\rsa_const[3] ),
    .B(net37));
 sg13g2_o21ai_1 _2330_ (.B1(_0438_),
    .Y(_0439_),
    .A1(_0029_),
    .A2(net31));
 sg13g2_nand2_1 _2331_ (.Y(_0440_),
    .A(net44),
    .B(_0439_));
 sg13g2_mux2_1 _2332_ (.A0(_0437_),
    .A1(_0440_),
    .S(net38),
    .X(_0441_));
 sg13g2_nand2_1 _2333_ (.Y(_0442_),
    .A(\rsa_unit_i.R_i[3] ),
    .B(net22));
 sg13g2_o21ai_1 _2334_ (.B1(_0442_),
    .Y(_0256_),
    .A1(net17),
    .A2(_0441_));
 sg13g2_buf_1 _2335_ (.A(_0045_),
    .X(_0443_));
 sg13g2_nand2_1 _2336_ (.Y(_0444_),
    .A(\rsa_const[4] ),
    .B(net37));
 sg13g2_o21ai_1 _2337_ (.B1(_0444_),
    .Y(_0445_),
    .A1(_0031_),
    .A2(net31));
 sg13g2_nand2_1 _2338_ (.Y(_0446_),
    .A(_0417_),
    .B(_0445_));
 sg13g2_mux2_1 _2339_ (.A0(_0443_),
    .A1(_0446_),
    .S(net38),
    .X(_0447_));
 sg13g2_nand2_1 _2340_ (.Y(_0448_),
    .A(\rsa_unit_i.R_i[4] ),
    .B(_0425_));
 sg13g2_o21ai_1 _2341_ (.B1(_0448_),
    .Y(_0257_),
    .A1(_0390_),
    .A2(_0447_));
 sg13g2_nand2_1 _2342_ (.Y(_0449_),
    .A(\rsa_const[5] ),
    .B(_0407_));
 sg13g2_o21ai_1 _2343_ (.B1(_0449_),
    .Y(_0450_),
    .A1(_0033_),
    .A2(net31));
 sg13g2_nand2_1 _2344_ (.Y(_0451_),
    .A(_0417_),
    .B(_0450_));
 sg13g2_mux2_1 _2345_ (.A0(_0046_),
    .A1(_0451_),
    .S(_0401_),
    .X(_0452_));
 sg13g2_nand2_1 _2346_ (.Y(_0453_),
    .A(\rsa_unit_i.R_i[5] ),
    .B(net22));
 sg13g2_o21ai_1 _2347_ (.B1(_0453_),
    .Y(_0258_),
    .A1(_0390_),
    .A2(_0452_));
 sg13g2_nand2_1 _2348_ (.Y(_0454_),
    .A(\rsa_const[6] ),
    .B(net37));
 sg13g2_o21ai_1 _2349_ (.B1(_0454_),
    .Y(_0455_),
    .A1(_0035_),
    .A2(net31));
 sg13g2_nand2_1 _2350_ (.Y(_0456_),
    .A(net44),
    .B(_0455_));
 sg13g2_mux2_1 _2351_ (.A0(_0047_),
    .A1(_0456_),
    .S(net38),
    .X(_0457_));
 sg13g2_nand2_1 _2352_ (.Y(_0458_),
    .A(\rsa_unit_i.R_i[6] ),
    .B(_0425_));
 sg13g2_o21ai_1 _2353_ (.B1(_0458_),
    .Y(_0259_),
    .A1(net17),
    .A2(_0457_));
 sg13g2_buf_1 _2354_ (.A(_0048_),
    .X(_0459_));
 sg13g2_nand2_1 _2355_ (.Y(_0460_),
    .A(\rsa_const[7] ),
    .B(net37));
 sg13g2_o21ai_1 _2356_ (.B1(_0460_),
    .Y(_0461_),
    .A1(_0037_),
    .A2(net31));
 sg13g2_nand2_1 _2357_ (.Y(_0462_),
    .A(net44),
    .B(_0461_));
 sg13g2_mux2_1 _2358_ (.A0(_0459_),
    .A1(_0462_),
    .S(net38),
    .X(_0463_));
 sg13g2_nand2_1 _2359_ (.Y(_0464_),
    .A(\rsa_unit_i.R_i[7] ),
    .B(net22));
 sg13g2_o21ai_1 _2360_ (.B1(_0464_),
    .Y(_0260_),
    .A1(net17),
    .A2(_0463_));
 sg13g2_buf_1 _2361_ (.A(_0049_),
    .X(_0465_));
 sg13g2_nand2b_1 _2362_ (.Y(_0466_),
    .B(net29),
    .A_N(_0039_));
 sg13g2_mux2_1 _2363_ (.A0(_0465_),
    .A1(_0466_),
    .S(_0400_),
    .X(_0467_));
 sg13g2_nand2_1 _2364_ (.Y(_0468_),
    .A(\rsa_unit_i.R_i[8] ),
    .B(net22));
 sg13g2_o21ai_1 _2365_ (.B1(_0468_),
    .Y(_0261_),
    .A1(net17),
    .A2(_0467_));
 sg13g2_nand3b_1 _2366_ (.B(net38),
    .C(net29),
    .Y(_0469_),
    .A_N(_0040_));
 sg13g2_nand2_1 _2367_ (.Y(_0470_),
    .A(\rsa_unit_i.R_i[9] ),
    .B(net22));
 sg13g2_o21ai_1 _2368_ (.B1(_0470_),
    .Y(_0262_),
    .A1(net17),
    .A2(_0469_));
 sg13g2_nor3_1 _2369_ (.A(net108),
    .B(_1391_),
    .C(_1396_),
    .Y(_0471_));
 sg13g2_buf_1 _2370_ (.A(_0471_),
    .X(_0472_));
 sg13g2_nand2_1 _2371_ (.Y(_0473_),
    .A(net61),
    .B(_0385_));
 sg13g2_buf_1 _2372_ (.A(_0473_),
    .X(_0474_));
 sg13g2_buf_1 _2373_ (.A(_0474_),
    .X(_0475_));
 sg13g2_inv_1 _2374_ (.Y(_0476_),
    .A(_0081_));
 sg13g2_a21oi_2 _2375_ (.B1(_0476_),
    .Y(_0477_),
    .A2(net61),
    .A1(net62));
 sg13g2_a21oi_1 _2376_ (.A1(_0082_),
    .A2(net32),
    .Y(_0478_),
    .B1(_0477_));
 sg13g2_nand2_1 _2377_ (.Y(_0479_),
    .A(_0106_),
    .B(_0474_));
 sg13g2_o21ai_1 _2378_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0475_),
    .A2(_0478_));
 sg13g2_buf_1 _2379_ (.A(_0424_),
    .X(_0481_));
 sg13g2_nand2_1 _2380_ (.Y(_0482_),
    .A(\rsa_unit_i.P_i[0] ),
    .B(net21));
 sg13g2_o21ai_1 _2381_ (.B1(_0482_),
    .Y(_0282_),
    .A1(net23),
    .A2(_0480_));
 sg13g2_inv_1 _2382_ (.Y(_0483_),
    .A(_0104_));
 sg13g2_mux2_1 _2383_ (.A0(_0084_),
    .A1(_0085_),
    .S(net32),
    .X(_0484_));
 sg13g2_nor2_1 _2384_ (.A(_0474_),
    .B(_0484_),
    .Y(_0485_));
 sg13g2_a21oi_1 _2385_ (.A1(_0483_),
    .A2(net36),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_buf_1 _2386_ (.A(\rsa_unit_i.P_i[1] ),
    .X(_0487_));
 sg13g2_nand2_1 _2387_ (.Y(_0488_),
    .A(net92),
    .B(net21));
 sg13g2_o21ai_1 _2388_ (.B1(_0488_),
    .Y(_0283_),
    .A1(net23),
    .A2(_0486_));
 sg13g2_inv_1 _2389_ (.Y(_0489_),
    .A(_0088_));
 sg13g2_nand2_1 _2390_ (.Y(_0490_),
    .A(net62),
    .B(net61));
 sg13g2_buf_1 _2391_ (.A(_0490_),
    .X(_0491_));
 sg13g2_buf_1 _2392_ (.A(net43),
    .X(_0492_));
 sg13g2_o21ai_1 _2393_ (.B1(_0087_),
    .Y(_0493_),
    .A1(_0378_),
    .A2(net64));
 sg13g2_buf_1 _2394_ (.A(_0493_),
    .X(_0494_));
 sg13g2_o21ai_1 _2395_ (.B1(_0494_),
    .Y(_0495_),
    .A1(_0489_),
    .A2(net35));
 sg13g2_mux2_1 _2396_ (.A0(_0495_),
    .A1(_0107_),
    .S(net36),
    .X(_0496_));
 sg13g2_nand2_1 _2397_ (.Y(_0497_),
    .A(\rsa_unit_i.P_i[2] ),
    .B(net21));
 sg13g2_o21ai_1 _2398_ (.B1(_0497_),
    .Y(_0284_),
    .A1(net23),
    .A2(_0496_));
 sg13g2_inv_1 _2399_ (.Y(_0498_),
    .A(_0090_));
 sg13g2_a21oi_1 _2400_ (.A1(net62),
    .A2(net61),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_a21o_1 _2401_ (.A2(_0384_),
    .A1(_0091_),
    .B1(_0499_),
    .X(_0500_));
 sg13g2_mux2_1 _2402_ (.A0(_0500_),
    .A1(_0109_),
    .S(net36),
    .X(_0501_));
 sg13g2_nand2_1 _2403_ (.Y(_0502_),
    .A(\rsa_unit_i.P_i[3] ),
    .B(net21));
 sg13g2_o21ai_1 _2404_ (.B1(_0502_),
    .Y(_0285_),
    .A1(net23),
    .A2(_0501_));
 sg13g2_buf_1 _2405_ (.A(_0111_),
    .X(_0503_));
 sg13g2_inv_1 _2406_ (.Y(_0504_),
    .A(_0503_));
 sg13g2_inv_1 _2407_ (.Y(_0505_),
    .A(_0093_));
 sg13g2_a21oi_1 _2408_ (.A1(net62),
    .A2(net61),
    .Y(_0506_),
    .B1(_0505_));
 sg13g2_a21o_1 _2409_ (.A2(_0384_),
    .A1(_0094_),
    .B1(_0506_),
    .X(_0507_));
 sg13g2_nor2_1 _2410_ (.A(_0474_),
    .B(_0507_),
    .Y(_0508_));
 sg13g2_a21oi_1 _2411_ (.A1(_0504_),
    .A2(net36),
    .Y(_0509_),
    .B1(_0508_));
 sg13g2_nand2_1 _2412_ (.Y(_0510_),
    .A(\rsa_unit_i.P_i[4] ),
    .B(_0481_));
 sg13g2_o21ai_1 _2413_ (.B1(_0510_),
    .Y(_0286_),
    .A1(net23),
    .A2(_0509_));
 sg13g2_mux2_1 _2414_ (.A0(_0096_),
    .A1(_0097_),
    .S(net32),
    .X(_0511_));
 sg13g2_buf_1 _2415_ (.A(_0113_),
    .X(_0512_));
 sg13g2_mux2_1 _2416_ (.A0(_0511_),
    .A1(_0512_),
    .S(_0475_),
    .X(_0513_));
 sg13g2_nand2_1 _2417_ (.Y(_0514_),
    .A(\rsa_unit_i.P_i[5] ),
    .B(_0481_));
 sg13g2_o21ai_1 _2418_ (.B1(_0514_),
    .Y(_0287_),
    .A1(_0389_),
    .A2(_0513_));
 sg13g2_and2_1 _2419_ (.A(_0099_),
    .B(net43),
    .X(_0515_));
 sg13g2_a21o_1 _2420_ (.A2(net32),
    .A1(_0100_),
    .B1(_0515_),
    .X(_0516_));
 sg13g2_mux2_1 _2421_ (.A0(_0516_),
    .A1(_0115_),
    .S(net36),
    .X(_0517_));
 sg13g2_nand2_1 _2422_ (.Y(_0518_),
    .A(\rsa_unit_i.P_i[6] ),
    .B(net21));
 sg13g2_o21ai_1 _2423_ (.B1(_0518_),
    .Y(_0288_),
    .A1(net23),
    .A2(_0517_));
 sg13g2_buf_1 _2424_ (.A(_0020_),
    .X(_0519_));
 sg13g2_inv_1 _2425_ (.Y(_0520_),
    .A(_0519_));
 sg13g2_and2_1 _2426_ (.A(_0102_),
    .B(net43),
    .X(_0521_));
 sg13g2_a21o_1 _2427_ (.A2(net32),
    .A1(_0103_),
    .B1(_0521_),
    .X(_0522_));
 sg13g2_nor2_1 _2428_ (.A(_0474_),
    .B(_0522_),
    .Y(_0523_));
 sg13g2_a21oi_1 _2429_ (.A1(_0520_),
    .A2(net36),
    .Y(_0524_),
    .B1(_0523_));
 sg13g2_nand2_1 _2430_ (.Y(_0525_),
    .A(\rsa_unit_i.P_i[7] ),
    .B(net21));
 sg13g2_o21ai_1 _2431_ (.B1(_0525_),
    .Y(_0289_),
    .A1(net23),
    .A2(_0524_));
 sg13g2_buf_2 _2432_ (.A(\rsa_unit_i.P_i[8] ),
    .X(_0526_));
 sg13g2_nand2_2 _2433_ (.Y(_0527_),
    .A(_0526_),
    .B(net43));
 sg13g2_nor2_1 _2434_ (.A(_0474_),
    .B(_0527_),
    .Y(_0528_));
 sg13g2_a21oi_1 _2435_ (.A1(\rsa_unit_i.mmm_square.adder2.gen_fa[8].fa.HA1.a ),
    .A2(net36),
    .Y(_0529_),
    .B1(_0528_));
 sg13g2_nand2_1 _2436_ (.Y(_0530_),
    .A(_0526_),
    .B(net21));
 sg13g2_o21ai_1 _2437_ (.B1(_0530_),
    .Y(_0290_),
    .A1(net23),
    .A2(_0529_));
 sg13g2_nor2_1 _2438_ (.A(net32),
    .B(net36),
    .Y(_0531_));
 sg13g2_buf_1 _2439_ (.A(\rsa_unit_i.P_i[9] ),
    .X(_0532_));
 sg13g2_o21ai_1 _2440_ (.B1(_0532_),
    .Y(_0533_),
    .A1(net21),
    .A2(_0531_));
 sg13g2_inv_1 _2441_ (.Y(_0291_),
    .A(_0533_));
 sg13g2_mux2_1 _2442_ (.A0(_0402_),
    .A1(\rsa_c[0] ),
    .S(_1372_),
    .X(_0292_));
 sg13g2_mux2_1 _2443_ (.A0(\rsa_unit_i.R_i[1] ),
    .A1(\rsa_c[1] ),
    .S(net40),
    .X(_0293_));
 sg13g2_mux2_1 _2444_ (.A0(\rsa_unit_i.R_i[2] ),
    .A1(\rsa_c[2] ),
    .S(net40),
    .X(_0294_));
 sg13g2_mux2_1 _2445_ (.A0(\rsa_unit_i.R_i[3] ),
    .A1(\rsa_c[3] ),
    .S(net40),
    .X(_0295_));
 sg13g2_mux2_1 _2446_ (.A0(\rsa_unit_i.R_i[4] ),
    .A1(\rsa_c[4] ),
    .S(net40),
    .X(_0296_));
 sg13g2_mux2_1 _2447_ (.A0(\rsa_unit_i.R_i[5] ),
    .A1(\rsa_c[5] ),
    .S(net40),
    .X(_0297_));
 sg13g2_mux2_1 _2448_ (.A0(\rsa_unit_i.R_i[6] ),
    .A1(\rsa_c[6] ),
    .S(net40),
    .X(_0298_));
 sg13g2_mux2_1 _2449_ (.A0(\rsa_unit_i.R_i[7] ),
    .A1(\rsa_c[7] ),
    .S(net40),
    .X(_0299_));
 sg13g2_nor2_1 _2450_ (.A(_1374_),
    .B(net109),
    .Y(_0534_));
 sg13g2_or2_1 _2451_ (.X(_0535_),
    .B(_0534_),
    .A(_1344_));
 sg13g2_buf_1 _2452_ (.A(_0535_),
    .X(_0536_));
 sg13g2_nor3_1 _2453_ (.A(net109),
    .B(_1379_),
    .C(_0536_),
    .Y(_0537_));
 sg13g2_a21o_1 _2454_ (.A2(_0536_),
    .A1(_1379_),
    .B1(_0537_),
    .X(_0300_));
 sg13g2_inv_1 _2455_ (.Y(_0538_),
    .A(_0055_));
 sg13g2_nor2_1 _2456_ (.A(_1375_),
    .B(_0534_),
    .Y(_0539_));
 sg13g2_o21ai_1 _2457_ (.B1(_0539_),
    .Y(_0540_),
    .A1(_1379_),
    .A2(_0538_));
 sg13g2_nor3_1 _2458_ (.A(_0538_),
    .B(_1380_),
    .C(_0536_),
    .Y(_0541_));
 sg13g2_a21o_1 _2459_ (.A2(_0540_),
    .A1(_1378_),
    .B1(_0541_),
    .X(_0301_));
 sg13g2_nand4_1 _2460_ (.B(_1378_),
    .C(_0055_),
    .A(_1379_),
    .Y(_0542_),
    .D(_0539_));
 sg13g2_a21oi_1 _2461_ (.A1(_1379_),
    .A2(_1378_),
    .Y(_0543_),
    .B1(_0538_));
 sg13g2_o21ai_1 _2462_ (.B1(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ),
    .Y(_0544_),
    .A1(_0536_),
    .A2(_0543_));
 sg13g2_o21ai_1 _2463_ (.B1(_0544_),
    .Y(_0302_),
    .A1(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ),
    .A2(_0542_));
 sg13g2_nand3_1 _2464_ (.B(_1378_),
    .C(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ),
    .A(_1379_),
    .Y(_0545_));
 sg13g2_nor3_1 _2465_ (.A(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ),
    .B(_0536_),
    .C(_0545_),
    .Y(_0546_));
 sg13g2_a21o_1 _2466_ (.A2(_0545_),
    .A1(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ),
    .B1(_0546_),
    .X(_0547_));
 sg13g2_a22oi_1 _2467_ (.Y(_0548_),
    .B1(_0547_),
    .B2(_0055_),
    .A2(_0536_),
    .A1(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ));
 sg13g2_inv_1 _2468_ (.Y(_0303_),
    .A(_0548_));
 sg13g2_nand2_1 _2469_ (.Y(_0549_),
    .A(_0051_),
    .B(_0534_));
 sg13g2_nor4_1 _2470_ (.A(_1328_),
    .B(\rsa_unit_i.rsa_control_fsm.state[3] ),
    .C(_1391_),
    .D(_0549_),
    .Y(_0550_));
 sg13g2_or2_1 _2471_ (.X(_0551_),
    .B(_0550_),
    .A(_1344_));
 sg13g2_buf_1 _2472_ (.A(_0551_),
    .X(_0552_));
 sg13g2_or2_1 _2473_ (.X(_0553_),
    .B(_0552_),
    .A(_0549_));
 sg13g2_buf_1 _2474_ (.A(_0553_),
    .X(_0554_));
 sg13g2_nand2_1 _2475_ (.Y(_0555_),
    .A(_1334_),
    .B(_0552_));
 sg13g2_o21ai_1 _2476_ (.B1(_0555_),
    .Y(_0304_),
    .A1(_1334_),
    .A2(_0554_));
 sg13g2_nor2_1 _2477_ (.A(_1334_),
    .B(_0549_),
    .Y(_0556_));
 sg13g2_o21ai_1 _2478_ (.B1(_1333_),
    .Y(_0557_),
    .A1(_0552_),
    .A2(_0556_));
 sg13g2_o21ai_1 _2479_ (.B1(_0557_),
    .Y(_0305_),
    .A1(_1335_),
    .A2(_0554_));
 sg13g2_nand3b_1 _2480_ (.B(_1333_),
    .C(_1334_),
    .Y(_0558_),
    .A_N(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ));
 sg13g2_a21oi_1 _2481_ (.A1(_1334_),
    .A2(_1333_),
    .Y(_0559_),
    .B1(_0549_));
 sg13g2_o21ai_1 _2482_ (.B1(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ),
    .Y(_0560_),
    .A1(_0552_),
    .A2(_0559_));
 sg13g2_o21ai_1 _2483_ (.B1(_0560_),
    .Y(_0306_),
    .A1(_0554_),
    .A2(_0558_));
 sg13g2_nand3_1 _2484_ (.B(_1333_),
    .C(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ),
    .A(_1334_),
    .Y(_0561_));
 sg13g2_nor3_1 _2485_ (.A(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ),
    .B(_0552_),
    .C(_0561_),
    .Y(_0562_));
 sg13g2_a21oi_1 _2486_ (.A1(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ),
    .A2(_0561_),
    .Y(_0563_),
    .B1(_0562_));
 sg13g2_nand2_1 _2487_ (.Y(_0564_),
    .A(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ),
    .B(_0552_));
 sg13g2_o21ai_1 _2488_ (.B1(_0564_),
    .Y(_0307_),
    .A1(_0549_),
    .A2(_0563_));
 sg13g2_nor2_1 _2489_ (.A(net108),
    .B(_0375_),
    .Y(_0565_));
 sg13g2_a21oi_1 _2490_ (.A1(_0492_),
    .A2(_0565_),
    .Y(_0566_),
    .B1(net57));
 sg13g2_buf_1 _2491_ (.A(_0566_),
    .X(_0567_));
 sg13g2_buf_1 _2492_ (.A(_0567_),
    .X(_0568_));
 sg13g2_buf_1 _2493_ (.A(net93),
    .X(_0569_));
 sg13g2_nor2b_1 _2494_ (.A(net77),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[1] ),
    .Y(_0570_));
 sg13g2_a22oi_1 _2495_ (.Y(_0571_),
    .B1(net35),
    .B2(_0570_),
    .A2(\rsa_e[0] ),
    .A1(net77));
 sg13g2_nor2_1 _2496_ (.A(\rsa_unit_i.rsa_control_fsm.exp[0] ),
    .B(net26),
    .Y(_0572_));
 sg13g2_a21oi_1 _2497_ (.A1(net26),
    .A2(_0571_),
    .Y(_0308_),
    .B1(_0572_));
 sg13g2_nor2b_1 _2498_ (.A(net77),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[2] ),
    .Y(_0573_));
 sg13g2_a22oi_1 _2499_ (.Y(_0574_),
    .B1(net35),
    .B2(_0573_),
    .A2(\rsa_e[1] ),
    .A1(net77));
 sg13g2_nor2_1 _2500_ (.A(\rsa_unit_i.rsa_control_fsm.exp[1] ),
    .B(net26),
    .Y(_0575_));
 sg13g2_a21oi_1 _2501_ (.A1(net26),
    .A2(_0574_),
    .Y(_0309_),
    .B1(_0575_));
 sg13g2_nor2b_1 _2502_ (.A(net93),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[3] ),
    .Y(_0576_));
 sg13g2_a22oi_1 _2503_ (.Y(_0577_),
    .B1(net35),
    .B2(_0576_),
    .A2(\rsa_e[2] ),
    .A1(net77));
 sg13g2_nor2_1 _2504_ (.A(\rsa_unit_i.rsa_control_fsm.exp[2] ),
    .B(_0567_),
    .Y(_0578_));
 sg13g2_a21oi_1 _2505_ (.A1(net26),
    .A2(_0577_),
    .Y(_0310_),
    .B1(_0578_));
 sg13g2_nor2b_1 _2506_ (.A(net93),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[4] ),
    .Y(_0579_));
 sg13g2_a22oi_1 _2507_ (.Y(_0580_),
    .B1(net35),
    .B2(_0579_),
    .A2(\rsa_e[3] ),
    .A1(net77));
 sg13g2_nor2_1 _2508_ (.A(\rsa_unit_i.rsa_control_fsm.exp[3] ),
    .B(_0567_),
    .Y(_0581_));
 sg13g2_a21oi_1 _2509_ (.A1(net26),
    .A2(_0580_),
    .Y(_0311_),
    .B1(_0581_));
 sg13g2_nor2b_1 _2510_ (.A(net93),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[5] ),
    .Y(_0582_));
 sg13g2_a22oi_1 _2511_ (.Y(_0583_),
    .B1(net35),
    .B2(_0582_),
    .A2(\rsa_e[4] ),
    .A1(net77));
 sg13g2_nor2_1 _2512_ (.A(\rsa_unit_i.rsa_control_fsm.exp[4] ),
    .B(_0567_),
    .Y(_0584_));
 sg13g2_a21oi_1 _2513_ (.A1(net26),
    .A2(_0583_),
    .Y(_0312_),
    .B1(_0584_));
 sg13g2_nor2b_1 _2514_ (.A(net93),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[6] ),
    .Y(_0585_));
 sg13g2_a22oi_1 _2515_ (.Y(_0586_),
    .B1(net35),
    .B2(_0585_),
    .A2(\rsa_e[5] ),
    .A1(_0569_));
 sg13g2_nor2_1 _2516_ (.A(\rsa_unit_i.rsa_control_fsm.exp[5] ),
    .B(_0567_),
    .Y(_0587_));
 sg13g2_a21oi_1 _2517_ (.A1(_0568_),
    .A2(_0586_),
    .Y(_0313_),
    .B1(_0587_));
 sg13g2_inv_1 _2518_ (.Y(_0588_),
    .A(\rsa_unit_i.rsa_control_fsm.exp[7] ));
 sg13g2_nor2_1 _2519_ (.A(net93),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_a22oi_1 _2520_ (.Y(_0590_),
    .B1(net35),
    .B2(_0589_),
    .A2(\rsa_e[6] ),
    .A1(_0569_));
 sg13g2_nor2_1 _2521_ (.A(\rsa_unit_i.rsa_control_fsm.exp[6] ),
    .B(_0567_),
    .Y(_0591_));
 sg13g2_a21oi_1 _2522_ (.A1(_0568_),
    .A2(_0590_),
    .Y(_0314_),
    .B1(_0591_));
 sg13g2_nand3_1 _2523_ (.B(\rsa_e[7] ),
    .C(net58),
    .A(net77),
    .Y(_0592_));
 sg13g2_o21ai_1 _2524_ (.B1(_0592_),
    .Y(_0315_),
    .A1(_0588_),
    .A2(net26));
 sg13g2_mux2_1 _2525_ (.A0(\synchronizer_spi_clk_inst.data_sync[1] ),
    .A1(net3),
    .S(net85),
    .X(_0316_));
 sg13g2_nand2_1 _2526_ (.Y(_0593_),
    .A(_1315_),
    .B(\synchronizer_spi_clk_inst.data_sync[1] ));
 sg13g2_o21ai_1 _2527_ (.B1(_0593_),
    .Y(_0317_),
    .A1(_1485_),
    .A2(net86));
 sg13g2_mux2_1 _2528_ (.A0(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .A1(net2),
    .S(net85),
    .X(_0318_));
 sg13g2_mux2_1 _2529_ (.A0(_1318_),
    .A1(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .S(_1417_),
    .X(_0319_));
 sg13g2_mux2_1 _2530_ (.A0(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .A1(net4),
    .S(net85),
    .X(_0320_));
 sg13g2_mux2_1 _2531_ (.A0(\rsa_spi_wrapper_i.spi_mosi ),
    .A1(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .S(_1417_),
    .X(_0321_));
 sg13g2_nand2_1 _2532_ (.Y(_0594_),
    .A(_1340_),
    .B(_1332_));
 sg13g2_o21ai_1 _2533_ (.B1(_0594_),
    .Y(_0595_),
    .A1(_0117_),
    .A2(_1342_));
 sg13g2_inv_1 _2534_ (.Y(_0120_),
    .A(_0595_));
 sg13g2_buf_1 _2535_ (.A(_0387_),
    .X(_0596_));
 sg13g2_buf_1 _2536_ (.A(net25),
    .X(_0597_));
 sg13g2_inv_1 _2537_ (.Y(_0598_),
    .A(_0052_));
 sg13g2_nor3_1 _2538_ (.A(_0598_),
    .B(_1396_),
    .C(\rsa_unit_i.rsa_control_fsm.state[6] ),
    .Y(_0599_));
 sg13g2_buf_1 _2539_ (.A(_0599_),
    .X(_0600_));
 sg13g2_buf_1 _2540_ (.A(_0600_),
    .X(_0601_));
 sg13g2_mux2_1 _2541_ (.A0(_0420_),
    .A1(_0023_),
    .S(net51),
    .X(_0602_));
 sg13g2_buf_1 _2542_ (.A(\rsa_unit_i.mmm_multiply.A_bit ),
    .X(_0603_));
 sg13g2_buf_1 _2543_ (.A(net91),
    .X(_0604_));
 sg13g2_nand2_1 _2544_ (.Y(_0605_),
    .A(_0604_),
    .B(net48));
 sg13g2_o21ai_1 _2545_ (.B1(_0605_),
    .Y(_0234_),
    .A1(_0597_),
    .A2(_0602_));
 sg13g2_mux2_1 _2546_ (.A0(_0429_),
    .A1(_0024_),
    .S(net51),
    .X(_0606_));
 sg13g2_nand2_1 _2547_ (.Y(_0607_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[1] ),
    .B(net48));
 sg13g2_o21ai_1 _2548_ (.B1(_0607_),
    .Y(_0235_),
    .A1(net20),
    .A2(_0606_));
 sg13g2_mux2_1 _2549_ (.A0(_0434_),
    .A1(_0026_),
    .S(net51),
    .X(_0608_));
 sg13g2_nand2_1 _2550_ (.Y(_0609_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[2] ),
    .B(net48));
 sg13g2_o21ai_1 _2551_ (.B1(_0609_),
    .Y(_0236_),
    .A1(net20),
    .A2(_0608_));
 sg13g2_mux2_1 _2552_ (.A0(_0440_),
    .A1(_0028_),
    .S(net51),
    .X(_0610_));
 sg13g2_nand2_1 _2553_ (.Y(_0611_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[3] ),
    .B(net48));
 sg13g2_o21ai_1 _2554_ (.B1(_0611_),
    .Y(_0237_),
    .A1(net20),
    .A2(_0610_));
 sg13g2_mux2_1 _2555_ (.A0(_0446_),
    .A1(_0030_),
    .S(net51),
    .X(_0612_));
 sg13g2_nand2_1 _2556_ (.Y(_0613_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[4] ),
    .B(net48));
 sg13g2_o21ai_1 _2557_ (.B1(_0613_),
    .Y(_0238_),
    .A1(net20),
    .A2(_0612_));
 sg13g2_mux2_1 _2558_ (.A0(_0451_),
    .A1(_0032_),
    .S(net51),
    .X(_0614_));
 sg13g2_nand2_1 _2559_ (.Y(_0615_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[5] ),
    .B(net48));
 sg13g2_o21ai_1 _2560_ (.B1(_0615_),
    .Y(_0239_),
    .A1(net20),
    .A2(_0614_));
 sg13g2_mux2_1 _2561_ (.A0(_0456_),
    .A1(_0034_),
    .S(net51),
    .X(_0616_));
 sg13g2_nand2_1 _2562_ (.Y(_0617_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[6] ),
    .B(_1401_));
 sg13g2_o21ai_1 _2563_ (.B1(_0617_),
    .Y(_0240_),
    .A1(net20),
    .A2(_0616_));
 sg13g2_buf_1 _2564_ (.A(_0600_),
    .X(_0618_));
 sg13g2_mux2_1 _2565_ (.A0(_0462_),
    .A1(_0036_),
    .S(net50),
    .X(_0619_));
 sg13g2_nand2_1 _2566_ (.Y(_0620_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[7] ),
    .B(net48));
 sg13g2_o21ai_1 _2567_ (.B1(_0620_),
    .Y(_0241_),
    .A1(net20),
    .A2(_0619_));
 sg13g2_mux2_1 _2568_ (.A0(_0466_),
    .A1(_0038_),
    .S(net50),
    .X(_0621_));
 sg13g2_buf_1 _2569_ (.A(net57),
    .X(_0622_));
 sg13g2_nand2_1 _2570_ (.Y(_0623_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[8] ),
    .B(net42));
 sg13g2_o21ai_1 _2571_ (.B1(_0623_),
    .Y(_0242_),
    .A1(net20),
    .A2(_0621_));
 sg13g2_inv_1 _2572_ (.Y(_0624_),
    .A(net29));
 sg13g2_nor4_1 _2573_ (.A(_0040_),
    .B(_0596_),
    .C(_0624_),
    .D(net51),
    .Y(_0625_));
 sg13g2_a21o_1 _2574_ (.A2(net48),
    .A1(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[9] ),
    .B1(_0625_),
    .X(_0243_));
 sg13g2_nand3_1 _2575_ (.B(_0386_),
    .C(_0600_),
    .A(_1342_),
    .Y(_0626_));
 sg13g2_buf_2 _2576_ (.A(_0626_),
    .X(_0627_));
 sg13g2_buf_1 _2577_ (.A(_0627_),
    .X(_0628_));
 sg13g2_buf_1 _2578_ (.A(_0061_),
    .X(_0629_));
 sg13g2_inv_1 _2579_ (.Y(_0630_),
    .A(net91));
 sg13g2_buf_1 _2580_ (.A(\rsa_unit_i.mmm_multiply.adder2.fa_bit0.HA1.a ),
    .X(_0631_));
 sg13g2_nand2_1 _2581_ (.Y(_0632_),
    .A(net75),
    .B(_0631_));
 sg13g2_buf_2 _2582_ (.A(_0632_),
    .X(_0633_));
 sg13g2_a21oi_1 _2583_ (.A1(_1398_),
    .A2(_0394_),
    .Y(_0634_),
    .B1(\rsa_unit_i.P_i[0] ));
 sg13g2_nand3_1 _2584_ (.B(_0408_),
    .C(_0410_),
    .A(_0391_),
    .Y(_0635_));
 sg13g2_and2_1 _2585_ (.A(_1398_),
    .B(_0402_),
    .X(_0636_));
 sg13g2_nand3_1 _2586_ (.B(net63),
    .C(_0636_),
    .A(_0391_),
    .Y(_0637_));
 sg13g2_o21ai_1 _2587_ (.B1(_0637_),
    .Y(_0638_),
    .A1(_0634_),
    .A2(_0635_));
 sg13g2_buf_1 _2588_ (.A(_0638_),
    .X(_0639_));
 sg13g2_nand3_1 _2589_ (.B(net98),
    .C(_0639_),
    .A(_1513_),
    .Y(_0640_));
 sg13g2_a21o_1 _2590_ (.A2(_0394_),
    .A1(net78),
    .B1(\rsa_unit_i.P_i[0] ),
    .X(_0641_));
 sg13g2_a221oi_1 _2591_ (.B2(_0641_),
    .C1(_0391_),
    .B1(net52),
    .A1(_0402_),
    .Y(_0642_),
    .A2(net37));
 sg13g2_buf_1 _2592_ (.A(_0642_),
    .X(_0643_));
 sg13g2_nor2_1 _2593_ (.A(_1513_),
    .B(net98),
    .Y(_0644_));
 sg13g2_a22oi_1 _2594_ (.Y(_0645_),
    .B1(_0639_),
    .B2(_0644_),
    .A2(_0643_),
    .A1(net98));
 sg13g2_inv_1 _2595_ (.Y(_0646_),
    .A(net92));
 sg13g2_a21oi_1 _2596_ (.A1(net78),
    .A2(_0395_),
    .Y(_0647_),
    .B1(_0646_));
 sg13g2_nor3_1 _2597_ (.A(net69),
    .B(_0025_),
    .C(net53),
    .Y(_0648_));
 sg13g2_mux2_1 _2598_ (.A0(_0647_),
    .A1(_0648_),
    .S(_0412_),
    .X(_0649_));
 sg13g2_buf_1 _2599_ (.A(_0649_),
    .X(_0650_));
 sg13g2_a21oi_1 _2600_ (.A1(_0640_),
    .A2(_0645_),
    .Y(_0651_),
    .B1(_0650_));
 sg13g2_and3_1 _2601_ (.X(_0652_),
    .A(_0640_),
    .B(_0645_),
    .C(_0650_));
 sg13g2_o21ai_1 _2602_ (.B1(_0603_),
    .Y(_0653_),
    .A1(_0651_),
    .A2(_0652_));
 sg13g2_o21ai_1 _2603_ (.B1(_0653_),
    .Y(_0654_),
    .A1(net90),
    .A2(_0633_));
 sg13g2_and2_1 _2604_ (.A(net63),
    .B(_0636_),
    .X(_0655_));
 sg13g2_nor2_1 _2605_ (.A(_0412_),
    .B(_0634_),
    .Y(_0656_));
 sg13g2_nor4_1 _2606_ (.A(_1459_),
    .B(_0630_),
    .C(_0655_),
    .D(_0656_),
    .Y(_0657_));
 sg13g2_a21oi_1 _2607_ (.A1(_1514_),
    .A2(_0631_),
    .Y(_0658_),
    .B1(net91));
 sg13g2_nor3_1 _2608_ (.A(_0391_),
    .B(_0657_),
    .C(_0658_),
    .Y(_0659_));
 sg13g2_nor2b_1 _2609_ (.A(_0659_),
    .B_N(_0041_),
    .Y(_0660_));
 sg13g2_nor4_1 _2610_ (.A(_0391_),
    .B(_0041_),
    .C(_0657_),
    .D(_0658_),
    .Y(_0661_));
 sg13g2_nor2_1 _2611_ (.A(_0660_),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_xnor2_1 _2612_ (.Y(_0663_),
    .A(_0654_),
    .B(_0662_));
 sg13g2_nand2_1 _2613_ (.Y(_0664_),
    .A(_0631_),
    .B(net42));
 sg13g2_o21ai_1 _2614_ (.B1(_0664_),
    .Y(_0244_),
    .A1(net19),
    .A2(_0663_));
 sg13g2_buf_1 _2615_ (.A(_0064_),
    .X(_0665_));
 sg13g2_nor4_1 _2616_ (.A(_1400_),
    .B(_1467_),
    .C(_0025_),
    .D(net53),
    .Y(_0666_));
 sg13g2_nand2_1 _2617_ (.Y(_0667_),
    .A(net92),
    .B(net98));
 sg13g2_a21oi_1 _2618_ (.A1(net78),
    .A2(net63),
    .Y(_0668_),
    .B1(_0667_));
 sg13g2_mux2_1 _2619_ (.A0(_0666_),
    .A1(_0668_),
    .S(net52),
    .X(_0669_));
 sg13g2_buf_2 _2620_ (.A(_0669_),
    .X(_0670_));
 sg13g2_inv_1 _2621_ (.Y(_0671_),
    .A(_0670_));
 sg13g2_nand2_1 _2622_ (.Y(_0672_),
    .A(_1513_),
    .B(_1467_));
 sg13g2_nor2_1 _2623_ (.A(_1513_),
    .B(_1467_),
    .Y(_0673_));
 sg13g2_a21oi_1 _2624_ (.A1(_0650_),
    .A2(_0672_),
    .Y(_0674_),
    .B1(_0673_));
 sg13g2_a221oi_1 _2625_ (.B2(_0639_),
    .C1(net89),
    .B1(_0674_),
    .A1(_0643_),
    .Y(_0675_),
    .A2(_0671_));
 sg13g2_nor3_1 _2626_ (.A(net69),
    .B(_0027_),
    .C(net53),
    .Y(_0676_));
 sg13g2_inv_1 _2627_ (.Y(_0677_),
    .A(\rsa_unit_i.P_i[2] ));
 sg13g2_a21oi_1 _2628_ (.A1(_0393_),
    .A2(_0394_),
    .Y(_0678_),
    .B1(_0677_));
 sg13g2_mux2_1 _2629_ (.A0(_0676_),
    .A1(_0678_),
    .S(net52),
    .X(_0679_));
 sg13g2_buf_2 _2630_ (.A(_0679_),
    .X(_0680_));
 sg13g2_nor4_1 _2631_ (.A(net89),
    .B(_0630_),
    .C(_0675_),
    .D(_0680_),
    .Y(_0681_));
 sg13g2_a21o_1 _2632_ (.A2(_0672_),
    .A1(_0650_),
    .B1(_0673_),
    .X(_0682_));
 sg13g2_a22oi_1 _2633_ (.Y(_0683_),
    .B1(_0682_),
    .B2(_0639_),
    .A2(_0670_),
    .A1(_0643_));
 sg13g2_and4_1 _2634_ (.A(net89),
    .B(_0603_),
    .C(_0680_),
    .D(_0683_),
    .X(_0684_));
 sg13g2_nor4_1 _2635_ (.A(net75),
    .B(_0675_),
    .C(_0680_),
    .D(_0683_),
    .Y(_0685_));
 sg13g2_and2_1 _2636_ (.A(net91),
    .B(_0680_),
    .X(_0686_));
 sg13g2_nor2_1 _2637_ (.A(net89),
    .B(_0633_),
    .Y(_0687_));
 sg13g2_a21o_1 _2638_ (.A2(_0686_),
    .A1(_0675_),
    .B1(_0687_),
    .X(_0688_));
 sg13g2_nor4_2 _2639_ (.A(_0681_),
    .B(_0684_),
    .C(_0685_),
    .Y(_0689_),
    .D(_0688_));
 sg13g2_nor2_1 _2640_ (.A(net90),
    .B(_0633_),
    .Y(_0690_));
 sg13g2_nor2_1 _2641_ (.A(_0690_),
    .B(_0661_),
    .Y(_0691_));
 sg13g2_a21o_1 _2642_ (.A2(_0691_),
    .A1(_0653_),
    .B1(_0660_),
    .X(_0692_));
 sg13g2_buf_1 _2643_ (.A(_0692_),
    .X(_0693_));
 sg13g2_xnor2_1 _2644_ (.Y(_0694_),
    .A(_0689_),
    .B(_0693_));
 sg13g2_xnor2_1 _2645_ (.Y(_0695_),
    .A(_0043_),
    .B(_0694_));
 sg13g2_nand2_1 _2646_ (.Y(_0696_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[1].fa.HA1.a ),
    .B(net42));
 sg13g2_o21ai_1 _2647_ (.B1(_0696_),
    .Y(_0245_),
    .A1(net19),
    .A2(_0695_));
 sg13g2_inv_1 _2648_ (.Y(_0697_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[2].fa.HA1.a ));
 sg13g2_inv_1 _2649_ (.Y(_0698_),
    .A(_0627_));
 sg13g2_nor2_1 _2650_ (.A(_0689_),
    .B(_0693_),
    .Y(_0699_));
 sg13g2_a21oi_2 _2651_ (.B1(_0043_),
    .Y(_0700_),
    .A2(_0693_),
    .A1(_0689_));
 sg13g2_buf_1 _2652_ (.A(net97),
    .X(_0701_));
 sg13g2_nor2_1 _2653_ (.A(net74),
    .B(_0633_),
    .Y(_0702_));
 sg13g2_nand3b_1 _2654_ (.B(net63),
    .C(net78),
    .Y(_0703_),
    .A_N(_0029_));
 sg13g2_o21ai_1 _2655_ (.B1(\rsa_unit_i.P_i[3] ),
    .Y(_0704_),
    .A1(net69),
    .A2(_0405_));
 sg13g2_mux2_1 _2656_ (.A0(_0703_),
    .A1(_0704_),
    .S(net52),
    .X(_0705_));
 sg13g2_buf_2 _2657_ (.A(_0705_),
    .X(_0706_));
 sg13g2_nor3_1 _2658_ (.A(net74),
    .B(net75),
    .C(_0706_),
    .Y(_0707_));
 sg13g2_nor3_1 _2659_ (.A(_1586_),
    .B(net75),
    .C(_0706_),
    .Y(_0708_));
 sg13g2_nor2b_1 _2660_ (.A(_1513_),
    .B_N(_0402_),
    .Y(_0709_));
 sg13g2_nand2b_1 _2661_ (.Y(_0710_),
    .B(_0025_),
    .A_N(net98));
 sg13g2_nand4_1 _2662_ (.B(_0394_),
    .C(_0709_),
    .A(_1398_),
    .Y(_0711_),
    .D(_0710_));
 sg13g2_nand2b_1 _2663_ (.Y(_0712_),
    .B(net98),
    .A_N(_1513_));
 sg13g2_and3_1 _2664_ (.X(_0713_),
    .A(_0408_),
    .B(_0410_),
    .C(_0712_));
 sg13g2_nor2b_1 _2665_ (.A(_1513_),
    .B_N(net92),
    .Y(_0714_));
 sg13g2_o21ai_1 _2666_ (.B1(_0714_),
    .Y(_0715_),
    .A1(net69),
    .A2(net53));
 sg13g2_a221oi_1 _2667_ (.B2(_0715_),
    .C1(_0634_),
    .B1(_0713_),
    .A1(_0412_),
    .Y(_0716_),
    .A2(_0711_));
 sg13g2_buf_1 _2668_ (.A(_0716_),
    .X(_0717_));
 sg13g2_o21ai_1 _2669_ (.B1(_0680_),
    .Y(_0718_),
    .A1(_0670_),
    .A2(_0717_));
 sg13g2_nor3_1 _2670_ (.A(_0670_),
    .B(_0680_),
    .C(_0717_),
    .Y(_0719_));
 sg13g2_a21o_1 _2671_ (.A2(_0718_),
    .A1(net89),
    .B1(_0719_),
    .X(_0720_));
 sg13g2_buf_1 _2672_ (.A(_0720_),
    .X(_0721_));
 sg13g2_mux2_1 _2673_ (.A0(_0707_),
    .A1(_0708_),
    .S(_0721_),
    .X(_0722_));
 sg13g2_and3_1 _2674_ (.X(_0723_),
    .A(net91),
    .B(_0408_),
    .C(_0410_));
 sg13g2_a221oi_1 _2675_ (.B2(_0723_),
    .C1(_0392_),
    .B1(_0641_),
    .A1(net91),
    .Y(_0724_),
    .A2(_0655_));
 sg13g2_nor2b_1 _2676_ (.A(_0391_),
    .B_N(\rsa_unit_i.mmm_multiply.A_bit ),
    .Y(_0725_));
 sg13g2_and3_1 _2677_ (.X(_0726_),
    .A(_0408_),
    .B(_0410_),
    .C(_0725_));
 sg13g2_a22oi_1 _2678_ (.Y(_0727_),
    .B1(_0726_),
    .B2(_0641_),
    .A2(_0725_),
    .A1(_0655_));
 sg13g2_nor2b_1 _2679_ (.A(_0724_),
    .B_N(_0727_),
    .Y(_0728_));
 sg13g2_buf_1 _2680_ (.A(_0728_),
    .X(_0729_));
 sg13g2_and4_1 _2681_ (.A(net74),
    .B(net91),
    .C(_0706_),
    .D(net30),
    .X(_0730_));
 sg13g2_and4_1 _2682_ (.A(_1586_),
    .B(net91),
    .C(_0706_),
    .D(net30),
    .X(_0731_));
 sg13g2_mux2_1 _2683_ (.A0(_0730_),
    .A1(_0731_),
    .S(_0721_),
    .X(_0732_));
 sg13g2_nor3_1 _2684_ (.A(net75),
    .B(_0706_),
    .C(_0729_),
    .Y(_0733_));
 sg13g2_nor4_2 _2685_ (.A(_0702_),
    .B(_0722_),
    .C(_0732_),
    .Y(_0734_),
    .D(_0733_));
 sg13g2_xor2_1 _2686_ (.B(_0734_),
    .A(_0437_),
    .X(_0735_));
 sg13g2_or3_1 _2687_ (.A(_0699_),
    .B(_0700_),
    .C(_0735_),
    .X(_0736_));
 sg13g2_o21ai_1 _2688_ (.B1(_0735_),
    .Y(_0737_),
    .A1(_0699_),
    .A2(_0700_));
 sg13g2_nand3_1 _2689_ (.B(_0736_),
    .C(_0737_),
    .A(_0698_),
    .Y(_0738_));
 sg13g2_o21ai_1 _2690_ (.B1(_0738_),
    .Y(_0246_),
    .A1(_0697_),
    .A2(net58));
 sg13g2_nand2_1 _2691_ (.Y(_0739_),
    .A(_0437_),
    .B(_0734_));
 sg13g2_o21ai_1 _2692_ (.B1(_0739_),
    .Y(_0740_),
    .A1(_0699_),
    .A2(_0700_));
 sg13g2_o21ai_1 _2693_ (.B1(_0740_),
    .Y(_0741_),
    .A1(_0437_),
    .A2(_0734_));
 sg13g2_buf_1 _2694_ (.A(_0741_),
    .X(_0742_));
 sg13g2_buf_1 _2695_ (.A(_1608_),
    .X(_0743_));
 sg13g2_nor2_1 _2696_ (.A(_0643_),
    .B(_0639_),
    .Y(_0744_));
 sg13g2_buf_1 _2697_ (.A(_0744_),
    .X(_0745_));
 sg13g2_nor2_1 _2698_ (.A(net73),
    .B(_0745_),
    .Y(_0746_));
 sg13g2_nor2_1 _2699_ (.A(_1609_),
    .B(_0745_),
    .Y(_0747_));
 sg13g2_and2_1 _2700_ (.A(net97),
    .B(_0706_),
    .X(_0748_));
 sg13g2_nand2b_1 _2701_ (.Y(_0749_),
    .B(\rsa_unit_i.P_i[3] ),
    .A_N(_0067_));
 sg13g2_a21oi_1 _2702_ (.A1(_0393_),
    .A2(_0395_),
    .Y(_0750_),
    .B1(_0749_));
 sg13g2_nor4_1 _2703_ (.A(net69),
    .B(net97),
    .C(_0029_),
    .D(_0405_),
    .Y(_0751_));
 sg13g2_mux2_1 _2704_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0412_),
    .X(_0752_));
 sg13g2_buf_1 _2705_ (.A(_0752_),
    .X(_0753_));
 sg13g2_nor4_1 _2706_ (.A(_0670_),
    .B(_0680_),
    .C(_0717_),
    .D(_0753_),
    .Y(_0754_));
 sg13g2_nor4_1 _2707_ (.A(_1564_),
    .B(_0670_),
    .C(_0717_),
    .D(_0753_),
    .Y(_0755_));
 sg13g2_nor3_1 _2708_ (.A(_1564_),
    .B(_0680_),
    .C(_0753_),
    .Y(_0756_));
 sg13g2_nor4_2 _2709_ (.A(_0748_),
    .B(_0754_),
    .C(_0755_),
    .Y(_0757_),
    .D(_0756_));
 sg13g2_mux2_1 _2710_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0757_),
    .X(_0758_));
 sg13g2_nand3b_1 _2711_ (.B(net63),
    .C(net78),
    .Y(_0759_),
    .A_N(_0031_));
 sg13g2_o21ai_1 _2712_ (.B1(\rsa_unit_i.P_i[4] ),
    .Y(_0760_),
    .A1(net69),
    .A2(net53));
 sg13g2_mux2_1 _2713_ (.A0(_0759_),
    .A1(_0760_),
    .S(net52),
    .X(_0761_));
 sg13g2_xnor2_1 _2714_ (.Y(_0762_),
    .A(_0758_),
    .B(_0761_));
 sg13g2_nor2_1 _2715_ (.A(net73),
    .B(_0633_),
    .Y(_0763_));
 sg13g2_a21o_1 _2716_ (.A2(_0762_),
    .A1(_0604_),
    .B1(_0763_),
    .X(_0764_));
 sg13g2_buf_1 _2717_ (.A(_0764_),
    .X(_0765_));
 sg13g2_xnor2_1 _2718_ (.Y(_0766_),
    .A(_0443_),
    .B(_0765_));
 sg13g2_xnor2_1 _2719_ (.Y(_0767_),
    .A(_0742_),
    .B(_0766_));
 sg13g2_nand2_1 _2720_ (.Y(_0768_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[3].fa.HA1.a ),
    .B(net42));
 sg13g2_o21ai_1 _2721_ (.B1(_0768_),
    .Y(_0247_),
    .A1(net19),
    .A2(_0767_));
 sg13g2_nand3_1 _2722_ (.B(net75),
    .C(_0631_),
    .A(_1625_),
    .Y(_0769_));
 sg13g2_nand2b_1 _2723_ (.Y(_0770_),
    .B(_0727_),
    .A_N(_0724_));
 sg13g2_nand3b_1 _2724_ (.B(net63),
    .C(net78),
    .Y(_0771_),
    .A_N(_0033_));
 sg13g2_o21ai_1 _2725_ (.B1(\rsa_unit_i.P_i[5] ),
    .Y(_0772_),
    .A1(net69),
    .A2(net53));
 sg13g2_mux2_1 _2726_ (.A0(_0771_),
    .A1(_0772_),
    .S(net52),
    .X(_0773_));
 sg13g2_buf_2 _2727_ (.A(_0773_),
    .X(_0774_));
 sg13g2_a21oi_1 _2728_ (.A1(_0770_),
    .A2(_0774_),
    .Y(_0775_),
    .B1(net75));
 sg13g2_nor2_1 _2729_ (.A(net44),
    .B(_0771_),
    .Y(_0776_));
 sg13g2_a21o_1 _2730_ (.A2(net29),
    .A1(\rsa_unit_i.P_i[5] ),
    .B1(_0776_),
    .X(_0777_));
 sg13g2_nor2_1 _2731_ (.A(_1608_),
    .B(_0761_),
    .Y(_0778_));
 sg13g2_nand4_1 _2732_ (.B(net30),
    .C(_0777_),
    .A(net96),
    .Y(_0779_),
    .D(_0778_));
 sg13g2_nor3_1 _2733_ (.A(net69),
    .B(_0031_),
    .C(net53),
    .Y(_0780_));
 sg13g2_inv_1 _2734_ (.Y(_0781_),
    .A(\rsa_unit_i.P_i[4] ));
 sg13g2_a21oi_1 _2735_ (.A1(net78),
    .A2(net63),
    .Y(_0782_),
    .B1(_0781_));
 sg13g2_mux2_1 _2736_ (.A0(_0780_),
    .A1(_0782_),
    .S(net52),
    .X(_0783_));
 sg13g2_nor2_1 _2737_ (.A(_1609_),
    .B(_0783_),
    .Y(_0784_));
 sg13g2_nand4_1 _2738_ (.B(net30),
    .C(_0777_),
    .A(_1625_),
    .Y(_0785_),
    .D(_0784_));
 sg13g2_and2_1 _2739_ (.A(net96),
    .B(_0774_),
    .X(_0786_));
 sg13g2_and2_1 _2740_ (.A(_1625_),
    .B(_0774_),
    .X(_0787_));
 sg13g2_a22oi_1 _2741_ (.Y(_0788_),
    .B1(_0787_),
    .B2(_0778_),
    .A2(_0784_),
    .A1(_0786_));
 sg13g2_nand4_1 _2742_ (.B(_0779_),
    .C(_0785_),
    .A(_0775_),
    .Y(_0789_),
    .D(_0788_));
 sg13g2_nor2_1 _2743_ (.A(net96),
    .B(_0774_),
    .Y(_0790_));
 sg13g2_nor2_1 _2744_ (.A(net96),
    .B(_0633_),
    .Y(_0791_));
 sg13g2_a21oi_1 _2745_ (.A1(net30),
    .A2(_0777_),
    .Y(_0792_),
    .B1(_1625_));
 sg13g2_nor4_1 _2746_ (.A(_0790_),
    .B(_0791_),
    .C(_0784_),
    .D(_0792_),
    .Y(_0793_));
 sg13g2_a21oi_1 _2747_ (.A1(net30),
    .A2(_0790_),
    .Y(_0794_),
    .B1(_0786_));
 sg13g2_nor4_1 _2748_ (.A(_0757_),
    .B(_0794_),
    .C(_0791_),
    .D(_0778_),
    .Y(_0795_));
 sg13g2_a221oi_1 _2749_ (.B2(_0757_),
    .C1(_0795_),
    .B1(_0793_),
    .A1(_0769_),
    .Y(_0796_),
    .A2(_0789_));
 sg13g2_nand2b_1 _2750_ (.Y(_0797_),
    .B(_0796_),
    .A_N(_0046_));
 sg13g2_nand2b_1 _2751_ (.Y(_0798_),
    .B(_0046_),
    .A_N(_0796_));
 sg13g2_nand2_1 _2752_ (.Y(_0799_),
    .A(_0797_),
    .B(_0798_));
 sg13g2_nor2_1 _2753_ (.A(_0437_),
    .B(_0734_),
    .Y(_0800_));
 sg13g2_nor3_1 _2754_ (.A(_0699_),
    .B(_0700_),
    .C(_0800_),
    .Y(_0801_));
 sg13g2_nand2b_1 _2755_ (.Y(_0802_),
    .B(_0739_),
    .A_N(_0443_));
 sg13g2_nand2b_1 _2756_ (.Y(_0803_),
    .B(_0765_),
    .A_N(_0443_));
 sg13g2_o21ai_1 _2757_ (.B1(_0803_),
    .Y(_0804_),
    .A1(_0801_),
    .A2(_0802_));
 sg13g2_a21oi_1 _2758_ (.A1(_0742_),
    .A2(_0765_),
    .Y(_0805_),
    .B1(_0804_));
 sg13g2_xnor2_1 _2759_ (.Y(_0806_),
    .A(_0799_),
    .B(_0805_));
 sg13g2_nand2_1 _2760_ (.Y(_0807_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[4].fa.HA1.a ),
    .B(net42));
 sg13g2_o21ai_1 _2761_ (.B1(_0807_),
    .Y(_0248_),
    .A1(net19),
    .A2(_0806_));
 sg13g2_nand2_1 _2762_ (.Y(_0808_),
    .A(_0803_),
    .B(_0797_));
 sg13g2_a21oi_1 _2763_ (.A1(net76),
    .A2(_0762_),
    .Y(_0809_),
    .B1(_0763_));
 sg13g2_nor2b_1 _2764_ (.A(_0796_),
    .B_N(_0046_),
    .Y(_0810_));
 sg13g2_a21oi_1 _2765_ (.A1(_0443_),
    .A2(_0809_),
    .Y(_0811_),
    .B1(_0810_));
 sg13g2_a22oi_1 _2766_ (.Y(_0812_),
    .B1(_0811_),
    .B2(_0742_),
    .A2(_0808_),
    .A1(_0798_));
 sg13g2_nor2_1 _2767_ (.A(_0774_),
    .B(_0784_),
    .Y(_0813_));
 sg13g2_nand2_1 _2768_ (.Y(_0814_),
    .A(_1609_),
    .B(_0783_));
 sg13g2_o21ai_1 _2769_ (.B1(net96),
    .Y(_0815_),
    .A1(_0774_),
    .A2(_0814_));
 sg13g2_a21oi_2 _2770_ (.B1(_0815_),
    .Y(_0816_),
    .A2(_0813_),
    .A1(_0757_));
 sg13g2_nor2b_1 _2771_ (.A(_0753_),
    .B_N(_0774_),
    .Y(_0817_));
 sg13g2_and2_1 _2772_ (.A(_0814_),
    .B(_0817_),
    .X(_0818_));
 sg13g2_nand2_1 _2773_ (.Y(_0819_),
    .A(_0416_),
    .B(_0704_));
 sg13g2_nand2_1 _2774_ (.Y(_0820_),
    .A(_0412_),
    .B(_0703_));
 sg13g2_a221oi_1 _2775_ (.B2(_1609_),
    .C1(_1586_),
    .B1(_0783_),
    .A1(_0819_),
    .Y(_0821_),
    .A2(_0820_));
 sg13g2_and3_1 _2776_ (.X(_0822_),
    .A(_1608_),
    .B(_0761_),
    .C(_0774_));
 sg13g2_a21o_1 _2777_ (.A2(_0821_),
    .A1(_0817_),
    .B1(_0822_),
    .X(_0823_));
 sg13g2_a21o_1 _2778_ (.A2(_0818_),
    .A1(_0721_),
    .B1(_0823_),
    .X(_0824_));
 sg13g2_buf_1 _2779_ (.A(_0824_),
    .X(_0825_));
 sg13g2_nand2_1 _2780_ (.Y(_0826_),
    .A(net37),
    .B(_0412_));
 sg13g2_nor2_1 _2781_ (.A(_0035_),
    .B(_0826_),
    .Y(_0827_));
 sg13g2_nand2_1 _2782_ (.Y(_0828_),
    .A(\rsa_unit_i.P_i[6] ),
    .B(net29));
 sg13g2_nand2b_1 _2783_ (.Y(_0829_),
    .B(_0828_),
    .A_N(_0827_));
 sg13g2_buf_2 _2784_ (.A(_0829_),
    .X(_0830_));
 sg13g2_nor3_1 _2785_ (.A(net95),
    .B(_0770_),
    .C(_0830_),
    .Y(_0831_));
 sg13g2_o21ai_1 _2786_ (.B1(_0831_),
    .Y(_0832_),
    .A1(_0816_),
    .A2(_0825_));
 sg13g2_nand2_1 _2787_ (.Y(_0833_),
    .A(_0770_),
    .B(_0830_));
 sg13g2_a21o_1 _2788_ (.A2(_0813_),
    .A1(_0757_),
    .B1(_0815_),
    .X(_0834_));
 sg13g2_buf_2 _2789_ (.A(_0834_),
    .X(_0835_));
 sg13g2_a21oi_1 _2790_ (.A1(_0721_),
    .A2(_0818_),
    .Y(_0836_),
    .B1(_0823_));
 sg13g2_buf_2 _2791_ (.A(_0836_),
    .X(_0837_));
 sg13g2_nor2b_1 _2792_ (.A(_0827_),
    .B_N(_0828_),
    .Y(_0838_));
 sg13g2_nor2_1 _2793_ (.A(net95),
    .B(_0838_),
    .Y(_0839_));
 sg13g2_nand3_1 _2794_ (.B(_0837_),
    .C(_0839_),
    .A(_0835_),
    .Y(_0840_));
 sg13g2_nand3_1 _2795_ (.B(_0833_),
    .C(_0840_),
    .A(_0832_),
    .Y(_0841_));
 sg13g2_nand3_1 _2796_ (.B(_0835_),
    .C(_0837_),
    .A(_0729_),
    .Y(_0842_));
 sg13g2_o21ai_1 _2797_ (.B1(_0830_),
    .Y(_0843_),
    .A1(_0816_),
    .A2(_0825_));
 sg13g2_o21ai_1 _2798_ (.B1(_0843_),
    .Y(_0844_),
    .A1(_0830_),
    .A2(_0842_));
 sg13g2_nor2_1 _2799_ (.A(_0334_),
    .B(net75),
    .Y(_0845_));
 sg13g2_buf_1 _2800_ (.A(net95),
    .X(_0846_));
 sg13g2_nor2_1 _2801_ (.A(net72),
    .B(_0633_),
    .Y(_0847_));
 sg13g2_a221oi_1 _2802_ (.B2(_0845_),
    .C1(_0847_),
    .B1(_0844_),
    .A1(net76),
    .Y(_0848_),
    .A2(_0841_));
 sg13g2_xnor2_1 _2803_ (.Y(_0849_),
    .A(_0047_),
    .B(_0848_));
 sg13g2_xnor2_1 _2804_ (.Y(_0850_),
    .A(_0812_),
    .B(_0849_));
 sg13g2_nand2_1 _2805_ (.Y(_0851_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[5].fa.HA1.a ),
    .B(net42));
 sg13g2_o21ai_1 _2806_ (.B1(_0851_),
    .Y(_0249_),
    .A1(net19),
    .A2(_0850_));
 sg13g2_a22oi_1 _2807_ (.Y(_0852_),
    .B1(_0844_),
    .B2(_0845_),
    .A2(_0841_),
    .A1(net76));
 sg13g2_nand2b_1 _2808_ (.Y(_0853_),
    .B(_0852_),
    .A_N(_0847_));
 sg13g2_a221oi_1 _2809_ (.B2(_0742_),
    .C1(_0853_),
    .B1(_0811_),
    .A1(_0798_),
    .Y(_0854_),
    .A2(_0808_));
 sg13g2_nand2_1 _2810_ (.Y(_0855_),
    .A(_0739_),
    .B(_0765_));
 sg13g2_and2_1 _2811_ (.A(_0047_),
    .B(_0797_),
    .X(_0856_));
 sg13g2_o21ai_1 _2812_ (.B1(_0856_),
    .Y(_0857_),
    .A1(_0801_),
    .A2(_0855_));
 sg13g2_o21ai_1 _2813_ (.B1(_0047_),
    .Y(_0858_),
    .A1(_0810_),
    .A2(_0848_));
 sg13g2_o21ai_1 _2814_ (.B1(_0858_),
    .Y(_0859_),
    .A1(_0804_),
    .A2(_0857_));
 sg13g2_nor2_1 _2815_ (.A(_0854_),
    .B(_0859_),
    .Y(_0860_));
 sg13g2_nor3_1 _2816_ (.A(_0037_),
    .B(_0396_),
    .C(net44),
    .Y(_0861_));
 sg13g2_a21oi_2 _2817_ (.B1(_0861_),
    .Y(_0862_),
    .A2(net29),
    .A1(\rsa_unit_i.P_i[7] ));
 sg13g2_xnor2_1 _2818_ (.Y(_0863_),
    .A(net94),
    .B(_0862_));
 sg13g2_nor4_1 _2819_ (.A(_0745_),
    .B(_0837_),
    .C(_0839_),
    .D(_0863_),
    .Y(_0864_));
 sg13g2_nor2_1 _2820_ (.A(_0745_),
    .B(_0863_),
    .Y(_0865_));
 sg13g2_nand3_1 _2821_ (.B(_0838_),
    .C(_0865_),
    .A(_0816_),
    .Y(_0866_));
 sg13g2_nor2_1 _2822_ (.A(net72),
    .B(_0745_),
    .Y(_0867_));
 sg13g2_nand3_1 _2823_ (.B(_0863_),
    .C(_0867_),
    .A(_0835_),
    .Y(_0868_));
 sg13g2_a21oi_1 _2824_ (.A1(_0866_),
    .A2(_0868_),
    .Y(_0869_),
    .B1(_0825_));
 sg13g2_nor2_1 _2825_ (.A(_0864_),
    .B(_0869_),
    .Y(_0870_));
 sg13g2_nor2_1 _2826_ (.A(_0745_),
    .B(_0838_),
    .Y(_0871_));
 sg13g2_nand3_1 _2827_ (.B(_0863_),
    .C(_0871_),
    .A(_0837_),
    .Y(_0872_));
 sg13g2_nand3_1 _2828_ (.B(_0816_),
    .C(_0865_),
    .A(net72),
    .Y(_0873_));
 sg13g2_o21ai_1 _2829_ (.B1(_0873_),
    .Y(_0874_),
    .A1(_0816_),
    .A2(_0872_));
 sg13g2_o21ai_1 _2830_ (.B1(net76),
    .Y(_0875_),
    .A1(net30),
    .A2(_0862_));
 sg13g2_nor2_1 _2831_ (.A(_0830_),
    .B(_0863_),
    .Y(_0876_));
 sg13g2_a22oi_1 _2832_ (.Y(_0877_),
    .B1(_0876_),
    .B2(net72),
    .A2(_0863_),
    .A1(_0839_));
 sg13g2_nor2_1 _2833_ (.A(_0745_),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_nor3_1 _2834_ (.A(_0874_),
    .B(_0875_),
    .C(_0878_),
    .Y(_0879_));
 sg13g2_a21oi_1 _2835_ (.A1(_0350_),
    .A2(_0631_),
    .Y(_0880_),
    .B1(net76));
 sg13g2_a21oi_1 _2836_ (.A1(_0870_),
    .A2(_0879_),
    .Y(_0881_),
    .B1(_0880_));
 sg13g2_xnor2_1 _2837_ (.Y(_0882_),
    .A(_0459_),
    .B(_0881_));
 sg13g2_xnor2_1 _2838_ (.Y(_0883_),
    .A(_0860_),
    .B(_0882_));
 sg13g2_nand2_1 _2839_ (.Y(_0884_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[6].fa.HA1.a ),
    .B(net42));
 sg13g2_o21ai_1 _2840_ (.B1(_0884_),
    .Y(_0250_),
    .A1(net19),
    .A2(_0883_));
 sg13g2_and2_1 _2841_ (.A(_0459_),
    .B(_0848_),
    .X(_0885_));
 sg13g2_nor2b_1 _2842_ (.A(_0881_),
    .B_N(_0459_),
    .Y(_0886_));
 sg13g2_a221oi_1 _2843_ (.B2(_0812_),
    .C1(_0886_),
    .B1(_0885_),
    .A1(_0459_),
    .Y(_0887_),
    .A2(_0859_));
 sg13g2_buf_2 _2844_ (.A(_0887_),
    .X(_0888_));
 sg13g2_inv_1 _2845_ (.Y(_0889_),
    .A(_0881_));
 sg13g2_o21ai_1 _2846_ (.B1(_0889_),
    .Y(_0890_),
    .A1(_0854_),
    .A2(_0859_));
 sg13g2_buf_1 _2847_ (.A(_0890_),
    .X(_0891_));
 sg13g2_nand2_1 _2848_ (.Y(_0892_),
    .A(_0888_),
    .B(_0891_));
 sg13g2_o21ai_1 _2849_ (.B1(_0838_),
    .Y(_0893_),
    .A1(_0816_),
    .A2(_0825_));
 sg13g2_nand3_1 _2850_ (.B(_0837_),
    .C(_0830_),
    .A(_0835_),
    .Y(_0894_));
 sg13g2_a21oi_1 _2851_ (.A1(net72),
    .A2(_0894_),
    .Y(_0895_),
    .B1(_0862_));
 sg13g2_nor2_1 _2852_ (.A(net72),
    .B(net94),
    .Y(_0896_));
 sg13g2_nor2_1 _2853_ (.A(net94),
    .B(_0862_),
    .Y(_0897_));
 sg13g2_a21oi_1 _2854_ (.A1(_0830_),
    .A2(_0896_),
    .Y(_0898_),
    .B1(_0897_));
 sg13g2_nand4_1 _2855_ (.B(_0835_),
    .C(_0837_),
    .A(_0350_),
    .Y(_0899_),
    .D(_0830_));
 sg13g2_nand3_1 _2856_ (.B(_0837_),
    .C(_0896_),
    .A(_0835_),
    .Y(_0900_));
 sg13g2_nand3_1 _2857_ (.B(_0899_),
    .C(_0900_),
    .A(_0898_),
    .Y(_0901_));
 sg13g2_a21o_1 _2858_ (.A2(_0895_),
    .A1(_0893_),
    .B1(_0901_),
    .X(_0902_));
 sg13g2_nor2_1 _2859_ (.A(_0039_),
    .B(_0826_),
    .Y(_0903_));
 sg13g2_a21oi_1 _2860_ (.A1(_0526_),
    .A2(net29),
    .Y(_0904_),
    .B1(_0903_));
 sg13g2_nor2_1 _2861_ (.A(_0770_),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_and2_1 _2862_ (.A(_0902_),
    .B(_0905_),
    .X(_0906_));
 sg13g2_buf_1 _2863_ (.A(_0906_),
    .X(_0907_));
 sg13g2_nand2_1 _2864_ (.Y(_0908_),
    .A(net30),
    .B(_0902_));
 sg13g2_nand2_1 _2865_ (.Y(_0909_),
    .A(_0904_),
    .B(_0908_));
 sg13g2_nand3b_1 _2866_ (.B(net76),
    .C(_0909_),
    .Y(_0910_),
    .A_N(_0907_));
 sg13g2_xnor2_1 _2867_ (.Y(_0911_),
    .A(_0465_),
    .B(_0910_));
 sg13g2_xnor2_1 _2868_ (.Y(_0912_),
    .A(_0892_),
    .B(_0911_));
 sg13g2_nand2_1 _2869_ (.Y(_0913_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[7].fa.HA1.a ),
    .B(net42));
 sg13g2_o21ai_1 _2870_ (.B1(_0913_),
    .Y(_0251_),
    .A1(net19),
    .A2(_0912_));
 sg13g2_nand2_1 _2871_ (.Y(_0914_),
    .A(net76),
    .B(_0698_));
 sg13g2_nor2_1 _2872_ (.A(_0040_),
    .B(_0826_),
    .Y(_0915_));
 sg13g2_nand2_1 _2873_ (.Y(_0916_),
    .A(_0532_),
    .B(net29));
 sg13g2_nand2b_1 _2874_ (.Y(_0917_),
    .B(_0916_),
    .A_N(_0915_));
 sg13g2_nand2_1 _2875_ (.Y(_0918_),
    .A(_0465_),
    .B(_0917_));
 sg13g2_nor2b_1 _2876_ (.A(_0915_),
    .B_N(_0916_),
    .Y(_0919_));
 sg13g2_and2_1 _2877_ (.A(_0465_),
    .B(_0919_),
    .X(_0920_));
 sg13g2_nand2_1 _2878_ (.Y(_0921_),
    .A(_0907_),
    .B(_0920_));
 sg13g2_o21ai_1 _2879_ (.B1(_0921_),
    .Y(_0922_),
    .A1(_0909_),
    .A2(_0918_));
 sg13g2_a221oi_1 _2880_ (.B2(_0905_),
    .C1(_0918_),
    .B1(_0902_),
    .A1(_0888_),
    .Y(_0923_),
    .A2(_0891_));
 sg13g2_and4_1 _2881_ (.A(_0888_),
    .B(_0891_),
    .C(_0909_),
    .D(_0920_),
    .X(_0924_));
 sg13g2_nand3b_1 _2882_ (.B(_0909_),
    .C(_0919_),
    .Y(_0925_),
    .A_N(_0465_));
 sg13g2_nand3_1 _2883_ (.B(_0908_),
    .C(_0917_),
    .A(_0904_),
    .Y(_0926_));
 sg13g2_a22oi_1 _2884_ (.Y(_0927_),
    .B1(_0925_),
    .B2(_0926_),
    .A2(_0891_),
    .A1(_0888_));
 sg13g2_nor4_1 _2885_ (.A(_0922_),
    .B(_0923_),
    .C(_0924_),
    .D(_0927_),
    .Y(_0928_));
 sg13g2_xnor2_1 _2886_ (.Y(_0929_),
    .A(_0907_),
    .B(_0919_));
 sg13g2_a21oi_1 _2887_ (.A1(net76),
    .A2(_0929_),
    .Y(_0930_),
    .B1(_0465_));
 sg13g2_and3_1 _2888_ (.X(_0931_),
    .A(_0888_),
    .B(_0891_),
    .C(_0930_));
 sg13g2_a22oi_1 _2889_ (.Y(_0932_),
    .B1(_0698_),
    .B2(_0931_),
    .A2(net57),
    .A1(\rsa_unit_i.mmm_multiply.adder2.gen_fa[8].fa.HA1.a ));
 sg13g2_o21ai_1 _2890_ (.B1(_0932_),
    .Y(_0252_),
    .A1(_0914_),
    .A2(_0928_));
 sg13g2_inv_1 _2891_ (.Y(_0933_),
    .A(_0478_));
 sg13g2_mux2_1 _2892_ (.A0(_0933_),
    .A1(_0080_),
    .S(net50),
    .X(_0934_));
 sg13g2_buf_1 _2893_ (.A(\rsa_unit_i.mmm_square.A_bit ),
    .X(_0935_));
 sg13g2_buf_1 _2894_ (.A(_0935_),
    .X(_0936_));
 sg13g2_buf_1 _2895_ (.A(net71),
    .X(_0937_));
 sg13g2_nand2_1 _2896_ (.Y(_0938_),
    .A(net60),
    .B(_0622_));
 sg13g2_o21ai_1 _2897_ (.B1(_0938_),
    .Y(_0263_),
    .A1(_0597_),
    .A2(_0934_));
 sg13g2_mux2_1 _2898_ (.A0(_0484_),
    .A1(_0083_),
    .S(net50),
    .X(_0939_));
 sg13g2_nand2_1 _2899_ (.Y(_0940_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[1] ),
    .B(_0622_));
 sg13g2_o21ai_1 _2900_ (.B1(_0940_),
    .Y(_0264_),
    .A1(net25),
    .A2(_0939_));
 sg13g2_mux2_1 _2901_ (.A0(_0495_),
    .A1(_0086_),
    .S(net50),
    .X(_0941_));
 sg13g2_buf_1 _2902_ (.A(net57),
    .X(_0942_));
 sg13g2_nand2_1 _2903_ (.Y(_0943_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[2] ),
    .B(net41));
 sg13g2_o21ai_1 _2904_ (.B1(_0943_),
    .Y(_0265_),
    .A1(net25),
    .A2(_0941_));
 sg13g2_mux2_1 _2905_ (.A0(_0500_),
    .A1(_0089_),
    .S(net50),
    .X(_0944_));
 sg13g2_nand2_1 _2906_ (.Y(_0945_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[3] ),
    .B(net41));
 sg13g2_o21ai_1 _2907_ (.B1(_0945_),
    .Y(_0266_),
    .A1(net25),
    .A2(_0944_));
 sg13g2_mux2_1 _2908_ (.A0(_0507_),
    .A1(_0092_),
    .S(net50),
    .X(_0946_));
 sg13g2_nand2_1 _2909_ (.Y(_0947_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[4] ),
    .B(net41));
 sg13g2_o21ai_1 _2910_ (.B1(_0947_),
    .Y(_0267_),
    .A1(net25),
    .A2(_0946_));
 sg13g2_mux2_1 _2911_ (.A0(_0511_),
    .A1(_0095_),
    .S(net50),
    .X(_0948_));
 sg13g2_nand2_1 _2912_ (.Y(_0949_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[5] ),
    .B(net41));
 sg13g2_o21ai_1 _2913_ (.B1(_0949_),
    .Y(_0268_),
    .A1(net25),
    .A2(_0948_));
 sg13g2_mux2_1 _2914_ (.A0(_0516_),
    .A1(_0098_),
    .S(_0618_),
    .X(_0950_));
 sg13g2_nand2_1 _2915_ (.Y(_0951_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[6] ),
    .B(net41));
 sg13g2_o21ai_1 _2916_ (.B1(_0951_),
    .Y(_0269_),
    .A1(net25),
    .A2(_0950_));
 sg13g2_mux2_1 _2917_ (.A0(_0522_),
    .A1(_0101_),
    .S(_0618_),
    .X(_0952_));
 sg13g2_nand2_1 _2918_ (.Y(_0953_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[7] ),
    .B(net41));
 sg13g2_o21ai_1 _2919_ (.B1(_0953_),
    .Y(_0270_),
    .A1(net25),
    .A2(_0952_));
 sg13g2_nor2_1 _2920_ (.A(_0527_),
    .B(_0600_),
    .Y(_0954_));
 sg13g2_a21oi_1 _2921_ (.A1(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[9] ),
    .A2(_0601_),
    .Y(_0955_),
    .B1(_0954_));
 sg13g2_nand2_1 _2922_ (.Y(_0956_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[8] ),
    .B(net41));
 sg13g2_o21ai_1 _2923_ (.B1(_0956_),
    .Y(_0271_),
    .A1(_0596_),
    .A2(_0955_));
 sg13g2_nor3_1 _2924_ (.A(net57),
    .B(net32),
    .C(_0601_),
    .Y(_0957_));
 sg13g2_a22oi_1 _2925_ (.Y(_0958_),
    .B1(_0957_),
    .B2(_0532_),
    .A2(net57),
    .A1(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[9] ));
 sg13g2_inv_1 _2926_ (.Y(_0272_),
    .A(_0958_));
 sg13g2_xor2_1 _2927_ (.B(_0105_),
    .A(net99),
    .X(_0959_));
 sg13g2_nor3_1 _2928_ (.A(net54),
    .B(net64),
    .C(_0959_),
    .Y(_0960_));
 sg13g2_xor2_1 _2929_ (.B(net92),
    .A(_0081_),
    .X(_0961_));
 sg13g2_a21oi_1 _2930_ (.A1(_0398_),
    .A2(_0472_),
    .Y(_0962_),
    .B1(_0961_));
 sg13g2_o21ai_1 _2931_ (.B1(_0935_),
    .Y(_0963_),
    .A1(_0960_),
    .A2(_0962_));
 sg13g2_inv_1 _2932_ (.Y(_0964_),
    .A(\rsa_unit_i.mmm_square.adder2.fa_bit0.HA1.a ));
 sg13g2_buf_1 _2933_ (.A(_0964_),
    .X(_0965_));
 sg13g2_nor2_1 _2934_ (.A(net90),
    .B(net70),
    .Y(_0966_));
 sg13g2_nor2_1 _2935_ (.A(net90),
    .B(_1460_),
    .Y(_0967_));
 sg13g2_mux2_1 _2936_ (.A0(net99),
    .A1(net92),
    .S(_0490_),
    .X(_0968_));
 sg13g2_nand2b_1 _2937_ (.Y(_0969_),
    .B(net90),
    .A_N(_1459_));
 sg13g2_a21oi_1 _2938_ (.A1(_0476_),
    .A2(_0969_),
    .Y(_0970_),
    .B1(net92));
 sg13g2_nor2_1 _2939_ (.A(_0383_),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_a21oi_1 _2940_ (.A1(_0646_),
    .A2(_1460_),
    .Y(_0972_),
    .B1(net90));
 sg13g2_nor3_1 _2941_ (.A(_0646_),
    .B(_1460_),
    .C(\rsa_unit_i.mmm_square.adder2.fa_bit0.HA1.a ),
    .Y(_0973_));
 sg13g2_o21ai_1 _2942_ (.B1(_0476_),
    .Y(_0974_),
    .A1(_0972_),
    .A2(_0973_));
 sg13g2_nand2b_1 _2943_ (.Y(_0975_),
    .B(net99),
    .A_N(_0105_));
 sg13g2_nand2b_1 _2944_ (.Y(_0976_),
    .B(_1459_),
    .A_N(net99));
 sg13g2_a21oi_1 _2945_ (.A1(_0975_),
    .A2(_0976_),
    .Y(_0977_),
    .B1(net90));
 sg13g2_inv_1 _2946_ (.Y(_0978_),
    .A(_0105_));
 sg13g2_a21oi_1 _2947_ (.A1(_0978_),
    .A2(_0969_),
    .Y(_0979_),
    .B1(net99));
 sg13g2_buf_1 _2948_ (.A(\rsa_unit_i.mmm_square.adder2.fa_bit0.HA1.a ),
    .X(_0980_));
 sg13g2_nor3_1 _2949_ (.A(_1460_),
    .B(net88),
    .C(_0975_),
    .Y(_0981_));
 sg13g2_nor4_1 _2950_ (.A(net43),
    .B(_0977_),
    .C(_0979_),
    .D(_0981_),
    .Y(_0982_));
 sg13g2_a221oi_1 _2951_ (.B2(_0974_),
    .C1(_0982_),
    .B1(_0971_),
    .A1(_0967_),
    .Y(_0983_),
    .A2(_0968_));
 sg13g2_and2_1 _2952_ (.A(net90),
    .B(\rsa_unit_i.P_i[1] ),
    .X(_0984_));
 sg13g2_o21ai_1 _2953_ (.B1(_0984_),
    .Y(_0985_),
    .A1(_0378_),
    .A2(net64));
 sg13g2_nand4_1 _2954_ (.B(net99),
    .C(_0397_),
    .A(_0629_),
    .Y(_0986_),
    .D(_0471_));
 sg13g2_nand2_1 _2955_ (.Y(_0987_),
    .A(_0985_),
    .B(_0986_));
 sg13g2_o21ai_1 _2956_ (.B1(net71),
    .Y(_0988_),
    .A1(net70),
    .A2(_0987_));
 sg13g2_nor2_1 _2957_ (.A(_0983_),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_a21oi_1 _2958_ (.A1(_0963_),
    .A2(_0966_),
    .Y(_0990_),
    .B1(_0989_));
 sg13g2_nor4_2 _2959_ (.A(_1391_),
    .B(_0978_),
    .C(_0379_),
    .Y(_0991_),
    .D(_0404_));
 sg13g2_nor2_2 _2960_ (.A(_0477_),
    .B(_0991_),
    .Y(_0992_));
 sg13g2_inv_1 _2961_ (.Y(_0993_),
    .A(_0935_));
 sg13g2_buf_1 _2962_ (.A(_0993_),
    .X(_0994_));
 sg13g2_nor3_1 _2963_ (.A(_1459_),
    .B(net59),
    .C(_0106_),
    .Y(_0995_));
 sg13g2_nand2_1 _2964_ (.Y(_0996_),
    .A(_1514_),
    .B(_0993_));
 sg13g2_nand2_1 _2965_ (.Y(_0997_),
    .A(_1459_),
    .B(_0935_));
 sg13g2_nand2b_1 _2966_ (.Y(_0998_),
    .B(net88),
    .A_N(_0106_));
 sg13g2_a21oi_1 _2967_ (.A1(_0996_),
    .A2(_0997_),
    .Y(_0999_),
    .B1(_0998_));
 sg13g2_a21o_1 _2968_ (.A2(_0995_),
    .A1(_0992_),
    .B1(_0999_),
    .X(_1000_));
 sg13g2_xnor2_1 _2969_ (.Y(_1001_),
    .A(_0483_),
    .B(_1000_));
 sg13g2_xnor2_1 _2970_ (.Y(_1002_),
    .A(_0990_),
    .B(_1001_));
 sg13g2_nand2_1 _2971_ (.Y(_1003_),
    .A(net88),
    .B(net41));
 sg13g2_o21ai_1 _2972_ (.B1(_1003_),
    .Y(_0273_),
    .A1(net19),
    .A2(_1002_));
 sg13g2_nand3_1 _2973_ (.B(_0397_),
    .C(_0471_),
    .A(_0108_),
    .Y(_1004_));
 sg13g2_buf_1 _2974_ (.A(_1004_),
    .X(_1005_));
 sg13g2_nand2_1 _2975_ (.Y(_1006_),
    .A(_0494_),
    .B(_1005_));
 sg13g2_nor4_1 _2976_ (.A(net89),
    .B(net88),
    .C(_0477_),
    .D(_0991_),
    .Y(_1007_));
 sg13g2_and2_1 _2977_ (.A(_1006_),
    .B(_1007_),
    .X(_1008_));
 sg13g2_and2_1 _2978_ (.A(_0494_),
    .B(_1005_),
    .X(_1009_));
 sg13g2_buf_1 _2979_ (.A(_1009_),
    .X(_1010_));
 sg13g2_o21ai_1 _2980_ (.B1(_0081_),
    .Y(_1011_),
    .A1(_0379_),
    .A2(net64));
 sg13g2_or4_1 _2981_ (.A(_1391_),
    .B(_0978_),
    .C(net54),
    .D(_0404_),
    .X(_1012_));
 sg13g2_buf_1 _2982_ (.A(_1012_),
    .X(_1013_));
 sg13g2_nand4_1 _2983_ (.B(_0964_),
    .C(_1011_),
    .A(net89),
    .Y(_1014_),
    .D(_1013_));
 sg13g2_nor2_1 _2984_ (.A(_1010_),
    .B(_1014_),
    .Y(_1015_));
 sg13g2_o21ai_1 _2985_ (.B1(_1467_),
    .Y(_1016_),
    .A1(_1540_),
    .A2(_1460_));
 sg13g2_mux2_1 _2986_ (.A0(_0967_),
    .A1(_1016_),
    .S(_0968_),
    .X(_1017_));
 sg13g2_mux2_1 _2987_ (.A0(_1008_),
    .A1(_1015_),
    .S(_1017_),
    .X(_1018_));
 sg13g2_nand4_1 _2988_ (.B(_1466_),
    .C(net62),
    .A(net99),
    .Y(_1019_),
    .D(net61));
 sg13g2_and2_1 _2989_ (.A(net92),
    .B(\rsa_spi_wrapper_i.config_regs[33] ),
    .X(_1020_));
 sg13g2_buf_1 _2990_ (.A(_1020_),
    .X(_1021_));
 sg13g2_o21ai_1 _2991_ (.B1(_1021_),
    .Y(_1022_),
    .A1(net54),
    .A2(net64));
 sg13g2_nand2_1 _2992_ (.Y(_1023_),
    .A(_1019_),
    .B(_1022_));
 sg13g2_nor3_2 _2993_ (.A(_1460_),
    .B(_0477_),
    .C(_0991_),
    .Y(_1024_));
 sg13g2_nor3_1 _2994_ (.A(_1564_),
    .B(_1023_),
    .C(_1024_),
    .Y(_1025_));
 sg13g2_nor2_1 _2995_ (.A(_0629_),
    .B(_0487_),
    .Y(_1026_));
 sg13g2_o21ai_1 _2996_ (.B1(_1026_),
    .Y(_1027_),
    .A1(net54),
    .A2(net64));
 sg13g2_nand4_1 _2997_ (.B(_1455_),
    .C(net62),
    .A(_1540_),
    .Y(_1028_),
    .D(net61));
 sg13g2_nand4_1 _2998_ (.B(_0986_),
    .C(_1027_),
    .A(_0985_),
    .Y(_1029_),
    .D(_1028_));
 sg13g2_buf_1 _2999_ (.A(_1029_),
    .X(_1030_));
 sg13g2_nand3_1 _3000_ (.B(_1024_),
    .C(_1030_),
    .A(_1564_),
    .Y(_1031_));
 sg13g2_nand2_1 _3001_ (.Y(_1032_),
    .A(_1011_),
    .B(_1013_));
 sg13g2_buf_2 _3002_ (.A(_1032_),
    .X(_1033_));
 sg13g2_and4_1 _3003_ (.A(_0985_),
    .B(_0986_),
    .C(_1027_),
    .D(_1028_),
    .X(_1034_));
 sg13g2_and3_1 _3004_ (.X(_1035_),
    .A(net89),
    .B(_1019_),
    .C(_1022_));
 sg13g2_a21oi_1 _3005_ (.A1(_1019_),
    .A2(_1022_),
    .Y(_1036_),
    .B1(_0665_));
 sg13g2_a221oi_1 _3006_ (.B2(_1035_),
    .C1(_1036_),
    .B1(_1034_),
    .A1(_0965_),
    .Y(_1037_),
    .A2(_1033_));
 sg13g2_nand3b_1 _3007_ (.B(_1031_),
    .C(_1037_),
    .Y(_1038_),
    .A_N(_1025_));
 sg13g2_nor2_1 _3008_ (.A(net59),
    .B(_1006_),
    .Y(_1039_));
 sg13g2_nand4_1 _3009_ (.B(_0108_),
    .C(net62),
    .A(_0105_),
    .Y(_1040_),
    .D(net61));
 sg13g2_and2_1 _3010_ (.A(_0081_),
    .B(_0087_),
    .X(_1041_));
 sg13g2_o21ai_1 _3011_ (.B1(_1041_),
    .Y(_1042_),
    .A1(net54),
    .A2(net64));
 sg13g2_a21oi_1 _3012_ (.A1(_1040_),
    .A2(_1042_),
    .Y(_1043_),
    .B1(_1564_));
 sg13g2_a22oi_1 _3013_ (.Y(_1044_),
    .B1(_1023_),
    .B2(_1043_),
    .A2(_1010_),
    .A1(_0992_));
 sg13g2_nand2_1 _3014_ (.Y(_1045_),
    .A(net71),
    .B(net88));
 sg13g2_nand2_1 _3015_ (.Y(_1046_),
    .A(_1454_),
    .B(net98));
 sg13g2_nor3_1 _3016_ (.A(net54),
    .B(_0381_),
    .C(_1046_),
    .Y(_1047_));
 sg13g2_a221oi_1 _3017_ (.B2(_1042_),
    .C1(_1047_),
    .B1(_1040_),
    .A1(_0491_),
    .Y(_1048_),
    .A2(_1021_));
 sg13g2_nor2_1 _3018_ (.A(_0665_),
    .B(_0965_),
    .Y(_1049_));
 sg13g2_o21ai_1 _3019_ (.B1(_1049_),
    .Y(_1050_),
    .A1(_0994_),
    .A2(_1048_));
 sg13g2_o21ai_1 _3020_ (.B1(_1050_),
    .Y(_1051_),
    .A1(_1044_),
    .A2(_1045_));
 sg13g2_a221oi_1 _3021_ (.B2(_1039_),
    .C1(_1051_),
    .B1(_1038_),
    .A1(net71),
    .Y(_1052_),
    .A2(_1018_));
 sg13g2_buf_1 _3022_ (.A(_1052_),
    .X(_1053_));
 sg13g2_a221oi_1 _3023_ (.B2(_0995_),
    .C1(_0999_),
    .B1(_0992_),
    .A1(_0963_),
    .Y(_1054_),
    .A2(_0966_));
 sg13g2_o21ai_1 _3024_ (.B1(_1054_),
    .Y(_1055_),
    .A1(_0983_),
    .A2(_0988_));
 sg13g2_nand2b_1 _3025_ (.Y(_1056_),
    .B(_0104_),
    .A_N(_1000_));
 sg13g2_a21oi_1 _3026_ (.A1(_0963_),
    .A2(_0966_),
    .Y(_1057_),
    .B1(_0483_));
 sg13g2_o21ai_1 _3027_ (.B1(_1057_),
    .Y(_1058_),
    .A1(_0983_),
    .A2(_0988_));
 sg13g2_nand3_1 _3028_ (.B(_1056_),
    .C(_1058_),
    .A(_1055_),
    .Y(_1059_));
 sg13g2_xnor2_1 _3029_ (.Y(_1060_),
    .A(_0107_),
    .B(_1059_));
 sg13g2_xnor2_1 _3030_ (.Y(_1061_),
    .A(_1053_),
    .B(_1060_));
 sg13g2_nand2_1 _3031_ (.Y(_1062_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[1].fa.HA1.a ),
    .B(_0942_));
 sg13g2_o21ai_1 _3032_ (.B1(_1062_),
    .Y(_0274_),
    .A1(_0628_),
    .A2(_1061_));
 sg13g2_nand2_1 _3033_ (.Y(_1063_),
    .A(_1053_),
    .B(_1059_));
 sg13g2_o21ai_1 _3034_ (.B1(_0107_),
    .Y(_1064_),
    .A1(_1053_),
    .A2(_1059_));
 sg13g2_nand2_1 _3035_ (.Y(_1065_),
    .A(_1063_),
    .B(_1064_));
 sg13g2_o21ai_1 _3036_ (.B1(net88),
    .Y(_1066_),
    .A1(_0477_),
    .A2(_0991_));
 sg13g2_buf_2 _3037_ (.A(_1066_),
    .X(_1067_));
 sg13g2_a21oi_1 _3038_ (.A1(_0110_),
    .A2(net39),
    .Y(_1068_),
    .B1(_0499_));
 sg13g2_buf_1 _3039_ (.A(_1068_),
    .X(_1069_));
 sg13g2_a221oi_1 _3040_ (.B2(_0494_),
    .C1(_1047_),
    .B1(_1005_),
    .A1(_0491_),
    .Y(_1070_),
    .A2(_1021_));
 sg13g2_nand3b_1 _3041_ (.B(_0487_),
    .C(net98),
    .Y(_1071_),
    .A_N(_0087_));
 sg13g2_a21oi_1 _3042_ (.A1(_0398_),
    .A2(_0472_),
    .Y(_1072_),
    .B1(_1071_));
 sg13g2_nor4_1 _3043_ (.A(_0108_),
    .B(net54),
    .C(_0381_),
    .D(_1046_),
    .Y(_1073_));
 sg13g2_nor3_2 _3044_ (.A(_1564_),
    .B(_1072_),
    .C(_1073_),
    .Y(_1074_));
 sg13g2_or4_1 _3045_ (.A(_1586_),
    .B(_1069_),
    .C(_1070_),
    .D(_1074_),
    .X(_1075_));
 sg13g2_nand3_1 _3046_ (.B(_1011_),
    .C(_1013_),
    .A(_0964_),
    .Y(_1076_));
 sg13g2_buf_2 _3047_ (.A(_1076_),
    .X(_1077_));
 sg13g2_nand3_1 _3048_ (.B(_1069_),
    .C(_1067_),
    .A(_1077_),
    .Y(_1078_));
 sg13g2_o21ai_1 _3049_ (.B1(_1078_),
    .Y(_1079_),
    .A1(_1067_),
    .A2(_1075_));
 sg13g2_nand2_1 _3050_ (.Y(_1080_),
    .A(_1024_),
    .B(_1030_));
 sg13g2_nand3_1 _3051_ (.B(_1024_),
    .C(_1030_),
    .A(_1010_),
    .Y(_1081_));
 sg13g2_buf_2 _3052_ (.A(_1081_),
    .X(_1082_));
 sg13g2_nand2_1 _3053_ (.Y(_1083_),
    .A(_1586_),
    .B(_1069_));
 sg13g2_a221oi_1 _3054_ (.B2(_1082_),
    .C1(_1083_),
    .B1(_1074_),
    .A1(_1080_),
    .Y(_1084_),
    .A2(_1070_));
 sg13g2_o21ai_1 _3055_ (.B1(net71),
    .Y(_1085_),
    .A1(_1079_),
    .A2(_1084_));
 sg13g2_nand3_1 _3056_ (.B(net71),
    .C(_1069_),
    .A(net74),
    .Y(_1086_));
 sg13g2_nor2_1 _3057_ (.A(_0980_),
    .B(_1033_),
    .Y(_1087_));
 sg13g2_a21o_1 _3058_ (.A2(net39),
    .A1(_0110_),
    .B1(_0499_),
    .X(_1088_));
 sg13g2_buf_1 _3059_ (.A(_1088_),
    .X(_1089_));
 sg13g2_nand4_1 _3060_ (.B(net71),
    .C(_1087_),
    .A(net74),
    .Y(_1090_),
    .D(net28));
 sg13g2_a221oi_1 _3061_ (.B2(_1030_),
    .C1(_1023_),
    .B1(_1024_),
    .A1(_0494_),
    .Y(_1091_),
    .A2(_1005_));
 sg13g2_a21oi_2 _3062_ (.B1(_1091_),
    .Y(_1092_),
    .A2(_1082_),
    .A1(_1074_));
 sg13g2_mux2_1 _3063_ (.A0(_1086_),
    .A1(_1090_),
    .S(_1092_),
    .X(_1093_));
 sg13g2_o21ai_1 _3064_ (.B1(net28),
    .Y(_1094_),
    .A1(_1070_),
    .A2(_1074_));
 sg13g2_o21ai_1 _3065_ (.B1(_0936_),
    .Y(_1095_),
    .A1(_0992_),
    .A2(_1094_));
 sg13g2_nor2_1 _3066_ (.A(net74),
    .B(net70),
    .Y(_1096_));
 sg13g2_nor4_1 _3067_ (.A(net97),
    .B(net59),
    .C(_1077_),
    .D(_1069_),
    .Y(_1097_));
 sg13g2_a21o_1 _3068_ (.A2(_1082_),
    .A1(_1074_),
    .B1(_1091_),
    .X(_1098_));
 sg13g2_a22oi_1 _3069_ (.Y(_1099_),
    .B1(_1097_),
    .B2(_1098_),
    .A2(_1096_),
    .A1(_1095_));
 sg13g2_nand3_1 _3070_ (.B(_1093_),
    .C(_1099_),
    .A(_1085_),
    .Y(_1100_));
 sg13g2_xor2_1 _3071_ (.B(_1100_),
    .A(_0109_),
    .X(_1101_));
 sg13g2_xnor2_1 _3072_ (.Y(_1102_),
    .A(_1065_),
    .B(_1101_));
 sg13g2_nand2_1 _3073_ (.Y(_1103_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[2].fa.HA1.a ),
    .B(_0942_));
 sg13g2_o21ai_1 _3074_ (.B1(_1103_),
    .Y(_0275_),
    .A1(_0628_),
    .A2(_1102_));
 sg13g2_nand4_1 _3075_ (.B(_1085_),
    .C(_1093_),
    .A(_0109_),
    .Y(_1104_),
    .D(_1099_));
 sg13g2_nand3_1 _3076_ (.B(_1064_),
    .C(_1104_),
    .A(_1063_),
    .Y(_1105_));
 sg13g2_buf_1 _3077_ (.A(_1105_),
    .X(_1106_));
 sg13g2_nand2b_1 _3078_ (.Y(_1107_),
    .B(_1100_),
    .A_N(_0109_));
 sg13g2_nand2_1 _3079_ (.Y(_1108_),
    .A(_1106_),
    .B(_1107_));
 sg13g2_a21oi_1 _3080_ (.A1(_0112_),
    .A2(net39),
    .Y(_1109_),
    .B1(_0506_));
 sg13g2_buf_1 _3081_ (.A(_1109_),
    .X(_1110_));
 sg13g2_nand3_1 _3082_ (.B(_1083_),
    .C(_1110_),
    .A(net73),
    .Y(_1111_));
 sg13g2_nand2_2 _3083_ (.Y(_1112_),
    .A(_1077_),
    .B(_1067_));
 sg13g2_nand2_1 _3084_ (.Y(_1113_),
    .A(net97),
    .B(_1089_));
 sg13g2_a21o_1 _3085_ (.A2(_0383_),
    .A1(_0112_),
    .B1(_0506_),
    .X(_1114_));
 sg13g2_buf_1 _3086_ (.A(_1114_),
    .X(_1115_));
 sg13g2_nand4_1 _3087_ (.B(_1112_),
    .C(_1113_),
    .A(_1608_),
    .Y(_1116_),
    .D(net27));
 sg13g2_mux2_1 _3088_ (.A0(_1111_),
    .A1(_1116_),
    .S(_1092_),
    .X(_1117_));
 sg13g2_and2_1 _3089_ (.A(_1077_),
    .B(_1067_),
    .X(_1118_));
 sg13g2_buf_1 _3090_ (.A(_1118_),
    .X(_1119_));
 sg13g2_nand3_1 _3091_ (.B(_1069_),
    .C(net27),
    .A(_1586_),
    .Y(_1120_));
 sg13g2_nand3_1 _3092_ (.B(net28),
    .C(_1110_),
    .A(net97),
    .Y(_1121_));
 sg13g2_o21ai_1 _3093_ (.B1(_1121_),
    .Y(_1122_),
    .A1(_1119_),
    .A2(_1120_));
 sg13g2_a22oi_1 _3094_ (.Y(_1123_),
    .B1(_1122_),
    .B2(net73),
    .A2(_1110_),
    .A1(_1119_));
 sg13g2_nand2_1 _3095_ (.Y(_1124_),
    .A(_1117_),
    .B(_1123_));
 sg13g2_nor2_1 _3096_ (.A(net73),
    .B(net70),
    .Y(_1125_));
 sg13g2_nor2_1 _3097_ (.A(net97),
    .B(net28),
    .Y(_1126_));
 sg13g2_buf_1 _3098_ (.A(_1126_),
    .X(_1127_));
 sg13g2_a221oi_1 _3099_ (.B2(_1082_),
    .C1(_1091_),
    .B1(_1074_),
    .A1(_1585_),
    .Y(_1128_),
    .A2(net28));
 sg13g2_buf_1 _3100_ (.A(_1128_),
    .X(_1129_));
 sg13g2_nor4_1 _3101_ (.A(_0992_),
    .B(net24),
    .C(_1110_),
    .D(net18),
    .Y(_1130_));
 sg13g2_nand2b_1 _3102_ (.Y(_1131_),
    .B(net71),
    .A_N(_1130_));
 sg13g2_or4_1 _3103_ (.A(_1077_),
    .B(net24),
    .C(_1110_),
    .D(net18),
    .X(_1132_));
 sg13g2_o21ai_1 _3104_ (.B1(_1110_),
    .Y(_1133_),
    .A1(net24),
    .A2(net18));
 sg13g2_nand2_1 _3105_ (.Y(_1134_),
    .A(_1609_),
    .B(_0936_));
 sg13g2_a21oi_1 _3106_ (.A1(_1132_),
    .A2(_1133_),
    .Y(_1135_),
    .B1(_1134_));
 sg13g2_a221oi_1 _3107_ (.B2(_1131_),
    .C1(_1135_),
    .B1(_1125_),
    .A1(_0937_),
    .Y(_1136_),
    .A2(_1124_));
 sg13g2_buf_2 _3108_ (.A(_1136_),
    .X(_1137_));
 sg13g2_xnor2_1 _3109_ (.Y(_1138_),
    .A(_0504_),
    .B(_1137_));
 sg13g2_xnor2_1 _3110_ (.Y(_1139_),
    .A(_1108_),
    .B(_1138_));
 sg13g2_nand2_1 _3111_ (.Y(_1140_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[3].fa.HA1.a ),
    .B(net49));
 sg13g2_o21ai_1 _3112_ (.B1(_1140_),
    .Y(_0276_),
    .A1(_0627_),
    .A2(_1139_));
 sg13g2_a22oi_1 _3113_ (.Y(_1141_),
    .B1(_1137_),
    .B2(_0503_),
    .A2(_1107_),
    .A1(_1106_));
 sg13g2_nor3_1 _3114_ (.A(net73),
    .B(net70),
    .C(_0503_),
    .Y(_1142_));
 sg13g2_nand2_1 _3115_ (.Y(_1143_),
    .A(net60),
    .B(_0504_));
 sg13g2_a21oi_1 _3116_ (.A1(_1117_),
    .A2(_1123_),
    .Y(_1144_),
    .B1(_1143_));
 sg13g2_a221oi_1 _3117_ (.B2(_1142_),
    .C1(_1144_),
    .B1(_1131_),
    .A1(_0504_),
    .Y(_1145_),
    .A2(_1135_));
 sg13g2_nor2b_1 _3118_ (.A(_1141_),
    .B_N(_1145_),
    .Y(_1146_));
 sg13g2_mux2_1 _3119_ (.A0(_0096_),
    .A1(_0114_),
    .S(_0382_),
    .X(_1147_));
 sg13g2_buf_2 _3120_ (.A(_1147_),
    .X(_1148_));
 sg13g2_nand2b_1 _3121_ (.Y(_1149_),
    .B(_1625_),
    .A_N(_1148_));
 sg13g2_buf_2 _3122_ (.A(_1149_),
    .X(_1150_));
 sg13g2_nand2_1 _3123_ (.Y(_1151_),
    .A(net96),
    .B(_1148_));
 sg13g2_nand2_1 _3124_ (.Y(_1152_),
    .A(_1150_),
    .B(_1151_));
 sg13g2_nor2_1 _3125_ (.A(net73),
    .B(net27),
    .Y(_1153_));
 sg13g2_or3_1 _3126_ (.A(net24),
    .B(net18),
    .C(_1153_),
    .X(_1154_));
 sg13g2_nor3_1 _3127_ (.A(net24),
    .B(net18),
    .C(_1152_),
    .Y(_1155_));
 sg13g2_nand2_1 _3128_ (.Y(_1156_),
    .A(net60),
    .B(_1112_));
 sg13g2_a221oi_1 _3129_ (.B2(_1115_),
    .C1(_1156_),
    .B1(_1155_),
    .A1(_1152_),
    .Y(_1157_),
    .A2(_1154_));
 sg13g2_or3_1 _3130_ (.A(net24),
    .B(net18),
    .C(_1152_),
    .X(_1158_));
 sg13g2_o21ai_1 _3131_ (.B1(_1115_),
    .Y(_1159_),
    .A1(_1127_),
    .A2(_1129_));
 sg13g2_a21o_1 _3132_ (.A2(_1159_),
    .A1(_1158_),
    .B1(_1609_),
    .X(_1160_));
 sg13g2_nor2_1 _3133_ (.A(net96),
    .B(_1148_),
    .Y(_1161_));
 sg13g2_o21ai_1 _3134_ (.B1(_1077_),
    .Y(_1162_),
    .A1(net59),
    .A2(_1067_));
 sg13g2_nand4_1 _3135_ (.B(net27),
    .C(_1161_),
    .A(net73),
    .Y(_1163_),
    .D(_1162_));
 sg13g2_nand2_1 _3136_ (.Y(_1164_),
    .A(_1608_),
    .B(net27));
 sg13g2_nor2b_1 _3137_ (.A(_1164_),
    .B_N(_1148_),
    .Y(_1165_));
 sg13g2_o21ai_1 _3138_ (.B1(_1624_),
    .Y(_1166_),
    .A1(net59),
    .A2(_1165_));
 sg13g2_nand4_1 _3139_ (.B(_0980_),
    .C(_0992_),
    .A(net60),
    .Y(_1167_),
    .D(_1148_));
 sg13g2_a21oi_1 _3140_ (.A1(_1033_),
    .A2(_1148_),
    .Y(_1168_),
    .B1(_0994_));
 sg13g2_or2_1 _3141_ (.X(_1169_),
    .B(_1168_),
    .A(net88));
 sg13g2_nand4_1 _3142_ (.B(_1166_),
    .C(_1167_),
    .A(_1163_),
    .Y(_1170_),
    .D(_1169_));
 sg13g2_a21o_1 _3143_ (.A2(_1160_),
    .A1(_1157_),
    .B1(_1170_),
    .X(_1171_));
 sg13g2_xnor2_1 _3144_ (.Y(_1172_),
    .A(_0512_),
    .B(_1171_));
 sg13g2_xnor2_1 _3145_ (.Y(_1173_),
    .A(_1146_),
    .B(_1172_));
 sg13g2_nand2_1 _3146_ (.Y(_1174_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[4].fa.HA1.a ),
    .B(net49));
 sg13g2_o21ai_1 _3147_ (.B1(_1174_),
    .Y(_0277_),
    .A1(_0627_),
    .A2(_1173_));
 sg13g2_a21oi_1 _3148_ (.A1(_0116_),
    .A2(net39),
    .Y(_1175_),
    .B1(_0515_));
 sg13g2_nand2_1 _3149_ (.Y(_1176_),
    .A(net95),
    .B(_1175_));
 sg13g2_a21o_1 _3150_ (.A2(net39),
    .A1(_0116_),
    .B1(_0515_),
    .X(_1177_));
 sg13g2_buf_2 _3151_ (.A(_1177_),
    .X(_1178_));
 sg13g2_nand3_1 _3152_ (.B(_1087_),
    .C(_1178_),
    .A(net95),
    .Y(_1179_));
 sg13g2_and2_1 _3153_ (.A(_1624_),
    .B(_1148_),
    .X(_1180_));
 sg13g2_buf_1 _3154_ (.A(_1180_),
    .X(_1181_));
 sg13g2_nand3_1 _3155_ (.B(net27),
    .C(_1150_),
    .A(net28),
    .Y(_1182_));
 sg13g2_nand3_1 _3156_ (.B(net27),
    .C(_1150_),
    .A(net74),
    .Y(_1183_));
 sg13g2_a21oi_1 _3157_ (.A1(_1182_),
    .A2(_1183_),
    .Y(_1184_),
    .B1(_1092_));
 sg13g2_nand3_1 _3158_ (.B(net28),
    .C(_1150_),
    .A(_0743_),
    .Y(_1185_));
 sg13g2_nand3_1 _3159_ (.B(_1608_),
    .C(_1150_),
    .A(net74),
    .Y(_1186_));
 sg13g2_a21oi_1 _3160_ (.A1(_1185_),
    .A2(_1186_),
    .Y(_1187_),
    .B1(_1092_));
 sg13g2_nor3_1 _3161_ (.A(_1069_),
    .B(_1110_),
    .C(_1161_),
    .Y(_1188_));
 sg13g2_nand3_1 _3162_ (.B(_1608_),
    .C(net28),
    .A(_1585_),
    .Y(_1189_));
 sg13g2_a21oi_1 _3163_ (.A1(_1164_),
    .A2(_1189_),
    .Y(_1190_),
    .B1(_1161_));
 sg13g2_a21o_1 _3164_ (.A2(_1188_),
    .A1(_0701_),
    .B1(_1190_),
    .X(_1191_));
 sg13g2_nor4_1 _3165_ (.A(_1181_),
    .B(_1184_),
    .C(_1187_),
    .D(_1191_),
    .Y(_1192_));
 sg13g2_mux2_1 _3166_ (.A0(_1176_),
    .A1(_1179_),
    .S(_1192_),
    .X(_1193_));
 sg13g2_a21o_1 _3167_ (.A2(_1183_),
    .A1(_1182_),
    .B1(_1092_),
    .X(_1194_));
 sg13g2_a21o_1 _3168_ (.A2(_1186_),
    .A1(_1185_),
    .B1(_1092_),
    .X(_1195_));
 sg13g2_a21oi_1 _3169_ (.A1(_0701_),
    .A2(_1188_),
    .Y(_1196_),
    .B1(_1190_));
 sg13g2_nor2_1 _3170_ (.A(_1181_),
    .B(_1178_),
    .Y(_1197_));
 sg13g2_and4_1 _3171_ (.A(_1194_),
    .B(_1195_),
    .C(_1196_),
    .D(_1197_),
    .X(_1198_));
 sg13g2_buf_2 _3172_ (.A(_1198_),
    .X(_1199_));
 sg13g2_nor2_1 _3173_ (.A(net72),
    .B(_1077_),
    .Y(_1200_));
 sg13g2_nand3_1 _3174_ (.B(_1150_),
    .C(_1178_),
    .A(net27),
    .Y(_1201_));
 sg13g2_nor3_2 _3175_ (.A(net24),
    .B(net18),
    .C(_1201_),
    .Y(_1202_));
 sg13g2_nand3_1 _3176_ (.B(_1150_),
    .C(_1178_),
    .A(_0743_),
    .Y(_1203_));
 sg13g2_nor3_2 _3177_ (.A(net24),
    .B(net18),
    .C(_1203_),
    .Y(_1204_));
 sg13g2_nand2_1 _3178_ (.Y(_1205_),
    .A(_1181_),
    .B(_1178_));
 sg13g2_o21ai_1 _3179_ (.B1(_1205_),
    .Y(_1206_),
    .A1(_1609_),
    .A2(_1201_));
 sg13g2_buf_1 _3180_ (.A(_1206_),
    .X(_1207_));
 sg13g2_or3_1 _3181_ (.A(_1202_),
    .B(_1204_),
    .C(_1207_),
    .X(_1208_));
 sg13g2_buf_1 _3182_ (.A(_1208_),
    .X(_1209_));
 sg13g2_a22oi_1 _3183_ (.Y(_1210_),
    .B1(_1200_),
    .B2(_1209_),
    .A2(_1199_),
    .A1(_0334_));
 sg13g2_nand3_1 _3184_ (.B(_1033_),
    .C(_1175_),
    .A(net70),
    .Y(_1211_));
 sg13g2_nand4_1 _3185_ (.B(_1033_),
    .C(_1151_),
    .A(net95),
    .Y(_1212_),
    .D(_1178_));
 sg13g2_nor4_1 _3186_ (.A(_1184_),
    .B(_1187_),
    .C(_1191_),
    .D(_1212_),
    .Y(_1213_));
 sg13g2_nor2_1 _3187_ (.A(_1033_),
    .B(_1178_),
    .Y(_1214_));
 sg13g2_o21ai_1 _3188_ (.B1(net88),
    .Y(_1215_),
    .A1(_1213_),
    .A2(_1214_));
 sg13g2_nand4_1 _3189_ (.B(_1210_),
    .C(_1211_),
    .A(_1193_),
    .Y(_1216_),
    .D(_1215_));
 sg13g2_a21oi_1 _3190_ (.A1(_1033_),
    .A2(_1209_),
    .Y(_1217_),
    .B1(net59));
 sg13g2_nor3_1 _3191_ (.A(net72),
    .B(net70),
    .C(_1217_),
    .Y(_1218_));
 sg13g2_a21oi_2 _3192_ (.B1(_1218_),
    .Y(_1219_),
    .A2(_1216_),
    .A1(net60));
 sg13g2_a221oi_1 _3193_ (.B2(_0503_),
    .C1(_1171_),
    .B1(_1137_),
    .A1(_1106_),
    .Y(_1220_),
    .A2(_1107_));
 sg13g2_a21oi_1 _3194_ (.A1(_0512_),
    .A2(_1145_),
    .Y(_1221_),
    .B1(_1171_));
 sg13g2_nor2_1 _3195_ (.A(_0512_),
    .B(_1145_),
    .Y(_1222_));
 sg13g2_a221oi_1 _3196_ (.B2(_0503_),
    .C1(_0512_),
    .B1(_1137_),
    .A1(_1106_),
    .Y(_1223_),
    .A2(_1107_));
 sg13g2_nor4_2 _3197_ (.A(_1220_),
    .B(_1221_),
    .C(_1222_),
    .Y(_1224_),
    .D(_1223_));
 sg13g2_xnor2_1 _3198_ (.Y(_1225_),
    .A(_1219_),
    .B(_1224_));
 sg13g2_xnor2_1 _3199_ (.Y(_1226_),
    .A(_0115_),
    .B(_1225_));
 sg13g2_nand2_1 _3200_ (.Y(_1227_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[5].fa.HA1.a ),
    .B(net49));
 sg13g2_o21ai_1 _3201_ (.B1(_1227_),
    .Y(_0278_),
    .A1(_0627_),
    .A2(_1226_));
 sg13g2_nand2_1 _3202_ (.Y(_1228_),
    .A(_1219_),
    .B(_1224_));
 sg13g2_o21ai_1 _3203_ (.B1(_0115_),
    .Y(_1229_),
    .A1(_1219_),
    .A2(_1224_));
 sg13g2_buf_1 _3204_ (.A(_1229_),
    .X(_1230_));
 sg13g2_nand2_1 _3205_ (.Y(_1231_),
    .A(_1228_),
    .B(_1230_));
 sg13g2_a21oi_1 _3206_ (.A1(_0021_),
    .A2(net39),
    .Y(_1232_),
    .B1(_0521_));
 sg13g2_buf_2 _3207_ (.A(_1232_),
    .X(_1233_));
 sg13g2_nand2_1 _3208_ (.Y(_1234_),
    .A(_1119_),
    .B(_1233_));
 sg13g2_nand4_1 _3209_ (.B(_1195_),
    .C(_1196_),
    .A(_1194_),
    .Y(_1235_),
    .D(_1197_));
 sg13g2_buf_1 _3210_ (.A(_1235_),
    .X(_1236_));
 sg13g2_or4_1 _3211_ (.A(net95),
    .B(_1202_),
    .C(_1204_),
    .D(_1207_),
    .X(_1237_));
 sg13g2_nand4_1 _3212_ (.B(_1236_),
    .C(_1237_),
    .A(net94),
    .Y(_1238_),
    .D(_1233_));
 sg13g2_nor4_2 _3213_ (.A(_0333_),
    .B(_1202_),
    .C(_1204_),
    .Y(_1239_),
    .D(_1207_));
 sg13g2_nor3_1 _3214_ (.A(_0350_),
    .B(_1119_),
    .C(_1233_),
    .Y(_1240_));
 sg13g2_o21ai_1 _3215_ (.B1(_1240_),
    .Y(_1241_),
    .A1(_1199_),
    .A2(_1239_));
 sg13g2_nand3_1 _3216_ (.B(_1238_),
    .C(_1241_),
    .A(_1234_),
    .Y(_1242_));
 sg13g2_nand3_1 _3217_ (.B(_1236_),
    .C(_1237_),
    .A(_1087_),
    .Y(_1243_));
 sg13g2_o21ai_1 _3218_ (.B1(_1233_),
    .Y(_1244_),
    .A1(_1199_),
    .A2(_1239_));
 sg13g2_o21ai_1 _3219_ (.B1(_1244_),
    .Y(_1245_),
    .A1(_1233_),
    .A2(_1243_));
 sg13g2_nor2_1 _3220_ (.A(net94),
    .B(net59),
    .Y(_1246_));
 sg13g2_nor2_1 _3221_ (.A(_1199_),
    .B(_1239_),
    .Y(_1247_));
 sg13g2_nor3_1 _3222_ (.A(net94),
    .B(_1067_),
    .C(_1233_),
    .Y(_1248_));
 sg13g2_nor3_1 _3223_ (.A(net94),
    .B(net60),
    .C(net70),
    .Y(_1249_));
 sg13g2_a21o_1 _3224_ (.A2(_1248_),
    .A1(_1247_),
    .B1(_1249_),
    .X(_1250_));
 sg13g2_a221oi_1 _3225_ (.B2(_1246_),
    .C1(_1250_),
    .B1(_1245_),
    .A1(net60),
    .Y(_1251_),
    .A2(_1242_));
 sg13g2_buf_2 _3226_ (.A(_1251_),
    .X(_1252_));
 sg13g2_xnor2_1 _3227_ (.Y(_1253_),
    .A(_0519_),
    .B(_1252_));
 sg13g2_xnor2_1 _3228_ (.Y(_1254_),
    .A(_1231_),
    .B(_1253_));
 sg13g2_nand2_1 _3229_ (.Y(_1255_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[6].fa.HA1.a ),
    .B(net49));
 sg13g2_o21ai_1 _3230_ (.B1(_1255_),
    .Y(_0279_),
    .A1(_0627_),
    .A2(_1254_));
 sg13g2_a21oi_1 _3231_ (.A1(_1219_),
    .A2(_1224_),
    .Y(_1256_),
    .B1(_1252_));
 sg13g2_a21oi_1 _3232_ (.A1(_1230_),
    .A2(_1256_),
    .Y(_1257_),
    .B1(_0520_));
 sg13g2_a21oi_1 _3233_ (.A1(_1231_),
    .A2(_1252_),
    .Y(_1258_),
    .B1(_1257_));
 sg13g2_buf_1 _3234_ (.A(_0022_),
    .X(_1259_));
 sg13g2_a21o_1 _3235_ (.A2(net39),
    .A1(_0021_),
    .B1(_0521_),
    .X(_1260_));
 sg13g2_buf_1 _3236_ (.A(_1260_),
    .X(_1261_));
 sg13g2_and2_1 _3237_ (.A(_0527_),
    .B(_1261_),
    .X(_1262_));
 sg13g2_nand3_1 _3238_ (.B(_1236_),
    .C(_1262_),
    .A(_0846_),
    .Y(_1263_));
 sg13g2_nand4_1 _3239_ (.B(net43),
    .C(_1112_),
    .A(_0526_),
    .Y(_1264_),
    .D(_1233_));
 sg13g2_nor4_1 _3240_ (.A(_1202_),
    .B(_1204_),
    .C(_1207_),
    .D(_1264_),
    .Y(_1265_));
 sg13g2_o21ai_1 _3241_ (.B1(_1265_),
    .Y(_1266_),
    .A1(_0334_),
    .A2(_1199_));
 sg13g2_nand4_1 _3242_ (.B(_0526_),
    .C(net43),
    .A(_0350_),
    .Y(_1267_),
    .D(_1112_));
 sg13g2_nor4_1 _3243_ (.A(_1202_),
    .B(_1204_),
    .C(_1207_),
    .D(_1267_),
    .Y(_1268_));
 sg13g2_o21ai_1 _3244_ (.B1(_1268_),
    .Y(_1269_),
    .A1(_0334_),
    .A2(_1199_));
 sg13g2_a21oi_1 _3245_ (.A1(_0526_),
    .A2(net43),
    .Y(_1270_),
    .B1(_0350_));
 sg13g2_nand3_1 _3246_ (.B(_1236_),
    .C(_1270_),
    .A(_0846_),
    .Y(_1271_));
 sg13g2_nand4_1 _3247_ (.B(_1266_),
    .C(_1269_),
    .A(_1263_),
    .Y(_1272_),
    .D(_1271_));
 sg13g2_o21ai_1 _3248_ (.B1(_1209_),
    .Y(_1273_),
    .A1(_1262_),
    .A2(_1270_));
 sg13g2_nor4_1 _3249_ (.A(_0349_),
    .B(_0527_),
    .C(_1119_),
    .D(_1261_),
    .Y(_1274_));
 sg13g2_a221oi_1 _3250_ (.B2(_1270_),
    .C1(_1274_),
    .B1(_1261_),
    .A1(_0527_),
    .Y(_1275_),
    .A2(_1119_));
 sg13g2_nand2_1 _3251_ (.Y(_1276_),
    .A(_1273_),
    .B(_1275_));
 sg13g2_nor3_2 _3252_ (.A(net59),
    .B(_1272_),
    .C(_1276_),
    .Y(_1277_));
 sg13g2_xnor2_1 _3253_ (.Y(_1278_),
    .A(_1259_),
    .B(_1277_));
 sg13g2_xnor2_1 _3254_ (.Y(_1279_),
    .A(_1258_),
    .B(_1278_));
 sg13g2_nand2_1 _3255_ (.Y(_1280_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[7].fa.HA1.a ),
    .B(net49));
 sg13g2_o21ai_1 _3256_ (.B1(_1280_),
    .Y(_0280_),
    .A1(_0627_),
    .A2(_1279_));
 sg13g2_nand2_1 _3257_ (.Y(_1281_),
    .A(_0937_),
    .B(_1242_));
 sg13g2_a21oi_1 _3258_ (.A1(_1245_),
    .A2(_1246_),
    .Y(_1282_),
    .B1(_1250_));
 sg13g2_nand2_1 _3259_ (.Y(_1283_),
    .A(_1281_),
    .B(_1282_));
 sg13g2_a221oi_1 _3260_ (.B2(_0520_),
    .C1(_1277_),
    .B1(_1283_),
    .A1(_1228_),
    .Y(_1284_),
    .A2(_1230_));
 sg13g2_nand2_1 _3261_ (.Y(_1285_),
    .A(_1259_),
    .B(_1252_));
 sg13g2_a21oi_1 _3262_ (.A1(_1228_),
    .A2(_1230_),
    .Y(_1286_),
    .B1(_1285_));
 sg13g2_nor2b_1 _3263_ (.A(_1277_),
    .B_N(_1259_),
    .Y(_1287_));
 sg13g2_nand3b_1 _3264_ (.B(_1252_),
    .C(_0519_),
    .Y(_1288_),
    .A_N(_1277_));
 sg13g2_nand3_1 _3265_ (.B(_1259_),
    .C(_1252_),
    .A(_0519_),
    .Y(_1289_));
 sg13g2_nand3b_1 _3266_ (.B(_1288_),
    .C(_1289_),
    .Y(_1290_),
    .A_N(_1287_));
 sg13g2_nand2_1 _3267_ (.Y(_1291_),
    .A(_0519_),
    .B(_1259_));
 sg13g2_a21oi_1 _3268_ (.A1(_1228_),
    .A2(_1230_),
    .Y(_1292_),
    .B1(_1291_));
 sg13g2_nor4_1 _3269_ (.A(_1284_),
    .B(_1286_),
    .C(_1290_),
    .D(_1292_),
    .Y(_1293_));
 sg13g2_a21o_1 _3270_ (.A2(_1261_),
    .A1(_1247_),
    .B1(_0349_),
    .X(_1294_));
 sg13g2_nand2_1 _3271_ (.Y(_1295_),
    .A(_0526_),
    .B(_1112_));
 sg13g2_a21oi_1 _3272_ (.A1(_1244_),
    .A2(_1294_),
    .Y(_1296_),
    .B1(_1295_));
 sg13g2_xnor2_1 _3273_ (.Y(_1297_),
    .A(_0532_),
    .B(_1296_));
 sg13g2_nand3b_1 _3274_ (.B(net60),
    .C(_0492_),
    .Y(_1298_),
    .A_N(_1297_));
 sg13g2_xor2_1 _3275_ (.B(_1298_),
    .A(_1293_),
    .X(_1299_));
 sg13g2_nand2_1 _3276_ (.Y(_1300_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[8].fa.HA1.a ),
    .B(net49));
 sg13g2_o21ai_1 _3277_ (.B1(_1300_),
    .Y(_0281_),
    .A1(_0627_),
    .A2(_1299_));
 sg13g2_nand2_1 _3278_ (.Y(_0118_),
    .A(_1308_),
    .B(\rsa_en_logic_i.state[0] ));
 sg13g2_nand2_1 _3279_ (.Y(_1301_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ),
    .B(_1325_));
 sg13g2_o21ai_1 _3280_ (.B1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ),
    .Y(_1302_),
    .A1(_1319_),
    .A2(_1355_));
 sg13g2_nand2_1 _3281_ (.Y(_1303_),
    .A(_1301_),
    .B(_1302_));
 sg13g2_nor2b_1 _3282_ (.A(_1355_),
    .B_N(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ),
    .Y(_1304_));
 sg13g2_nand3_1 _3283_ (.B(_1314_),
    .C(_1304_),
    .A(_1318_),
    .Y(_1305_));
 sg13g2_a21oi_1 _3284_ (.A1(_1359_),
    .A2(_1305_),
    .Y(_1306_),
    .B1(_1317_));
 sg13g2_a221oi_1 _3285_ (.B2(net86),
    .C1(_1306_),
    .B1(_1303_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0] ),
    .Y(_0119_),
    .A2(_1360_));
 sg13g2_dfrbp_1 _3286_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(_0120_),
    .Q_N(\rsa_unit_i.rsa_control_fsm.state[0] ),
    .Q(_0117_));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _3289__156 (.L_HI(net156));
 sg13g2_buf_1 _3289_ (.A(net156),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3290_ (.A(net157),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3291_ (.A(net158),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3292_ (.A(net159),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3293_ (.A(net160),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3294_ (.A(net161),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3295_ (.A(net162),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3296_ (.A(net163),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3297_ (.A(\rsa_spi_wrapper_i.config_regs[56] ),
    .X(net7));
 sg13g2_buf_1 _3298_ (.A(\rsa_spi_wrapper_i.config_regs[57] ),
    .X(net8));
 sg13g2_buf_1 _3299_ (.A(\rsa_spi_wrapper_i.config_regs[58] ),
    .X(net9));
 sg13g2_buf_1 _3300_ (.A(\rsa_spi_wrapper_i.config_regs[59] ),
    .X(net10));
 sg13g2_buf_1 _3301_ (.A(\rsa_spi_wrapper_i.config_regs[60] ),
    .X(net11));
 sg13g2_buf_1 _3302_ (.A(\rsa_spi_wrapper_i.config_regs[61] ),
    .X(net12));
 sg13g2_buf_1 _3303_ (.A(\rsa_spi_wrapper_i.config_regs[62] ),
    .X(net13));
 sg13g2_buf_1 _3304_ (.A(\rsa_spi_wrapper_i.config_regs[63] ),
    .X(net14));
 sg13g2_buf_1 _3305_ (.A(net150),
    .X(uo_out[0]));
 sg13g2_buf_1 _3306_ (.A(net151),
    .X(uo_out[1]));
 sg13g2_buf_1 _3307_ (.A(net152),
    .X(uo_out[2]));
 sg13g2_buf_1 _3308_ (.A(\rsa_spi_wrapper_i.spi_miso ),
    .X(net15));
 sg13g2_buf_1 _3309_ (.A(irq),
    .X(net16));
 sg13g2_buf_1 _3310_ (.A(net153),
    .X(uo_out[5]));
 sg13g2_buf_1 _3311_ (.A(net154),
    .X(uo_out[6]));
 sg13g2_buf_1 _3312_ (.A(net155),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \gpio_wrapper_i.gpio_start_cmd_i.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net142),
    .D(_0121_),
    .Q_N(_1736_),
    .Q(\gpio_wrapper_i.gpio_start_cmd_i.data_dly ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.gpio_stop_cmd_i.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0122_),
    .Q_N(_1735_),
    .Q(\gpio_wrapper_i.gpio_stop_cmd_i.data_dly ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.sync_gpio_start.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0123_),
    .Q_N(_1734_),
    .Q(\gpio_wrapper_i.sync_gpio_start.data_sync[1] ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.sync_gpio_start.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0124_),
    .Q_N(_1733_),
    .Q(\gpio_wrapper_i.gpio_start_cmd_i.data ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.sync_gpio_stop.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net145),
    .D(_0125_),
    .Q_N(_1732_),
    .Q(\gpio_wrapper_i.sync_gpio_stop.data_sync[1] ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.sync_gpio_stop.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0126_),
    .Q_N(_1731_),
    .Q(\gpio_wrapper_i.gpio_stop_cmd_i.data ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.irq_reg$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net147),
    .D(_0127_),
    .Q_N(_0058_),
    .Q(irq));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[0]$_DFF_PN1_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net136),
    .D(_0118_),
    .Q_N(\rsa_en_logic_i.state[0] ),
    .Q(_1752_));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net142),
    .D(_0000_),
    .Q_N(_1737_),
    .Q(\rsa_en_logic_i.state[1] ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[2]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(_0001_),
    .Q_N(_1738_),
    .Q(\rsa_en_logic_i.state[2] ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[3]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net147),
    .D(_0002_),
    .Q_N(_1739_),
    .Q(\rsa_en_logic_i.state[3] ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[4]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net144),
    .D(_0003_),
    .Q_N(_1740_),
    .Q(\rsa_en_logic_i.state[4] ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[5]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(_0004_),
    .Q_N(_0053_),
    .Q(\rsa_en_logic_i.state[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_start_cmd_i.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net142),
    .D(_0128_),
    .Q_N(_1730_),
    .Q(\rsa_spi_wrapper_i.spi_start_cmd_i.data_dly ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net143),
    .D(_0129_),
    .Q_N(_1729_),
    .Q(\rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net128),
    .D(_0130_),
    .Q_N(_0056_),
    .Q(\rsa_spi_wrapper_i.config_regs[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net139),
    .D(_0131_),
    .Q_N(_0060_),
    .Q(\rsa_spi_wrapper_i.config_regs[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net128),
    .D(_0132_),
    .Q_N(_0063_),
    .Q(\rsa_spi_wrapper_i.config_regs[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0133_),
    .Q_N(_0066_),
    .Q(\rsa_spi_wrapper_i.config_regs[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net127),
    .D(_0134_),
    .Q_N(_0069_),
    .Q(\rsa_spi_wrapper_i.config_regs[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net128),
    .D(_0135_),
    .Q_N(_0072_),
    .Q(\rsa_spi_wrapper_i.config_regs[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0136_),
    .Q_N(_0075_),
    .Q(\rsa_spi_wrapper_i.config_regs[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net124),
    .D(_0137_),
    .Q_N(_0078_),
    .Q(\rsa_spi_wrapper_i.config_regs[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net136),
    .D(_0138_),
    .Q_N(_1728_),
    .Q(\rsa_spi_wrapper_i.config_regs[8] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net136),
    .D(_0139_),
    .Q_N(_1727_),
    .Q(\rsa_spi_wrapper_i.config_regs[9] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net120),
    .D(_0140_),
    .Q_N(_1726_),
    .Q(\rsa_spi_wrapper_i.config_regs[10] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net124),
    .D(_0141_),
    .Q_N(_1725_),
    .Q(\rsa_spi_wrapper_i.config_regs[11] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net120),
    .D(_0142_),
    .Q_N(_1724_),
    .Q(\rsa_spi_wrapper_i.config_regs[12] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net124),
    .D(_0143_),
    .Q_N(_1723_),
    .Q(\rsa_spi_wrapper_i.config_regs[13] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net124),
    .D(_0144_),
    .Q_N(_1722_),
    .Q(\rsa_spi_wrapper_i.config_regs[14] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net121),
    .D(_0145_),
    .Q_N(_1721_),
    .Q(\rsa_spi_wrapper_i.config_regs[15] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net136),
    .D(_0146_),
    .Q_N(_0105_),
    .Q(\rsa_p[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net136),
    .D(_0147_),
    .Q_N(_1720_),
    .Q(\rsa_p[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net136),
    .D(_0148_),
    .Q_N(_0108_),
    .Q(\rsa_p[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net137),
    .D(_0149_),
    .Q_N(_0110_),
    .Q(\rsa_p[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net138),
    .D(_0150_),
    .Q_N(_0112_),
    .Q(\rsa_p[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net137),
    .D(_0151_),
    .Q_N(_0114_),
    .Q(\rsa_p[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net137),
    .D(_0152_),
    .Q_N(_0116_),
    .Q(\rsa_p[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net137),
    .D(_0153_),
    .Q_N(_0021_),
    .Q(\rsa_p[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net119),
    .D(_0154_),
    .Q_N(_1719_),
    .Q(\rsa_e[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net124),
    .D(_0155_),
    .Q_N(_1718_),
    .Q(\rsa_e[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net124),
    .D(_0156_),
    .Q_N(_1717_),
    .Q(\rsa_e[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net122),
    .D(_0157_),
    .Q_N(_1716_),
    .Q(\rsa_e[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net122),
    .D(_0158_),
    .Q_N(_1715_),
    .Q(\rsa_e[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net122),
    .D(_0159_),
    .Q_N(_1714_),
    .Q(\rsa_e[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net122),
    .D(_0160_),
    .Q_N(_1713_),
    .Q(\rsa_e[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net119),
    .D(_0161_),
    .Q_N(_1712_),
    .Q(\rsa_e[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net132),
    .D(_0162_),
    .Q_N(_0057_),
    .Q(\rsa_spi_wrapper_i.config_regs[32] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net133),
    .D(_0163_),
    .Q_N(_0061_),
    .Q(\rsa_spi_wrapper_i.config_regs[33] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net126),
    .D(_0164_),
    .Q_N(_0064_),
    .Q(\rsa_spi_wrapper_i.config_regs[34] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net117),
    .D(_0165_),
    .Q_N(_0067_),
    .Q(\rsa_spi_wrapper_i.config_regs[35] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net126),
    .D(_0166_),
    .Q_N(_0070_),
    .Q(\rsa_spi_wrapper_i.config_regs[36] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net118),
    .D(_0167_),
    .Q_N(_0073_),
    .Q(\rsa_spi_wrapper_i.config_regs[37] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net118),
    .D(_0168_),
    .Q_N(_0076_),
    .Q(\rsa_spi_wrapper_i.config_regs[38] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net126),
    .D(_0169_),
    .Q_N(_0079_),
    .Q(\rsa_spi_wrapper_i.config_regs[39] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net132),
    .D(_0170_),
    .Q_N(_0082_),
    .Q(\rsa_const[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net132),
    .D(_0171_),
    .Q_N(_0085_),
    .Q(\rsa_const[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net126),
    .D(_0172_),
    .Q_N(_0088_),
    .Q(\rsa_const[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net118),
    .D(_0173_),
    .Q_N(_0091_),
    .Q(\rsa_const[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net137),
    .D(_0174_),
    .Q_N(_0094_),
    .Q(\rsa_const[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net118),
    .D(_0175_),
    .Q_N(_0097_),
    .Q(\rsa_const[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net132),
    .D(_0176_),
    .Q_N(_0100_),
    .Q(\rsa_const[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net137),
    .D(_0177_),
    .Q_N(_0103_),
    .Q(\rsa_const[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net121),
    .D(_0178_),
    .Q_N(_1711_),
    .Q(\rsa_spi_wrapper_i.config_regs[48] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net137),
    .D(_0179_),
    .Q_N(_1710_),
    .Q(\rsa_spi_wrapper_i.config_regs[49] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net126),
    .D(_0180_),
    .Q_N(_1709_),
    .Q(\rsa_spi_wrapper_i.config_regs[50] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net121),
    .D(_0181_),
    .Q_N(_1708_),
    .Q(\rsa_spi_wrapper_i.config_regs[51] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net126),
    .D(_0182_),
    .Q_N(_1707_),
    .Q(\rsa_spi_wrapper_i.config_regs[52] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net129),
    .D(_0183_),
    .Q_N(_1706_),
    .Q(\rsa_spi_wrapper_i.config_regs[53] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net126),
    .D(_0184_),
    .Q_N(_1705_),
    .Q(\rsa_spi_wrapper_i.config_regs[54] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net120),
    .D(_0185_),
    .Q_N(_1704_),
    .Q(\rsa_spi_wrapper_i.config_regs[55] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net128),
    .D(_0186_),
    .Q_N(_1703_),
    .Q(\rsa_spi_wrapper_i.config_regs[56] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net128),
    .D(_0187_),
    .Q_N(_1702_),
    .Q(\rsa_spi_wrapper_i.config_regs[57] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0188_),
    .Q_N(_1701_),
    .Q(\rsa_spi_wrapper_i.config_regs[58] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net127),
    .D(_0189_),
    .Q_N(_1700_),
    .Q(\rsa_spi_wrapper_i.config_regs[59] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net127),
    .D(_0190_),
    .Q_N(_1699_),
    .Q(\rsa_spi_wrapper_i.config_regs[60] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net127),
    .D(_0191_),
    .Q_N(_1698_),
    .Q(\rsa_spi_wrapper_i.config_regs[61] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0192_),
    .Q_N(_1697_),
    .Q(\rsa_spi_wrapper_i.config_regs[62] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net128),
    .D(_0193_),
    .Q_N(_1696_),
    .Q(\rsa_spi_wrapper_i.config_regs[63] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.addr[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net129),
    .D(_0194_),
    .Q_N(_1695_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.addr[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net139),
    .D(_0195_),
    .Q_N(_1694_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.addr[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net139),
    .D(_0196_),
    .Q_N(_0050_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.addr[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net128),
    .D(_0197_),
    .Q_N(_1693_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net139),
    .D(_0198_),
    .Q_N(_1692_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net139),
    .D(_0199_),
    .Q_N(_1691_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net124),
    .D(_0200_),
    .Q_N(_1690_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net123),
    .D(_0201_),
    .Q_N(_1689_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net123),
    .D(_0202_),
    .Q_N(_1688_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net123),
    .D(_0203_),
    .Q_N(_1687_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net123),
    .D(_0204_),
    .Q_N(_1686_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net124),
    .D(_0205_),
    .Q_N(_1685_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.dv$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net140),
    .D(_0206_),
    .Q_N(_1684_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o_vld ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net140),
    .D(_0207_),
    .Q_N(_1683_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rising_edge_detector_eof.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0208_),
    .Q_N(_1682_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rising_edge_detector_spi_clk.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net145),
    .D(_0209_),
    .Q_N(_1681_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net140),
    .D(_0210_),
    .Q_N(_1680_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net129),
    .D(_0211_),
    .Q_N(_1679_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net129),
    .D(_0212_),
    .Q_N(_1678_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net125),
    .D(_0213_),
    .Q_N(_1677_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net123),
    .D(_0214_),
    .Q_N(_1676_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net123),
    .D(_0215_),
    .Q_N(_1675_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net123),
    .D(_0216_),
    .Q_N(_1674_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net125),
    .D(_0217_),
    .Q_N(_1673_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net147),
    .D(_0218_),
    .Q_N(_1672_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net147),
    .D(_0219_),
    .Q_N(_1671_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net147),
    .D(_0220_),
    .Q_N(_1670_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net145),
    .D(_0221_),
    .Q_N(_1669_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0]$_DFF_PN1_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net147),
    .D(_0119_),
    .Q_N(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0] ),
    .Q(_1753_));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net140),
    .D(_0005_),
    .Q_N(_1741_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net147),
    .D(_0006_),
    .Q_N(_1742_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3]$_DFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net145),
    .D(_0007_),
    .Q_N(_1743_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4]$_DFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net140),
    .D(_0008_),
    .Q_N(_1668_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net140),
    .D(_0222_),
    .Q_N(_0059_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net140),
    .D(_0223_),
    .Q_N(_0062_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net138),
    .D(_0224_),
    .Q_N(_0065_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net138),
    .D(_0225_),
    .Q_N(_0068_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net137),
    .D(_0226_),
    .Q_N(_0071_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net139),
    .D(_0227_),
    .Q_N(_0074_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net139),
    .D(_0228_),
    .Q_N(_0077_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net139),
    .D(_0229_),
    .Q_N(_1667_),
    .Q(\rsa_spi_wrapper_i.spi_miso ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net141),
    .D(_0230_),
    .Q_N(_1666_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net141),
    .D(_0231_),
    .Q_N(_1665_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net147),
    .D(_0232_),
    .Q_N(_1664_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net141),
    .D(_0233_),
    .Q_N(_1663_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net115),
    .D(_0234_),
    .Q_N(_1662_),
    .Q(\rsa_unit_i.mmm_multiply.A_bit ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net113),
    .D(_0235_),
    .Q_N(_0023_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net113),
    .D(_0236_),
    .Q_N(_0024_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(_0237_),
    .Q_N(_0026_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(_0238_),
    .Q_N(_0028_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(_0239_),
    .Q_N(_0030_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net113),
    .D(_0240_),
    .Q_N(_0032_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net113),
    .D(_0241_),
    .Q_N(_0034_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net113),
    .D(_0242_),
    .Q_N(_0036_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net112),
    .D(_0243_),
    .Q_N(_0038_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[9] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net112),
    .D(_0244_),
    .Q_N(_0042_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.fa_bit0.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net115),
    .D(_0245_),
    .Q_N(_0041_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[1].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net113),
    .D(_0246_),
    .Q_N(_0043_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[2].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net112),
    .D(_0247_),
    .Q_N(_0044_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[3].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net112),
    .D(_0248_),
    .Q_N(_0045_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[4].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net112),
    .D(_0249_),
    .Q_N(_0046_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[5].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net112),
    .D(_0250_),
    .Q_N(_0047_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[6].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net112),
    .D(_0251_),
    .Q_N(_0048_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[7].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net112),
    .D(_0252_),
    .Q_N(_0049_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[8].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net120),
    .D(_0253_),
    .Q_N(_1661_),
    .Q(\rsa_unit_i.R_i[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net115),
    .D(_0254_),
    .Q_N(_0025_),
    .Q(\rsa_unit_i.R_i[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net119),
    .D(_0255_),
    .Q_N(_0027_),
    .Q(\rsa_unit_i.R_i[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net119),
    .D(_0256_),
    .Q_N(_0029_),
    .Q(\rsa_unit_i.R_i[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net120),
    .D(_0257_),
    .Q_N(_0031_),
    .Q(\rsa_unit_i.R_i[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(_0258_),
    .Q_N(_0033_),
    .Q(\rsa_unit_i.R_i[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net113),
    .D(_0259_),
    .Q_N(_0035_),
    .Q(\rsa_unit_i.R_i[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net113),
    .D(_0260_),
    .Q_N(_0037_),
    .Q(\rsa_unit_i.R_i[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net116),
    .D(_0261_),
    .Q_N(_0039_),
    .Q(\rsa_unit_i.R_i[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net116),
    .D(_0262_),
    .Q_N(_0040_),
    .Q(\rsa_unit_i.R_i[9] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net131),
    .D(_0263_),
    .Q_N(_1660_),
    .Q(\rsa_unit_i.mmm_square.A_bit ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net131),
    .D(_0264_),
    .Q_N(_0080_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net131),
    .D(_0265_),
    .Q_N(_0083_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net117),
    .D(_0266_),
    .Q_N(_0086_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net117),
    .D(_0267_),
    .Q_N(_0089_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net117),
    .D(_0268_),
    .Q_N(_0092_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net117),
    .D(_0269_),
    .Q_N(_0095_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0270_),
    .Q_N(_0098_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net117),
    .D(_0271_),
    .Q_N(_0101_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net117),
    .D(_0272_),
    .Q_N(_1659_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[9] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net132),
    .D(_0273_),
    .Q_N(_0106_),
    .Q(\rsa_unit_i.mmm_square.adder2.fa_bit0.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0274_),
    .Q_N(_0104_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[1].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0275_),
    .Q_N(_0107_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[2].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net135),
    .D(_0276_),
    .Q_N(_0109_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[3].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net135),
    .D(_0277_),
    .Q_N(_0111_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[4].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net135),
    .D(_0278_),
    .Q_N(_0113_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[5].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net135),
    .D(_0279_),
    .Q_N(_0115_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[6].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net135),
    .D(_0280_),
    .Q_N(_0020_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[7].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net135),
    .D(_0281_),
    .Q_N(_0022_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[8].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net132),
    .D(_0282_),
    .Q_N(_0081_),
    .Q(\rsa_unit_i.P_i[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net132),
    .D(_0283_),
    .Q_N(_0084_),
    .Q(\rsa_unit_i.P_i[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net132),
    .D(_0284_),
    .Q_N(_0087_),
    .Q(\rsa_unit_i.P_i[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net118),
    .D(_0285_),
    .Q_N(_0090_),
    .Q(\rsa_unit_i.P_i[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net131),
    .D(_0286_),
    .Q_N(_0093_),
    .Q(\rsa_unit_i.P_i[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net117),
    .D(_0287_),
    .Q_N(_0096_),
    .Q(\rsa_unit_i.P_i[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0288_),
    .Q_N(_0099_),
    .Q(\rsa_unit_i.P_i[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0289_),
    .Q_N(_0102_),
    .Q(\rsa_unit_i.P_i[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0290_),
    .Q_N(_1658_),
    .Q(\rsa_unit_i.P_i[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net133),
    .D(_0291_),
    .Q_N(_1657_),
    .Q(\rsa_unit_i.P_i[9] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net129),
    .D(_0292_),
    .Q_N(_1656_),
    .Q(\rsa_c[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net126),
    .D(_0293_),
    .Q_N(_1655_),
    .Q(\rsa_c[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net119),
    .D(_0294_),
    .Q_N(_1654_),
    .Q(\rsa_c[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net119),
    .D(_0295_),
    .Q_N(_1653_),
    .Q(\rsa_c[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net120),
    .D(_0296_),
    .Q_N(_1652_),
    .Q(\rsa_c[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net120),
    .D(_0297_),
    .Q_N(_1651_),
    .Q(\rsa_c[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net119),
    .D(_0298_),
    .Q_N(_1650_),
    .Q(\rsa_c[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net120),
    .D(_0299_),
    .Q_N(_1649_),
    .Q(\rsa_c[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_rounds[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net143),
    .D(_0300_),
    .Q_N(_1648_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_rounds[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_rounds[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net143),
    .D(_0301_),
    .Q_N(_1647_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_rounds[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_rounds[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net142),
    .D(_0302_),
    .Q_N(_1646_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_rounds[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net143),
    .D(_0303_),
    .Q_N(_1645_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_steps[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0304_),
    .Q_N(_1644_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_steps[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_steps[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0305_),
    .Q_N(_1643_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_steps[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_steps[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0306_),
    .Q_N(_1642_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_steps[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0307_),
    .Q_N(_1641_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net119),
    .D(_0308_),
    .Q_N(_1640_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net121),
    .D(_0309_),
    .Q_N(_1639_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net121),
    .D(_0310_),
    .Q_N(_1638_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net122),
    .D(_0311_),
    .Q_N(_1637_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net122),
    .D(_0312_),
    .Q_N(_1636_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net122),
    .D(_0313_),
    .Q_N(_1635_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net122),
    .D(_0314_),
    .Q_N(_1634_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net121),
    .D(_0315_),
    .Q_N(_1744_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[10]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net136),
    .D(_0009_),
    .Q_N(_1745_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[10] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[11]$_DFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net136),
    .D(_0010_),
    .Q_N(_0052_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[11] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net134),
    .D(_0011_),
    .Q_N(_1746_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[2]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net142),
    .D(_0012_),
    .Q_N(_1747_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[3]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net142),
    .D(_0013_),
    .Q_N(_1748_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[4]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(_0014_),
    .Q_N(_0055_),
    .Q(eoc_rsa));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[5]$_DFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0015_),
    .Q_N(_1749_),
    .Q(\rsa_unit_i.rsa_control_fsm.increment_rounds ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[6]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net144),
    .D(_0016_),
    .Q_N(_1750_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[7]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net142),
    .D(_0017_),
    .Q_N(_1751_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[8]$_DFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net135),
    .D(_0018_),
    .Q_N(_0054_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[9]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net142),
    .D(_0019_),
    .Q_N(_0051_),
    .Q(\rsa_unit_i.rsa_control_fsm.load_exp ));
 sg13g2_dfrbp_1 \synchronizer_spi_clk_inst.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net145),
    .D(_0316_),
    .Q_N(_1633_),
    .Q(\synchronizer_spi_clk_inst.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_clk_inst.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0317_),
    .Q_N(_1632_),
    .Q(\rsa_spi_wrapper_i.spi_clk ));
 sg13g2_dfrbp_1 \synchronizer_spi_cs_n_inst.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net145),
    .D(_0318_),
    .Q_N(_1631_),
    .Q(\synchronizer_spi_cs_n_inst.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_cs_n_inst.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net145),
    .D(_0319_),
    .Q_N(_1630_),
    .Q(\rsa_spi_wrapper_i.spi_cs_n ));
 sg13g2_dfrbp_1 \synchronizer_spi_mosi_inst.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net145),
    .D(_0320_),
    .Q_N(_1629_),
    .Q(\synchronizer_spi_mosi_inst.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_mosi_inst.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net146),
    .D(_0321_),
    .Q_N(_1628_),
    .Q(\rsa_spi_wrapper_i.spi_mosi ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[1]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[2]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[3]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[4]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[5]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[6]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[7]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[4]));
 sg13g2_buf_2 fanout17 (.A(_0390_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_1129_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0628_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0597_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0481_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0425_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0389_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1127_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0596_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0568_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1115_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1089_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0414_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0729_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0419_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0384_),
    .X(net32));
 sg13g2_buf_4 fanout33 (.X(net33),
    .A(_1483_));
 sg13g2_buf_2 fanout34 (.A(_1464_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0492_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0475_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0407_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0401_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0383_),
    .X(net39));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(_1372_));
 sg13g2_buf_2 fanout41 (.A(_0942_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0622_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0491_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0417_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1533_),
    .X(net45));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(_1488_));
 sg13g2_buf_2 fanout47 (.A(_1453_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1401_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1390_),
    .X(net49));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(_0618_));
 sg13g2_buf_2 fanout51 (.A(_0601_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0416_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0405_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0379_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1479_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1445_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1375_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1342_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0994_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0937_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0472_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0398_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0395_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0381_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1470_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1462_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1444_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1431_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1400_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0965_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0936_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0846_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0743_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0701_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0630_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0604_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0569_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0393_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1525_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1481_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1447_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1430_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1427_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1425_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1417_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1364_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1315_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0980_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0665_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0629_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0603_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0487_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0375_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0349_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0333_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_1624_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1585_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1466_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_1454_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1443_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_1442_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_1441_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_1440_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_1439_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_1438_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_1437_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_1423_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1374_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1370_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1314_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_1307_),
    .X(net111));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(net116));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(net115));
 sg13g2_buf_2 fanout114 (.A(net115),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(net116),
    .X(net115));
 sg13g2_buf_1 fanout116 (.A(net130),
    .X(net116));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(net130));
 sg13g2_buf_2 fanout118 (.A(net130),
    .X(net118));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(net121));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(net121));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(net130));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(net125));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(net125));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(net125));
 sg13g2_buf_2 fanout125 (.A(net130),
    .X(net125));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(net129));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(net128));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(net129));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(net130));
 sg13g2_buf_2 fanout130 (.A(net149),
    .X(net130));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(net133));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(net133));
 sg13g2_buf_2 fanout133 (.A(net149),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net135));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net149));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(net138));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net141));
 sg13g2_buf_2 fanout138 (.A(net141),
    .X(net138));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net140));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(net141));
 sg13g2_buf_2 fanout141 (.A(net148),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net144));
 sg13g2_buf_2 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net148));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net146));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net148));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(net148));
 sg13g2_buf_1 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_1 fanout149 (.A(net1),
    .X(net149));
 sg13g2_tielo _3305__150 (.L_LO(net150));
 sg13g2_tielo _3306__151 (.L_LO(net151));
 sg13g2_tielo _3307__152 (.L_LO(net152));
 sg13g2_tielo _3310__153 (.L_LO(net153));
 sg13g2_tielo _3311__154 (.L_LO(net154));
 sg13g2_tielo _3312__155 (.L_LO(net155));
 sg13g2_tiehi _3290__157 (.L_HI(net157));
 sg13g2_tiehi _3291__158 (.L_HI(net158));
 sg13g2_tiehi _3292__159 (.L_HI(net159));
 sg13g2_tiehi _3293__160 (.L_HI(net160));
 sg13g2_tiehi _3294__161 (.L_HI(net161));
 sg13g2_tiehi _3295__162 (.L_HI(net162));
 sg13g2_tiehi _3296__163 (.L_HI(net163));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload2 (.A(clknet_leaf_29_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_leaf_2_clk));
 sg13g2_buf_16 clkload4 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_12_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_25_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_24_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_fill_1 FILLER_0_21 ();
 sg13g2_fill_2 FILLER_0_86 ();
 sg13g2_fill_1 FILLER_0_88 ();
 sg13g2_fill_2 FILLER_0_115 ();
 sg13g2_fill_1 FILLER_0_117 ();
 sg13g2_fill_2 FILLER_0_156 ();
 sg13g2_fill_2 FILLER_0_308 ();
 sg13g2_fill_1 FILLER_0_318 ();
 sg13g2_fill_1 FILLER_0_328 ();
 sg13g2_fill_1 FILLER_0_379 ();
 sg13g2_fill_2 FILLER_0_396 ();
 sg13g2_fill_1 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_4 FILLER_1_7 ();
 sg13g2_fill_1 FILLER_1_11 ();
 sg13g2_fill_1 FILLER_1_56 ();
 sg13g2_fill_2 FILLER_1_83 ();
 sg13g2_fill_2 FILLER_1_101 ();
 sg13g2_fill_2 FILLER_1_232 ();
 sg13g2_fill_2 FILLER_1_239 ();
 sg13g2_fill_1 FILLER_1_241 ();
 sg13g2_fill_1 FILLER_1_260 ();
 sg13g2_fill_2 FILLER_1_271 ();
 sg13g2_fill_1 FILLER_1_285 ();
 sg13g2_fill_1 FILLER_1_330 ();
 sg13g2_fill_1 FILLER_1_336 ();
 sg13g2_fill_1 FILLER_1_356 ();
 sg13g2_fill_2 FILLER_1_361 ();
 sg13g2_fill_2 FILLER_1_375 ();
 sg13g2_fill_1 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_fill_1 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_108 ();
 sg13g2_fill_1 FILLER_2_115 ();
 sg13g2_fill_1 FILLER_2_121 ();
 sg13g2_fill_1 FILLER_2_127 ();
 sg13g2_fill_2 FILLER_2_160 ();
 sg13g2_fill_1 FILLER_2_162 ();
 sg13g2_decap_4 FILLER_2_223 ();
 sg13g2_fill_2 FILLER_2_267 ();
 sg13g2_fill_2 FILLER_2_275 ();
 sg13g2_fill_2 FILLER_2_284 ();
 sg13g2_fill_1 FILLER_2_300 ();
 sg13g2_fill_2 FILLER_2_384 ();
 sg13g2_fill_2 FILLER_2_391 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_27 ();
 sg13g2_fill_2 FILLER_3_36 ();
 sg13g2_fill_1 FILLER_3_51 ();
 sg13g2_fill_1 FILLER_3_101 ();
 sg13g2_fill_2 FILLER_3_157 ();
 sg13g2_fill_1 FILLER_3_177 ();
 sg13g2_fill_2 FILLER_3_224 ();
 sg13g2_fill_2 FILLER_3_230 ();
 sg13g2_fill_2 FILLER_3_259 ();
 sg13g2_fill_1 FILLER_3_266 ();
 sg13g2_fill_1 FILLER_3_272 ();
 sg13g2_fill_1 FILLER_3_277 ();
 sg13g2_fill_1 FILLER_3_283 ();
 sg13g2_fill_2 FILLER_3_289 ();
 sg13g2_fill_1 FILLER_3_296 ();
 sg13g2_fill_2 FILLER_3_302 ();
 sg13g2_fill_2 FILLER_3_334 ();
 sg13g2_fill_1 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_fill_2 FILLER_4_64 ();
 sg13g2_fill_1 FILLER_4_93 ();
 sg13g2_fill_1 FILLER_4_117 ();
 sg13g2_fill_1 FILLER_4_123 ();
 sg13g2_fill_1 FILLER_4_133 ();
 sg13g2_fill_1 FILLER_4_138 ();
 sg13g2_fill_1 FILLER_4_165 ();
 sg13g2_fill_1 FILLER_4_205 ();
 sg13g2_decap_4 FILLER_4_211 ();
 sg13g2_fill_2 FILLER_4_215 ();
 sg13g2_fill_1 FILLER_4_221 ();
 sg13g2_fill_1 FILLER_4_226 ();
 sg13g2_fill_1 FILLER_4_265 ();
 sg13g2_fill_2 FILLER_4_273 ();
 sg13g2_fill_1 FILLER_4_275 ();
 sg13g2_fill_1 FILLER_4_280 ();
 sg13g2_fill_1 FILLER_4_286 ();
 sg13g2_fill_1 FILLER_4_295 ();
 sg13g2_fill_1 FILLER_4_336 ();
 sg13g2_fill_1 FILLER_4_342 ();
 sg13g2_fill_1 FILLER_4_353 ();
 sg13g2_fill_1 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_9 ();
 sg13g2_fill_1 FILLER_5_41 ();
 sg13g2_fill_1 FILLER_5_93 ();
 sg13g2_fill_1 FILLER_5_134 ();
 sg13g2_decap_4 FILLER_5_176 ();
 sg13g2_fill_2 FILLER_5_206 ();
 sg13g2_fill_1 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_223 ();
 sg13g2_decap_4 FILLER_5_230 ();
 sg13g2_fill_1 FILLER_5_238 ();
 sg13g2_decap_4 FILLER_5_250 ();
 sg13g2_fill_2 FILLER_5_380 ();
 sg13g2_fill_1 FILLER_5_382 ();
 sg13g2_fill_2 FILLER_5_387 ();
 sg13g2_fill_1 FILLER_5_389 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_fill_2 FILLER_6_94 ();
 sg13g2_fill_1 FILLER_6_154 ();
 sg13g2_fill_1 FILLER_6_162 ();
 sg13g2_fill_1 FILLER_6_172 ();
 sg13g2_decap_4 FILLER_6_178 ();
 sg13g2_fill_1 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_251 ();
 sg13g2_fill_1 FILLER_6_258 ();
 sg13g2_fill_1 FILLER_6_264 ();
 sg13g2_fill_1 FILLER_6_281 ();
 sg13g2_fill_1 FILLER_6_293 ();
 sg13g2_fill_1 FILLER_6_300 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_fill_2 FILLER_6_311 ();
 sg13g2_fill_1 FILLER_6_323 ();
 sg13g2_fill_1 FILLER_6_359 ();
 sg13g2_fill_1 FILLER_6_367 ();
 sg13g2_fill_2 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_6_419 ();
 sg13g2_decap_4 FILLER_6_426 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_31 ();
 sg13g2_fill_2 FILLER_7_89 ();
 sg13g2_fill_1 FILLER_7_127 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_251 ();
 sg13g2_fill_1 FILLER_7_256 ();
 sg13g2_fill_1 FILLER_7_262 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_fill_2 FILLER_7_303 ();
 sg13g2_fill_1 FILLER_7_305 ();
 sg13g2_fill_1 FILLER_7_311 ();
 sg13g2_fill_1 FILLER_7_329 ();
 sg13g2_fill_2 FILLER_7_335 ();
 sg13g2_fill_1 FILLER_7_337 ();
 sg13g2_fill_2 FILLER_7_357 ();
 sg13g2_fill_1 FILLER_7_364 ();
 sg13g2_fill_2 FILLER_7_402 ();
 sg13g2_fill_2 FILLER_8_94 ();
 sg13g2_fill_1 FILLER_8_96 ();
 sg13g2_fill_1 FILLER_8_120 ();
 sg13g2_fill_2 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_138 ();
 sg13g2_fill_2 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_185 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_fill_2 FILLER_8_244 ();
 sg13g2_fill_2 FILLER_8_272 ();
 sg13g2_fill_2 FILLER_8_283 ();
 sg13g2_fill_2 FILLER_8_344 ();
 sg13g2_fill_1 FILLER_8_346 ();
 sg13g2_fill_1 FILLER_8_352 ();
 sg13g2_fill_1 FILLER_8_377 ();
 sg13g2_fill_2 FILLER_8_382 ();
 sg13g2_fill_2 FILLER_8_415 ();
 sg13g2_fill_1 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_426 ();
 sg13g2_fill_1 FILLER_9_62 ();
 sg13g2_fill_1 FILLER_9_68 ();
 sg13g2_fill_1 FILLER_9_108 ();
 sg13g2_fill_2 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_167 ();
 sg13g2_fill_2 FILLER_9_187 ();
 sg13g2_fill_1 FILLER_9_273 ();
 sg13g2_fill_1 FILLER_9_298 ();
 sg13g2_fill_1 FILLER_9_309 ();
 sg13g2_fill_1 FILLER_9_320 ();
 sg13g2_fill_1 FILLER_9_340 ();
 sg13g2_fill_2 FILLER_9_380 ();
 sg13g2_fill_1 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_149 ();
 sg13g2_fill_1 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_170 ();
 sg13g2_fill_2 FILLER_10_228 ();
 sg13g2_fill_2 FILLER_10_284 ();
 sg13g2_fill_2 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_fill_1 FILLER_10_339 ();
 sg13g2_fill_2 FILLER_10_371 ();
 sg13g2_fill_1 FILLER_10_378 ();
 sg13g2_decap_4 FILLER_10_384 ();
 sg13g2_fill_1 FILLER_10_388 ();
 sg13g2_fill_1 FILLER_10_397 ();
 sg13g2_fill_1 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_79 ();
 sg13g2_fill_2 FILLER_11_104 ();
 sg13g2_fill_2 FILLER_11_117 ();
 sg13g2_fill_1 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_135 ();
 sg13g2_fill_1 FILLER_11_137 ();
 sg13g2_fill_2 FILLER_11_176 ();
 sg13g2_decap_4 FILLER_11_197 ();
 sg13g2_fill_2 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_fill_1 FILLER_11_250 ();
 sg13g2_fill_1 FILLER_11_344 ();
 sg13g2_fill_1 FILLER_11_369 ();
 sg13g2_fill_1 FILLER_11_378 ();
 sg13g2_fill_1 FILLER_11_384 ();
 sg13g2_fill_1 FILLER_11_393 ();
 sg13g2_fill_1 FILLER_11_420 ();
 sg13g2_decap_4 FILLER_11_425 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_fill_1 FILLER_12_26 ();
 sg13g2_fill_1 FILLER_12_37 ();
 sg13g2_fill_1 FILLER_12_77 ();
 sg13g2_fill_2 FILLER_12_104 ();
 sg13g2_fill_1 FILLER_12_116 ();
 sg13g2_fill_2 FILLER_12_123 ();
 sg13g2_fill_1 FILLER_12_164 ();
 sg13g2_fill_1 FILLER_12_201 ();
 sg13g2_fill_1 FILLER_12_212 ();
 sg13g2_fill_1 FILLER_12_217 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_fill_1 FILLER_12_234 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_256 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_fill_1 FILLER_12_297 ();
 sg13g2_fill_2 FILLER_12_391 ();
 sg13g2_fill_2 FILLER_12_398 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_27 ();
 sg13g2_fill_2 FILLER_13_39 ();
 sg13g2_fill_2 FILLER_13_67 ();
 sg13g2_fill_1 FILLER_13_69 ();
 sg13g2_fill_2 FILLER_13_96 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_108 ();
 sg13g2_fill_2 FILLER_13_125 ();
 sg13g2_fill_2 FILLER_13_199 ();
 sg13g2_fill_1 FILLER_13_218 ();
 sg13g2_fill_1 FILLER_13_223 ();
 sg13g2_fill_1 FILLER_13_250 ();
 sg13g2_fill_2 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_292 ();
 sg13g2_fill_2 FILLER_13_306 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_fill_1 FILLER_13_357 ();
 sg13g2_decap_4 FILLER_13_381 ();
 sg13g2_fill_2 FILLER_13_390 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_fill_2 FILLER_14_26 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_64 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_fill_2 FILLER_14_85 ();
 sg13g2_fill_1 FILLER_14_87 ();
 sg13g2_fill_1 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_191 ();
 sg13g2_fill_1 FILLER_14_197 ();
 sg13g2_fill_1 FILLER_14_203 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_fill_2 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_378 ();
 sg13g2_fill_2 FILLER_14_384 ();
 sg13g2_fill_1 FILLER_14_386 ();
 sg13g2_fill_2 FILLER_14_396 ();
 sg13g2_fill_1 FILLER_14_398 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_15_26 ();
 sg13g2_fill_1 FILLER_15_47 ();
 sg13g2_fill_1 FILLER_15_74 ();
 sg13g2_fill_1 FILLER_15_85 ();
 sg13g2_fill_1 FILLER_15_90 ();
 sg13g2_fill_2 FILLER_15_97 ();
 sg13g2_fill_2 FILLER_15_108 ();
 sg13g2_fill_1 FILLER_15_144 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_189 ();
 sg13g2_fill_2 FILLER_15_205 ();
 sg13g2_fill_1 FILLER_15_212 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_276 ();
 sg13g2_fill_1 FILLER_15_326 ();
 sg13g2_fill_1 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_342 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_fill_1 FILLER_15_365 ();
 sg13g2_fill_2 FILLER_15_370 ();
 sg13g2_fill_2 FILLER_15_377 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_5 ();
 sg13g2_decap_4 FILLER_16_13 ();
 sg13g2_decap_4 FILLER_16_32 ();
 sg13g2_fill_1 FILLER_16_89 ();
 sg13g2_fill_1 FILLER_16_95 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_142 ();
 sg13g2_decap_8 FILLER_16_194 ();
 sg13g2_decap_8 FILLER_16_201 ();
 sg13g2_fill_2 FILLER_16_208 ();
 sg13g2_fill_2 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_263 ();
 sg13g2_fill_2 FILLER_16_269 ();
 sg13g2_fill_1 FILLER_16_318 ();
 sg13g2_fill_1 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_349 ();
 sg13g2_decap_4 FILLER_16_410 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_2 FILLER_17_128 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_fill_2 FILLER_17_313 ();
 sg13g2_fill_1 FILLER_17_321 ();
 sg13g2_fill_2 FILLER_17_342 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_2 FILLER_17_387 ();
 sg13g2_fill_1 FILLER_17_402 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_27 ();
 sg13g2_fill_1 FILLER_18_38 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_69 ();
 sg13g2_fill_2 FILLER_18_144 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_fill_1 FILLER_18_194 ();
 sg13g2_decap_4 FILLER_18_217 ();
 sg13g2_fill_2 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_fill_1 FILLER_18_347 ();
 sg13g2_fill_1 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_decap_4 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_5 ();
 sg13g2_fill_1 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_fill_1 FILLER_19_105 ();
 sg13g2_decap_4 FILLER_19_111 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_194 ();
 sg13g2_fill_2 FILLER_19_206 ();
 sg13g2_fill_1 FILLER_19_208 ();
 sg13g2_decap_4 FILLER_19_223 ();
 sg13g2_decap_4 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_281 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_fill_2 FILLER_19_292 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_decap_4 FILLER_19_336 ();
 sg13g2_fill_2 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_385 ();
 sg13g2_decap_4 FILLER_19_425 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_33 ();
 sg13g2_fill_1 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_66 ();
 sg13g2_fill_1 FILLER_20_85 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_fill_2 FILLER_20_128 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_decap_4 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_268 ();
 sg13g2_fill_2 FILLER_20_295 ();
 sg13g2_fill_2 FILLER_20_301 ();
 sg13g2_fill_2 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_354 ();
 sg13g2_fill_1 FILLER_20_395 ();
 sg13g2_fill_2 FILLER_20_427 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_fill_1 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_87 ();
 sg13g2_decap_4 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_136 ();
 sg13g2_fill_1 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_202 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_fill_2 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_243 ();
 sg13g2_decap_8 FILLER_21_255 ();
 sg13g2_fill_2 FILLER_21_281 ();
 sg13g2_decap_8 FILLER_21_286 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_fill_2 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_415 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_27 ();
 sg13g2_fill_1 FILLER_22_32 ();
 sg13g2_fill_2 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_fill_2 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_232 ();
 sg13g2_decap_4 FILLER_22_296 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_fill_1 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_fill_1 FILLER_23_80 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_fill_2 FILLER_23_200 ();
 sg13g2_decap_4 FILLER_23_228 ();
 sg13g2_fill_2 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_274 ();
 sg13g2_fill_2 FILLER_23_301 ();
 sg13g2_fill_1 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_409 ();
 sg13g2_fill_1 FILLER_23_416 ();
 sg13g2_fill_2 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_fill_2 FILLER_24_153 ();
 sg13g2_fill_1 FILLER_24_160 ();
 sg13g2_fill_2 FILLER_24_167 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_decap_8 FILLER_24_255 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_fill_2 FILLER_24_292 ();
 sg13g2_decap_4 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_323 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_356 ();
 sg13g2_fill_1 FILLER_24_365 ();
 sg13g2_fill_2 FILLER_25_36 ();
 sg13g2_fill_1 FILLER_25_43 ();
 sg13g2_fill_2 FILLER_25_71 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_123 ();
 sg13g2_fill_1 FILLER_25_128 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_295 ();
 sg13g2_fill_1 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_374 ();
 sg13g2_fill_1 FILLER_25_379 ();
 sg13g2_decap_4 FILLER_26_212 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_352 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_390 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_27_40 ();
 sg13g2_fill_1 FILLER_27_42 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_fill_1 FILLER_27_62 ();
 sg13g2_fill_2 FILLER_27_138 ();
 sg13g2_fill_2 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_fill_1 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_73 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_fill_2 FILLER_28_224 ();
 sg13g2_fill_1 FILLER_28_388 ();
 sg13g2_fill_1 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_29_41 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_decap_4 FILLER_29_236 ();
 sg13g2_fill_1 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_263 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_fill_1 FILLER_29_359 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_51 ();
 sg13g2_fill_1 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_74 ();
 sg13g2_fill_1 FILLER_30_76 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_240 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_fill_1 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_27 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_decap_4 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_243 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_32_26 ();
 sg13g2_fill_1 FILLER_32_34 ();
 sg13g2_fill_1 FILLER_32_71 ();
 sg13g2_fill_2 FILLER_32_164 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_fill_2 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_82 ();
 sg13g2_fill_1 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_fill_2 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_167 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_2 FILLER_33_228 ();
 sg13g2_fill_1 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_315 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_348 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_fill_2 FILLER_33_392 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_1 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_140 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_315 ();
 sg13g2_fill_1 FILLER_35_36 ();
 sg13g2_fill_2 FILLER_35_73 ();
 sg13g2_fill_2 FILLER_35_162 ();
 sg13g2_fill_2 FILLER_35_174 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_272 ();
 sg13g2_fill_1 FILLER_35_343 ();
 sg13g2_fill_1 FILLER_35_424 ();
 sg13g2_fill_1 FILLER_36_5 ();
 sg13g2_fill_1 FILLER_36_77 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_2 FILLER_36_122 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_297 ();
 sg13g2_fill_2 FILLER_36_402 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_2 FILLER_37_91 ();
 sg13g2_fill_2 FILLER_37_258 ();
 sg13g2_fill_1 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_279 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_fill_1 FILLER_37_321 ();
 sg13g2_fill_1 FILLER_37_377 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_93 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_2 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_2 FILLER_38_183 ();
 sg13g2_fill_1 FILLER_38_189 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_241 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_382 ();
 sg13g2_fill_1 FILLER_38_399 ();
 sg13g2_fill_1 FILLER_38_410 ();
 sg13g2_fill_1 FILLER_38_419 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
