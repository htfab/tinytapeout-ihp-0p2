module tt_um_ccattuto_conway (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire _4601_;
 wire _4602_;
 wire _4603_;
 wire _4604_;
 wire _4605_;
 wire _4606_;
 wire _4607_;
 wire _4608_;
 wire _4609_;
 wire _4610_;
 wire _4611_;
 wire _4612_;
 wire _4613_;
 wire _4614_;
 wire _4615_;
 wire _4616_;
 wire _4617_;
 wire _4618_;
 wire _4619_;
 wire _4620_;
 wire _4621_;
 wire _4622_;
 wire _4623_;
 wire _4624_;
 wire _4625_;
 wire _4626_;
 wire _4627_;
 wire _4628_;
 wire _4629_;
 wire _4630_;
 wire _4631_;
 wire _4632_;
 wire _4633_;
 wire _4634_;
 wire _4635_;
 wire _4636_;
 wire _4637_;
 wire _4638_;
 wire _4639_;
 wire _4640_;
 wire _4641_;
 wire _4642_;
 wire _4643_;
 wire _4644_;
 wire _4645_;
 wire _4646_;
 wire _4647_;
 wire _4648_;
 wire _4649_;
 wire _4650_;
 wire _4651_;
 wire _4652_;
 wire _4653_;
 wire _4654_;
 wire _4655_;
 wire _4656_;
 wire _4657_;
 wire _4658_;
 wire _4659_;
 wire _4660_;
 wire _4661_;
 wire _4662_;
 wire _4663_;
 wire _4664_;
 wire _4665_;
 wire _4666_;
 wire _4667_;
 wire _4668_;
 wire _4669_;
 wire _4670_;
 wire _4671_;
 wire _4672_;
 wire _4673_;
 wire _4674_;
 wire _4675_;
 wire _4676_;
 wire _4677_;
 wire _4678_;
 wire _4679_;
 wire _4680_;
 wire _4681_;
 wire _4682_;
 wire _4683_;
 wire _4684_;
 wire _4685_;
 wire _4686_;
 wire _4687_;
 wire _4688_;
 wire _4689_;
 wire _4690_;
 wire _4691_;
 wire _4692_;
 wire _4693_;
 wire _4694_;
 wire _4695_;
 wire _4696_;
 wire _4697_;
 wire _4698_;
 wire _4699_;
 wire _4700_;
 wire _4701_;
 wire _4702_;
 wire _4703_;
 wire _4704_;
 wire _4705_;
 wire _4706_;
 wire _4707_;
 wire _4708_;
 wire _4709_;
 wire _4710_;
 wire _4711_;
 wire _4712_;
 wire _4713_;
 wire _4714_;
 wire _4715_;
 wire _4716_;
 wire _4717_;
 wire _4718_;
 wire _4719_;
 wire _4720_;
 wire _4721_;
 wire _4722_;
 wire _4723_;
 wire _4724_;
 wire _4725_;
 wire _4726_;
 wire _4727_;
 wire _4728_;
 wire _4729_;
 wire _4730_;
 wire _4731_;
 wire _4732_;
 wire _4733_;
 wire _4734_;
 wire _4735_;
 wire _4736_;
 wire _4737_;
 wire _4738_;
 wire _4739_;
 wire _4740_;
 wire _4741_;
 wire _4742_;
 wire _4743_;
 wire _4744_;
 wire _4745_;
 wire _4746_;
 wire _4747_;
 wire _4748_;
 wire _4749_;
 wire _4750_;
 wire _4751_;
 wire _4752_;
 wire _4753_;
 wire _4754_;
 wire _4755_;
 wire _4756_;
 wire _4757_;
 wire _4758_;
 wire _4759_;
 wire _4760_;
 wire _4761_;
 wire _4762_;
 wire _4763_;
 wire _4764_;
 wire _4765_;
 wire _4766_;
 wire _4767_;
 wire _4768_;
 wire _4769_;
 wire _4770_;
 wire _4771_;
 wire _4772_;
 wire _4773_;
 wire _4774_;
 wire _4775_;
 wire _4776_;
 wire _4777_;
 wire _4778_;
 wire _4779_;
 wire _4780_;
 wire _4781_;
 wire _4782_;
 wire _4783_;
 wire _4784_;
 wire _4785_;
 wire _4786_;
 wire _4787_;
 wire _4788_;
 wire _4789_;
 wire _4790_;
 wire _4791_;
 wire _4792_;
 wire _4793_;
 wire _4794_;
 wire _4795_;
 wire _4796_;
 wire _4797_;
 wire _4798_;
 wire _4799_;
 wire _4800_;
 wire _4801_;
 wire _4802_;
 wire _4803_;
 wire _4804_;
 wire _4805_;
 wire _4806_;
 wire _4807_;
 wire _4808_;
 wire _4809_;
 wire _4810_;
 wire _4811_;
 wire _4812_;
 wire _4813_;
 wire _4814_;
 wire _4815_;
 wire _4816_;
 wire _4817_;
 wire _4818_;
 wire _4819_;
 wire _4820_;
 wire _4821_;
 wire _4822_;
 wire _4823_;
 wire _4824_;
 wire _4825_;
 wire _4826_;
 wire _4827_;
 wire _4828_;
 wire _4829_;
 wire _4830_;
 wire _4831_;
 wire _4832_;
 wire _4833_;
 wire _4834_;
 wire _4835_;
 wire _4836_;
 wire _4837_;
 wire _4838_;
 wire _4839_;
 wire _4840_;
 wire _4841_;
 wire _4842_;
 wire _4843_;
 wire _4844_;
 wire _4845_;
 wire _4846_;
 wire _4847_;
 wire _4848_;
 wire _4849_;
 wire _4850_;
 wire _4851_;
 wire _4852_;
 wire _4853_;
 wire _4854_;
 wire _4855_;
 wire _4856_;
 wire _4857_;
 wire _4858_;
 wire _4859_;
 wire _4860_;
 wire _4861_;
 wire _4862_;
 wire _4863_;
 wire _4864_;
 wire _4865_;
 wire _4866_;
 wire _4867_;
 wire _4868_;
 wire _4869_;
 wire _4870_;
 wire _4871_;
 wire _4872_;
 wire _4873_;
 wire _4874_;
 wire _4875_;
 wire _4876_;
 wire _4877_;
 wire _4878_;
 wire _4879_;
 wire _4880_;
 wire _4881_;
 wire _4882_;
 wire _4883_;
 wire _4884_;
 wire _4885_;
 wire _4886_;
 wire _4887_;
 wire _4888_;
 wire _4889_;
 wire _4890_;
 wire _4891_;
 wire _4892_;
 wire _4893_;
 wire _4894_;
 wire _4895_;
 wire _4896_;
 wire _4897_;
 wire _4898_;
 wire _4899_;
 wire _4900_;
 wire _4901_;
 wire _4902_;
 wire _4903_;
 wire _4904_;
 wire _4905_;
 wire _4906_;
 wire _4907_;
 wire _4908_;
 wire _4909_;
 wire _4910_;
 wire _4911_;
 wire _4912_;
 wire _4913_;
 wire _4914_;
 wire _4915_;
 wire _4916_;
 wire _4917_;
 wire _4918_;
 wire _4919_;
 wire _4920_;
 wire _4921_;
 wire _4922_;
 wire _4923_;
 wire _4924_;
 wire _4925_;
 wire _4926_;
 wire _4927_;
 wire _4928_;
 wire _4929_;
 wire _4930_;
 wire _4931_;
 wire _4932_;
 wire _4933_;
 wire _4934_;
 wire _4935_;
 wire _4936_;
 wire _4937_;
 wire _4938_;
 wire _4939_;
 wire _4940_;
 wire _4941_;
 wire _4942_;
 wire _4943_;
 wire _4944_;
 wire _4945_;
 wire _4946_;
 wire _4947_;
 wire _4948_;
 wire _4949_;
 wire _4950_;
 wire _4951_;
 wire _4952_;
 wire _4953_;
 wire _4954_;
 wire _4955_;
 wire _4956_;
 wire _4957_;
 wire _4958_;
 wire _4959_;
 wire _4960_;
 wire _4961_;
 wire _4962_;
 wire _4963_;
 wire _4964_;
 wire _4965_;
 wire _4966_;
 wire _4967_;
 wire _4968_;
 wire _4969_;
 wire _4970_;
 wire _4971_;
 wire _4972_;
 wire _4973_;
 wire _4974_;
 wire _4975_;
 wire _4976_;
 wire _4977_;
 wire _4978_;
 wire _4979_;
 wire _4980_;
 wire _4981_;
 wire _4982_;
 wire _4983_;
 wire _4984_;
 wire _4985_;
 wire _4986_;
 wire _4987_;
 wire _4988_;
 wire _4989_;
 wire _4990_;
 wire _4991_;
 wire _4992_;
 wire _4993_;
 wire _4994_;
 wire _4995_;
 wire _4996_;
 wire _4997_;
 wire _4998_;
 wire _4999_;
 wire _5000_;
 wire _5001_;
 wire _5002_;
 wire _5003_;
 wire _5004_;
 wire _5005_;
 wire _5006_;
 wire _5007_;
 wire _5008_;
 wire _5009_;
 wire _5010_;
 wire _5011_;
 wire _5012_;
 wire _5013_;
 wire _5014_;
 wire _5015_;
 wire _5016_;
 wire _5017_;
 wire _5018_;
 wire _5019_;
 wire _5020_;
 wire _5021_;
 wire _5022_;
 wire _5023_;
 wire _5024_;
 wire _5025_;
 wire _5026_;
 wire _5027_;
 wire _5028_;
 wire _5029_;
 wire _5030_;
 wire _5031_;
 wire _5032_;
 wire _5033_;
 wire _5034_;
 wire _5035_;
 wire _5036_;
 wire _5037_;
 wire _5038_;
 wire _5039_;
 wire _5040_;
 wire _5041_;
 wire _5042_;
 wire _5043_;
 wire _5044_;
 wire _5045_;
 wire _5046_;
 wire _5047_;
 wire _5048_;
 wire _5049_;
 wire _5050_;
 wire _5051_;
 wire _5052_;
 wire _5053_;
 wire _5054_;
 wire _5055_;
 wire _5056_;
 wire _5057_;
 wire _5058_;
 wire _5059_;
 wire _5060_;
 wire _5061_;
 wire _5062_;
 wire _5063_;
 wire _5064_;
 wire _5065_;
 wire _5066_;
 wire _5067_;
 wire _5068_;
 wire _5069_;
 wire _5070_;
 wire _5071_;
 wire _5072_;
 wire _5073_;
 wire _5074_;
 wire _5075_;
 wire _5076_;
 wire _5077_;
 wire _5078_;
 wire _5079_;
 wire _5080_;
 wire _5081_;
 wire _5082_;
 wire _5083_;
 wire _5084_;
 wire _5085_;
 wire _5086_;
 wire _5087_;
 wire _5088_;
 wire _5089_;
 wire _5090_;
 wire _5091_;
 wire _5092_;
 wire _5093_;
 wire _5094_;
 wire _5095_;
 wire _5096_;
 wire _5097_;
 wire _5098_;
 wire _5099_;
 wire _5100_;
 wire _5101_;
 wire _5102_;
 wire _5103_;
 wire _5104_;
 wire _5105_;
 wire _5106_;
 wire _5107_;
 wire _5108_;
 wire _5109_;
 wire _5110_;
 wire _5111_;
 wire _5112_;
 wire _5113_;
 wire _5114_;
 wire _5115_;
 wire _5116_;
 wire _5117_;
 wire _5118_;
 wire _5119_;
 wire _5120_;
 wire _5121_;
 wire _5122_;
 wire _5123_;
 wire _5124_;
 wire _5125_;
 wire _5126_;
 wire _5127_;
 wire _5128_;
 wire _5129_;
 wire _5130_;
 wire _5131_;
 wire _5132_;
 wire _5133_;
 wire _5134_;
 wire _5135_;
 wire _5136_;
 wire _5137_;
 wire _5138_;
 wire _5139_;
 wire _5140_;
 wire _5141_;
 wire _5142_;
 wire _5143_;
 wire _5144_;
 wire _5145_;
 wire _5146_;
 wire _5147_;
 wire _5148_;
 wire _5149_;
 wire _5150_;
 wire _5151_;
 wire _5152_;
 wire _5153_;
 wire _5154_;
 wire _5155_;
 wire _5156_;
 wire _5157_;
 wire _5158_;
 wire _5159_;
 wire _5160_;
 wire _5161_;
 wire _5162_;
 wire _5163_;
 wire _5164_;
 wire _5165_;
 wire _5166_;
 wire _5167_;
 wire _5168_;
 wire _5169_;
 wire _5170_;
 wire _5171_;
 wire _5172_;
 wire _5173_;
 wire _5174_;
 wire _5175_;
 wire _5176_;
 wire _5177_;
 wire _5178_;
 wire _5179_;
 wire _5180_;
 wire _5181_;
 wire _5182_;
 wire _5183_;
 wire _5184_;
 wire _5185_;
 wire _5186_;
 wire _5187_;
 wire _5188_;
 wire _5189_;
 wire _5190_;
 wire _5191_;
 wire _5192_;
 wire _5193_;
 wire _5194_;
 wire _5195_;
 wire _5196_;
 wire _5197_;
 wire _5198_;
 wire _5199_;
 wire _5200_;
 wire _5201_;
 wire _5202_;
 wire _5203_;
 wire _5204_;
 wire _5205_;
 wire _5206_;
 wire _5207_;
 wire _5208_;
 wire _5209_;
 wire _5210_;
 wire _5211_;
 wire _5212_;
 wire _5213_;
 wire _5214_;
 wire _5215_;
 wire _5216_;
 wire _5217_;
 wire _5218_;
 wire _5219_;
 wire _5220_;
 wire _5221_;
 wire _5222_;
 wire _5223_;
 wire _5224_;
 wire _5225_;
 wire _5226_;
 wire _5227_;
 wire _5228_;
 wire _5229_;
 wire _5230_;
 wire _5231_;
 wire _5232_;
 wire _5233_;
 wire _5234_;
 wire _5235_;
 wire _5236_;
 wire _5237_;
 wire _5238_;
 wire _5239_;
 wire _5240_;
 wire _5241_;
 wire _5242_;
 wire _5243_;
 wire _5244_;
 wire _5245_;
 wire _5246_;
 wire _5247_;
 wire _5248_;
 wire _5249_;
 wire _5250_;
 wire _5251_;
 wire _5252_;
 wire _5253_;
 wire _5254_;
 wire _5255_;
 wire _5256_;
 wire _5257_;
 wire _5258_;
 wire _5259_;
 wire _5260_;
 wire _5261_;
 wire _5262_;
 wire _5263_;
 wire _5264_;
 wire _5265_;
 wire _5266_;
 wire _5267_;
 wire _5268_;
 wire _5269_;
 wire _5270_;
 wire _5271_;
 wire _5272_;
 wire _5273_;
 wire _5274_;
 wire _5275_;
 wire _5276_;
 wire _5277_;
 wire _5278_;
 wire _5279_;
 wire _5280_;
 wire _5281_;
 wire _5282_;
 wire _5283_;
 wire _5284_;
 wire _5285_;
 wire _5286_;
 wire _5287_;
 wire _5288_;
 wire _5289_;
 wire _5290_;
 wire _5291_;
 wire _5292_;
 wire _5293_;
 wire _5294_;
 wire _5295_;
 wire _5296_;
 wire _5297_;
 wire _5298_;
 wire _5299_;
 wire _5300_;
 wire _5301_;
 wire _5302_;
 wire _5303_;
 wire _5304_;
 wire _5305_;
 wire _5306_;
 wire _5307_;
 wire _5308_;
 wire _5309_;
 wire _5310_;
 wire _5311_;
 wire _5312_;
 wire _5313_;
 wire _5314_;
 wire _5315_;
 wire _5316_;
 wire _5317_;
 wire _5318_;
 wire _5319_;
 wire _5320_;
 wire _5321_;
 wire _5322_;
 wire _5323_;
 wire _5324_;
 wire _5325_;
 wire _5326_;
 wire _5327_;
 wire _5328_;
 wire _5329_;
 wire _5330_;
 wire _5331_;
 wire _5332_;
 wire _5333_;
 wire _5334_;
 wire _5335_;
 wire _5336_;
 wire _5337_;
 wire _5338_;
 wire _5339_;
 wire _5340_;
 wire _5341_;
 wire _5342_;
 wire _5343_;
 wire _5344_;
 wire _5345_;
 wire _5346_;
 wire _5347_;
 wire _5348_;
 wire _5349_;
 wire _5350_;
 wire _5351_;
 wire _5352_;
 wire _5353_;
 wire _5354_;
 wire _5355_;
 wire _5356_;
 wire _5357_;
 wire _5358_;
 wire _5359_;
 wire _5360_;
 wire _5361_;
 wire _5362_;
 wire _5363_;
 wire _5364_;
 wire _5365_;
 wire _5366_;
 wire _5367_;
 wire _5368_;
 wire _5369_;
 wire _5370_;
 wire _5371_;
 wire _5372_;
 wire _5373_;
 wire _5374_;
 wire _5375_;
 wire _5376_;
 wire _5377_;
 wire _5378_;
 wire _5379_;
 wire _5380_;
 wire _5381_;
 wire _5382_;
 wire _5383_;
 wire _5384_;
 wire _5385_;
 wire _5386_;
 wire _5387_;
 wire _5388_;
 wire _5389_;
 wire _5390_;
 wire _5391_;
 wire _5392_;
 wire _5393_;
 wire _5394_;
 wire _5395_;
 wire _5396_;
 wire _5397_;
 wire _5398_;
 wire _5399_;
 wire _5400_;
 wire _5401_;
 wire _5402_;
 wire _5403_;
 wire _5404_;
 wire _5405_;
 wire _5406_;
 wire _5407_;
 wire _5408_;
 wire _5409_;
 wire _5410_;
 wire _5411_;
 wire _5412_;
 wire _5413_;
 wire _5414_;
 wire _5415_;
 wire _5416_;
 wire _5417_;
 wire _5418_;
 wire clknet_leaf_0_clk;
 wire net417;
 wire \action[0] ;
 wire \action[1] ;
 wire \action[2] ;
 wire \action[3] ;
 wire \action[4] ;
 wire \action[5] ;
 wire \action[6] ;
 wire \action[7] ;
 wire \board_state[0] ;
 wire \board_state[100] ;
 wire \board_state[101] ;
 wire \board_state[102] ;
 wire \board_state[103] ;
 wire \board_state[104] ;
 wire \board_state[105] ;
 wire \board_state[106] ;
 wire \board_state[107] ;
 wire \board_state[108] ;
 wire \board_state[109] ;
 wire \board_state[10] ;
 wire \board_state[110] ;
 wire \board_state[111] ;
 wire \board_state[112] ;
 wire \board_state[113] ;
 wire \board_state[114] ;
 wire \board_state[115] ;
 wire \board_state[116] ;
 wire \board_state[117] ;
 wire \board_state[118] ;
 wire \board_state[119] ;
 wire \board_state[11] ;
 wire \board_state[120] ;
 wire \board_state[121] ;
 wire \board_state[122] ;
 wire \board_state[123] ;
 wire \board_state[124] ;
 wire \board_state[125] ;
 wire \board_state[126] ;
 wire \board_state[127] ;
 wire \board_state[128] ;
 wire \board_state[129] ;
 wire \board_state[12] ;
 wire \board_state[130] ;
 wire \board_state[131] ;
 wire \board_state[132] ;
 wire \board_state[133] ;
 wire \board_state[134] ;
 wire \board_state[135] ;
 wire \board_state[136] ;
 wire \board_state[137] ;
 wire \board_state[138] ;
 wire \board_state[139] ;
 wire \board_state[13] ;
 wire \board_state[140] ;
 wire \board_state[141] ;
 wire \board_state[142] ;
 wire \board_state[143] ;
 wire \board_state[144] ;
 wire \board_state[145] ;
 wire \board_state[146] ;
 wire \board_state[147] ;
 wire \board_state[148] ;
 wire \board_state[149] ;
 wire \board_state[14] ;
 wire \board_state[150] ;
 wire \board_state[151] ;
 wire \board_state[152] ;
 wire \board_state[153] ;
 wire \board_state[154] ;
 wire \board_state[155] ;
 wire \board_state[156] ;
 wire \board_state[157] ;
 wire \board_state[158] ;
 wire \board_state[159] ;
 wire \board_state[15] ;
 wire \board_state[160] ;
 wire \board_state[161] ;
 wire \board_state[162] ;
 wire \board_state[163] ;
 wire \board_state[164] ;
 wire \board_state[165] ;
 wire \board_state[166] ;
 wire \board_state[167] ;
 wire \board_state[168] ;
 wire \board_state[169] ;
 wire \board_state[16] ;
 wire \board_state[170] ;
 wire \board_state[171] ;
 wire \board_state[172] ;
 wire \board_state[173] ;
 wire \board_state[174] ;
 wire \board_state[175] ;
 wire \board_state[176] ;
 wire \board_state[177] ;
 wire \board_state[178] ;
 wire \board_state[179] ;
 wire \board_state[17] ;
 wire \board_state[180] ;
 wire \board_state[181] ;
 wire \board_state[182] ;
 wire \board_state[183] ;
 wire \board_state[184] ;
 wire \board_state[185] ;
 wire \board_state[186] ;
 wire \board_state[187] ;
 wire \board_state[188] ;
 wire \board_state[189] ;
 wire \board_state[18] ;
 wire \board_state[190] ;
 wire \board_state[191] ;
 wire \board_state[192] ;
 wire \board_state[193] ;
 wire \board_state[194] ;
 wire \board_state[195] ;
 wire \board_state[196] ;
 wire \board_state[197] ;
 wire \board_state[198] ;
 wire \board_state[199] ;
 wire \board_state[19] ;
 wire \board_state[1] ;
 wire \board_state[200] ;
 wire \board_state[201] ;
 wire \board_state[202] ;
 wire \board_state[203] ;
 wire \board_state[204] ;
 wire \board_state[205] ;
 wire \board_state[206] ;
 wire \board_state[207] ;
 wire \board_state[208] ;
 wire \board_state[209] ;
 wire \board_state[20] ;
 wire \board_state[210] ;
 wire \board_state[211] ;
 wire \board_state[212] ;
 wire \board_state[213] ;
 wire \board_state[214] ;
 wire \board_state[215] ;
 wire \board_state[216] ;
 wire \board_state[217] ;
 wire \board_state[218] ;
 wire \board_state[219] ;
 wire \board_state[21] ;
 wire \board_state[220] ;
 wire \board_state[221] ;
 wire \board_state[222] ;
 wire \board_state[223] ;
 wire \board_state[224] ;
 wire \board_state[225] ;
 wire \board_state[226] ;
 wire \board_state[227] ;
 wire \board_state[228] ;
 wire \board_state[229] ;
 wire \board_state[22] ;
 wire \board_state[230] ;
 wire \board_state[231] ;
 wire \board_state[232] ;
 wire \board_state[233] ;
 wire \board_state[234] ;
 wire \board_state[235] ;
 wire \board_state[236] ;
 wire \board_state[237] ;
 wire \board_state[238] ;
 wire \board_state[239] ;
 wire \board_state[23] ;
 wire \board_state[240] ;
 wire \board_state[241] ;
 wire \board_state[242] ;
 wire \board_state[243] ;
 wire \board_state[244] ;
 wire \board_state[245] ;
 wire \board_state[246] ;
 wire \board_state[247] ;
 wire \board_state[248] ;
 wire \board_state[249] ;
 wire \board_state[24] ;
 wire \board_state[250] ;
 wire \board_state[251] ;
 wire \board_state[252] ;
 wire \board_state[253] ;
 wire \board_state[254] ;
 wire \board_state[255] ;
 wire \board_state[256] ;
 wire \board_state[257] ;
 wire \board_state[258] ;
 wire \board_state[259] ;
 wire \board_state[25] ;
 wire \board_state[260] ;
 wire \board_state[261] ;
 wire \board_state[262] ;
 wire \board_state[263] ;
 wire \board_state[264] ;
 wire \board_state[265] ;
 wire \board_state[266] ;
 wire \board_state[267] ;
 wire \board_state[268] ;
 wire \board_state[269] ;
 wire \board_state[26] ;
 wire \board_state[270] ;
 wire \board_state[271] ;
 wire \board_state[272] ;
 wire \board_state[273] ;
 wire \board_state[274] ;
 wire \board_state[275] ;
 wire \board_state[276] ;
 wire \board_state[277] ;
 wire \board_state[278] ;
 wire \board_state[279] ;
 wire \board_state[27] ;
 wire \board_state[280] ;
 wire \board_state[281] ;
 wire \board_state[282] ;
 wire \board_state[283] ;
 wire \board_state[284] ;
 wire \board_state[285] ;
 wire \board_state[286] ;
 wire \board_state[287] ;
 wire \board_state[288] ;
 wire \board_state[289] ;
 wire \board_state[28] ;
 wire \board_state[290] ;
 wire \board_state[291] ;
 wire \board_state[292] ;
 wire \board_state[293] ;
 wire \board_state[294] ;
 wire \board_state[295] ;
 wire \board_state[296] ;
 wire \board_state[297] ;
 wire \board_state[298] ;
 wire \board_state[299] ;
 wire \board_state[29] ;
 wire \board_state[2] ;
 wire \board_state[300] ;
 wire \board_state[301] ;
 wire \board_state[302] ;
 wire \board_state[303] ;
 wire \board_state[304] ;
 wire \board_state[305] ;
 wire \board_state[306] ;
 wire \board_state[307] ;
 wire \board_state[308] ;
 wire \board_state[309] ;
 wire \board_state[30] ;
 wire \board_state[310] ;
 wire \board_state[311] ;
 wire \board_state[312] ;
 wire \board_state[313] ;
 wire \board_state[314] ;
 wire \board_state[315] ;
 wire \board_state[316] ;
 wire \board_state[317] ;
 wire \board_state[318] ;
 wire \board_state[319] ;
 wire \board_state[31] ;
 wire \board_state[320] ;
 wire \board_state[321] ;
 wire \board_state[322] ;
 wire \board_state[323] ;
 wire \board_state[324] ;
 wire \board_state[325] ;
 wire \board_state[326] ;
 wire \board_state[327] ;
 wire \board_state[328] ;
 wire \board_state[329] ;
 wire \board_state[32] ;
 wire \board_state[330] ;
 wire \board_state[331] ;
 wire \board_state[332] ;
 wire \board_state[333] ;
 wire \board_state[334] ;
 wire \board_state[335] ;
 wire \board_state[336] ;
 wire \board_state[337] ;
 wire \board_state[338] ;
 wire \board_state[339] ;
 wire \board_state[33] ;
 wire \board_state[340] ;
 wire \board_state[341] ;
 wire \board_state[342] ;
 wire \board_state[343] ;
 wire \board_state[344] ;
 wire \board_state[345] ;
 wire \board_state[346] ;
 wire \board_state[347] ;
 wire \board_state[348] ;
 wire \board_state[349] ;
 wire \board_state[34] ;
 wire \board_state[350] ;
 wire \board_state[351] ;
 wire \board_state[352] ;
 wire \board_state[353] ;
 wire \board_state[354] ;
 wire \board_state[355] ;
 wire \board_state[356] ;
 wire \board_state[357] ;
 wire \board_state[358] ;
 wire \board_state[359] ;
 wire \board_state[35] ;
 wire \board_state[360] ;
 wire \board_state[361] ;
 wire \board_state[362] ;
 wire \board_state[363] ;
 wire \board_state[364] ;
 wire \board_state[365] ;
 wire \board_state[366] ;
 wire \board_state[367] ;
 wire \board_state[368] ;
 wire \board_state[369] ;
 wire \board_state[36] ;
 wire \board_state[370] ;
 wire \board_state[371] ;
 wire \board_state[372] ;
 wire \board_state[373] ;
 wire \board_state[374] ;
 wire \board_state[375] ;
 wire \board_state[376] ;
 wire \board_state[377] ;
 wire \board_state[378] ;
 wire \board_state[379] ;
 wire \board_state[37] ;
 wire \board_state[380] ;
 wire \board_state[381] ;
 wire \board_state[382] ;
 wire \board_state[383] ;
 wire \board_state[384] ;
 wire \board_state[385] ;
 wire \board_state[386] ;
 wire \board_state[387] ;
 wire \board_state[388] ;
 wire \board_state[389] ;
 wire \board_state[38] ;
 wire \board_state[390] ;
 wire \board_state[391] ;
 wire \board_state[392] ;
 wire \board_state[393] ;
 wire \board_state[394] ;
 wire \board_state[395] ;
 wire \board_state[396] ;
 wire \board_state[397] ;
 wire \board_state[398] ;
 wire \board_state[399] ;
 wire \board_state[39] ;
 wire \board_state[3] ;
 wire \board_state[400] ;
 wire \board_state[401] ;
 wire \board_state[402] ;
 wire \board_state[403] ;
 wire \board_state[404] ;
 wire \board_state[405] ;
 wire \board_state[406] ;
 wire \board_state[407] ;
 wire \board_state[408] ;
 wire \board_state[409] ;
 wire \board_state[40] ;
 wire \board_state[410] ;
 wire \board_state[411] ;
 wire \board_state[412] ;
 wire \board_state[413] ;
 wire \board_state[414] ;
 wire \board_state[415] ;
 wire \board_state[416] ;
 wire \board_state[417] ;
 wire \board_state[418] ;
 wire \board_state[419] ;
 wire \board_state[41] ;
 wire \board_state[420] ;
 wire \board_state[421] ;
 wire \board_state[422] ;
 wire \board_state[423] ;
 wire \board_state[424] ;
 wire \board_state[425] ;
 wire \board_state[426] ;
 wire \board_state[427] ;
 wire \board_state[428] ;
 wire \board_state[429] ;
 wire \board_state[42] ;
 wire \board_state[430] ;
 wire \board_state[431] ;
 wire \board_state[432] ;
 wire \board_state[433] ;
 wire \board_state[434] ;
 wire \board_state[435] ;
 wire \board_state[436] ;
 wire \board_state[437] ;
 wire \board_state[438] ;
 wire \board_state[439] ;
 wire \board_state[43] ;
 wire \board_state[440] ;
 wire \board_state[441] ;
 wire \board_state[442] ;
 wire \board_state[443] ;
 wire \board_state[444] ;
 wire \board_state[445] ;
 wire \board_state[446] ;
 wire \board_state[447] ;
 wire \board_state[448] ;
 wire \board_state[449] ;
 wire \board_state[44] ;
 wire \board_state[450] ;
 wire \board_state[451] ;
 wire \board_state[452] ;
 wire \board_state[453] ;
 wire \board_state[454] ;
 wire \board_state[455] ;
 wire \board_state[456] ;
 wire \board_state[457] ;
 wire \board_state[458] ;
 wire \board_state[459] ;
 wire \board_state[45] ;
 wire \board_state[460] ;
 wire \board_state[461] ;
 wire \board_state[462] ;
 wire \board_state[463] ;
 wire \board_state[464] ;
 wire \board_state[465] ;
 wire \board_state[466] ;
 wire \board_state[467] ;
 wire \board_state[468] ;
 wire \board_state[469] ;
 wire \board_state[46] ;
 wire \board_state[470] ;
 wire \board_state[471] ;
 wire \board_state[472] ;
 wire \board_state[473] ;
 wire \board_state[474] ;
 wire \board_state[475] ;
 wire \board_state[476] ;
 wire \board_state[477] ;
 wire \board_state[478] ;
 wire \board_state[479] ;
 wire \board_state[47] ;
 wire \board_state[480] ;
 wire \board_state[481] ;
 wire \board_state[482] ;
 wire \board_state[483] ;
 wire \board_state[484] ;
 wire \board_state[485] ;
 wire \board_state[486] ;
 wire \board_state[487] ;
 wire \board_state[488] ;
 wire \board_state[489] ;
 wire \board_state[48] ;
 wire \board_state[490] ;
 wire \board_state[491] ;
 wire \board_state[492] ;
 wire \board_state[493] ;
 wire \board_state[494] ;
 wire \board_state[495] ;
 wire \board_state[496] ;
 wire \board_state[497] ;
 wire \board_state[498] ;
 wire \board_state[499] ;
 wire \board_state[49] ;
 wire \board_state[4] ;
 wire \board_state[500] ;
 wire \board_state[501] ;
 wire \board_state[502] ;
 wire \board_state[503] ;
 wire \board_state[504] ;
 wire \board_state[505] ;
 wire \board_state[506] ;
 wire \board_state[507] ;
 wire \board_state[508] ;
 wire \board_state[509] ;
 wire \board_state[50] ;
 wire \board_state[510] ;
 wire \board_state[511] ;
 wire \board_state[51] ;
 wire \board_state[52] ;
 wire \board_state[53] ;
 wire \board_state[54] ;
 wire \board_state[55] ;
 wire \board_state[56] ;
 wire \board_state[57] ;
 wire \board_state[58] ;
 wire \board_state[59] ;
 wire \board_state[5] ;
 wire \board_state[60] ;
 wire \board_state[61] ;
 wire \board_state[62] ;
 wire \board_state[63] ;
 wire \board_state[64] ;
 wire \board_state[65] ;
 wire \board_state[66] ;
 wire \board_state[67] ;
 wire \board_state[68] ;
 wire \board_state[69] ;
 wire \board_state[6] ;
 wire \board_state[70] ;
 wire \board_state[71] ;
 wire \board_state[72] ;
 wire \board_state[73] ;
 wire \board_state[74] ;
 wire \board_state[75] ;
 wire \board_state[76] ;
 wire \board_state[77] ;
 wire \board_state[78] ;
 wire \board_state[79] ;
 wire \board_state[7] ;
 wire \board_state[80] ;
 wire \board_state[81] ;
 wire \board_state[82] ;
 wire \board_state[83] ;
 wire \board_state[84] ;
 wire \board_state[85] ;
 wire \board_state[86] ;
 wire \board_state[87] ;
 wire \board_state[88] ;
 wire \board_state[89] ;
 wire \board_state[8] ;
 wire \board_state[90] ;
 wire \board_state[91] ;
 wire \board_state[92] ;
 wire \board_state[93] ;
 wire \board_state[94] ;
 wire \board_state[95] ;
 wire \board_state[96] ;
 wire \board_state[97] ;
 wire \board_state[98] ;
 wire \board_state[99] ;
 wire \board_state[9] ;
 wire \board_state_next[0] ;
 wire \board_state_next[100] ;
 wire \board_state_next[101] ;
 wire \board_state_next[102] ;
 wire \board_state_next[103] ;
 wire \board_state_next[104] ;
 wire \board_state_next[105] ;
 wire \board_state_next[106] ;
 wire \board_state_next[107] ;
 wire \board_state_next[108] ;
 wire \board_state_next[109] ;
 wire \board_state_next[10] ;
 wire \board_state_next[110] ;
 wire \board_state_next[111] ;
 wire \board_state_next[112] ;
 wire \board_state_next[113] ;
 wire \board_state_next[114] ;
 wire \board_state_next[115] ;
 wire \board_state_next[116] ;
 wire \board_state_next[117] ;
 wire \board_state_next[118] ;
 wire \board_state_next[119] ;
 wire \board_state_next[11] ;
 wire \board_state_next[120] ;
 wire \board_state_next[121] ;
 wire \board_state_next[122] ;
 wire \board_state_next[123] ;
 wire \board_state_next[124] ;
 wire \board_state_next[125] ;
 wire \board_state_next[126] ;
 wire \board_state_next[127] ;
 wire \board_state_next[128] ;
 wire \board_state_next[129] ;
 wire \board_state_next[12] ;
 wire \board_state_next[130] ;
 wire \board_state_next[131] ;
 wire \board_state_next[132] ;
 wire \board_state_next[133] ;
 wire \board_state_next[134] ;
 wire \board_state_next[135] ;
 wire \board_state_next[136] ;
 wire \board_state_next[137] ;
 wire \board_state_next[138] ;
 wire \board_state_next[139] ;
 wire \board_state_next[13] ;
 wire \board_state_next[140] ;
 wire \board_state_next[141] ;
 wire \board_state_next[142] ;
 wire \board_state_next[143] ;
 wire \board_state_next[144] ;
 wire \board_state_next[145] ;
 wire \board_state_next[146] ;
 wire \board_state_next[147] ;
 wire \board_state_next[148] ;
 wire \board_state_next[149] ;
 wire \board_state_next[14] ;
 wire \board_state_next[150] ;
 wire \board_state_next[151] ;
 wire \board_state_next[152] ;
 wire \board_state_next[153] ;
 wire \board_state_next[154] ;
 wire \board_state_next[155] ;
 wire \board_state_next[156] ;
 wire \board_state_next[157] ;
 wire \board_state_next[158] ;
 wire \board_state_next[159] ;
 wire \board_state_next[15] ;
 wire \board_state_next[160] ;
 wire \board_state_next[161] ;
 wire \board_state_next[162] ;
 wire \board_state_next[163] ;
 wire \board_state_next[164] ;
 wire \board_state_next[165] ;
 wire \board_state_next[166] ;
 wire \board_state_next[167] ;
 wire \board_state_next[168] ;
 wire \board_state_next[169] ;
 wire \board_state_next[16] ;
 wire \board_state_next[170] ;
 wire \board_state_next[171] ;
 wire \board_state_next[172] ;
 wire \board_state_next[173] ;
 wire \board_state_next[174] ;
 wire \board_state_next[175] ;
 wire \board_state_next[176] ;
 wire \board_state_next[177] ;
 wire \board_state_next[178] ;
 wire \board_state_next[179] ;
 wire \board_state_next[17] ;
 wire \board_state_next[180] ;
 wire \board_state_next[181] ;
 wire \board_state_next[182] ;
 wire \board_state_next[183] ;
 wire \board_state_next[184] ;
 wire \board_state_next[185] ;
 wire \board_state_next[186] ;
 wire \board_state_next[187] ;
 wire \board_state_next[188] ;
 wire \board_state_next[189] ;
 wire \board_state_next[18] ;
 wire \board_state_next[190] ;
 wire \board_state_next[191] ;
 wire \board_state_next[192] ;
 wire \board_state_next[193] ;
 wire \board_state_next[194] ;
 wire \board_state_next[195] ;
 wire \board_state_next[196] ;
 wire \board_state_next[197] ;
 wire \board_state_next[198] ;
 wire \board_state_next[199] ;
 wire \board_state_next[19] ;
 wire \board_state_next[1] ;
 wire \board_state_next[200] ;
 wire \board_state_next[201] ;
 wire \board_state_next[202] ;
 wire \board_state_next[203] ;
 wire \board_state_next[204] ;
 wire \board_state_next[205] ;
 wire \board_state_next[206] ;
 wire \board_state_next[207] ;
 wire \board_state_next[208] ;
 wire \board_state_next[209] ;
 wire \board_state_next[20] ;
 wire \board_state_next[210] ;
 wire \board_state_next[211] ;
 wire \board_state_next[212] ;
 wire \board_state_next[213] ;
 wire \board_state_next[214] ;
 wire \board_state_next[215] ;
 wire \board_state_next[216] ;
 wire \board_state_next[217] ;
 wire \board_state_next[218] ;
 wire \board_state_next[219] ;
 wire \board_state_next[21] ;
 wire \board_state_next[220] ;
 wire \board_state_next[221] ;
 wire \board_state_next[222] ;
 wire \board_state_next[223] ;
 wire \board_state_next[224] ;
 wire \board_state_next[225] ;
 wire \board_state_next[226] ;
 wire \board_state_next[227] ;
 wire \board_state_next[228] ;
 wire \board_state_next[229] ;
 wire \board_state_next[22] ;
 wire \board_state_next[230] ;
 wire \board_state_next[231] ;
 wire \board_state_next[232] ;
 wire \board_state_next[233] ;
 wire \board_state_next[234] ;
 wire \board_state_next[235] ;
 wire \board_state_next[236] ;
 wire \board_state_next[237] ;
 wire \board_state_next[238] ;
 wire \board_state_next[239] ;
 wire \board_state_next[23] ;
 wire \board_state_next[240] ;
 wire \board_state_next[241] ;
 wire \board_state_next[242] ;
 wire \board_state_next[243] ;
 wire \board_state_next[244] ;
 wire \board_state_next[245] ;
 wire \board_state_next[246] ;
 wire \board_state_next[247] ;
 wire \board_state_next[248] ;
 wire \board_state_next[249] ;
 wire \board_state_next[24] ;
 wire \board_state_next[250] ;
 wire \board_state_next[251] ;
 wire \board_state_next[252] ;
 wire \board_state_next[253] ;
 wire \board_state_next[254] ;
 wire \board_state_next[255] ;
 wire \board_state_next[256] ;
 wire \board_state_next[257] ;
 wire \board_state_next[258] ;
 wire \board_state_next[259] ;
 wire \board_state_next[25] ;
 wire \board_state_next[260] ;
 wire \board_state_next[261] ;
 wire \board_state_next[262] ;
 wire \board_state_next[263] ;
 wire \board_state_next[264] ;
 wire \board_state_next[265] ;
 wire \board_state_next[266] ;
 wire \board_state_next[267] ;
 wire \board_state_next[268] ;
 wire \board_state_next[269] ;
 wire \board_state_next[26] ;
 wire \board_state_next[270] ;
 wire \board_state_next[271] ;
 wire \board_state_next[272] ;
 wire \board_state_next[273] ;
 wire \board_state_next[274] ;
 wire \board_state_next[275] ;
 wire \board_state_next[276] ;
 wire \board_state_next[277] ;
 wire \board_state_next[278] ;
 wire \board_state_next[279] ;
 wire \board_state_next[27] ;
 wire \board_state_next[280] ;
 wire \board_state_next[281] ;
 wire \board_state_next[282] ;
 wire \board_state_next[283] ;
 wire \board_state_next[284] ;
 wire \board_state_next[285] ;
 wire \board_state_next[286] ;
 wire \board_state_next[287] ;
 wire \board_state_next[288] ;
 wire \board_state_next[289] ;
 wire \board_state_next[28] ;
 wire \board_state_next[290] ;
 wire \board_state_next[291] ;
 wire \board_state_next[292] ;
 wire \board_state_next[293] ;
 wire \board_state_next[294] ;
 wire \board_state_next[295] ;
 wire \board_state_next[296] ;
 wire \board_state_next[297] ;
 wire \board_state_next[298] ;
 wire \board_state_next[299] ;
 wire \board_state_next[29] ;
 wire \board_state_next[2] ;
 wire \board_state_next[300] ;
 wire \board_state_next[301] ;
 wire \board_state_next[302] ;
 wire \board_state_next[303] ;
 wire \board_state_next[304] ;
 wire \board_state_next[305] ;
 wire \board_state_next[306] ;
 wire \board_state_next[307] ;
 wire \board_state_next[308] ;
 wire \board_state_next[309] ;
 wire \board_state_next[30] ;
 wire \board_state_next[310] ;
 wire \board_state_next[311] ;
 wire \board_state_next[312] ;
 wire \board_state_next[313] ;
 wire \board_state_next[314] ;
 wire \board_state_next[315] ;
 wire \board_state_next[316] ;
 wire \board_state_next[317] ;
 wire \board_state_next[318] ;
 wire \board_state_next[319] ;
 wire \board_state_next[31] ;
 wire \board_state_next[320] ;
 wire \board_state_next[321] ;
 wire \board_state_next[322] ;
 wire \board_state_next[323] ;
 wire \board_state_next[324] ;
 wire \board_state_next[325] ;
 wire \board_state_next[326] ;
 wire \board_state_next[327] ;
 wire \board_state_next[328] ;
 wire \board_state_next[329] ;
 wire \board_state_next[32] ;
 wire \board_state_next[330] ;
 wire \board_state_next[331] ;
 wire \board_state_next[332] ;
 wire \board_state_next[333] ;
 wire \board_state_next[334] ;
 wire \board_state_next[335] ;
 wire \board_state_next[336] ;
 wire \board_state_next[337] ;
 wire \board_state_next[338] ;
 wire \board_state_next[339] ;
 wire \board_state_next[33] ;
 wire \board_state_next[340] ;
 wire \board_state_next[341] ;
 wire \board_state_next[342] ;
 wire \board_state_next[343] ;
 wire \board_state_next[344] ;
 wire \board_state_next[345] ;
 wire \board_state_next[346] ;
 wire \board_state_next[347] ;
 wire \board_state_next[348] ;
 wire \board_state_next[349] ;
 wire \board_state_next[34] ;
 wire \board_state_next[350] ;
 wire \board_state_next[351] ;
 wire \board_state_next[352] ;
 wire \board_state_next[353] ;
 wire \board_state_next[354] ;
 wire \board_state_next[355] ;
 wire \board_state_next[356] ;
 wire \board_state_next[357] ;
 wire \board_state_next[358] ;
 wire \board_state_next[359] ;
 wire \board_state_next[35] ;
 wire \board_state_next[360] ;
 wire \board_state_next[361] ;
 wire \board_state_next[362] ;
 wire \board_state_next[363] ;
 wire \board_state_next[364] ;
 wire \board_state_next[365] ;
 wire \board_state_next[366] ;
 wire \board_state_next[367] ;
 wire \board_state_next[368] ;
 wire \board_state_next[369] ;
 wire \board_state_next[36] ;
 wire \board_state_next[370] ;
 wire \board_state_next[371] ;
 wire \board_state_next[372] ;
 wire \board_state_next[373] ;
 wire \board_state_next[374] ;
 wire \board_state_next[375] ;
 wire \board_state_next[376] ;
 wire \board_state_next[377] ;
 wire \board_state_next[378] ;
 wire \board_state_next[379] ;
 wire \board_state_next[37] ;
 wire \board_state_next[380] ;
 wire \board_state_next[381] ;
 wire \board_state_next[382] ;
 wire \board_state_next[383] ;
 wire \board_state_next[384] ;
 wire \board_state_next[385] ;
 wire \board_state_next[386] ;
 wire \board_state_next[387] ;
 wire \board_state_next[388] ;
 wire \board_state_next[389] ;
 wire \board_state_next[38] ;
 wire \board_state_next[390] ;
 wire \board_state_next[391] ;
 wire \board_state_next[392] ;
 wire \board_state_next[393] ;
 wire \board_state_next[394] ;
 wire \board_state_next[395] ;
 wire \board_state_next[396] ;
 wire \board_state_next[397] ;
 wire \board_state_next[398] ;
 wire \board_state_next[399] ;
 wire \board_state_next[39] ;
 wire \board_state_next[3] ;
 wire \board_state_next[400] ;
 wire \board_state_next[401] ;
 wire \board_state_next[402] ;
 wire \board_state_next[403] ;
 wire \board_state_next[404] ;
 wire \board_state_next[405] ;
 wire \board_state_next[406] ;
 wire \board_state_next[407] ;
 wire \board_state_next[408] ;
 wire \board_state_next[409] ;
 wire \board_state_next[40] ;
 wire \board_state_next[410] ;
 wire \board_state_next[411] ;
 wire \board_state_next[412] ;
 wire \board_state_next[413] ;
 wire \board_state_next[414] ;
 wire \board_state_next[415] ;
 wire \board_state_next[416] ;
 wire \board_state_next[417] ;
 wire \board_state_next[418] ;
 wire \board_state_next[419] ;
 wire \board_state_next[41] ;
 wire \board_state_next[420] ;
 wire \board_state_next[421] ;
 wire \board_state_next[422] ;
 wire \board_state_next[423] ;
 wire \board_state_next[424] ;
 wire \board_state_next[425] ;
 wire \board_state_next[426] ;
 wire \board_state_next[427] ;
 wire \board_state_next[428] ;
 wire \board_state_next[429] ;
 wire \board_state_next[42] ;
 wire \board_state_next[430] ;
 wire \board_state_next[431] ;
 wire \board_state_next[432] ;
 wire \board_state_next[433] ;
 wire \board_state_next[434] ;
 wire \board_state_next[435] ;
 wire \board_state_next[436] ;
 wire \board_state_next[437] ;
 wire \board_state_next[438] ;
 wire \board_state_next[439] ;
 wire \board_state_next[43] ;
 wire \board_state_next[440] ;
 wire \board_state_next[441] ;
 wire \board_state_next[442] ;
 wire \board_state_next[443] ;
 wire \board_state_next[444] ;
 wire \board_state_next[445] ;
 wire \board_state_next[446] ;
 wire \board_state_next[447] ;
 wire \board_state_next[448] ;
 wire \board_state_next[449] ;
 wire \board_state_next[44] ;
 wire \board_state_next[450] ;
 wire \board_state_next[451] ;
 wire \board_state_next[452] ;
 wire \board_state_next[453] ;
 wire \board_state_next[454] ;
 wire \board_state_next[455] ;
 wire \board_state_next[456] ;
 wire \board_state_next[457] ;
 wire \board_state_next[458] ;
 wire \board_state_next[459] ;
 wire \board_state_next[45] ;
 wire \board_state_next[460] ;
 wire \board_state_next[461] ;
 wire \board_state_next[462] ;
 wire \board_state_next[463] ;
 wire \board_state_next[464] ;
 wire \board_state_next[465] ;
 wire \board_state_next[466] ;
 wire \board_state_next[467] ;
 wire \board_state_next[468] ;
 wire \board_state_next[469] ;
 wire \board_state_next[46] ;
 wire \board_state_next[470] ;
 wire \board_state_next[471] ;
 wire \board_state_next[472] ;
 wire \board_state_next[473] ;
 wire \board_state_next[474] ;
 wire \board_state_next[475] ;
 wire \board_state_next[476] ;
 wire \board_state_next[477] ;
 wire \board_state_next[478] ;
 wire \board_state_next[479] ;
 wire \board_state_next[47] ;
 wire \board_state_next[480] ;
 wire \board_state_next[481] ;
 wire \board_state_next[482] ;
 wire \board_state_next[483] ;
 wire \board_state_next[484] ;
 wire \board_state_next[485] ;
 wire \board_state_next[486] ;
 wire \board_state_next[487] ;
 wire \board_state_next[488] ;
 wire \board_state_next[489] ;
 wire \board_state_next[48] ;
 wire \board_state_next[490] ;
 wire \board_state_next[491] ;
 wire \board_state_next[492] ;
 wire \board_state_next[493] ;
 wire \board_state_next[494] ;
 wire \board_state_next[495] ;
 wire \board_state_next[496] ;
 wire \board_state_next[497] ;
 wire \board_state_next[498] ;
 wire \board_state_next[499] ;
 wire \board_state_next[49] ;
 wire \board_state_next[4] ;
 wire \board_state_next[500] ;
 wire \board_state_next[501] ;
 wire \board_state_next[502] ;
 wire \board_state_next[503] ;
 wire \board_state_next[504] ;
 wire \board_state_next[505] ;
 wire \board_state_next[506] ;
 wire \board_state_next[507] ;
 wire \board_state_next[508] ;
 wire \board_state_next[509] ;
 wire \board_state_next[50] ;
 wire \board_state_next[510] ;
 wire \board_state_next[511] ;
 wire \board_state_next[51] ;
 wire \board_state_next[52] ;
 wire \board_state_next[53] ;
 wire \board_state_next[54] ;
 wire \board_state_next[55] ;
 wire \board_state_next[56] ;
 wire \board_state_next[57] ;
 wire \board_state_next[58] ;
 wire \board_state_next[59] ;
 wire \board_state_next[5] ;
 wire \board_state_next[60] ;
 wire \board_state_next[61] ;
 wire \board_state_next[62] ;
 wire \board_state_next[63] ;
 wire \board_state_next[64] ;
 wire \board_state_next[65] ;
 wire \board_state_next[66] ;
 wire \board_state_next[67] ;
 wire \board_state_next[68] ;
 wire \board_state_next[69] ;
 wire \board_state_next[6] ;
 wire \board_state_next[70] ;
 wire \board_state_next[71] ;
 wire \board_state_next[72] ;
 wire \board_state_next[73] ;
 wire \board_state_next[74] ;
 wire \board_state_next[75] ;
 wire \board_state_next[76] ;
 wire \board_state_next[77] ;
 wire \board_state_next[78] ;
 wire \board_state_next[79] ;
 wire \board_state_next[7] ;
 wire \board_state_next[80] ;
 wire \board_state_next[81] ;
 wire \board_state_next[82] ;
 wire \board_state_next[83] ;
 wire \board_state_next[84] ;
 wire \board_state_next[85] ;
 wire \board_state_next[86] ;
 wire \board_state_next[87] ;
 wire \board_state_next[88] ;
 wire \board_state_next[89] ;
 wire \board_state_next[8] ;
 wire \board_state_next[90] ;
 wire \board_state_next[91] ;
 wire \board_state_next[92] ;
 wire \board_state_next[93] ;
 wire \board_state_next[94] ;
 wire \board_state_next[95] ;
 wire \board_state_next[96] ;
 wire \board_state_next[97] ;
 wire \board_state_next[98] ;
 wire \board_state_next[99] ;
 wire \board_state_next[9] ;
 wire \cell_index[0] ;
 wire \cell_index[1] ;
 wire \cell_index[2] ;
 wire \cell_index[3] ;
 wire \cell_index[4] ;
 wire \cell_index[5] ;
 wire \cell_index[6] ;
 wire \cell_index[7] ;
 wire \cell_index[8] ;
 wire \cell_x[0] ;
 wire \cell_x[1] ;
 wire \cell_x[2] ;
 wire \cell_x[3] ;
 wire \cell_x[4] ;
 wire \cell_y[0] ;
 wire \cell_y[1] ;
 wire \cell_y[2] ;
 wire \cell_y[3] ;
 wire \colindex[0] ;
 wire \colindex[1] ;
 wire \colindex[2] ;
 wire \colindex[3] ;
 wire \colindex[4] ;
 wire \colindex[5] ;
 wire hsync;
 wire \hvsync_inst.hpos[0] ;
 wire \hvsync_inst.hpos[1] ;
 wire \hvsync_inst.hpos[2] ;
 wire \hvsync_inst.hpos[3] ;
 wire \hvsync_inst.hpos[9] ;
 wire \hvsync_inst.vpos[0] ;
 wire \hvsync_inst.vpos[1] ;
 wire \hvsync_inst.vpos[2] ;
 wire \hvsync_inst.vpos[3] ;
 wire \hvsync_inst.vpos[8] ;
 wire \hvsync_inst.vpos[9] ;
 wire \hvsync_inst.vsync ;
 wire \lfsr.lfsr_reg[0] ;
 wire \lfsr.lfsr_reg[10] ;
 wire \lfsr.lfsr_reg[11] ;
 wire \lfsr.lfsr_reg[12] ;
 wire \lfsr.lfsr_reg[13] ;
 wire \lfsr.lfsr_reg[14] ;
 wire \lfsr.lfsr_reg[15] ;
 wire \lfsr.lfsr_reg[1] ;
 wire \lfsr.lfsr_reg[2] ;
 wire \lfsr.lfsr_reg[3] ;
 wire \lfsr.lfsr_reg[4] ;
 wire \lfsr.lfsr_reg[5] ;
 wire \lfsr.lfsr_reg[6] ;
 wire \lfsr.lfsr_reg[7] ;
 wire \lfsr.lfsr_reg[8] ;
 wire \lfsr.lfsr_reg[9] ;
 wire \neigh_index[0] ;
 wire \neigh_index[1] ;
 wire \neigh_index[2] ;
 wire \neigh_index[3] ;
 wire \num_neighbors[0] ;
 wire \num_neighbors[1] ;
 wire \num_neighbors[2] ;
 wire \num_neighbors[3] ;
 wire running;
 wire \timer[0] ;
 wire \timer[10] ;
 wire \timer[11] ;
 wire \timer[12] ;
 wire \timer[13] ;
 wire \timer[14] ;
 wire \timer[15] ;
 wire \timer[16] ;
 wire \timer[17] ;
 wire \timer[18] ;
 wire \timer[19] ;
 wire \timer[1] ;
 wire \timer[20] ;
 wire \timer[21] ;
 wire \timer[22] ;
 wire \timer[23] ;
 wire \timer[24] ;
 wire \timer[25] ;
 wire \timer[26] ;
 wire \timer[27] ;
 wire \timer[28] ;
 wire \timer[29] ;
 wire \timer[2] ;
 wire \timer[30] ;
 wire \timer[31] ;
 wire \timer[3] ;
 wire \timer[4] ;
 wire \timer[5] ;
 wire \timer[6] ;
 wire \timer[7] ;
 wire \timer[8] ;
 wire \timer[9] ;
 wire \txindex[0] ;
 wire \txindex[1] ;
 wire \txindex[2] ;
 wire \txindex[3] ;
 wire \txindex[4] ;
 wire \txindex[5] ;
 wire \txstate[0] ;
 wire \txstate[2] ;
 wire \txstate[3] ;
 wire \txstate[4] ;
 wire \txstate[5] ;
 wire \txstate[6] ;
 wire \txstate[7] ;
 wire \txstate[8] ;
 wire \uart_rx_data[0] ;
 wire \uart_rx_data[1] ;
 wire \uart_rx_data[2] ;
 wire \uart_rx_data[3] ;
 wire \uart_rx_data[4] ;
 wire \uart_rx_data[5] ;
 wire \uart_rx_data[6] ;
 wire \uart_rx_data[7] ;
 wire \uart_rx_inst.bitIndex[0] ;
 wire \uart_rx_inst.bitIndex[1] ;
 wire \uart_rx_inst.bitIndex[2] ;
 wire \uart_rx_inst.data[0] ;
 wire \uart_rx_inst.data[1] ;
 wire \uart_rx_inst.data[2] ;
 wire \uart_rx_inst.data[3] ;
 wire \uart_rx_inst.data[4] ;
 wire \uart_rx_inst.data[5] ;
 wire \uart_rx_inst.data[6] ;
 wire \uart_rx_inst.data[7] ;
 wire \uart_rx_inst.inputReg[0] ;
 wire \uart_rx_inst.inputReg[1] ;
 wire \uart_rx_inst.inputReg[2] ;
 wire \uart_rx_inst.out_latched ;
 wire \uart_rx_inst.ready ;
 wire \uart_rx_inst.rxCounter[0] ;
 wire \uart_rx_inst.rxCounter[1] ;
 wire \uart_rx_inst.rxCounter[2] ;
 wire \uart_rx_inst.rxCounter[3] ;
 wire \uart_rx_inst.sampleCount[0] ;
 wire \uart_rx_inst.sampleCount[1] ;
 wire \uart_rx_inst.sampleCount[2] ;
 wire \uart_rx_inst.sampleCount[3] ;
 wire \uart_rx_inst.state[0] ;
 wire \uart_rx_inst.state[1] ;
 wire \uart_rx_inst.state[2] ;
 wire \uart_rx_inst.state[3] ;
 wire \uart_rx_inst.valid ;
 wire uart_tx;
 wire \uart_tx_data[0] ;
 wire \uart_tx_data[1] ;
 wire \uart_tx_data[2] ;
 wire \uart_tx_data[3] ;
 wire \uart_tx_data[4] ;
 wire \uart_tx_data[5] ;
 wire \uart_tx_data[6] ;
 wire \uart_tx_inst.bitIndex[0] ;
 wire \uart_tx_inst.bitIndex[1] ;
 wire \uart_tx_inst.bitIndex[2] ;
 wire \uart_tx_inst.data[0] ;
 wire \uart_tx_inst.data[1] ;
 wire \uart_tx_inst.data[2] ;
 wire \uart_tx_inst.data[3] ;
 wire \uart_tx_inst.data[4] ;
 wire \uart_tx_inst.data[5] ;
 wire \uart_tx_inst.data[6] ;
 wire \uart_tx_inst.ready ;
 wire \uart_tx_inst.state[0] ;
 wire \uart_tx_inst.state[1] ;
 wire \uart_tx_inst.state[2] ;
 wire \uart_tx_inst.state[3] ;
 wire \uart_tx_inst.txCounter[0] ;
 wire \uart_tx_inst.txCounter[1] ;
 wire \uart_tx_inst.txCounter[2] ;
 wire \uart_tx_inst.txCounter[3] ;
 wire \uart_tx_inst.txCounter[4] ;
 wire \uart_tx_inst.txCounter[5] ;
 wire \uart_tx_inst.txCounter[6] ;
 wire \uart_tx_inst.txCounter[7] ;
 wire \uart_tx_inst.valid ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _5421_ (.A(\txstate[2] ),
    .X(_1783_));
 sg13g2_nor2_1 _5422_ (.A(\hvsync_inst.vsync ),
    .B(_0055_),
    .Y(_1784_));
 sg13g2_buf_2 _5423_ (.A(\action[3] ),
    .X(_1785_));
 sg13g2_buf_1 _5424_ (.A(\action[2] ),
    .X(_1786_));
 sg13g2_nor2_1 _5425_ (.A(_1785_),
    .B(net400),
    .Y(_1787_));
 sg13g2_buf_1 _5426_ (.A(\action[6] ),
    .X(_1788_));
 sg13g2_buf_1 _5427_ (.A(\action[7] ),
    .X(_1789_));
 sg13g2_buf_1 _5428_ (.A(_1789_),
    .X(_1790_));
 sg13g2_nor2_2 _5429_ (.A(_1788_),
    .B(net382),
    .Y(_1791_));
 sg13g2_and2_1 _5430_ (.A(_1787_),
    .B(_1791_),
    .X(_1792_));
 sg13g2_buf_1 _5431_ (.A(net1),
    .X(_1793_));
 sg13g2_o21ai_1 _5432_ (.B1(net401),
    .Y(_1794_),
    .A1(_1784_),
    .A2(_1792_));
 sg13g2_buf_1 _5433_ (.A(_1788_),
    .X(_1795_));
 sg13g2_buf_1 _5434_ (.A(net401),
    .X(_1796_));
 sg13g2_nand2_1 _5435_ (.Y(_1797_),
    .A(net381),
    .B(net399));
 sg13g2_buf_1 _5436_ (.A(net399),
    .X(_1798_));
 sg13g2_buf_1 _5437_ (.A(\uart_tx_inst.valid ),
    .X(_1799_));
 sg13g2_buf_1 _5438_ (.A(\uart_tx_inst.ready ),
    .X(_1800_));
 sg13g2_nand2b_1 _5439_ (.Y(_1801_),
    .B(net397),
    .A_N(net398));
 sg13g2_nand2b_1 _5440_ (.Y(_1802_),
    .B(net398),
    .A_N(net397));
 sg13g2_nand4_1 _5441_ (.B(net382),
    .C(_1801_),
    .A(net380),
    .Y(_1803_),
    .D(_1802_));
 sg13g2_and2_1 _5442_ (.A(_1785_),
    .B(\hvsync_inst.vsync ),
    .X(_1804_));
 sg13g2_o21ai_1 _5443_ (.B1(net399),
    .Y(_1805_),
    .A1(net400),
    .A2(_1804_));
 sg13g2_buf_1 _5444_ (.A(_0054_),
    .X(_1806_));
 sg13g2_buf_1 _5445_ (.A(\cell_x[4] ),
    .X(_1807_));
 sg13g2_buf_2 _5446_ (.A(\cell_x[3] ),
    .X(_1808_));
 sg13g2_buf_1 _5447_ (.A(_1808_),
    .X(_1809_));
 sg13g2_nand2_2 _5448_ (.Y(_1810_),
    .A(_1807_),
    .B(_1809_));
 sg13g2_buf_2 _5449_ (.A(\cell_x[2] ),
    .X(_1811_));
 sg13g2_buf_1 _5450_ (.A(_1811_),
    .X(_1812_));
 sg13g2_buf_1 _5451_ (.A(net378),
    .X(_1813_));
 sg13g2_buf_2 _5452_ (.A(\cell_x[1] ),
    .X(_1814_));
 sg13g2_buf_1 _5453_ (.A(_1814_),
    .X(_1815_));
 sg13g2_buf_1 _5454_ (.A(net377),
    .X(_1816_));
 sg13g2_buf_1 _5455_ (.A(_1816_),
    .X(_1817_));
 sg13g2_nand2_1 _5456_ (.Y(_1818_),
    .A(_1813_),
    .B(net276));
 sg13g2_buf_1 _5457_ (.A(\cell_y[2] ),
    .X(_1819_));
 sg13g2_buf_1 _5458_ (.A(\cell_y[3] ),
    .X(_1820_));
 sg13g2_buf_1 _5459_ (.A(\cell_y[1] ),
    .X(_1821_));
 sg13g2_buf_1 _5460_ (.A(_1821_),
    .X(_1822_));
 sg13g2_buf_1 _5461_ (.A(\cell_y[0] ),
    .X(_1823_));
 sg13g2_buf_1 _5462_ (.A(net393),
    .X(_1824_));
 sg13g2_nand4_1 _5463_ (.B(_1820_),
    .C(net376),
    .A(_1819_),
    .Y(_1825_),
    .D(net375));
 sg13g2_or4_1 _5464_ (.A(net396),
    .B(_1810_),
    .C(_1818_),
    .D(_1825_),
    .X(_1826_));
 sg13g2_buf_2 _5465_ (.A(_1826_),
    .X(_1827_));
 sg13g2_nand2b_1 _5466_ (.Y(_1828_),
    .B(_1827_),
    .A_N(_1805_));
 sg13g2_nand4_1 _5467_ (.B(_1797_),
    .C(_1803_),
    .A(_1794_),
    .Y(_1829_),
    .D(_1828_));
 sg13g2_inv_1 _5468_ (.Y(_1830_),
    .A(net401));
 sg13g2_buf_1 _5469_ (.A(_1830_),
    .X(_1831_));
 sg13g2_buf_1 _5470_ (.A(net374),
    .X(_1832_));
 sg13g2_buf_1 _5471_ (.A(\txstate[0] ),
    .X(_1833_));
 sg13g2_buf_1 _5472_ (.A(\txindex[1] ),
    .X(_1834_));
 sg13g2_buf_1 _5473_ (.A(\txindex[0] ),
    .X(_1835_));
 sg13g2_nor2b_1 _5474_ (.A(net392),
    .B_N(net391),
    .Y(_1836_));
 sg13g2_buf_1 _5475_ (.A(\txindex[2] ),
    .X(_1837_));
 sg13g2_nand2b_1 _5476_ (.Y(_1838_),
    .B(_0056_),
    .A_N(_1837_));
 sg13g2_buf_1 _5477_ (.A(\txindex[5] ),
    .X(_1839_));
 sg13g2_buf_1 _5478_ (.A(\txindex[4] ),
    .X(_1840_));
 sg13g2_buf_1 _5479_ (.A(\txindex[3] ),
    .X(_1841_));
 sg13g2_and3_1 _5480_ (.X(_1842_),
    .A(_1839_),
    .B(_1840_),
    .C(_1841_));
 sg13g2_o21ai_1 _5481_ (.B1(_1842_),
    .Y(_1843_),
    .A1(_1836_),
    .A2(_1838_));
 sg13g2_buf_1 _5482_ (.A(_1843_),
    .X(_1844_));
 sg13g2_nor2b_1 _5483_ (.A(net398),
    .B_N(net397),
    .Y(_1845_));
 sg13g2_a22oi_1 _5484_ (.Y(_1846_),
    .B1(_1845_),
    .B2(_1783_),
    .A2(_1844_),
    .A1(_1833_));
 sg13g2_nor3_1 _5485_ (.A(net330),
    .B(_0053_),
    .C(_1846_),
    .Y(_1847_));
 sg13g2_a21o_1 _5486_ (.A2(_1829_),
    .A1(_1783_),
    .B1(_1847_),
    .X(_0029_));
 sg13g2_buf_1 _5487_ (.A(\uart_tx_inst.txCounter[1] ),
    .X(_1848_));
 sg13g2_buf_2 _5488_ (.A(\uart_tx_inst.txCounter[0] ),
    .X(_1849_));
 sg13g2_nand4_1 _5489_ (.B(\uart_tx_inst.txCounter[2] ),
    .C(_1848_),
    .A(\uart_tx_inst.txCounter[3] ),
    .Y(_1850_),
    .D(_1849_));
 sg13g2_buf_1 _5490_ (.A(_1850_),
    .X(_1851_));
 sg13g2_nor2_1 _5491_ (.A(\uart_tx_inst.txCounter[5] ),
    .B(\uart_tx_inst.txCounter[4] ),
    .Y(_1852_));
 sg13g2_nand2_1 _5492_ (.Y(_1853_),
    .A(\uart_tx_inst.txCounter[7] ),
    .B(\uart_tx_inst.txCounter[6] ));
 sg13g2_a21oi_1 _5493_ (.A1(_1851_),
    .A2(_1852_),
    .Y(_1854_),
    .B1(_1853_));
 sg13g2_buf_1 _5494_ (.A(_1854_),
    .X(_1855_));
 sg13g2_nand2_1 _5495_ (.Y(_1856_),
    .A(net397),
    .B(_1799_));
 sg13g2_buf_2 _5496_ (.A(_1856_),
    .X(_1857_));
 sg13g2_nand2_1 _5497_ (.Y(_1858_),
    .A(net401),
    .B(_1857_));
 sg13g2_nor2_1 _5498_ (.A(net262),
    .B(_1858_),
    .Y(_1859_));
 sg13g2_nor2_1 _5499_ (.A(net374),
    .B(_1857_),
    .Y(_1860_));
 sg13g2_buf_1 _5500_ (.A(_1860_),
    .X(_1861_));
 sg13g2_a21o_1 _5501_ (.A2(_1859_),
    .A1(\uart_tx_inst.state[2] ),
    .B1(_1861_),
    .X(_0042_));
 sg13g2_buf_2 _5502_ (.A(\uart_tx_inst.bitIndex[1] ),
    .X(_1862_));
 sg13g2_buf_1 _5503_ (.A(\uart_tx_inst.bitIndex[0] ),
    .X(_1863_));
 sg13g2_nand2_1 _5504_ (.Y(_1864_),
    .A(_1862_),
    .B(net390));
 sg13g2_nor2_1 _5505_ (.A(_0057_),
    .B(_1864_),
    .Y(_1865_));
 sg13g2_nand2_1 _5506_ (.Y(_1866_),
    .A(net262),
    .B(_1865_));
 sg13g2_buf_1 _5507_ (.A(\uart_tx_inst.state[1] ),
    .X(_1867_));
 sg13g2_a22oi_1 _5508_ (.Y(_1868_),
    .B1(_1866_),
    .B2(_1867_),
    .A2(_1855_),
    .A1(\uart_tx_inst.state[2] ));
 sg13g2_nor2_1 _5509_ (.A(_1858_),
    .B(_1868_),
    .Y(_0041_));
 sg13g2_buf_1 _5510_ (.A(net330),
    .X(_1869_));
 sg13g2_buf_2 _5511_ (.A(\uart_rx_inst.state[1] ),
    .X(_1870_));
 sg13g2_buf_1 _5512_ (.A(_1870_),
    .X(_1871_));
 sg13g2_buf_1 _5513_ (.A(\uart_rx_inst.sampleCount[3] ),
    .X(_1872_));
 sg13g2_buf_2 _5514_ (.A(\uart_rx_inst.sampleCount[2] ),
    .X(_1873_));
 sg13g2_buf_2 _5515_ (.A(\uart_rx_inst.sampleCount[1] ),
    .X(_1874_));
 sg13g2_buf_1 _5516_ (.A(\uart_rx_inst.sampleCount[0] ),
    .X(_1875_));
 sg13g2_nand4_1 _5517_ (.B(_1873_),
    .C(_1874_),
    .A(_1872_),
    .Y(_1876_),
    .D(net389));
 sg13g2_buf_1 _5518_ (.A(_1876_),
    .X(_1877_));
 sg13g2_buf_1 _5519_ (.A(\uart_rx_inst.rxCounter[2] ),
    .X(_1878_));
 sg13g2_nand2_1 _5520_ (.Y(_1879_),
    .A(\uart_rx_inst.rxCounter[3] ),
    .B(_1878_));
 sg13g2_buf_1 _5521_ (.A(_1879_),
    .X(_1880_));
 sg13g2_buf_1 _5522_ (.A(\uart_rx_inst.bitIndex[1] ),
    .X(_1881_));
 sg13g2_buf_2 _5523_ (.A(\uart_rx_inst.bitIndex[0] ),
    .X(_1882_));
 sg13g2_nand2_1 _5524_ (.Y(_1883_),
    .A(_1881_),
    .B(_1882_));
 sg13g2_or4_1 _5525_ (.A(_0059_),
    .B(_1877_),
    .C(_1880_),
    .D(_1883_),
    .X(_1884_));
 sg13g2_o21ai_1 _5526_ (.B1(_1873_),
    .Y(_1885_),
    .A1(_1874_),
    .A2(net389));
 sg13g2_nand2b_1 _5527_ (.Y(_1886_),
    .B(_1885_),
    .A_N(_1872_));
 sg13g2_buf_1 _5528_ (.A(\uart_rx_inst.state[2] ),
    .X(_1887_));
 sg13g2_inv_1 _5529_ (.Y(_1888_),
    .A(_1887_));
 sg13g2_buf_1 _5530_ (.A(_1880_),
    .X(_1889_));
 sg13g2_nor2_1 _5531_ (.A(_1888_),
    .B(net274),
    .Y(_1890_));
 sg13g2_a22oi_1 _5532_ (.Y(_1891_),
    .B1(_1886_),
    .B2(_1890_),
    .A2(_1884_),
    .A1(net373));
 sg13g2_nor2_1 _5533_ (.A(_1869_),
    .B(_1891_),
    .Y(_0037_));
 sg13g2_inv_1 _5534_ (.Y(_1892_),
    .A(net381));
 sg13g2_or2_1 _5535_ (.X(_1893_),
    .B(net398),
    .A(net397));
 sg13g2_nand2_1 _5536_ (.Y(_1894_),
    .A(net398),
    .B(_1892_));
 sg13g2_nand2b_1 _5537_ (.Y(_1895_),
    .B(_0058_),
    .A_N(net398));
 sg13g2_nand3_1 _5538_ (.B(_1894_),
    .C(_1895_),
    .A(net397),
    .Y(_1896_));
 sg13g2_o21ai_1 _5539_ (.B1(_1896_),
    .Y(_1897_),
    .A1(_1892_),
    .A2(_1893_));
 sg13g2_nand2_1 _5540_ (.Y(_1898_),
    .A(net401),
    .B(net382));
 sg13g2_nand3_1 _5541_ (.B(_1804_),
    .C(_1827_),
    .A(net401),
    .Y(_1899_));
 sg13g2_nand3_1 _5542_ (.B(_1898_),
    .C(_1899_),
    .A(_1794_),
    .Y(_1900_));
 sg13g2_a21o_1 _5543_ (.A2(_1897_),
    .A1(net399),
    .B1(_1900_),
    .X(_1901_));
 sg13g2_nand3_1 _5544_ (.B(_1786_),
    .C(_1827_),
    .A(net399),
    .Y(_1902_));
 sg13g2_buf_1 _5545_ (.A(_1902_),
    .X(_1903_));
 sg13g2_nand2b_1 _5546_ (.Y(_1904_),
    .B(_1903_),
    .A_N(_1901_));
 sg13g2_nand2_1 _5547_ (.Y(_1905_),
    .A(\txstate[3] ),
    .B(_1904_));
 sg13g2_buf_2 _5548_ (.A(\txstate[8] ),
    .X(_1906_));
 sg13g2_or4_1 _5549_ (.A(_1839_),
    .B(_1840_),
    .C(_1841_),
    .D(_1837_),
    .X(_1907_));
 sg13g2_buf_1 _5550_ (.A(_1907_),
    .X(_1908_));
 sg13g2_nor2_1 _5551_ (.A(net392),
    .B(_1908_),
    .Y(_1909_));
 sg13g2_nor2_1 _5552_ (.A(net374),
    .B(_0058_),
    .Y(_1910_));
 sg13g2_nand3_1 _5553_ (.B(_1909_),
    .C(_1910_),
    .A(_1906_),
    .Y(_1911_));
 sg13g2_nand2_1 _5554_ (.Y(_0030_),
    .A(_1905_),
    .B(_1911_));
 sg13g2_buf_1 _5555_ (.A(net399),
    .X(_1912_));
 sg13g2_buf_1 _5556_ (.A(net372),
    .X(_1913_));
 sg13g2_buf_1 _5557_ (.A(\uart_rx_inst.state[0] ),
    .X(_1914_));
 sg13g2_and2_1 _5558_ (.A(\uart_rx_inst.rxCounter[3] ),
    .B(_1878_),
    .X(_1915_));
 sg13g2_buf_2 _5559_ (.A(_1915_),
    .X(_1916_));
 sg13g2_buf_2 _5560_ (.A(\uart_rx_inst.state[3] ),
    .X(_1917_));
 sg13g2_inv_1 _5561_ (.Y(_1918_),
    .A(_1877_));
 sg13g2_buf_1 _5562_ (.A(\uart_rx_inst.inputReg[1] ),
    .X(_1919_));
 sg13g2_buf_1 _5563_ (.A(\uart_rx_inst.inputReg[0] ),
    .X(_1920_));
 sg13g2_buf_1 _5564_ (.A(\uart_rx_inst.inputReg[2] ),
    .X(_1921_));
 sg13g2_nand3_1 _5565_ (.B(_1920_),
    .C(_1921_),
    .A(_1919_),
    .Y(_1922_));
 sg13g2_nand3_1 _5566_ (.B(_1918_),
    .C(_1922_),
    .A(_1917_),
    .Y(_1923_));
 sg13g2_or3_1 _5567_ (.A(_1873_),
    .B(_1874_),
    .C(net389),
    .X(_1924_));
 sg13g2_buf_1 _5568_ (.A(_1924_),
    .X(_1925_));
 sg13g2_nand2b_1 _5569_ (.Y(_1926_),
    .B(_1887_),
    .A_N(_1872_));
 sg13g2_nor3_1 _5570_ (.A(_1919_),
    .B(_1920_),
    .C(_1921_),
    .Y(_1927_));
 sg13g2_nor2_1 _5571_ (.A(_1926_),
    .B(_1927_),
    .Y(_1928_));
 sg13g2_nand3_1 _5572_ (.B(_1925_),
    .C(_1928_),
    .A(_1885_),
    .Y(_1929_));
 sg13g2_nand3_1 _5573_ (.B(_1923_),
    .C(_1929_),
    .A(_1916_),
    .Y(_1930_));
 sg13g2_o21ai_1 _5574_ (.B1(_1930_),
    .Y(_1931_),
    .A1(_1914_),
    .A2(_1916_));
 sg13g2_nand2_1 _5575_ (.Y(_0036_),
    .A(net329),
    .B(_1931_));
 sg13g2_inv_1 _5576_ (.Y(_1932_),
    .A(net3));
 sg13g2_buf_2 _5577_ (.A(\action[1] ),
    .X(_1933_));
 sg13g2_nand2_1 _5578_ (.Y(_1934_),
    .A(net380),
    .B(_1933_));
 sg13g2_buf_2 _5579_ (.A(\uart_rx_inst.valid ),
    .X(_1935_));
 sg13g2_buf_1 _5580_ (.A(running),
    .X(_1936_));
 sg13g2_inv_1 _5581_ (.Y(_1937_),
    .A(_1936_));
 sg13g2_buf_1 _5582_ (.A(\timer[22] ),
    .X(_1938_));
 sg13g2_buf_1 _5583_ (.A(\timer[19] ),
    .X(_1939_));
 sg13g2_inv_1 _5584_ (.Y(_1940_),
    .A(\timer[16] ));
 sg13g2_buf_1 _5585_ (.A(\timer[15] ),
    .X(_1941_));
 sg13g2_buf_1 _5586_ (.A(\timer[14] ),
    .X(_1942_));
 sg13g2_buf_1 _5587_ (.A(\timer[10] ),
    .X(_1943_));
 sg13g2_and4_1 _5588_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .C(\timer[11] ),
    .D(_1943_),
    .X(_1944_));
 sg13g2_nor2b_1 _5589_ (.A(_0060_),
    .B_N(_1944_),
    .Y(_1945_));
 sg13g2_nor3_1 _5590_ (.A(_1941_),
    .B(_1942_),
    .C(_1945_),
    .Y(_1946_));
 sg13g2_buf_1 _5591_ (.A(\timer[17] ),
    .X(_1947_));
 sg13g2_nor2_1 _5592_ (.A(\timer[18] ),
    .B(_1947_),
    .Y(_1948_));
 sg13g2_o21ai_1 _5593_ (.B1(_1948_),
    .Y(_1949_),
    .A1(_1940_),
    .A2(_1946_));
 sg13g2_buf_1 _5594_ (.A(\timer[20] ),
    .X(_1950_));
 sg13g2_or2_1 _5595_ (.X(_1951_),
    .B(_1950_),
    .A(\timer[21] ));
 sg13g2_a21o_1 _5596_ (.A2(_1949_),
    .A1(_1939_),
    .B1(_1951_),
    .X(_1952_));
 sg13g2_buf_1 _5597_ (.A(\timer[9] ),
    .X(_1953_));
 sg13g2_and2_1 _5598_ (.A(_1953_),
    .B(_1944_),
    .X(_1954_));
 sg13g2_buf_1 _5599_ (.A(_1954_),
    .X(_1955_));
 sg13g2_nor4_1 _5600_ (.A(\timer[18] ),
    .B(_1947_),
    .C(_1941_),
    .D(_1942_),
    .Y(_1956_));
 sg13g2_buf_1 _5601_ (.A(\timer[3] ),
    .X(_1957_));
 sg13g2_nor3_1 _5602_ (.A(\timer[8] ),
    .B(_1957_),
    .C(_1951_),
    .Y(_1958_));
 sg13g2_buf_1 _5603_ (.A(\timer[7] ),
    .X(_1959_));
 sg13g2_buf_1 _5604_ (.A(\timer[4] ),
    .X(_1960_));
 sg13g2_nor4_1 _5605_ (.A(_1959_),
    .B(\timer[6] ),
    .C(\timer[5] ),
    .D(_1960_),
    .Y(_1961_));
 sg13g2_buf_1 _5606_ (.A(\timer[2] ),
    .X(_1962_));
 sg13g2_buf_1 _5607_ (.A(\timer[1] ),
    .X(_1963_));
 sg13g2_buf_2 _5608_ (.A(\timer[0] ),
    .X(_1964_));
 sg13g2_nor4_1 _5609_ (.A(_1940_),
    .B(_1962_),
    .C(_1963_),
    .D(_1964_),
    .Y(_1965_));
 sg13g2_buf_1 _5610_ (.A(\timer[23] ),
    .X(_1966_));
 sg13g2_nor2b_1 _5611_ (.A(_1966_),
    .B_N(_1938_),
    .Y(_1967_));
 sg13g2_and4_1 _5612_ (.A(_1939_),
    .B(_1961_),
    .C(_1965_),
    .D(_1967_),
    .X(_1968_));
 sg13g2_nand4_1 _5613_ (.B(_1956_),
    .C(_1958_),
    .A(_1955_),
    .Y(_1969_),
    .D(_1968_));
 sg13g2_nor2_1 _5614_ (.A(\timer[31] ),
    .B(\timer[30] ),
    .Y(_1970_));
 sg13g2_nor4_1 _5615_ (.A(\timer[26] ),
    .B(\timer[25] ),
    .C(\timer[24] ),
    .D(_1966_),
    .Y(_1971_));
 sg13g2_nor3_1 _5616_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .C(\timer[27] ),
    .Y(_1972_));
 sg13g2_nand4_1 _5617_ (.B(_1970_),
    .C(_1971_),
    .A(_1969_),
    .Y(_1973_),
    .D(_1972_));
 sg13g2_a21oi_1 _5618_ (.A1(_1938_),
    .A2(_1952_),
    .Y(_1974_),
    .B1(_1973_));
 sg13g2_nor3_1 _5619_ (.A(_1935_),
    .B(_1937_),
    .C(_1974_),
    .Y(_1975_));
 sg13g2_nand2b_1 _5620_ (.Y(_1976_),
    .B(_1975_),
    .A_N(_1934_));
 sg13g2_or2_1 _5621_ (.X(_1977_),
    .B(\uart_rx_data[3] ),
    .A(\uart_rx_data[1] ));
 sg13g2_nand2b_1 _5622_ (.Y(_1978_),
    .B(\uart_rx_data[5] ),
    .A_N(\uart_rx_data[2] ));
 sg13g2_nor4_2 _5623_ (.A(\uart_rx_data[7] ),
    .B(\uart_rx_data[6] ),
    .C(_1977_),
    .Y(_1979_),
    .D(_1978_));
 sg13g2_buf_1 _5624_ (.A(\uart_rx_inst.ready ),
    .X(_1980_));
 sg13g2_nand2_1 _5625_ (.Y(_1981_),
    .A(_1980_),
    .B(_1935_));
 sg13g2_inv_1 _5626_ (.Y(_1982_),
    .A(_1981_));
 sg13g2_and4_1 _5627_ (.A(net399),
    .B(_1933_),
    .C(_1979_),
    .D(_1982_),
    .X(_1983_));
 sg13g2_buf_1 _5628_ (.A(_1983_),
    .X(_1984_));
 sg13g2_buf_1 _5629_ (.A(\uart_rx_data[0] ),
    .X(_1985_));
 sg13g2_buf_1 _5630_ (.A(\uart_rx_data[4] ),
    .X(_1986_));
 sg13g2_nor2b_1 _5631_ (.A(_1985_),
    .B_N(_1986_),
    .Y(_1987_));
 sg13g2_and3_1 _5632_ (.X(_1988_),
    .A(net380),
    .B(net400),
    .C(_1827_));
 sg13g2_a21oi_1 _5633_ (.A1(_1984_),
    .A2(_1987_),
    .Y(_1989_),
    .B1(_1988_));
 sg13g2_o21ai_1 _5634_ (.B1(_1989_),
    .Y(_0022_),
    .A1(_1932_),
    .A2(_1976_));
 sg13g2_buf_1 _5635_ (.A(\action[4] ),
    .X(_1990_));
 sg13g2_nor4_2 _5636_ (.A(net396),
    .B(_1810_),
    .C(_1818_),
    .Y(_1991_),
    .D(_1825_));
 sg13g2_inv_1 _5637_ (.Y(_1992_),
    .A(_1844_));
 sg13g2_o21ai_1 _5638_ (.B1(_1833_),
    .Y(_1993_),
    .A1(_0061_),
    .A2(_1992_));
 sg13g2_buf_1 _5639_ (.A(_1790_),
    .X(_1994_));
 sg13g2_a22oi_1 _5640_ (.Y(_1995_),
    .B1(_1993_),
    .B2(net328),
    .A2(_1991_),
    .A1(_1990_));
 sg13g2_nor2_1 _5641_ (.A(net275),
    .B(_1995_),
    .Y(_0027_));
 sg13g2_buf_1 _5642_ (.A(\colindex[5] ),
    .X(_1996_));
 sg13g2_inv_1 _5643_ (.Y(_1997_),
    .A(_1996_));
 sg13g2_buf_1 _5644_ (.A(\txstate[6] ),
    .X(_1998_));
 sg13g2_and2_1 _5645_ (.A(_1998_),
    .B(_1910_),
    .X(_1999_));
 sg13g2_nand2_1 _5646_ (.Y(_2000_),
    .A(_1997_),
    .B(_1999_));
 sg13g2_o21ai_1 _5647_ (.B1(_2000_),
    .Y(_2001_),
    .A1(_0063_),
    .A2(_1903_));
 sg13g2_a21o_1 _5648_ (.A2(_1901_),
    .A1(\txstate[4] ),
    .B1(_2001_),
    .X(_0031_));
 sg13g2_nand2b_1 _5649_ (.Y(_2002_),
    .B(_1988_),
    .A_N(_0061_));
 sg13g2_nor2b_1 _5650_ (.A(net397),
    .B_N(net398),
    .Y(_2003_));
 sg13g2_nand3_1 _5651_ (.B(_1783_),
    .C(_2003_),
    .A(net328),
    .Y(_2004_));
 sg13g2_nand2_1 _5652_ (.Y(_2005_),
    .A(_1794_),
    .B(_1899_));
 sg13g2_o21ai_1 _5653_ (.B1(_1833_),
    .Y(_2006_),
    .A1(net381),
    .A2(_2005_));
 sg13g2_nand4_1 _5654_ (.B(_2002_),
    .C(_2004_),
    .A(net329),
    .Y(_0028_),
    .D(_2006_));
 sg13g2_inv_1 _5655_ (.Y(_2007_),
    .A(\hvsync_inst.vsync ));
 sg13g2_inv_1 _5656_ (.Y(_2008_),
    .A(_0055_));
 sg13g2_nand2_1 _5657_ (.Y(_2009_),
    .A(_2007_),
    .B(_2008_));
 sg13g2_nor2b_1 _5658_ (.A(_0064_),
    .B_N(_1785_),
    .Y(_2010_));
 sg13g2_buf_1 _5659_ (.A(\action[5] ),
    .X(_2011_));
 sg13g2_buf_2 _5660_ (.A(\neigh_index[3] ),
    .X(_2012_));
 sg13g2_buf_1 _5661_ (.A(_2012_),
    .X(_2013_));
 sg13g2_buf_1 _5662_ (.A(\neigh_index[2] ),
    .X(_2014_));
 sg13g2_buf_1 _5663_ (.A(_2014_),
    .X(_2015_));
 sg13g2_buf_1 _5664_ (.A(net370),
    .X(_2016_));
 sg13g2_buf_1 _5665_ (.A(\neigh_index[0] ),
    .X(_2017_));
 sg13g2_buf_1 _5666_ (.A(\neigh_index[1] ),
    .X(_2018_));
 sg13g2_or2_1 _5667_ (.X(_2019_),
    .B(net386),
    .A(_2017_));
 sg13g2_buf_1 _5668_ (.A(_2019_),
    .X(_2020_));
 sg13g2_nor2_1 _5669_ (.A(net327),
    .B(_2020_),
    .Y(_2021_));
 sg13g2_nand3_1 _5670_ (.B(net371),
    .C(_2021_),
    .A(net387),
    .Y(_2022_));
 sg13g2_nand2_1 _5671_ (.Y(_2023_),
    .A(_1991_),
    .B(_2022_));
 sg13g2_o21ai_1 _5672_ (.B1(_2023_),
    .Y(_2024_),
    .A1(_1991_),
    .A2(_2010_));
 sg13g2_buf_1 _5673_ (.A(net330),
    .X(_2025_));
 sg13g2_a21oi_1 _5674_ (.A1(_2009_),
    .A2(_2024_),
    .Y(_0023_),
    .B1(net273));
 sg13g2_inv_1 _5675_ (.Y(_2026_),
    .A(\txstate[4] ));
 sg13g2_buf_1 _5676_ (.A(\cell_x[0] ),
    .X(_2027_));
 sg13g2_buf_8 _5677_ (.A(_2027_),
    .X(_2028_));
 sg13g2_nor4_2 _5678_ (.A(_1808_),
    .B(_1811_),
    .C(_1814_),
    .Y(_2029_),
    .D(_2028_));
 sg13g2_nor2_1 _5679_ (.A(net393),
    .B(net395),
    .Y(_2030_));
 sg13g2_buf_1 _5680_ (.A(_2030_),
    .X(_2031_));
 sg13g2_nor2_2 _5681_ (.A(net394),
    .B(_1821_),
    .Y(_2032_));
 sg13g2_nand4_1 _5682_ (.B(_2029_),
    .C(net326),
    .A(_0065_),
    .Y(_2033_),
    .D(_2032_));
 sg13g2_nand2b_1 _5683_ (.Y(_2034_),
    .B(_2033_),
    .A_N(_0063_));
 sg13g2_a22oi_1 _5684_ (.Y(_2035_),
    .B1(_2003_),
    .B2(_2034_),
    .A2(_1845_),
    .A1(_0063_));
 sg13g2_o21ai_1 _5685_ (.B1(_1795_),
    .Y(_2036_),
    .A1(_2026_),
    .A2(_2035_));
 sg13g2_o21ai_1 _5686_ (.B1(_1991_),
    .Y(_2037_),
    .A1(net400),
    .A2(_2010_));
 sg13g2_buf_1 _5687_ (.A(net330),
    .X(_2038_));
 sg13g2_a21oi_1 _5688_ (.A1(_2036_),
    .A2(_2037_),
    .Y(_0026_),
    .B1(net272));
 sg13g2_a22oi_1 _5689_ (.Y(_2039_),
    .B1(_1982_),
    .B2(\action[0] ),
    .A2(_1827_),
    .A1(_1990_));
 sg13g2_nor2_1 _5690_ (.A(net275),
    .B(_2039_),
    .Y(_0024_));
 sg13g2_buf_2 _5691_ (.A(\txstate[7] ),
    .X(_2040_));
 sg13g2_nor4_1 _5692_ (.A(_1839_),
    .B(_1840_),
    .C(_1841_),
    .D(_1837_),
    .Y(_2041_));
 sg13g2_and2_1 _5693_ (.A(_2040_),
    .B(_2041_),
    .X(_2042_));
 sg13g2_buf_2 _5694_ (.A(_2042_),
    .X(_2043_));
 sg13g2_a22oi_1 _5695_ (.Y(_2044_),
    .B1(_1910_),
    .B2(_2043_),
    .A2(_1904_),
    .A1(\txstate[5] ));
 sg13g2_inv_1 _5696_ (.Y(_0032_),
    .A(_2044_));
 sg13g2_nor2_1 _5697_ (.A(_1797_),
    .B(_1802_),
    .Y(_2045_));
 sg13g2_a22oi_1 _5698_ (.Y(_2046_),
    .B1(_2045_),
    .B2(\txstate[3] ),
    .A2(_1999_),
    .A1(_1996_));
 sg13g2_o21ai_1 _5699_ (.B1(_2046_),
    .Y(_2047_),
    .A1(_0066_),
    .A2(_1903_));
 sg13g2_a21o_1 _5700_ (.A2(_1900_),
    .A1(_1906_),
    .B1(_2047_),
    .X(_0035_));
 sg13g2_a21oi_1 _5701_ (.A1(_2040_),
    .A2(_1908_),
    .Y(_2048_),
    .B1(_1906_));
 sg13g2_nand3_1 _5702_ (.B(_2003_),
    .C(_2033_),
    .A(\txstate[4] ),
    .Y(_2049_));
 sg13g2_o21ai_1 _5703_ (.B1(_2049_),
    .Y(_2050_),
    .A1(_1909_),
    .A2(_2048_));
 sg13g2_nand2b_1 _5704_ (.Y(_2051_),
    .B(_1903_),
    .A_N(_1900_));
 sg13g2_a22oi_1 _5705_ (.Y(_2052_),
    .B1(_2051_),
    .B2(_1998_),
    .A2(_2050_),
    .A1(_1910_));
 sg13g2_inv_1 _5706_ (.Y(_0033_),
    .A(_2052_));
 sg13g2_nand2b_1 _5707_ (.Y(_2053_),
    .B(_1985_),
    .A_N(_1986_));
 sg13g2_nand3_1 _5708_ (.B(_1982_),
    .C(_2053_),
    .A(_1979_),
    .Y(_2054_));
 sg13g2_nand2b_1 _5709_ (.Y(_2055_),
    .B(_2054_),
    .A_N(_1934_));
 sg13g2_nor2_1 _5710_ (.A(_0061_),
    .B(_1898_),
    .Y(_2056_));
 sg13g2_buf_1 _5711_ (.A(_0062_),
    .X(_2057_));
 sg13g2_nand2_1 _5712_ (.Y(_2058_),
    .A(_1985_),
    .B(_1986_));
 sg13g2_or2_1 _5713_ (.X(_2059_),
    .B(_1986_),
    .A(_1985_));
 sg13g2_buf_1 _5714_ (.A(_2059_),
    .X(_2060_));
 sg13g2_o21ai_1 _5715_ (.B1(_2060_),
    .Y(_2061_),
    .A1(_2057_),
    .A2(_2058_));
 sg13g2_nor4_1 _5716_ (.A(_0063_),
    .B(_1797_),
    .C(_1802_),
    .D(_2033_),
    .Y(_2062_));
 sg13g2_a221oi_1 _5717_ (.B2(_1984_),
    .C1(_2062_),
    .B1(_2061_),
    .A1(_1992_),
    .Y(_2063_),
    .A2(_2056_));
 sg13g2_o21ai_1 _5718_ (.B1(_2063_),
    .Y(_0021_),
    .A1(_1975_),
    .A2(_2055_));
 sg13g2_inv_1 _5719_ (.Y(_2064_),
    .A(_0068_));
 sg13g2_inv_1 _5720_ (.Y(_2065_),
    .A(_1917_));
 sg13g2_nor2_1 _5721_ (.A(_2065_),
    .B(_1880_),
    .Y(_2066_));
 sg13g2_inv_1 _5722_ (.Y(_2067_),
    .A(_1870_));
 sg13g2_nor2_1 _5723_ (.A(_2067_),
    .B(_1884_),
    .Y(_2068_));
 sg13g2_a221oi_1 _5724_ (.B2(_1877_),
    .C1(_2068_),
    .B1(_2066_),
    .A1(_2064_),
    .Y(_2069_),
    .A2(net274));
 sg13g2_nor2_1 _5725_ (.A(_1869_),
    .B(_2069_),
    .Y(_0039_));
 sg13g2_buf_1 _5726_ (.A(\uart_tx_inst.state[0] ),
    .X(_2070_));
 sg13g2_a21o_1 _5727_ (.A2(net262),
    .A1(\uart_tx_inst.state[3] ),
    .B1(_2070_),
    .X(_2071_));
 sg13g2_buf_1 _5728_ (.A(_1832_),
    .X(_2072_));
 sg13g2_a21o_1 _5729_ (.A2(_2071_),
    .A1(_1857_),
    .B1(net271),
    .X(_0040_));
 sg13g2_a21o_1 _5730_ (.A2(_1981_),
    .A1(\action[0] ),
    .B1(net271),
    .X(_0020_));
 sg13g2_nor2b_1 _5731_ (.A(_1789_),
    .B_N(_1788_),
    .Y(_2073_));
 sg13g2_nand2_1 _5732_ (.Y(_2074_),
    .A(_2040_),
    .B(net380));
 sg13g2_a21oi_1 _5733_ (.A1(_1787_),
    .A2(_2073_),
    .Y(_2075_),
    .B1(_2074_));
 sg13g2_a21oi_1 _5734_ (.A1(\txstate[5] ),
    .A2(_2045_),
    .Y(_2076_),
    .B1(_2075_));
 sg13g2_o21ai_1 _5735_ (.B1(_2076_),
    .Y(_0034_),
    .A1(_1805_),
    .A2(_1827_));
 sg13g2_nand2b_1 _5736_ (.Y(_2077_),
    .B(\uart_tx_inst.state[3] ),
    .A_N(net262));
 sg13g2_nand3_1 _5737_ (.B(net262),
    .C(_1865_),
    .A(_1867_),
    .Y(_2078_));
 sg13g2_a21oi_1 _5738_ (.A1(_2077_),
    .A2(_2078_),
    .Y(_0043_),
    .B1(_1858_));
 sg13g2_and2_1 _5739_ (.A(_0067_),
    .B(net274),
    .X(_2079_));
 sg13g2_nand2_1 _5740_ (.Y(_2080_),
    .A(_1885_),
    .B(_1927_));
 sg13g2_a21oi_1 _5741_ (.A1(_1925_),
    .A2(_2080_),
    .Y(_2081_),
    .B1(_1926_));
 sg13g2_nor3_1 _5742_ (.A(_2065_),
    .B(_1877_),
    .C(_1922_),
    .Y(_2082_));
 sg13g2_nor4_1 _5743_ (.A(net388),
    .B(net274),
    .C(_2081_),
    .D(_2082_),
    .Y(_2083_));
 sg13g2_nor3_1 _5744_ (.A(_2072_),
    .B(_2079_),
    .C(_2083_),
    .Y(_0038_));
 sg13g2_nor2_1 _5745_ (.A(_1936_),
    .B(_2058_),
    .Y(_2084_));
 sg13g2_inv_2 _5746_ (.Y(_2085_),
    .A(net387));
 sg13g2_nand2_1 _5747_ (.Y(_2086_),
    .A(net371),
    .B(_2021_));
 sg13g2_nor2_1 _5748_ (.A(_1827_),
    .B(_2086_),
    .Y(_2087_));
 sg13g2_nor3_1 _5749_ (.A(net374),
    .B(_2085_),
    .C(_2087_),
    .Y(_2088_));
 sg13g2_a21oi_1 _5750_ (.A1(_1984_),
    .A2(_2084_),
    .Y(_2089_),
    .B1(_2088_));
 sg13g2_o21ai_1 _5751_ (.B1(_2089_),
    .Y(_0025_),
    .A1(net3),
    .A2(_1976_));
 sg13g2_buf_1 _5752_ (.A(\hvsync_inst.vpos[8] ),
    .X(_2090_));
 sg13g2_nand2b_1 _5753_ (.Y(_2091_),
    .B(_2090_),
    .A_N(\hvsync_inst.vpos[9] ));
 sg13g2_buf_4 _5754_ (.X(_2092_),
    .A(\cell_index[6] ));
 sg13g2_buf_2 _5755_ (.A(\cell_index[7] ),
    .X(_2093_));
 sg13g2_nand2_1 _5756_ (.Y(_2094_),
    .A(_2092_),
    .B(_2093_));
 sg13g2_buf_1 _5757_ (.A(\cell_index[5] ),
    .X(_2095_));
 sg13g2_nand2b_1 _5758_ (.Y(_2096_),
    .B(\hvsync_inst.vpos[3] ),
    .A_N(_2095_));
 sg13g2_buf_1 _5759_ (.A(\hvsync_inst.vpos[1] ),
    .X(_2097_));
 sg13g2_inv_1 _5760_ (.Y(_2098_),
    .A(\hvsync_inst.vpos[2] ));
 sg13g2_buf_2 _5761_ (.A(\cell_index[8] ),
    .X(_2099_));
 sg13g2_nand3_1 _5762_ (.B(_2098_),
    .C(_2099_),
    .A(_2097_),
    .Y(_2100_));
 sg13g2_nor4_1 _5763_ (.A(_2091_),
    .B(_2094_),
    .C(_2096_),
    .D(_2100_),
    .Y(_0045_));
 sg13g2_buf_2 _5764_ (.A(\cell_index[0] ),
    .X(_2101_));
 sg13g2_buf_1 _5765_ (.A(_2101_),
    .X(_2102_));
 sg13g2_buf_2 _5766_ (.A(_2102_),
    .X(_2103_));
 sg13g2_buf_1 _5767_ (.A(\cell_index[1] ),
    .X(_2104_));
 sg13g2_buf_1 _5768_ (.A(_2104_),
    .X(_2105_));
 sg13g2_buf_1 _5769_ (.A(_2105_),
    .X(_2106_));
 sg13g2_buf_1 _5770_ (.A(\cell_index[2] ),
    .X(_2107_));
 sg13g2_buf_1 _5771_ (.A(_2107_),
    .X(_2108_));
 sg13g2_buf_1 _5772_ (.A(net367),
    .X(_2109_));
 sg13g2_nor3_1 _5773_ (.A(net325),
    .B(net324),
    .C(net323),
    .Y(_2110_));
 sg13g2_and3_1 _5774_ (.X(_2111_),
    .A(net325),
    .B(net324),
    .C(net323));
 sg13g2_buf_1 _5775_ (.A(\cell_index[3] ),
    .X(_2112_));
 sg13g2_buf_2 _5776_ (.A(net385),
    .X(_2113_));
 sg13g2_buf_1 _5777_ (.A(\hvsync_inst.hpos[9] ),
    .X(_2114_));
 sg13g2_nand2_1 _5778_ (.Y(_2115_),
    .A(net366),
    .B(_2114_));
 sg13g2_nor4_1 _5779_ (.A(\cell_index[4] ),
    .B(_2110_),
    .C(_2111_),
    .D(_2115_),
    .Y(_0044_));
 sg13g2_inv_1 _5780_ (.Y(_2116_),
    .A(\cell_index[0] ));
 sg13g2_buf_2 _5781_ (.A(\hvsync_inst.hpos[2] ),
    .X(_2117_));
 sg13g2_buf_1 _5782_ (.A(\hvsync_inst.hpos[3] ),
    .X(_2118_));
 sg13g2_buf_1 _5783_ (.A(\hvsync_inst.hpos[1] ),
    .X(_2119_));
 sg13g2_buf_1 _5784_ (.A(\hvsync_inst.hpos[0] ),
    .X(_2120_));
 sg13g2_and2_1 _5785_ (.A(_2119_),
    .B(_2120_),
    .X(_2121_));
 sg13g2_buf_1 _5786_ (.A(_2121_),
    .X(_2122_));
 sg13g2_nand3_1 _5787_ (.B(_2118_),
    .C(_2122_),
    .A(_2117_),
    .Y(_2123_));
 sg13g2_nor2_2 _5788_ (.A(_2116_),
    .B(_2123_),
    .Y(_2124_));
 sg13g2_inv_1 _5789_ (.Y(_2125_),
    .A(\cell_index[4] ));
 sg13g2_nor4_1 _5790_ (.A(_2104_),
    .B(_2112_),
    .C(_2107_),
    .D(_2125_),
    .Y(_2126_));
 sg13g2_and3_1 _5791_ (.X(_2127_),
    .A(_2114_),
    .B(_2124_),
    .C(_2126_));
 sg13g2_buf_1 _5792_ (.A(_2127_),
    .X(_2128_));
 sg13g2_nand2b_1 _5793_ (.Y(_2129_),
    .B(\hvsync_inst.vpos[9] ),
    .A_N(_2090_));
 sg13g2_nor4_1 _5794_ (.A(_2097_),
    .B(_2093_),
    .C(_2096_),
    .D(_2129_),
    .Y(_2130_));
 sg13g2_buf_1 _5795_ (.A(\hvsync_inst.vpos[0] ),
    .X(_2131_));
 sg13g2_nor4_1 _5796_ (.A(_2131_),
    .B(_2098_),
    .C(_2092_),
    .D(_2099_),
    .Y(_2132_));
 sg13g2_a21oi_1 _5797_ (.A1(_2130_),
    .A2(_2132_),
    .Y(_2133_),
    .B1(_1830_));
 sg13g2_buf_1 _5798_ (.A(_2133_),
    .X(_2134_));
 sg13g2_and2_1 _5799_ (.A(_2128_),
    .B(_2134_),
    .X(_2135_));
 sg13g2_buf_2 _5800_ (.A(_2135_),
    .X(_2136_));
 sg13g2_nand3_1 _5801_ (.B(_2131_),
    .C(\hvsync_inst.vpos[2] ),
    .A(_2097_),
    .Y(_2137_));
 sg13g2_buf_1 _5802_ (.A(_2137_),
    .X(_2138_));
 sg13g2_nor2_1 _5803_ (.A(net374),
    .B(_2128_),
    .Y(_2139_));
 sg13g2_buf_1 _5804_ (.A(_2139_),
    .X(_2140_));
 sg13g2_a21o_1 _5805_ (.A2(_2138_),
    .A1(_2136_),
    .B1(net213),
    .X(_2141_));
 sg13g2_nand2_1 _5806_ (.Y(_2142_),
    .A(_2128_),
    .B(_2134_));
 sg13g2_o21ai_1 _5807_ (.B1(_0070_),
    .Y(_2143_),
    .A1(_2142_),
    .A2(_2138_));
 sg13g2_o21ai_1 _5808_ (.B1(_2143_),
    .Y(_2144_),
    .A1(_0070_),
    .A2(_2141_));
 sg13g2_buf_1 _5809_ (.A(_2144_),
    .X(_2145_));
 sg13g2_nand2_1 _5810_ (.Y(_2146_),
    .A(_2131_),
    .B(_2128_));
 sg13g2_xor2_1 _5811_ (.B(_2146_),
    .A(_2097_),
    .X(_2147_));
 sg13g2_nor2_1 _5812_ (.A(net374),
    .B(_2147_),
    .Y(_2148_));
 sg13g2_buf_1 _5813_ (.A(_2148_),
    .X(_1650_));
 sg13g2_nand2b_1 _5814_ (.Y(_2149_),
    .B(net401),
    .A_N(_2128_));
 sg13g2_buf_2 _5815_ (.A(_2149_),
    .X(_2150_));
 sg13g2_nand2_1 _5816_ (.Y(_2151_),
    .A(_2097_),
    .B(_2131_));
 sg13g2_xor2_1 _5817_ (.B(_2151_),
    .A(_0069_),
    .X(_2152_));
 sg13g2_nand2_1 _5818_ (.Y(_2153_),
    .A(_2136_),
    .B(_2152_));
 sg13g2_o21ai_1 _5819_ (.B1(_2153_),
    .Y(_2154_),
    .A1(_0069_),
    .A2(_2150_));
 sg13g2_buf_1 _5820_ (.A(_2154_),
    .X(_2155_));
 sg13g2_nand3_1 _5821_ (.B(_1650_),
    .C(_2155_),
    .A(_2145_),
    .Y(_2156_));
 sg13g2_nor2_1 _5822_ (.A(_1650_),
    .B(_2155_),
    .Y(_2157_));
 sg13g2_nand2b_1 _5823_ (.Y(_2158_),
    .B(_2157_),
    .A_N(_2145_));
 sg13g2_nand2_1 _5824_ (.Y(_0009_),
    .A(_2156_),
    .B(_2158_));
 sg13g2_xnor2_1 _5825_ (.Y(_0010_),
    .A(_2145_),
    .B(_2155_));
 sg13g2_inv_1 _5826_ (.Y(_2159_),
    .A(_0597_));
 sg13g2_nand2_1 _5827_ (.Y(_2160_),
    .A(_2131_),
    .B(net213));
 sg13g2_o21ai_1 _5828_ (.B1(_2160_),
    .Y(_1649_),
    .A1(_2159_),
    .A2(_2142_));
 sg13g2_a21oi_1 _5829_ (.A1(_1650_),
    .A2(_1649_),
    .Y(_2161_),
    .B1(_2155_));
 sg13g2_or2_1 _5830_ (.X(_2162_),
    .B(_1649_),
    .A(_1650_));
 sg13g2_nor2b_1 _5831_ (.A(_2145_),
    .B_N(_2155_),
    .Y(_2163_));
 sg13g2_a22oi_1 _5832_ (.Y(_0011_),
    .B1(_2162_),
    .B2(_2163_),
    .A2(_2161_),
    .A1(_2145_));
 sg13g2_a22oi_1 _5833_ (.Y(_0012_),
    .B1(_2163_),
    .B2(_1650_),
    .A2(_2157_),
    .A1(_2145_));
 sg13g2_nor3_1 _5834_ (.A(_2040_),
    .B(_1906_),
    .C(_0058_),
    .Y(_2164_));
 sg13g2_a21oi_1 _5835_ (.A1(_1789_),
    .A2(_1833_),
    .Y(_2165_),
    .B1(_2073_));
 sg13g2_or2_1 _5836_ (.X(_2166_),
    .B(_2165_),
    .A(_2164_));
 sg13g2_buf_2 _5837_ (.A(_2166_),
    .X(_2167_));
 sg13g2_nor2b_1 _5838_ (.A(_2040_),
    .B_N(_1834_),
    .Y(_2168_));
 sg13g2_nor3_1 _5839_ (.A(_1789_),
    .B(_1908_),
    .C(_2168_),
    .Y(_2169_));
 sg13g2_a21oi_2 _5840_ (.B1(_2169_),
    .Y(_2170_),
    .A2(_1844_),
    .A1(_1789_));
 sg13g2_nor2_1 _5841_ (.A(_2167_),
    .B(_2170_),
    .Y(_2171_));
 sg13g2_buf_2 _5842_ (.A(_2171_),
    .X(_2172_));
 sg13g2_and2_1 _5843_ (.A(net392),
    .B(net391),
    .X(_2173_));
 sg13g2_buf_1 _5844_ (.A(_2173_),
    .X(_2174_));
 sg13g2_nand3_1 _5845_ (.B(_1837_),
    .C(_2174_),
    .A(_1841_),
    .Y(_2175_));
 sg13g2_nor2_1 _5846_ (.A(_1840_),
    .B(_2175_),
    .Y(_2176_));
 sg13g2_a21o_1 _5847_ (.A2(_1844_),
    .A1(net382),
    .B1(_2169_),
    .X(_2177_));
 sg13g2_a21oi_1 _5848_ (.A1(_2177_),
    .A2(_2175_),
    .Y(_2178_),
    .B1(_2167_));
 sg13g2_nor2b_1 _5849_ (.A(_2178_),
    .B_N(_1840_),
    .Y(_2179_));
 sg13g2_a21oi_1 _5850_ (.A1(_2172_),
    .A2(_2176_),
    .Y(_2180_),
    .B1(_2179_));
 sg13g2_buf_1 _5851_ (.A(_0080_),
    .X(_2181_));
 sg13g2_inv_1 _5852_ (.Y(_2182_),
    .A(_2181_));
 sg13g2_nor2_2 _5853_ (.A(_2164_),
    .B(_2165_),
    .Y(_2183_));
 sg13g2_nand4_1 _5854_ (.B(net392),
    .C(_2182_),
    .A(_1837_),
    .Y(_2184_),
    .D(_2183_));
 sg13g2_xor2_1 _5855_ (.B(_2184_),
    .A(_1841_),
    .X(_2185_));
 sg13g2_inv_1 _5856_ (.Y(_2186_),
    .A(_2185_));
 sg13g2_nor2_1 _5857_ (.A(_2180_),
    .B(_2186_),
    .Y(_2187_));
 sg13g2_nand2_1 _5858_ (.Y(_2188_),
    .A(_0056_),
    .B(_2167_));
 sg13g2_xnor2_1 _5859_ (.Y(_2189_),
    .A(net392),
    .B(net391));
 sg13g2_o21ai_1 _5860_ (.B1(_2183_),
    .Y(_2190_),
    .A1(_2170_),
    .A2(_2189_));
 sg13g2_and2_1 _5861_ (.A(_2188_),
    .B(_2190_),
    .X(_2191_));
 sg13g2_buf_1 _5862_ (.A(_2191_),
    .X(_2192_));
 sg13g2_inv_1 _5863_ (.Y(_2193_),
    .A(_0081_));
 sg13g2_o21ai_1 _5864_ (.B1(_2183_),
    .Y(_2194_),
    .A1(_2170_),
    .A2(_2174_));
 sg13g2_nand2_1 _5865_ (.Y(_2195_),
    .A(_2193_),
    .B(_2194_));
 sg13g2_nand3_1 _5866_ (.B(_2174_),
    .C(_2172_),
    .A(_0081_),
    .Y(_2196_));
 sg13g2_and2_1 _5867_ (.A(_2195_),
    .B(_2196_),
    .X(_2197_));
 sg13g2_buf_1 _5868_ (.A(_2197_),
    .X(_2198_));
 sg13g2_nor2_1 _5869_ (.A(_2181_),
    .B(_2183_),
    .Y(_2199_));
 sg13g2_a21oi_2 _5870_ (.B1(_2199_),
    .Y(_2200_),
    .A2(_2172_),
    .A1(_2181_));
 sg13g2_nand2_1 _5871_ (.Y(_2201_),
    .A(_2198_),
    .B(_2200_));
 sg13g2_buf_2 _5872_ (.A(_2201_),
    .X(_2202_));
 sg13g2_a21o_1 _5873_ (.A2(_2172_),
    .A1(_2181_),
    .B1(_2199_),
    .X(_2203_));
 sg13g2_buf_1 _5874_ (.A(_2203_),
    .X(_2204_));
 sg13g2_nand2_1 _5875_ (.Y(_2205_),
    .A(_2204_),
    .B(net240));
 sg13g2_o21ai_1 _5876_ (.B1(_2205_),
    .Y(_2206_),
    .A1(net240),
    .A2(_2202_));
 sg13g2_nand2_1 _5877_ (.Y(_2207_),
    .A(_2188_),
    .B(_2190_));
 sg13g2_buf_2 _5878_ (.A(_2207_),
    .X(_2208_));
 sg13g2_buf_1 _5879_ (.A(_2208_),
    .X(_2209_));
 sg13g2_buf_1 _5880_ (.A(_2198_),
    .X(_2210_));
 sg13g2_o21ai_1 _5881_ (.B1(net401),
    .Y(_2211_),
    .A1(_2167_),
    .A2(_2177_));
 sg13g2_or2_1 _5882_ (.X(_2212_),
    .B(_2185_),
    .A(_2211_));
 sg13g2_buf_2 _5883_ (.A(_2212_),
    .X(_2213_));
 sg13g2_inv_1 _5884_ (.Y(_2214_),
    .A(_2213_));
 sg13g2_nand2_1 _5885_ (.Y(_2215_),
    .A(net103),
    .B(_2214_));
 sg13g2_nor2_1 _5886_ (.A(_2202_),
    .B(_2214_),
    .Y(_2216_));
 sg13g2_nor2_1 _5887_ (.A(_2200_),
    .B(_2213_),
    .Y(_2217_));
 sg13g2_o21ai_1 _5888_ (.B1(_2209_),
    .Y(_2218_),
    .A1(_2216_),
    .A2(_2217_));
 sg13g2_o21ai_1 _5889_ (.B1(_2218_),
    .Y(_2219_),
    .A1(net212),
    .A2(_2215_));
 sg13g2_buf_1 _5890_ (.A(_2180_),
    .X(_2220_));
 sg13g2_buf_1 _5891_ (.A(_2204_),
    .X(_2221_));
 sg13g2_nor2_1 _5892_ (.A(_2204_),
    .B(_2208_),
    .Y(_2222_));
 sg13g2_a22oi_1 _5893_ (.Y(_2223_),
    .B1(_2222_),
    .B2(net211),
    .A2(_2187_),
    .A1(net171));
 sg13g2_nor2_1 _5894_ (.A(net103),
    .B(_2223_),
    .Y(_2224_));
 sg13g2_a221oi_1 _5895_ (.B2(net211),
    .C1(_2224_),
    .B1(_2219_),
    .A1(_2187_),
    .Y(_2225_),
    .A2(_2206_));
 sg13g2_buf_1 _5896_ (.A(_2213_),
    .X(_2226_));
 sg13g2_nand2_1 _5897_ (.Y(_2227_),
    .A(_2195_),
    .B(_2196_));
 sg13g2_buf_1 _5898_ (.A(_2227_),
    .X(_2228_));
 sg13g2_nor2_1 _5899_ (.A(net170),
    .B(net240),
    .Y(_2229_));
 sg13g2_a21o_1 _5900_ (.A2(_2176_),
    .A1(_2172_),
    .B1(_2179_),
    .X(_2230_));
 sg13g2_buf_1 _5901_ (.A(_2230_),
    .X(_2231_));
 sg13g2_nand2_2 _5902_ (.Y(_2232_),
    .A(_1793_),
    .B(net209));
 sg13g2_inv_1 _5903_ (.Y(_1720_),
    .A(_2232_));
 sg13g2_a21oi_1 _5904_ (.A1(net170),
    .A2(_1720_),
    .Y(_2233_),
    .B1(_2204_));
 sg13g2_a22oi_1 _5905_ (.Y(_2234_),
    .B1(_2233_),
    .B2(net240),
    .A2(_2229_),
    .A1(net171));
 sg13g2_nor2_1 _5906_ (.A(_2204_),
    .B(_2192_),
    .Y(_2235_));
 sg13g2_nor2_1 _5907_ (.A(net209),
    .B(_2213_),
    .Y(_2236_));
 sg13g2_nand2_1 _5908_ (.Y(_2237_),
    .A(net170),
    .B(_2204_));
 sg13g2_nor2_1 _5909_ (.A(_2236_),
    .B(_2237_),
    .Y(_2238_));
 sg13g2_a21oi_1 _5910_ (.A1(_2187_),
    .A2(_2235_),
    .Y(_2239_),
    .B1(_2238_));
 sg13g2_o21ai_1 _5911_ (.B1(_2239_),
    .Y(_2240_),
    .A1(net210),
    .A2(_2234_));
 sg13g2_nand2_1 _5912_ (.Y(_2241_),
    .A(_1840_),
    .B(_1841_));
 sg13g2_nor2_1 _5913_ (.A(_2241_),
    .B(_2184_),
    .Y(_2242_));
 sg13g2_xnor2_1 _5914_ (.Y(_2243_),
    .A(_1839_),
    .B(_2242_));
 sg13g2_or2_1 _5915_ (.X(_2244_),
    .B(_2243_),
    .A(_2211_));
 sg13g2_buf_1 _5916_ (.A(_2244_),
    .X(_2245_));
 sg13g2_mux2_1 _5917_ (.A0(_2225_),
    .A1(_2240_),
    .S(_2245_),
    .X(_2246_));
 sg13g2_nand2_1 _5918_ (.Y(_0013_),
    .A(net329),
    .B(_2246_));
 sg13g2_buf_1 _5919_ (.A(_2245_),
    .X(_2247_));
 sg13g2_o21ai_1 _5920_ (.B1(net103),
    .Y(_2248_),
    .A1(net209),
    .A2(net212));
 sg13g2_nor2_2 _5921_ (.A(net103),
    .B(_2208_),
    .Y(_2249_));
 sg13g2_o21ai_1 _5922_ (.B1(net211),
    .Y(_2250_),
    .A1(net210),
    .A2(_2249_));
 sg13g2_nand2_1 _5923_ (.Y(_2251_),
    .A(_2248_),
    .B(_2250_));
 sg13g2_nand2_2 _5924_ (.Y(_2252_),
    .A(_2227_),
    .B(_2208_));
 sg13g2_o21ai_1 _5925_ (.B1(net211),
    .Y(_2253_),
    .A1(net171),
    .A2(_2252_));
 sg13g2_buf_1 _5926_ (.A(_2214_),
    .X(_1719_));
 sg13g2_a22oi_1 _5927_ (.Y(_2254_),
    .B1(_2253_),
    .B2(net168),
    .A2(_2251_),
    .A1(net171));
 sg13g2_nand4_1 _5928_ (.B(_2228_),
    .C(_2220_),
    .A(_1796_),
    .Y(_2255_),
    .D(net210));
 sg13g2_a21o_1 _5929_ (.A2(_2255_),
    .A1(_2215_),
    .B1(net171),
    .X(_2256_));
 sg13g2_o21ai_1 _5930_ (.B1(_2213_),
    .Y(_2257_),
    .A1(net209),
    .A2(_2249_));
 sg13g2_o21ai_1 _5931_ (.B1(_2257_),
    .Y(_2258_),
    .A1(net103),
    .A2(net211));
 sg13g2_nand3_1 _5932_ (.B(net171),
    .C(_2258_),
    .A(net372),
    .Y(_2259_));
 sg13g2_nor3_1 _5933_ (.A(net170),
    .B(net168),
    .C(_2232_),
    .Y(_2260_));
 sg13g2_o21ai_1 _5934_ (.B1(net212),
    .Y(_2261_),
    .A1(_2236_),
    .A2(_2260_));
 sg13g2_nand4_1 _5935_ (.B(_2256_),
    .C(_2259_),
    .A(net169),
    .Y(_2262_),
    .D(_2261_));
 sg13g2_o21ai_1 _5936_ (.B1(_2262_),
    .Y(_0014_),
    .A1(net169),
    .A2(_2254_));
 sg13g2_buf_1 _5937_ (.A(_2200_),
    .X(_2263_));
 sg13g2_nor2_1 _5938_ (.A(net103),
    .B(net240),
    .Y(_2264_));
 sg13g2_nor2_1 _5939_ (.A(_2209_),
    .B(_1719_),
    .Y(_2265_));
 sg13g2_a21oi_1 _5940_ (.A1(_1719_),
    .A2(_2264_),
    .Y(_2266_),
    .B1(_2265_));
 sg13g2_nand3_1 _5941_ (.B(net168),
    .C(_2237_),
    .A(net240),
    .Y(_2267_));
 sg13g2_o21ai_1 _5942_ (.B1(_2267_),
    .Y(_2268_),
    .A1(_2263_),
    .A2(_2266_));
 sg13g2_nand2_1 _5943_ (.Y(_2269_),
    .A(net399),
    .B(net170));
 sg13g2_nor4_1 _5944_ (.A(_2245_),
    .B(_2186_),
    .C(_2222_),
    .D(_2269_),
    .Y(_2270_));
 sg13g2_a21oi_1 _5945_ (.A1(net169),
    .A2(_2268_),
    .Y(_2271_),
    .B1(_2270_));
 sg13g2_nand4_1 _5946_ (.B(net170),
    .C(_2222_),
    .A(net380),
    .Y(_2272_),
    .D(net210));
 sg13g2_inv_1 _5947_ (.Y(_1721_),
    .A(_2245_));
 sg13g2_a21oi_1 _5948_ (.A1(_2215_),
    .A2(_2272_),
    .Y(_2273_),
    .B1(_1721_));
 sg13g2_nor2_1 _5949_ (.A(_2245_),
    .B(_2202_),
    .Y(_2274_));
 sg13g2_o21ai_1 _5950_ (.B1(net212),
    .Y(_2275_),
    .A1(_2217_),
    .A2(_2274_));
 sg13g2_nor2_1 _5951_ (.A(_2204_),
    .B(_2213_),
    .Y(_2276_));
 sg13g2_nor3_1 _5952_ (.A(_2210_),
    .B(_2263_),
    .C(net168),
    .Y(_2277_));
 sg13g2_nor2_1 _5953_ (.A(_2245_),
    .B(net212),
    .Y(_2278_));
 sg13g2_o21ai_1 _5954_ (.B1(_2278_),
    .Y(_2279_),
    .A1(_2276_),
    .A2(_2277_));
 sg13g2_nand2_1 _5955_ (.Y(_2280_),
    .A(_2275_),
    .B(_2279_));
 sg13g2_nor3_1 _5956_ (.A(_1720_),
    .B(_2273_),
    .C(_2280_),
    .Y(_2281_));
 sg13g2_a21oi_1 _5957_ (.A1(_1720_),
    .A2(_2271_),
    .Y(_0015_),
    .B1(_2281_));
 sg13g2_nor2_1 _5958_ (.A(_1831_),
    .B(_2236_),
    .Y(_2282_));
 sg13g2_a21oi_1 _5959_ (.A1(_2221_),
    .A2(_2282_),
    .Y(_2283_),
    .B1(_2276_));
 sg13g2_nor2_1 _5960_ (.A(net103),
    .B(_2213_),
    .Y(_2284_));
 sg13g2_a221oi_1 _5961_ (.B2(net171),
    .C1(net212),
    .B1(_2284_),
    .A1(_2185_),
    .Y(_2285_),
    .A2(_1720_));
 sg13g2_a21o_1 _5962_ (.A2(_2283_),
    .A1(net212),
    .B1(_2285_),
    .X(_2286_));
 sg13g2_o21ai_1 _5963_ (.B1(_2286_),
    .Y(_2287_),
    .A1(_2202_),
    .A2(_2232_));
 sg13g2_nand2_1 _5964_ (.Y(_2288_),
    .A(net103),
    .B(_2208_));
 sg13g2_nand3_1 _5965_ (.B(_2213_),
    .C(_2288_),
    .A(net208),
    .Y(_2289_));
 sg13g2_o21ai_1 _5966_ (.B1(_2289_),
    .Y(_2290_),
    .A1(net208),
    .A2(_2252_));
 sg13g2_a221oi_1 _5967_ (.B2(net380),
    .C1(_1720_),
    .B1(_2290_),
    .A1(_2229_),
    .Y(_2291_),
    .A2(_2276_));
 sg13g2_nand2_1 _5968_ (.Y(_2292_),
    .A(_2198_),
    .B(net240));
 sg13g2_nand4_1 _5969_ (.B(net171),
    .C(_2292_),
    .A(net380),
    .Y(_2293_),
    .D(_2252_));
 sg13g2_a21oi_1 _5970_ (.A1(_2185_),
    .A2(_2293_),
    .Y(_2294_),
    .B1(_2232_));
 sg13g2_nor3_1 _5971_ (.A(net169),
    .B(_2291_),
    .C(_2294_),
    .Y(_2295_));
 sg13g2_a21oi_1 _5972_ (.A1(net169),
    .A2(_2287_),
    .Y(_0016_),
    .B1(_2295_));
 sg13g2_a21oi_1 _5973_ (.A1(_2292_),
    .A2(_2252_),
    .Y(_2296_),
    .B1(net209));
 sg13g2_a221oi_1 _5974_ (.B2(net209),
    .C1(_2296_),
    .B1(_2249_),
    .A1(net208),
    .Y(_2297_),
    .A2(net212));
 sg13g2_inv_1 _5975_ (.Y(_2298_),
    .A(_2205_));
 sg13g2_xnor2_1 _5976_ (.Y(_2299_),
    .A(_2208_),
    .B(_2202_));
 sg13g2_a221oi_1 _5977_ (.B2(net209),
    .C1(_2226_),
    .B1(_2299_),
    .A1(_2228_),
    .Y(_2300_),
    .A2(_2298_));
 sg13g2_a21oi_1 _5978_ (.A1(net210),
    .A2(_2297_),
    .Y(_2301_),
    .B1(_2300_));
 sg13g2_nor2_1 _5979_ (.A(net330),
    .B(_2301_),
    .Y(_2302_));
 sg13g2_nand3_1 _5980_ (.B(_2236_),
    .C(_2264_),
    .A(net208),
    .Y(_2303_));
 sg13g2_nor2_1 _5981_ (.A(_2227_),
    .B(net208),
    .Y(_2304_));
 sg13g2_a21oi_1 _5982_ (.A1(net208),
    .A2(_2292_),
    .Y(_2305_),
    .B1(_2304_));
 sg13g2_o21ai_1 _5983_ (.B1(_2292_),
    .Y(_2306_),
    .A1(_2200_),
    .A2(_2252_));
 sg13g2_nand2_1 _5984_ (.Y(_2307_),
    .A(net211),
    .B(_2306_));
 sg13g2_o21ai_1 _5985_ (.B1(_2307_),
    .Y(_2308_),
    .A1(net211),
    .A2(_2305_));
 sg13g2_nand3_1 _5986_ (.B(_2226_),
    .C(_2308_),
    .A(_1912_),
    .Y(_2309_));
 sg13g2_and3_1 _5987_ (.X(_2310_),
    .A(_1721_),
    .B(_2303_),
    .C(_2309_));
 sg13g2_a21oi_1 _5988_ (.A1(net169),
    .A2(_2302_),
    .Y(_0017_),
    .B1(_2310_));
 sg13g2_nand3_1 _5989_ (.B(_2205_),
    .C(_2202_),
    .A(_1798_),
    .Y(_2311_));
 sg13g2_xnor2_1 _5990_ (.Y(_2312_),
    .A(net208),
    .B(net240));
 sg13g2_a22oi_1 _5991_ (.Y(_2313_),
    .B1(_2312_),
    .B2(_2284_),
    .A2(_2311_),
    .A1(net210));
 sg13g2_a21oi_1 _5992_ (.A1(net169),
    .A2(_2313_),
    .Y(_2314_),
    .B1(_1720_));
 sg13g2_nand3_1 _5993_ (.B(_2221_),
    .C(_2249_),
    .A(_1912_),
    .Y(_2315_));
 sg13g2_a21oi_1 _5994_ (.A1(_2185_),
    .A2(_2315_),
    .Y(_2316_),
    .B1(_2247_));
 sg13g2_a21oi_1 _5995_ (.A1(net168),
    .A2(_2249_),
    .Y(_2317_),
    .B1(net209));
 sg13g2_nand2b_1 _5996_ (.Y(_2318_),
    .B(_1798_),
    .A_N(_2317_));
 sg13g2_o21ai_1 _5997_ (.B1(net210),
    .Y(_2319_),
    .A1(_1831_),
    .A2(_2229_));
 sg13g2_nand3_1 _5998_ (.B(_2318_),
    .C(_2319_),
    .A(_1721_),
    .Y(_2320_));
 sg13g2_o21ai_1 _5999_ (.B1(_2320_),
    .Y(_0018_),
    .A1(_2314_),
    .A2(_2316_));
 sg13g2_o21ai_1 _6000_ (.B1(net210),
    .Y(_2321_),
    .A1(_2235_),
    .A2(_2269_));
 sg13g2_xnor2_1 _6001_ (.Y(_2322_),
    .A(net170),
    .B(_2205_));
 sg13g2_nor2_1 _6002_ (.A(_2186_),
    .B(_2232_),
    .Y(_2323_));
 sg13g2_a22oi_1 _6003_ (.Y(_2324_),
    .B1(_2322_),
    .B2(_2323_),
    .A2(_2321_),
    .A1(_2318_));
 sg13g2_buf_1 _6004_ (.A(net372),
    .X(_2325_));
 sg13g2_nand3_1 _6005_ (.B(net208),
    .C(net211),
    .A(net170),
    .Y(_2326_));
 sg13g2_nand3_1 _6006_ (.B(_2231_),
    .C(_2298_),
    .A(_2210_),
    .Y(_2327_));
 sg13g2_nand3_1 _6007_ (.B(_2326_),
    .C(_2327_),
    .A(net168),
    .Y(_2328_));
 sg13g2_o21ai_1 _6008_ (.B1(_2328_),
    .Y(_2329_),
    .A1(net168),
    .A2(_2264_));
 sg13g2_o21ai_1 _6009_ (.B1(_2220_),
    .Y(_2330_),
    .A1(_2216_),
    .A2(_2264_));
 sg13g2_nand4_1 _6010_ (.B(_2247_),
    .C(_2329_),
    .A(net322),
    .Y(_2331_),
    .D(_2330_));
 sg13g2_o21ai_1 _6011_ (.B1(_2331_),
    .Y(_0019_),
    .A1(net169),
    .A2(_2324_));
 sg13g2_nor2_1 _6012_ (.A(_1933_),
    .B(\action[0] ),
    .Y(_2332_));
 sg13g2_nand4_1 _6013_ (.B(_2085_),
    .C(_1791_),
    .A(net1),
    .Y(_2333_),
    .D(_2332_));
 sg13g2_nor3_1 _6014_ (.A(net400),
    .B(_1990_),
    .C(_0064_),
    .Y(_2334_));
 sg13g2_nor2b_1 _6015_ (.A(_2333_),
    .B_N(_2334_),
    .Y(_2335_));
 sg13g2_buf_1 _6016_ (.A(net332),
    .X(_2336_));
 sg13g2_inv_1 _6017_ (.Y(_2337_),
    .A(_1810_));
 sg13g2_buf_1 _6018_ (.A(net369),
    .X(_2338_));
 sg13g2_nor2b_1 _6019_ (.A(net321),
    .B_N(_1815_),
    .Y(_2339_));
 sg13g2_buf_1 _6020_ (.A(_2339_),
    .X(_2340_));
 sg13g2_inv_2 _6021_ (.Y(_2341_),
    .A(net369));
 sg13g2_nor2_1 _6022_ (.A(_1815_),
    .B(net320),
    .Y(_2342_));
 sg13g2_buf_2 _6023_ (.A(_2342_),
    .X(_2343_));
 sg13g2_a22oi_1 _6024_ (.Y(_2344_),
    .B1(_2343_),
    .B2(net375),
    .A2(net260),
    .A1(_2337_));
 sg13g2_inv_1 _6025_ (.Y(_2345_),
    .A(_1808_));
 sg13g2_buf_1 _6026_ (.A(_2338_),
    .X(_2346_));
 sg13g2_nand2b_1 _6027_ (.Y(_2347_),
    .B(net269),
    .A_N(net331));
 sg13g2_inv_1 _6028_ (.Y(_2348_),
    .A(net395));
 sg13g2_buf_1 _6029_ (.A(_2348_),
    .X(_2349_));
 sg13g2_o21ai_1 _6030_ (.B1(net319),
    .Y(_2350_),
    .A1(net365),
    .A2(_2347_));
 sg13g2_and3_1 _6031_ (.X(_2351_),
    .A(_1811_),
    .B(net377),
    .C(net369));
 sg13g2_buf_2 _6032_ (.A(_2351_),
    .X(_2352_));
 sg13g2_nor2b_1 _6033_ (.A(_1810_),
    .B_N(_2352_),
    .Y(_2353_));
 sg13g2_a21oi_1 _6034_ (.A1(net375),
    .A2(_2350_),
    .Y(_2354_),
    .B1(_2353_));
 sg13g2_o21ai_1 _6035_ (.B1(_2354_),
    .Y(_2355_),
    .A1(net270),
    .A2(_2344_));
 sg13g2_nor2_1 _6036_ (.A(net377),
    .B(net369),
    .Y(_2356_));
 sg13g2_buf_1 _6037_ (.A(_2356_),
    .X(_2357_));
 sg13g2_nand3_1 _6038_ (.B(net270),
    .C(net268),
    .A(net375),
    .Y(_2358_));
 sg13g2_nand2_1 _6039_ (.Y(_2359_),
    .A(net377),
    .B(net369));
 sg13g2_buf_2 _6040_ (.A(_2359_),
    .X(_2360_));
 sg13g2_nand2b_1 _6041_ (.Y(_2361_),
    .B(net378),
    .A_N(net377));
 sg13g2_o21ai_1 _6042_ (.B1(_2361_),
    .Y(_2362_),
    .A1(net332),
    .A2(_2360_));
 sg13g2_inv_1 _6043_ (.Y(_2363_),
    .A(net378));
 sg13g2_buf_1 _6044_ (.A(_2363_),
    .X(_2364_));
 sg13g2_nor2_1 _6045_ (.A(_2363_),
    .B(net320),
    .Y(_2365_));
 sg13g2_inv_1 _6046_ (.Y(_2366_),
    .A(\cell_y[0] ));
 sg13g2_buf_1 _6047_ (.A(_2366_),
    .X(_2367_));
 sg13g2_a22oi_1 _6048_ (.Y(_2368_),
    .B1(_2365_),
    .B2(net364),
    .A2(net260),
    .A1(net267));
 sg13g2_nand2_1 _6049_ (.Y(_2369_),
    .A(net319),
    .B(_2368_));
 sg13g2_o21ai_1 _6050_ (.B1(_2369_),
    .Y(_2370_),
    .A1(net319),
    .A2(_2362_));
 sg13g2_buf_1 _6051_ (.A(net379),
    .X(_2371_));
 sg13g2_a21oi_1 _6052_ (.A1(_2358_),
    .A2(_2370_),
    .Y(_2372_),
    .B1(net318));
 sg13g2_nor2_1 _6053_ (.A(net364),
    .B(net319),
    .Y(_2373_));
 sg13g2_buf_1 _6054_ (.A(_2373_),
    .X(_2374_));
 sg13g2_nand2_1 _6055_ (.Y(_2375_),
    .A(net331),
    .B(net320));
 sg13g2_nor2b_1 _6056_ (.A(net332),
    .B_N(net331),
    .Y(_2376_));
 sg13g2_a21oi_1 _6057_ (.A1(net332),
    .A2(_2375_),
    .Y(_2377_),
    .B1(_2376_));
 sg13g2_buf_1 _6058_ (.A(_0073_),
    .X(_2378_));
 sg13g2_nor2_2 _6059_ (.A(net365),
    .B(net321),
    .Y(_2379_));
 sg13g2_nand3b_1 _6060_ (.B(net384),
    .C(_2379_),
    .Y(_2380_),
    .A_N(net331));
 sg13g2_o21ai_1 _6061_ (.B1(_2380_),
    .Y(_2381_),
    .A1(net318),
    .A2(_2377_));
 sg13g2_a21oi_1 _6062_ (.A1(_2374_),
    .A2(_2381_),
    .Y(_2382_),
    .B1(_1820_));
 sg13g2_o21ai_1 _6063_ (.B1(_2382_),
    .Y(_2383_),
    .A1(_2355_),
    .A2(_2372_));
 sg13g2_nand2_1 _6064_ (.Y(_2384_),
    .A(net365),
    .B(net321));
 sg13g2_and2_1 _6065_ (.A(_1808_),
    .B(_1811_),
    .X(_2385_));
 sg13g2_buf_1 _6066_ (.A(_2385_),
    .X(_2386_));
 sg13g2_buf_1 _6067_ (.A(_2386_),
    .X(_2387_));
 sg13g2_nand2_1 _6068_ (.Y(_2388_),
    .A(net364),
    .B(net266));
 sg13g2_o21ai_1 _6069_ (.B1(_2388_),
    .Y(_2389_),
    .A1(net270),
    .A2(_2384_));
 sg13g2_inv_1 _6070_ (.Y(_2390_),
    .A(_1820_));
 sg13g2_a21oi_1 _6071_ (.A1(net319),
    .A2(_2389_),
    .Y(_2391_),
    .B1(_2390_));
 sg13g2_nand2_1 _6072_ (.Y(_2392_),
    .A(net378),
    .B(net321));
 sg13g2_nor2_1 _6073_ (.A(_2348_),
    .B(net320),
    .Y(_2393_));
 sg13g2_nor3_1 _6074_ (.A(net395),
    .B(net378),
    .C(net321),
    .Y(_2394_));
 sg13g2_o21ai_1 _6075_ (.B1(net379),
    .Y(_2395_),
    .A1(_2393_),
    .A2(_2394_));
 sg13g2_a21oi_1 _6076_ (.A1(_2392_),
    .A2(_2395_),
    .Y(_2396_),
    .B1(net276));
 sg13g2_nand2_1 _6077_ (.Y(_2397_),
    .A(net267),
    .B(net260));
 sg13g2_nand2_1 _6078_ (.Y(_2398_),
    .A(_2397_),
    .B(_2392_));
 sg13g2_o21ai_1 _6079_ (.B1(_1807_),
    .Y(_2399_),
    .A1(net379),
    .A2(net269));
 sg13g2_nor2_1 _6080_ (.A(_2398_),
    .B(_2399_),
    .Y(_2400_));
 sg13g2_nor2_1 _6081_ (.A(net395),
    .B(net331),
    .Y(_2401_));
 sg13g2_buf_1 _6082_ (.A(net395),
    .X(_2402_));
 sg13g2_buf_1 _6083_ (.A(net365),
    .X(_2403_));
 sg13g2_xor2_1 _6084_ (.B(net321),
    .A(net378),
    .X(_2404_));
 sg13g2_nor3_1 _6085_ (.A(net363),
    .B(net317),
    .C(_2404_),
    .Y(_2405_));
 sg13g2_nor3_1 _6086_ (.A(_2400_),
    .B(_2401_),
    .C(_2405_),
    .Y(_2406_));
 sg13g2_o21ai_1 _6087_ (.B1(net375),
    .Y(_2407_),
    .A1(_2396_),
    .A2(_2406_));
 sg13g2_a21oi_1 _6088_ (.A1(net270),
    .A2(_2360_),
    .Y(_2408_),
    .B1(net317));
 sg13g2_inv_1 _6089_ (.Y(_2409_),
    .A(net268));
 sg13g2_o21ai_1 _6090_ (.B1(_2409_),
    .Y(_2410_),
    .A1(net332),
    .A2(_2360_));
 sg13g2_nor2_1 _6091_ (.A(net393),
    .B(net319),
    .Y(_2411_));
 sg13g2_buf_1 _6092_ (.A(_2411_),
    .X(_2412_));
 sg13g2_o21ai_1 _6093_ (.B1(_2412_),
    .Y(_2413_),
    .A1(_2408_),
    .A2(_2410_));
 sg13g2_nand3_1 _6094_ (.B(_2407_),
    .C(_2413_),
    .A(_2391_),
    .Y(_2414_));
 sg13g2_nand4_1 _6095_ (.B(net376),
    .C(_2383_),
    .A(net394),
    .Y(_2415_),
    .D(_2414_));
 sg13g2_mux2_1 _6096_ (.A0(_0084_),
    .A1(net396),
    .S(net332),
    .X(_2416_));
 sg13g2_o21ai_1 _6097_ (.B1(_2031_),
    .Y(_2417_),
    .A1(net318),
    .A2(_2416_));
 sg13g2_mux2_1 _6098_ (.A0(net396),
    .A1(net384),
    .S(net276),
    .X(_2418_));
 sg13g2_nor2_1 _6099_ (.A(net317),
    .B(_2418_),
    .Y(_2419_));
 sg13g2_nor2_1 _6100_ (.A(net379),
    .B(net267),
    .Y(_2420_));
 sg13g2_buf_1 _6101_ (.A(_2420_),
    .X(_2421_));
 sg13g2_a21oi_1 _6102_ (.A1(net318),
    .A2(net276),
    .Y(_2422_),
    .B1(net257));
 sg13g2_nand2_1 _6103_ (.Y(_2423_),
    .A(net393),
    .B(net395));
 sg13g2_nor2_2 _6104_ (.A(net378),
    .B(net377),
    .Y(_2424_));
 sg13g2_nor2_1 _6105_ (.A(_2423_),
    .B(_2424_),
    .Y(_2425_));
 sg13g2_o21ai_1 _6106_ (.B1(_2425_),
    .Y(_2426_),
    .A1(net396),
    .A2(_2422_));
 sg13g2_o21ai_1 _6107_ (.B1(_2426_),
    .Y(_2427_),
    .A1(_2417_),
    .A2(_2419_));
 sg13g2_o21ai_1 _6108_ (.B1(net363),
    .Y(_2428_),
    .A1(net318),
    .A2(_2375_));
 sg13g2_nor2_1 _6109_ (.A(_1808_),
    .B(net378),
    .Y(_2429_));
 sg13g2_buf_1 _6110_ (.A(_2429_),
    .X(_2430_));
 sg13g2_o21ai_1 _6111_ (.B1(_2361_),
    .Y(_2431_),
    .A1(net364),
    .A2(_2430_));
 sg13g2_or3_1 _6112_ (.A(_1811_),
    .B(net377),
    .C(_2028_),
    .X(_2432_));
 sg13g2_buf_1 _6113_ (.A(_2432_),
    .X(_2433_));
 sg13g2_nand2_1 _6114_ (.Y(_2434_),
    .A(_2423_),
    .B(_2433_));
 sg13g2_a221oi_1 _6115_ (.B2(net269),
    .C1(_2434_),
    .B1(_2431_),
    .A1(net364),
    .Y(_2435_),
    .A2(_2428_));
 sg13g2_nand2_1 _6116_ (.Y(_2436_),
    .A(net394),
    .B(_2390_));
 sg13g2_nor2_2 _6117_ (.A(net376),
    .B(_2436_),
    .Y(_2437_));
 sg13g2_o21ai_1 _6118_ (.B1(_2437_),
    .Y(_2438_),
    .A1(_2427_),
    .A2(_2435_));
 sg13g2_nor3_1 _6119_ (.A(_1785_),
    .B(net400),
    .C(_2333_),
    .Y(_2439_));
 sg13g2_nor2_1 _6120_ (.A(net365),
    .B(net320),
    .Y(_2440_));
 sg13g2_nand2_1 _6121_ (.Y(_2441_),
    .A(_2349_),
    .B(_2424_));
 sg13g2_nand2_1 _6122_ (.Y(_2442_),
    .A(_1818_),
    .B(_2441_));
 sg13g2_nor2_1 _6123_ (.A(_1813_),
    .B(_2409_),
    .Y(_2443_));
 sg13g2_a21o_1 _6124_ (.A2(net266),
    .A1(net269),
    .B1(_2443_),
    .X(_2444_));
 sg13g2_nor2_1 _6125_ (.A(net267),
    .B(net331),
    .Y(_2445_));
 sg13g2_nand2_1 _6126_ (.Y(_2446_),
    .A(_1809_),
    .B(net267));
 sg13g2_a22oi_1 _6127_ (.Y(_2447_),
    .B1(_2446_),
    .B2(net320),
    .A2(_2445_),
    .A1(_2403_));
 sg13g2_a21oi_1 _6128_ (.A1(_2403_),
    .A2(_2340_),
    .Y(_2448_),
    .B1(_2367_));
 sg13g2_o21ai_1 _6129_ (.B1(_2448_),
    .Y(_2449_),
    .A1(net363),
    .A2(_2447_));
 sg13g2_a221oi_1 _6130_ (.B2(net363),
    .C1(_2449_),
    .B1(_2444_),
    .A1(_2440_),
    .Y(_2450_),
    .A2(_2442_));
 sg13g2_a21oi_1 _6131_ (.A1(net321),
    .A2(_2361_),
    .Y(_2451_),
    .B1(net379));
 sg13g2_o21ai_1 _6132_ (.B1(_2412_),
    .Y(_2452_),
    .A1(_2376_),
    .A2(_2451_));
 sg13g2_nor2_1 _6133_ (.A(_2347_),
    .B(_2446_),
    .Y(_2453_));
 sg13g2_a21oi_1 _6134_ (.A1(_2417_),
    .A2(_2452_),
    .Y(_2454_),
    .B1(_2453_));
 sg13g2_nand2_1 _6135_ (.Y(_2455_),
    .A(\cell_y[2] ),
    .B(_1820_));
 sg13g2_nor2_2 _6136_ (.A(net376),
    .B(_2455_),
    .Y(_2456_));
 sg13g2_o21ai_1 _6137_ (.B1(_2456_),
    .Y(_2457_),
    .A1(_2450_),
    .A2(_2454_));
 sg13g2_and4_1 _6138_ (.A(_2415_),
    .B(_2438_),
    .C(_2439_),
    .D(_2457_),
    .X(_2458_));
 sg13g2_nand2_1 _6139_ (.Y(_2459_),
    .A(net364),
    .B(_2349_));
 sg13g2_mux2_1 _6140_ (.A0(net384),
    .A1(_0084_),
    .S(net321),
    .X(_2460_));
 sg13g2_nor2_1 _6141_ (.A(_2366_),
    .B(\cell_x[4] ),
    .Y(_2461_));
 sg13g2_buf_1 _6142_ (.A(_2461_),
    .X(_2462_));
 sg13g2_o21ai_1 _6143_ (.B1(_2462_),
    .Y(_2463_),
    .A1(_2345_),
    .A2(_2460_));
 sg13g2_buf_1 _6144_ (.A(_2463_),
    .X(_2464_));
 sg13g2_a21oi_1 _6145_ (.A1(net331),
    .A2(_2464_),
    .Y(_2465_),
    .B1(_2356_));
 sg13g2_nand2_1 _6146_ (.Y(_2466_),
    .A(_2440_),
    .B(_2464_));
 sg13g2_o21ai_1 _6147_ (.B1(_2466_),
    .Y(_2467_),
    .A1(_2371_),
    .A2(_2465_));
 sg13g2_nor2_1 _6148_ (.A(_1816_),
    .B(_2384_),
    .Y(_2468_));
 sg13g2_a22oi_1 _6149_ (.Y(_2469_),
    .B1(_2468_),
    .B2(_2459_),
    .A2(_2464_),
    .A1(net320));
 sg13g2_nor2_1 _6150_ (.A(net270),
    .B(_2469_),
    .Y(_2470_));
 sg13g2_a221oi_1 _6151_ (.B2(_2336_),
    .C1(_2470_),
    .B1(_2467_),
    .A1(_2459_),
    .Y(_2471_),
    .A2(_2464_));
 sg13g2_nand2_1 _6152_ (.Y(_2472_),
    .A(net267),
    .B(net269));
 sg13g2_nand2_1 _6153_ (.Y(_2473_),
    .A(_1812_),
    .B(_2340_));
 sg13g2_o21ai_1 _6154_ (.B1(_2473_),
    .Y(_2474_),
    .A1(_2472_),
    .A2(_2411_));
 sg13g2_nor2_1 _6155_ (.A(_1812_),
    .B(_2338_),
    .Y(_2475_));
 sg13g2_xnor2_1 _6156_ (.Y(_2476_),
    .A(net365),
    .B(_2475_));
 sg13g2_o21ai_1 _6157_ (.B1(_2411_),
    .Y(_2477_),
    .A1(net276),
    .A2(_2476_));
 sg13g2_inv_1 _6158_ (.Y(_2478_),
    .A(net257));
 sg13g2_o21ai_1 _6159_ (.B1(_2425_),
    .Y(_2479_),
    .A1(net396),
    .A2(_2478_));
 sg13g2_a22oi_1 _6160_ (.Y(_2480_),
    .B1(_2477_),
    .B2(_2479_),
    .A2(_2474_),
    .A1(net318));
 sg13g2_buf_1 _6161_ (.A(_1820_),
    .X(_2481_));
 sg13g2_o21ai_1 _6162_ (.B1(net362),
    .Y(_2482_),
    .A1(_2471_),
    .A2(_2480_));
 sg13g2_and2_1 _6163_ (.A(_1814_),
    .B(net369),
    .X(_2483_));
 sg13g2_buf_2 _6164_ (.A(_2483_),
    .X(_2484_));
 sg13g2_a22oi_1 _6165_ (.Y(_2485_),
    .B1(_2430_),
    .B2(_2484_),
    .A2(net268),
    .A1(net332));
 sg13g2_o21ai_1 _6166_ (.B1(net363),
    .Y(_2486_),
    .A1(_2357_),
    .A2(_2365_));
 sg13g2_nor2_1 _6167_ (.A(net319),
    .B(net267),
    .Y(_2487_));
 sg13g2_o21ai_1 _6168_ (.B1(net318),
    .Y(_2488_),
    .A1(_2401_),
    .A2(_2487_));
 sg13g2_nand4_1 _6169_ (.B(_2485_),
    .C(_2486_),
    .A(_1824_),
    .Y(_2489_),
    .D(_2488_));
 sg13g2_a22oi_1 _6170_ (.Y(_2490_),
    .B1(_2387_),
    .B2(_0084_),
    .A2(_2343_),
    .A1(_2364_));
 sg13g2_nor2_1 _6171_ (.A(net269),
    .B(_2424_),
    .Y(_2491_));
 sg13g2_o21ai_1 _6172_ (.B1(net363),
    .Y(_2492_),
    .A1(_2451_),
    .A2(_2491_));
 sg13g2_o21ai_1 _6173_ (.B1(_2492_),
    .Y(_2493_),
    .A1(net363),
    .A2(_2490_));
 sg13g2_nand2_1 _6174_ (.Y(_2494_),
    .A(net364),
    .B(_2493_));
 sg13g2_a21o_1 _6175_ (.A2(_2494_),
    .A1(_2489_),
    .B1(net362),
    .X(_2495_));
 sg13g2_and3_1 _6176_ (.X(_2496_),
    .A(_1822_),
    .B(_2482_),
    .C(_2495_));
 sg13g2_nand3_1 _6177_ (.B(_2371_),
    .C(_2445_),
    .A(net393),
    .Y(_2497_));
 sg13g2_a21oi_1 _6178_ (.A1(_2397_),
    .A2(_2497_),
    .Y(_2498_),
    .B1(_2402_));
 sg13g2_nand2_1 _6179_ (.Y(_2499_),
    .A(net395),
    .B(net365));
 sg13g2_nor2_1 _6180_ (.A(_2347_),
    .B(_2499_),
    .Y(_2500_));
 sg13g2_a21oi_1 _6181_ (.A1(net267),
    .A2(_2343_),
    .Y(_2501_),
    .B1(net260));
 sg13g2_and4_1 _6182_ (.A(_1808_),
    .B(_1811_),
    .C(_1814_),
    .D(_2027_),
    .X(_2502_));
 sg13g2_buf_2 _6183_ (.A(_2502_),
    .X(_2503_));
 sg13g2_o21ai_1 _6184_ (.B1(net395),
    .Y(_2504_),
    .A1(_2430_),
    .A2(_2503_));
 sg13g2_o21ai_1 _6185_ (.B1(_2504_),
    .Y(_2505_),
    .A1(net379),
    .A2(_2501_));
 sg13g2_a21oi_1 _6186_ (.A1(_2357_),
    .A2(_2387_),
    .Y(_2506_),
    .B1(_2505_));
 sg13g2_nor2b_1 _6187_ (.A(_1808_),
    .B_N(net377),
    .Y(_2507_));
 sg13g2_o21ai_1 _6188_ (.B1(_2348_),
    .Y(_2508_),
    .A1(_2341_),
    .A2(_2507_));
 sg13g2_o21ai_1 _6189_ (.B1(_2508_),
    .Y(_2509_),
    .A1(net331),
    .A2(_1810_));
 sg13g2_a21oi_1 _6190_ (.A1(_2384_),
    .A2(_2473_),
    .Y(_2510_),
    .B1(net319));
 sg13g2_a221oi_1 _6191_ (.B2(_2364_),
    .C1(_2510_),
    .B1(_2509_),
    .A1(net365),
    .Y(_2511_),
    .A2(_2445_));
 sg13g2_or2_1 _6192_ (.X(_2512_),
    .B(_2511_),
    .A(net375));
 sg13g2_o21ai_1 _6193_ (.B1(_2512_),
    .Y(_2513_),
    .A1(net364),
    .A2(_2506_));
 sg13g2_nor4_1 _6194_ (.A(_2390_),
    .B(_2498_),
    .C(_2500_),
    .D(_2513_),
    .Y(_2514_));
 sg13g2_nor2_1 _6195_ (.A(net379),
    .B(net269),
    .Y(_2515_));
 sg13g2_o21ai_1 _6196_ (.B1(net317),
    .Y(_2516_),
    .A1(net393),
    .A2(net332));
 sg13g2_a221oi_1 _6197_ (.B2(_2393_),
    .C1(net266),
    .B1(_2516_),
    .A1(_1823_),
    .Y(_2517_),
    .A2(_2515_));
 sg13g2_nand2_1 _6198_ (.Y(_2518_),
    .A(net269),
    .B(_2499_));
 sg13g2_nand3_1 _6199_ (.B(_2376_),
    .C(_2518_),
    .A(_1824_),
    .Y(_2519_));
 sg13g2_o21ai_1 _6200_ (.B1(_2519_),
    .Y(_2520_),
    .A1(net276),
    .A2(_2517_));
 sg13g2_o21ai_1 _6201_ (.B1(_1817_),
    .Y(_2521_),
    .A1(_2421_),
    .A2(_2440_));
 sg13g2_a21oi_1 _6202_ (.A1(net379),
    .A2(net268),
    .Y(_2522_),
    .B1(_2365_));
 sg13g2_a21oi_1 _6203_ (.A1(net317),
    .A2(_2424_),
    .Y(_2523_),
    .B1(net266));
 sg13g2_mux2_1 _6204_ (.A0(_2522_),
    .A1(_2523_),
    .S(_1823_),
    .X(_2524_));
 sg13g2_a21oi_1 _6205_ (.A1(_2521_),
    .A2(_2524_),
    .Y(_2525_),
    .B1(_2402_));
 sg13g2_nor3_1 _6206_ (.A(net362),
    .B(_2520_),
    .C(_2525_),
    .Y(_2526_));
 sg13g2_nor3_1 _6207_ (.A(_1822_),
    .B(_2514_),
    .C(_2526_),
    .Y(_2527_));
 sg13g2_or3_1 _6208_ (.A(_1819_),
    .B(_2496_),
    .C(_2527_),
    .X(_2528_));
 sg13g2_nand2b_1 _6209_ (.Y(_2529_),
    .B(_2439_),
    .A_N(_2334_));
 sg13g2_nand2b_1 _6210_ (.Y(_2530_),
    .B(\lfsr.lfsr_reg[0] ),
    .A_N(_2335_));
 sg13g2_a22oi_1 _6211_ (.Y(_2531_),
    .B1(_2529_),
    .B2(_2530_),
    .A2(_2528_),
    .A1(_2458_));
 sg13g2_a21o_1 _6212_ (.A2(_2335_),
    .A1(\board_state_next[511] ),
    .B1(_2531_),
    .X(_2532_));
 sg13g2_buf_2 _6213_ (.A(_2532_),
    .X(_2533_));
 sg13g2_buf_1 _6214_ (.A(_2533_),
    .X(_2534_));
 sg13g2_buf_1 _6215_ (.A(_2534_),
    .X(_2535_));
 sg13g2_inv_1 _6216_ (.Y(_2536_),
    .A(_2032_));
 sg13g2_nor2_2 _6217_ (.A(_2481_),
    .B(_2536_),
    .Y(_2537_));
 sg13g2_nand2_1 _6218_ (.Y(_2538_),
    .A(net326),
    .B(_2537_));
 sg13g2_buf_2 _6219_ (.A(_2538_),
    .X(_2539_));
 sg13g2_buf_1 _6220_ (.A(_2539_),
    .X(_2540_));
 sg13g2_a21oi_1 _6221_ (.A1(net400),
    .A2(_1990_),
    .Y(_2541_),
    .B1(_1785_));
 sg13g2_nor2_1 _6222_ (.A(_2334_),
    .B(_2541_),
    .Y(_2542_));
 sg13g2_nor2_1 _6223_ (.A(_2333_),
    .B(_2542_),
    .Y(_2543_));
 sg13g2_buf_2 _6224_ (.A(_2543_),
    .X(_2544_));
 sg13g2_nand2_1 _6225_ (.Y(_2545_),
    .A(_2029_),
    .B(_2544_));
 sg13g2_buf_1 _6226_ (.A(_2545_),
    .X(_2546_));
 sg13g2_buf_1 _6227_ (.A(_2546_),
    .X(_2547_));
 sg13g2_nor2_1 _6228_ (.A(net247),
    .B(_2547_),
    .Y(_2548_));
 sg13g2_mux2_1 _6229_ (.A0(\board_state[0] ),
    .A1(net59),
    .S(_2548_),
    .X(_0609_));
 sg13g2_buf_1 _6230_ (.A(net67),
    .X(_2549_));
 sg13g2_inv_1 _6231_ (.Y(_2550_),
    .A(_2544_));
 sg13g2_buf_2 _6232_ (.A(_0077_),
    .X(_2551_));
 sg13g2_nor3_2 _6233_ (.A(net394),
    .B(_2481_),
    .C(_2551_),
    .Y(_2552_));
 sg13g2_nand2_1 _6234_ (.Y(_2553_),
    .A(net316),
    .B(_2552_));
 sg13g2_buf_1 _6235_ (.A(_2553_),
    .X(_2554_));
 sg13g2_nor2_1 _6236_ (.A(_2550_),
    .B(_2554_),
    .Y(_2555_));
 sg13g2_buf_1 _6237_ (.A(_2555_),
    .X(_2556_));
 sg13g2_nand3_1 _6238_ (.B(net257),
    .C(net206),
    .A(net268),
    .Y(_2557_));
 sg13g2_mux2_1 _6239_ (.A0(net58),
    .A1(\board_state[100] ),
    .S(_2557_),
    .X(_0610_));
 sg13g2_nand3_1 _6240_ (.B(net257),
    .C(net206),
    .A(_2343_),
    .Y(_2558_));
 sg13g2_mux2_1 _6241_ (.A0(net58),
    .A1(\board_state[101] ),
    .S(_2558_),
    .X(_0611_));
 sg13g2_nand3_1 _6242_ (.B(net257),
    .C(net206),
    .A(net260),
    .Y(_2559_));
 sg13g2_mux2_1 _6243_ (.A0(_2549_),
    .A1(\board_state[102] ),
    .S(_2559_),
    .X(_0612_));
 sg13g2_nand3_1 _6244_ (.B(_2352_),
    .C(net206),
    .A(net317),
    .Y(_2560_));
 sg13g2_mux2_1 _6245_ (.A0(net58),
    .A1(\board_state[103] ),
    .S(_2560_),
    .X(_0613_));
 sg13g2_nand3_1 _6246_ (.B(_2424_),
    .C(net206),
    .A(_2379_),
    .Y(_2561_));
 sg13g2_mux2_1 _6247_ (.A0(net58),
    .A1(\board_state[104] ),
    .S(_2561_),
    .X(_0614_));
 sg13g2_nand2_1 _6248_ (.Y(_2562_),
    .A(_2453_),
    .B(net206));
 sg13g2_mux2_1 _6249_ (.A0(net58),
    .A1(\board_state[105] ),
    .S(_2562_),
    .X(_0615_));
 sg13g2_nand3_1 _6250_ (.B(_2379_),
    .C(_2556_),
    .A(_2376_),
    .Y(_2563_));
 sg13g2_mux2_1 _6251_ (.A0(net58),
    .A1(\board_state[106] ),
    .S(_2563_),
    .X(_0616_));
 sg13g2_nor2_1 _6252_ (.A(net317),
    .B(net270),
    .Y(_2564_));
 sg13g2_nand3_1 _6253_ (.B(_2564_),
    .C(_2556_),
    .A(_2484_),
    .Y(_2565_));
 sg13g2_mux2_1 _6254_ (.A0(net58),
    .A1(\board_state[107] ),
    .S(_2565_),
    .X(_0617_));
 sg13g2_nand3_1 _6255_ (.B(net266),
    .C(net206),
    .A(net268),
    .Y(_2566_));
 sg13g2_mux2_1 _6256_ (.A0(_2549_),
    .A1(\board_state[108] ),
    .S(_2566_),
    .X(_0618_));
 sg13g2_nand3_1 _6257_ (.B(net266),
    .C(net206),
    .A(_2343_),
    .Y(_2567_));
 sg13g2_mux2_1 _6258_ (.A0(net58),
    .A1(\board_state[109] ),
    .S(_2567_),
    .X(_0619_));
 sg13g2_buf_1 _6259_ (.A(_2544_),
    .X(_2568_));
 sg13g2_nand3_1 _6260_ (.B(net260),
    .C(_2564_),
    .A(_2568_),
    .Y(_2569_));
 sg13g2_buf_1 _6261_ (.A(_2569_),
    .X(_2570_));
 sg13g2_buf_1 _6262_ (.A(_2570_),
    .X(_2571_));
 sg13g2_nor2_1 _6263_ (.A(net247),
    .B(net167),
    .Y(_2572_));
 sg13g2_mux2_1 _6264_ (.A0(\board_state[10] ),
    .A1(net59),
    .S(_2572_),
    .X(_0620_));
 sg13g2_nand4_1 _6265_ (.B(net276),
    .C(_2379_),
    .A(net270),
    .Y(_2573_),
    .D(_2555_));
 sg13g2_mux2_1 _6266_ (.A0(net59),
    .A1(\board_state[110] ),
    .S(_2573_),
    .X(_0621_));
 sg13g2_nand2_1 _6267_ (.Y(_2574_),
    .A(_2484_),
    .B(_2386_));
 sg13g2_nor3_1 _6268_ (.A(_2550_),
    .B(_2574_),
    .C(_2554_),
    .Y(_2575_));
 sg13g2_mux2_1 _6269_ (.A0(\board_state[111] ),
    .A1(_2535_),
    .S(_2575_),
    .X(_0622_));
 sg13g2_nand2_1 _6270_ (.Y(_2576_),
    .A(net259),
    .B(_2552_));
 sg13g2_buf_2 _6271_ (.A(_2576_),
    .X(_2577_));
 sg13g2_buf_1 _6272_ (.A(_2577_),
    .X(_2578_));
 sg13g2_nor2_1 _6273_ (.A(_2547_),
    .B(net239),
    .Y(_2579_));
 sg13g2_mux2_1 _6274_ (.A0(\board_state[112] ),
    .A1(net59),
    .S(_2579_),
    .X(_0623_));
 sg13g2_nand3_1 _6275_ (.B(_2544_),
    .C(_2343_),
    .A(_2430_),
    .Y(_2580_));
 sg13g2_buf_1 _6276_ (.A(_2580_),
    .X(_2581_));
 sg13g2_buf_1 _6277_ (.A(_2581_),
    .X(_2582_));
 sg13g2_nor2_1 _6278_ (.A(net239),
    .B(_2582_),
    .Y(_2583_));
 sg13g2_mux2_1 _6279_ (.A0(\board_state[113] ),
    .A1(net59),
    .S(_2583_),
    .X(_0624_));
 sg13g2_nand3_1 _6280_ (.B(_2544_),
    .C(net260),
    .A(_2430_),
    .Y(_2584_));
 sg13g2_buf_1 _6281_ (.A(_2584_),
    .X(_2585_));
 sg13g2_buf_1 _6282_ (.A(_2585_),
    .X(_2586_));
 sg13g2_nor2_1 _6283_ (.A(_2578_),
    .B(_2586_),
    .Y(_2587_));
 sg13g2_mux2_1 _6284_ (.A0(\board_state[114] ),
    .A1(net59),
    .S(_2587_),
    .X(_0625_));
 sg13g2_nand3_1 _6285_ (.B(_2544_),
    .C(_2484_),
    .A(_2430_),
    .Y(_2588_));
 sg13g2_buf_1 _6286_ (.A(_2588_),
    .X(_2589_));
 sg13g2_buf_1 _6287_ (.A(_2589_),
    .X(_2590_));
 sg13g2_nor2_1 _6288_ (.A(_2578_),
    .B(_2590_),
    .Y(_2591_));
 sg13g2_mux2_1 _6289_ (.A0(\board_state[115] ),
    .A1(net59),
    .S(_2591_),
    .X(_0626_));
 sg13g2_nand3_1 _6290_ (.B(net246),
    .C(net257),
    .A(net268),
    .Y(_2592_));
 sg13g2_buf_1 _6291_ (.A(_2592_),
    .X(_2593_));
 sg13g2_buf_1 _6292_ (.A(_2593_),
    .X(_2594_));
 sg13g2_nor2_1 _6293_ (.A(net239),
    .B(_2594_),
    .Y(_2595_));
 sg13g2_mux2_1 _6294_ (.A0(\board_state[116] ),
    .A1(_2535_),
    .S(_2595_),
    .X(_0627_));
 sg13g2_nand3_1 _6295_ (.B(_2343_),
    .C(net257),
    .A(net246),
    .Y(_2596_));
 sg13g2_buf_1 _6296_ (.A(_2596_),
    .X(_2597_));
 sg13g2_buf_1 _6297_ (.A(_2597_),
    .X(_2598_));
 sg13g2_nor2_1 _6298_ (.A(net239),
    .B(_2598_),
    .Y(_2599_));
 sg13g2_mux2_1 _6299_ (.A0(\board_state[117] ),
    .A1(net59),
    .S(_2599_),
    .X(_0628_));
 sg13g2_buf_1 _6300_ (.A(_2534_),
    .X(_2600_));
 sg13g2_nand3_1 _6301_ (.B(net260),
    .C(net257),
    .A(net246),
    .Y(_2601_));
 sg13g2_buf_1 _6302_ (.A(_2601_),
    .X(_2602_));
 sg13g2_buf_1 _6303_ (.A(_2602_),
    .X(_2603_));
 sg13g2_nor2_1 _6304_ (.A(net239),
    .B(net164),
    .Y(_2604_));
 sg13g2_mux2_1 _6305_ (.A0(\board_state[118] ),
    .A1(_2600_),
    .S(_2604_),
    .X(_0629_));
 sg13g2_nand3_1 _6306_ (.B(_2568_),
    .C(_2352_),
    .A(net317),
    .Y(_2605_));
 sg13g2_buf_1 _6307_ (.A(_2605_),
    .X(_2606_));
 sg13g2_buf_1 _6308_ (.A(_2606_),
    .X(_2607_));
 sg13g2_nor2_1 _6309_ (.A(net239),
    .B(net163),
    .Y(_2608_));
 sg13g2_mux2_1 _6310_ (.A0(\board_state[119] ),
    .A1(net57),
    .S(_2608_),
    .X(_0630_));
 sg13g2_nand3_1 _6311_ (.B(_2484_),
    .C(_2564_),
    .A(net246),
    .Y(_2609_));
 sg13g2_buf_1 _6312_ (.A(_2609_),
    .X(_2610_));
 sg13g2_buf_1 _6313_ (.A(_2610_),
    .X(_2611_));
 sg13g2_nor2_1 _6314_ (.A(net247),
    .B(net162),
    .Y(_2612_));
 sg13g2_mux2_1 _6315_ (.A0(\board_state[11] ),
    .A1(net57),
    .S(_2612_),
    .X(_0631_));
 sg13g2_nand3_1 _6316_ (.B(_2379_),
    .C(_2424_),
    .A(net246),
    .Y(_2613_));
 sg13g2_buf_1 _6317_ (.A(_2613_),
    .X(_2614_));
 sg13g2_buf_1 _6318_ (.A(_2614_),
    .X(_2615_));
 sg13g2_nor2_1 _6319_ (.A(net239),
    .B(net161),
    .Y(_2616_));
 sg13g2_mux2_1 _6320_ (.A0(\board_state[120] ),
    .A1(net57),
    .S(_2616_),
    .X(_0632_));
 sg13g2_nand2_1 _6321_ (.Y(_2617_),
    .A(net246),
    .B(_2453_));
 sg13g2_buf_1 _6322_ (.A(_2617_),
    .X(_2618_));
 sg13g2_buf_1 _6323_ (.A(_2618_),
    .X(_2619_));
 sg13g2_nor2_1 _6324_ (.A(_2577_),
    .B(net160),
    .Y(_2620_));
 sg13g2_mux2_1 _6325_ (.A0(\board_state[121] ),
    .A1(net57),
    .S(_2620_),
    .X(_0633_));
 sg13g2_nor2_1 _6326_ (.A(net167),
    .B(net239),
    .Y(_2621_));
 sg13g2_mux2_1 _6327_ (.A0(\board_state[122] ),
    .A1(_2600_),
    .S(_2621_),
    .X(_0634_));
 sg13g2_nor2_1 _6328_ (.A(_2577_),
    .B(net162),
    .Y(_2622_));
 sg13g2_mux2_1 _6329_ (.A0(\board_state[123] ),
    .A1(net57),
    .S(_2622_),
    .X(_0635_));
 sg13g2_nand3_1 _6330_ (.B(_2544_),
    .C(net266),
    .A(net268),
    .Y(_2623_));
 sg13g2_buf_1 _6331_ (.A(_2623_),
    .X(_2624_));
 sg13g2_buf_1 _6332_ (.A(_2624_),
    .X(_2625_));
 sg13g2_nor2_1 _6333_ (.A(_2577_),
    .B(net202),
    .Y(_2626_));
 sg13g2_mux2_1 _6334_ (.A0(\board_state[124] ),
    .A1(net57),
    .S(_2626_),
    .X(_0636_));
 sg13g2_nand3_1 _6335_ (.B(_2343_),
    .C(net266),
    .A(net246),
    .Y(_2627_));
 sg13g2_buf_1 _6336_ (.A(_2627_),
    .X(_2628_));
 sg13g2_buf_1 _6337_ (.A(_2628_),
    .X(_2629_));
 sg13g2_nor2_1 _6338_ (.A(_2577_),
    .B(net159),
    .Y(_2630_));
 sg13g2_mux2_1 _6339_ (.A0(\board_state[125] ),
    .A1(net57),
    .S(_2630_),
    .X(_0637_));
 sg13g2_nand4_1 _6340_ (.B(net276),
    .C(_2544_),
    .A(net270),
    .Y(_2631_),
    .D(_2379_));
 sg13g2_buf_1 _6341_ (.A(_2631_),
    .X(_2632_));
 sg13g2_buf_1 _6342_ (.A(_2632_),
    .X(_2633_));
 sg13g2_nor2_1 _6343_ (.A(_2577_),
    .B(net201),
    .Y(_2634_));
 sg13g2_mux2_1 _6344_ (.A0(\board_state[126] ),
    .A1(net57),
    .S(_2634_),
    .X(_0638_));
 sg13g2_buf_1 _6345_ (.A(net67),
    .X(_2635_));
 sg13g2_nand2_1 _6346_ (.Y(_2636_),
    .A(net246),
    .B(_2503_));
 sg13g2_buf_1 _6347_ (.A(_2636_),
    .X(_2637_));
 sg13g2_buf_1 _6348_ (.A(_2637_),
    .X(_2638_));
 sg13g2_nor2_1 _6349_ (.A(_2577_),
    .B(net158),
    .Y(_2639_));
 sg13g2_mux2_1 _6350_ (.A0(\board_state[127] ),
    .A1(_2635_),
    .S(_2639_),
    .X(_0639_));
 sg13g2_nand2_1 _6351_ (.Y(_2640_),
    .A(net326),
    .B(_2437_));
 sg13g2_buf_2 _6352_ (.A(_2640_),
    .X(_2641_));
 sg13g2_buf_1 _6353_ (.A(_2641_),
    .X(_2642_));
 sg13g2_nor2_1 _6354_ (.A(net207),
    .B(net245),
    .Y(_2643_));
 sg13g2_mux2_1 _6355_ (.A0(\board_state[128] ),
    .A1(net56),
    .S(_2643_),
    .X(_0640_));
 sg13g2_nor2_1 _6356_ (.A(net205),
    .B(net245),
    .Y(_2644_));
 sg13g2_mux2_1 _6357_ (.A0(\board_state[129] ),
    .A1(net56),
    .S(_2644_),
    .X(_0641_));
 sg13g2_nor2_1 _6358_ (.A(net247),
    .B(net202),
    .Y(_2645_));
 sg13g2_mux2_1 _6359_ (.A0(\board_state[12] ),
    .A1(_2635_),
    .S(_2645_),
    .X(_0642_));
 sg13g2_nor2_1 _6360_ (.A(net204),
    .B(net245),
    .Y(_2646_));
 sg13g2_mux2_1 _6361_ (.A0(\board_state[130] ),
    .A1(net56),
    .S(_2646_),
    .X(_0643_));
 sg13g2_nor2_1 _6362_ (.A(net203),
    .B(net245),
    .Y(_2647_));
 sg13g2_mux2_1 _6363_ (.A0(\board_state[131] ),
    .A1(net56),
    .S(_2647_),
    .X(_0644_));
 sg13g2_nor2_1 _6364_ (.A(net166),
    .B(net245),
    .Y(_2648_));
 sg13g2_mux2_1 _6365_ (.A0(\board_state[132] ),
    .A1(net56),
    .S(_2648_),
    .X(_0645_));
 sg13g2_nor2_1 _6366_ (.A(net165),
    .B(net245),
    .Y(_2649_));
 sg13g2_mux2_1 _6367_ (.A0(\board_state[133] ),
    .A1(net56),
    .S(_2649_),
    .X(_0646_));
 sg13g2_nor2_1 _6368_ (.A(net164),
    .B(_2642_),
    .Y(_2650_));
 sg13g2_mux2_1 _6369_ (.A0(\board_state[134] ),
    .A1(net56),
    .S(_2650_),
    .X(_0647_));
 sg13g2_nor2_1 _6370_ (.A(net163),
    .B(_2642_),
    .Y(_2651_));
 sg13g2_mux2_1 _6371_ (.A0(\board_state[135] ),
    .A1(net56),
    .S(_2651_),
    .X(_0648_));
 sg13g2_buf_1 _6372_ (.A(net67),
    .X(_2652_));
 sg13g2_nor2_1 _6373_ (.A(net161),
    .B(net245),
    .Y(_2653_));
 sg13g2_mux2_1 _6374_ (.A0(\board_state[136] ),
    .A1(net55),
    .S(_2653_),
    .X(_0649_));
 sg13g2_nor2_1 _6375_ (.A(net160),
    .B(net245),
    .Y(_2654_));
 sg13g2_mux2_1 _6376_ (.A0(\board_state[137] ),
    .A1(net55),
    .S(_2654_),
    .X(_0650_));
 sg13g2_nor2_1 _6377_ (.A(net167),
    .B(_2641_),
    .Y(_2655_));
 sg13g2_mux2_1 _6378_ (.A0(\board_state[138] ),
    .A1(net55),
    .S(_2655_),
    .X(_0651_));
 sg13g2_nor2_1 _6379_ (.A(net162),
    .B(_2641_),
    .Y(_2656_));
 sg13g2_mux2_1 _6380_ (.A0(\board_state[139] ),
    .A1(net55),
    .S(_2656_),
    .X(_0652_));
 sg13g2_nor2_1 _6381_ (.A(net247),
    .B(net159),
    .Y(_2657_));
 sg13g2_mux2_1 _6382_ (.A0(\board_state[13] ),
    .A1(_2652_),
    .S(_2657_),
    .X(_0653_));
 sg13g2_nor2_1 _6383_ (.A(net202),
    .B(_2641_),
    .Y(_2658_));
 sg13g2_mux2_1 _6384_ (.A0(\board_state[140] ),
    .A1(net55),
    .S(_2658_),
    .X(_0654_));
 sg13g2_nor2_1 _6385_ (.A(net159),
    .B(_2641_),
    .Y(_2659_));
 sg13g2_mux2_1 _6386_ (.A0(\board_state[141] ),
    .A1(net55),
    .S(_2659_),
    .X(_0655_));
 sg13g2_nor2_1 _6387_ (.A(net201),
    .B(_2641_),
    .Y(_2660_));
 sg13g2_mux2_1 _6388_ (.A0(\board_state[142] ),
    .A1(net55),
    .S(_2660_),
    .X(_0656_));
 sg13g2_nor2_1 _6389_ (.A(net158),
    .B(_2641_),
    .Y(_2661_));
 sg13g2_mux2_1 _6390_ (.A0(\board_state[143] ),
    .A1(net55),
    .S(_2661_),
    .X(_0657_));
 sg13g2_nand2_1 _6391_ (.Y(_2662_),
    .A(net258),
    .B(_2437_));
 sg13g2_buf_1 _6392_ (.A(_2662_),
    .X(_2663_));
 sg13g2_buf_1 _6393_ (.A(_2663_),
    .X(_2664_));
 sg13g2_nor2_1 _6394_ (.A(net207),
    .B(net238),
    .Y(_2665_));
 sg13g2_mux2_1 _6395_ (.A0(\board_state[144] ),
    .A1(_2652_),
    .S(_2665_),
    .X(_0658_));
 sg13g2_buf_1 _6396_ (.A(net67),
    .X(_2666_));
 sg13g2_nor2_1 _6397_ (.A(net205),
    .B(net238),
    .Y(_2667_));
 sg13g2_mux2_1 _6398_ (.A0(\board_state[145] ),
    .A1(net54),
    .S(_2667_),
    .X(_0659_));
 sg13g2_nor2_1 _6399_ (.A(net204),
    .B(net238),
    .Y(_2668_));
 sg13g2_mux2_1 _6400_ (.A0(\board_state[146] ),
    .A1(net54),
    .S(_2668_),
    .X(_0660_));
 sg13g2_nor2_1 _6401_ (.A(net203),
    .B(net238),
    .Y(_2669_));
 sg13g2_mux2_1 _6402_ (.A0(\board_state[147] ),
    .A1(net54),
    .S(_2669_),
    .X(_0661_));
 sg13g2_nor2_1 _6403_ (.A(net166),
    .B(net238),
    .Y(_2670_));
 sg13g2_mux2_1 _6404_ (.A0(\board_state[148] ),
    .A1(net54),
    .S(_2670_),
    .X(_0662_));
 sg13g2_nor2_1 _6405_ (.A(net165),
    .B(net238),
    .Y(_2671_));
 sg13g2_mux2_1 _6406_ (.A0(\board_state[149] ),
    .A1(net54),
    .S(_2671_),
    .X(_0663_));
 sg13g2_nor2_1 _6407_ (.A(_2540_),
    .B(net201),
    .Y(_2672_));
 sg13g2_mux2_1 _6408_ (.A0(\board_state[14] ),
    .A1(_2666_),
    .S(_2672_),
    .X(_0664_));
 sg13g2_nor2_1 _6409_ (.A(net164),
    .B(net238),
    .Y(_2673_));
 sg13g2_mux2_1 _6410_ (.A0(\board_state[150] ),
    .A1(net54),
    .S(_2673_),
    .X(_0665_));
 sg13g2_nor2_1 _6411_ (.A(net163),
    .B(_2664_),
    .Y(_2674_));
 sg13g2_mux2_1 _6412_ (.A0(\board_state[151] ),
    .A1(_2666_),
    .S(_2674_),
    .X(_0666_));
 sg13g2_nor2_1 _6413_ (.A(net161),
    .B(_2664_),
    .Y(_2675_));
 sg13g2_mux2_1 _6414_ (.A0(\board_state[152] ),
    .A1(net54),
    .S(_2675_),
    .X(_0667_));
 sg13g2_nor2_1 _6415_ (.A(net160),
    .B(net238),
    .Y(_2676_));
 sg13g2_mux2_1 _6416_ (.A0(\board_state[153] ),
    .A1(net54),
    .S(_2676_),
    .X(_0668_));
 sg13g2_buf_1 _6417_ (.A(net67),
    .X(_2677_));
 sg13g2_nor2_1 _6418_ (.A(net167),
    .B(_2663_),
    .Y(_2678_));
 sg13g2_mux2_1 _6419_ (.A0(\board_state[154] ),
    .A1(net53),
    .S(_2678_),
    .X(_0669_));
 sg13g2_nor2_1 _6420_ (.A(net162),
    .B(_2663_),
    .Y(_2679_));
 sg13g2_mux2_1 _6421_ (.A0(\board_state[155] ),
    .A1(net53),
    .S(_2679_),
    .X(_0670_));
 sg13g2_nor2_1 _6422_ (.A(net202),
    .B(_2663_),
    .Y(_2680_));
 sg13g2_mux2_1 _6423_ (.A0(\board_state[156] ),
    .A1(net53),
    .S(_2680_),
    .X(_0671_));
 sg13g2_nor2_1 _6424_ (.A(net159),
    .B(_2663_),
    .Y(_2681_));
 sg13g2_mux2_1 _6425_ (.A0(\board_state[157] ),
    .A1(net53),
    .S(_2681_),
    .X(_0672_));
 sg13g2_nor2_1 _6426_ (.A(net201),
    .B(_2663_),
    .Y(_2682_));
 sg13g2_mux2_1 _6427_ (.A0(\board_state[158] ),
    .A1(net53),
    .S(_2682_),
    .X(_0673_));
 sg13g2_nor2_1 _6428_ (.A(net158),
    .B(_2663_),
    .Y(_2683_));
 sg13g2_mux2_1 _6429_ (.A0(\board_state[159] ),
    .A1(net53),
    .S(_2683_),
    .X(_0674_));
 sg13g2_nor2_1 _6430_ (.A(_2540_),
    .B(_2638_),
    .Y(_2684_));
 sg13g2_mux2_1 _6431_ (.A0(\board_state[15] ),
    .A1(_2677_),
    .S(_2684_),
    .X(_0675_));
 sg13g2_nand2_1 _6432_ (.Y(_2685_),
    .A(_2437_),
    .B(net316));
 sg13g2_buf_1 _6433_ (.A(_2685_),
    .X(_2686_));
 sg13g2_buf_1 _6434_ (.A(_2686_),
    .X(_2687_));
 sg13g2_nor2_1 _6435_ (.A(net207),
    .B(net244),
    .Y(_2688_));
 sg13g2_mux2_1 _6436_ (.A0(\board_state[160] ),
    .A1(net53),
    .S(_2688_),
    .X(_0676_));
 sg13g2_nor2_1 _6437_ (.A(net205),
    .B(net244),
    .Y(_2689_));
 sg13g2_mux2_1 _6438_ (.A0(\board_state[161] ),
    .A1(_2677_),
    .S(_2689_),
    .X(_0677_));
 sg13g2_nor2_1 _6439_ (.A(net204),
    .B(net244),
    .Y(_2690_));
 sg13g2_mux2_1 _6440_ (.A0(\board_state[162] ),
    .A1(net53),
    .S(_2690_),
    .X(_0678_));
 sg13g2_buf_1 _6441_ (.A(net67),
    .X(_2691_));
 sg13g2_nor2_1 _6442_ (.A(net203),
    .B(net244),
    .Y(_2692_));
 sg13g2_mux2_1 _6443_ (.A0(\board_state[163] ),
    .A1(net52),
    .S(_2692_),
    .X(_0679_));
 sg13g2_nor2_1 _6444_ (.A(net166),
    .B(net244),
    .Y(_2693_));
 sg13g2_mux2_1 _6445_ (.A0(\board_state[164] ),
    .A1(net52),
    .S(_2693_),
    .X(_0680_));
 sg13g2_nor2_1 _6446_ (.A(net165),
    .B(_2687_),
    .Y(_2694_));
 sg13g2_mux2_1 _6447_ (.A0(\board_state[165] ),
    .A1(net52),
    .S(_2694_),
    .X(_0681_));
 sg13g2_nor2_1 _6448_ (.A(net164),
    .B(net244),
    .Y(_2695_));
 sg13g2_mux2_1 _6449_ (.A0(\board_state[166] ),
    .A1(net52),
    .S(_2695_),
    .X(_0682_));
 sg13g2_nor2_1 _6450_ (.A(net163),
    .B(_2687_),
    .Y(_2696_));
 sg13g2_mux2_1 _6451_ (.A0(\board_state[167] ),
    .A1(net52),
    .S(_2696_),
    .X(_0683_));
 sg13g2_nor2_1 _6452_ (.A(net161),
    .B(net244),
    .Y(_2697_));
 sg13g2_mux2_1 _6453_ (.A0(\board_state[168] ),
    .A1(net52),
    .S(_2697_),
    .X(_0684_));
 sg13g2_nor2_1 _6454_ (.A(net160),
    .B(net244),
    .Y(_2698_));
 sg13g2_mux2_1 _6455_ (.A0(\board_state[169] ),
    .A1(_2691_),
    .S(_2698_),
    .X(_0685_));
 sg13g2_nand2_1 _6456_ (.Y(_2699_),
    .A(_2537_),
    .B(net258));
 sg13g2_buf_1 _6457_ (.A(_2699_),
    .X(_2700_));
 sg13g2_buf_1 _6458_ (.A(_2700_),
    .X(_2701_));
 sg13g2_nor2_1 _6459_ (.A(net207),
    .B(net237),
    .Y(_2702_));
 sg13g2_mux2_1 _6460_ (.A0(\board_state[16] ),
    .A1(_2691_),
    .S(_2702_),
    .X(_0686_));
 sg13g2_nor2_1 _6461_ (.A(net167),
    .B(_2686_),
    .Y(_2703_));
 sg13g2_mux2_1 _6462_ (.A0(\board_state[170] ),
    .A1(net52),
    .S(_2703_),
    .X(_0687_));
 sg13g2_nor2_1 _6463_ (.A(net162),
    .B(_2686_),
    .Y(_2704_));
 sg13g2_mux2_1 _6464_ (.A0(\board_state[171] ),
    .A1(net52),
    .S(_2704_),
    .X(_0688_));
 sg13g2_buf_1 _6465_ (.A(_2533_),
    .X(_2705_));
 sg13g2_buf_1 _6466_ (.A(net66),
    .X(_2706_));
 sg13g2_nor2_1 _6467_ (.A(_2625_),
    .B(_2686_),
    .Y(_2707_));
 sg13g2_mux2_1 _6468_ (.A0(\board_state[172] ),
    .A1(net51),
    .S(_2707_),
    .X(_0689_));
 sg13g2_nor2_1 _6469_ (.A(_2629_),
    .B(_2686_),
    .Y(_2708_));
 sg13g2_mux2_1 _6470_ (.A0(\board_state[173] ),
    .A1(net51),
    .S(_2708_),
    .X(_0690_));
 sg13g2_nor2_1 _6471_ (.A(_2633_),
    .B(_2686_),
    .Y(_2709_));
 sg13g2_mux2_1 _6472_ (.A0(\board_state[174] ),
    .A1(_2706_),
    .S(_2709_),
    .X(_0691_));
 sg13g2_nor2_1 _6473_ (.A(_2638_),
    .B(_2686_),
    .Y(_2710_));
 sg13g2_mux2_1 _6474_ (.A0(\board_state[175] ),
    .A1(_2706_),
    .S(_2710_),
    .X(_0692_));
 sg13g2_nand2_1 _6475_ (.Y(_2711_),
    .A(net259),
    .B(_2437_));
 sg13g2_buf_2 _6476_ (.A(_2711_),
    .X(_2712_));
 sg13g2_buf_1 _6477_ (.A(_2712_),
    .X(_2713_));
 sg13g2_nor2_1 _6478_ (.A(net207),
    .B(net236),
    .Y(_2714_));
 sg13g2_mux2_1 _6479_ (.A0(\board_state[176] ),
    .A1(net51),
    .S(_2714_),
    .X(_0693_));
 sg13g2_nor2_1 _6480_ (.A(_2582_),
    .B(net236),
    .Y(_2715_));
 sg13g2_mux2_1 _6481_ (.A0(\board_state[177] ),
    .A1(net51),
    .S(_2715_),
    .X(_0694_));
 sg13g2_nor2_1 _6482_ (.A(net204),
    .B(net236),
    .Y(_2716_));
 sg13g2_mux2_1 _6483_ (.A0(\board_state[178] ),
    .A1(net51),
    .S(_2716_),
    .X(_0695_));
 sg13g2_nor2_1 _6484_ (.A(net203),
    .B(net236),
    .Y(_2717_));
 sg13g2_mux2_1 _6485_ (.A0(\board_state[179] ),
    .A1(net51),
    .S(_2717_),
    .X(_0696_));
 sg13g2_nor2_1 _6486_ (.A(net205),
    .B(net237),
    .Y(_2718_));
 sg13g2_mux2_1 _6487_ (.A0(\board_state[17] ),
    .A1(net51),
    .S(_2718_),
    .X(_0697_));
 sg13g2_nor2_1 _6488_ (.A(net166),
    .B(net236),
    .Y(_2719_));
 sg13g2_mux2_1 _6489_ (.A0(\board_state[180] ),
    .A1(net51),
    .S(_2719_),
    .X(_0698_));
 sg13g2_buf_1 _6490_ (.A(net66),
    .X(_2720_));
 sg13g2_nor2_1 _6491_ (.A(net165),
    .B(net236),
    .Y(_2721_));
 sg13g2_mux2_1 _6492_ (.A0(\board_state[181] ),
    .A1(net50),
    .S(_2721_),
    .X(_0699_));
 sg13g2_nor2_1 _6493_ (.A(_2603_),
    .B(net236),
    .Y(_2722_));
 sg13g2_mux2_1 _6494_ (.A0(\board_state[182] ),
    .A1(net50),
    .S(_2722_),
    .X(_0700_));
 sg13g2_nor2_1 _6495_ (.A(net163),
    .B(net236),
    .Y(_2723_));
 sg13g2_mux2_1 _6496_ (.A0(\board_state[183] ),
    .A1(net50),
    .S(_2723_),
    .X(_0701_));
 sg13g2_nor2_1 _6497_ (.A(_2615_),
    .B(_2713_),
    .Y(_2724_));
 sg13g2_mux2_1 _6498_ (.A0(\board_state[184] ),
    .A1(net50),
    .S(_2724_),
    .X(_0702_));
 sg13g2_nor2_1 _6499_ (.A(net160),
    .B(_2713_),
    .Y(_2725_));
 sg13g2_mux2_1 _6500_ (.A0(\board_state[185] ),
    .A1(net50),
    .S(_2725_),
    .X(_0703_));
 sg13g2_nor2_1 _6501_ (.A(_2571_),
    .B(_2712_),
    .Y(_2726_));
 sg13g2_mux2_1 _6502_ (.A0(\board_state[186] ),
    .A1(net50),
    .S(_2726_),
    .X(_0704_));
 sg13g2_nor2_1 _6503_ (.A(_2611_),
    .B(_2712_),
    .Y(_2727_));
 sg13g2_mux2_1 _6504_ (.A0(\board_state[187] ),
    .A1(_2720_),
    .S(_2727_),
    .X(_0705_));
 sg13g2_nor2_1 _6505_ (.A(_2625_),
    .B(_2712_),
    .Y(_2728_));
 sg13g2_mux2_1 _6506_ (.A0(\board_state[188] ),
    .A1(_2720_),
    .S(_2728_),
    .X(_0706_));
 sg13g2_nor2_1 _6507_ (.A(_2629_),
    .B(_2712_),
    .Y(_2729_));
 sg13g2_mux2_1 _6508_ (.A0(\board_state[189] ),
    .A1(net50),
    .S(_2729_),
    .X(_0707_));
 sg13g2_nor2_1 _6509_ (.A(net204),
    .B(net237),
    .Y(_2730_));
 sg13g2_mux2_1 _6510_ (.A0(\board_state[18] ),
    .A1(net50),
    .S(_2730_),
    .X(_0708_));
 sg13g2_buf_1 _6511_ (.A(_2705_),
    .X(_2731_));
 sg13g2_nor2_1 _6512_ (.A(_2633_),
    .B(_2712_),
    .Y(_2732_));
 sg13g2_mux2_1 _6513_ (.A0(\board_state[190] ),
    .A1(_2731_),
    .S(_2732_),
    .X(_0709_));
 sg13g2_nor2_1 _6514_ (.A(net158),
    .B(_2712_),
    .Y(_2733_));
 sg13g2_mux2_1 _6515_ (.A0(\board_state[191] ),
    .A1(_2731_),
    .S(_2733_),
    .X(_0710_));
 sg13g2_nor2_2 _6516_ (.A(_2551_),
    .B(_2436_),
    .Y(_2734_));
 sg13g2_nand2_1 _6517_ (.Y(_2735_),
    .A(net326),
    .B(_2734_));
 sg13g2_buf_1 _6518_ (.A(_2735_),
    .X(_2736_));
 sg13g2_buf_1 _6519_ (.A(_2736_),
    .X(_2737_));
 sg13g2_nor2_1 _6520_ (.A(net207),
    .B(net243),
    .Y(_2738_));
 sg13g2_mux2_1 _6521_ (.A0(\board_state[192] ),
    .A1(net49),
    .S(_2738_),
    .X(_0711_));
 sg13g2_nor2_1 _6522_ (.A(net205),
    .B(net243),
    .Y(_2739_));
 sg13g2_mux2_1 _6523_ (.A0(\board_state[193] ),
    .A1(net49),
    .S(_2739_),
    .X(_0712_));
 sg13g2_nor2_1 _6524_ (.A(net204),
    .B(net243),
    .Y(_2740_));
 sg13g2_mux2_1 _6525_ (.A0(\board_state[194] ),
    .A1(net49),
    .S(_2740_),
    .X(_0713_));
 sg13g2_nor2_1 _6526_ (.A(net203),
    .B(net243),
    .Y(_2741_));
 sg13g2_mux2_1 _6527_ (.A0(\board_state[195] ),
    .A1(net49),
    .S(_2741_),
    .X(_0714_));
 sg13g2_nor2_1 _6528_ (.A(net166),
    .B(_2737_),
    .Y(_2742_));
 sg13g2_mux2_1 _6529_ (.A0(\board_state[196] ),
    .A1(net49),
    .S(_2742_),
    .X(_0715_));
 sg13g2_nor2_1 _6530_ (.A(net165),
    .B(net243),
    .Y(_2743_));
 sg13g2_mux2_1 _6531_ (.A0(\board_state[197] ),
    .A1(net49),
    .S(_2743_),
    .X(_0716_));
 sg13g2_nor2_1 _6532_ (.A(net164),
    .B(net243),
    .Y(_2744_));
 sg13g2_mux2_1 _6533_ (.A0(\board_state[198] ),
    .A1(net49),
    .S(_2744_),
    .X(_0717_));
 sg13g2_nor2_1 _6534_ (.A(net163),
    .B(_2737_),
    .Y(_2745_));
 sg13g2_mux2_1 _6535_ (.A0(\board_state[199] ),
    .A1(net49),
    .S(_2745_),
    .X(_0718_));
 sg13g2_buf_1 _6536_ (.A(_2705_),
    .X(_2746_));
 sg13g2_nor2_1 _6537_ (.A(net203),
    .B(net237),
    .Y(_2747_));
 sg13g2_mux2_1 _6538_ (.A0(\board_state[19] ),
    .A1(_2746_),
    .S(_2747_),
    .X(_0719_));
 sg13g2_nor2_1 _6539_ (.A(net247),
    .B(net205),
    .Y(_2748_));
 sg13g2_mux2_1 _6540_ (.A0(\board_state[1] ),
    .A1(_2746_),
    .S(_2748_),
    .X(_0720_));
 sg13g2_nor2_1 _6541_ (.A(net161),
    .B(net243),
    .Y(_2749_));
 sg13g2_mux2_1 _6542_ (.A0(\board_state[200] ),
    .A1(net48),
    .S(_2749_),
    .X(_0721_));
 sg13g2_nor2_1 _6543_ (.A(net160),
    .B(net243),
    .Y(_2750_));
 sg13g2_mux2_1 _6544_ (.A0(\board_state[201] ),
    .A1(net48),
    .S(_2750_),
    .X(_0722_));
 sg13g2_nor2_1 _6545_ (.A(net167),
    .B(_2736_),
    .Y(_2751_));
 sg13g2_mux2_1 _6546_ (.A0(\board_state[202] ),
    .A1(net48),
    .S(_2751_),
    .X(_0723_));
 sg13g2_nor2_1 _6547_ (.A(net162),
    .B(_2736_),
    .Y(_2752_));
 sg13g2_mux2_1 _6548_ (.A0(\board_state[203] ),
    .A1(net48),
    .S(_2752_),
    .X(_0724_));
 sg13g2_nor2_1 _6549_ (.A(net202),
    .B(_2736_),
    .Y(_2753_));
 sg13g2_mux2_1 _6550_ (.A0(\board_state[204] ),
    .A1(net48),
    .S(_2753_),
    .X(_0725_));
 sg13g2_nor2_1 _6551_ (.A(net159),
    .B(_2736_),
    .Y(_2754_));
 sg13g2_mux2_1 _6552_ (.A0(\board_state[205] ),
    .A1(net48),
    .S(_2754_),
    .X(_0726_));
 sg13g2_nor2_1 _6553_ (.A(net201),
    .B(_2736_),
    .Y(_2755_));
 sg13g2_mux2_1 _6554_ (.A0(\board_state[206] ),
    .A1(net48),
    .S(_2755_),
    .X(_0727_));
 sg13g2_nor2_1 _6555_ (.A(net158),
    .B(_2736_),
    .Y(_2756_));
 sg13g2_mux2_1 _6556_ (.A0(\board_state[207] ),
    .A1(net48),
    .S(_2756_),
    .X(_0728_));
 sg13g2_buf_1 _6557_ (.A(net66),
    .X(_2757_));
 sg13g2_nand2_1 _6558_ (.Y(_2758_),
    .A(net258),
    .B(_2734_));
 sg13g2_buf_1 _6559_ (.A(_2758_),
    .X(_2759_));
 sg13g2_buf_1 _6560_ (.A(_2759_),
    .X(_2760_));
 sg13g2_nor2_1 _6561_ (.A(net207),
    .B(_2760_),
    .Y(_2761_));
 sg13g2_mux2_1 _6562_ (.A0(\board_state[208] ),
    .A1(net47),
    .S(_2761_),
    .X(_0729_));
 sg13g2_nor2_1 _6563_ (.A(net205),
    .B(net235),
    .Y(_2762_));
 sg13g2_mux2_1 _6564_ (.A0(\board_state[209] ),
    .A1(_2757_),
    .S(_2762_),
    .X(_0730_));
 sg13g2_nor2_1 _6565_ (.A(net166),
    .B(net237),
    .Y(_2763_));
 sg13g2_mux2_1 _6566_ (.A0(\board_state[20] ),
    .A1(_2757_),
    .S(_2763_),
    .X(_0731_));
 sg13g2_nor2_1 _6567_ (.A(net204),
    .B(net235),
    .Y(_2764_));
 sg13g2_mux2_1 _6568_ (.A0(\board_state[210] ),
    .A1(net47),
    .S(_2764_),
    .X(_0732_));
 sg13g2_nor2_1 _6569_ (.A(net203),
    .B(net235),
    .Y(_2765_));
 sg13g2_mux2_1 _6570_ (.A0(\board_state[211] ),
    .A1(net47),
    .S(_2765_),
    .X(_0733_));
 sg13g2_nor2_1 _6571_ (.A(net166),
    .B(net235),
    .Y(_2766_));
 sg13g2_mux2_1 _6572_ (.A0(\board_state[212] ),
    .A1(net47),
    .S(_2766_),
    .X(_0734_));
 sg13g2_nor2_1 _6573_ (.A(net165),
    .B(_2760_),
    .Y(_2767_));
 sg13g2_mux2_1 _6574_ (.A0(\board_state[213] ),
    .A1(net47),
    .S(_2767_),
    .X(_0735_));
 sg13g2_nor2_1 _6575_ (.A(net164),
    .B(net235),
    .Y(_2768_));
 sg13g2_mux2_1 _6576_ (.A0(\board_state[214] ),
    .A1(net47),
    .S(_2768_),
    .X(_0736_));
 sg13g2_nor2_1 _6577_ (.A(net163),
    .B(net235),
    .Y(_2769_));
 sg13g2_mux2_1 _6578_ (.A0(\board_state[215] ),
    .A1(net47),
    .S(_2769_),
    .X(_0737_));
 sg13g2_nor2_1 _6579_ (.A(net161),
    .B(net235),
    .Y(_2770_));
 sg13g2_mux2_1 _6580_ (.A0(\board_state[216] ),
    .A1(net47),
    .S(_2770_),
    .X(_0738_));
 sg13g2_buf_1 _6581_ (.A(net66),
    .X(_2771_));
 sg13g2_nor2_1 _6582_ (.A(net160),
    .B(net235),
    .Y(_2772_));
 sg13g2_mux2_1 _6583_ (.A0(\board_state[217] ),
    .A1(net46),
    .S(_2772_),
    .X(_0739_));
 sg13g2_nor2_1 _6584_ (.A(net167),
    .B(_2759_),
    .Y(_2773_));
 sg13g2_mux2_1 _6585_ (.A0(\board_state[218] ),
    .A1(net46),
    .S(_2773_),
    .X(_0740_));
 sg13g2_nor2_1 _6586_ (.A(net162),
    .B(_2759_),
    .Y(_2774_));
 sg13g2_mux2_1 _6587_ (.A0(\board_state[219] ),
    .A1(net46),
    .S(_2774_),
    .X(_0741_));
 sg13g2_nor2_1 _6588_ (.A(net165),
    .B(net237),
    .Y(_2775_));
 sg13g2_mux2_1 _6589_ (.A0(\board_state[21] ),
    .A1(net46),
    .S(_2775_),
    .X(_0742_));
 sg13g2_nor2_1 _6590_ (.A(net202),
    .B(_2759_),
    .Y(_2776_));
 sg13g2_mux2_1 _6591_ (.A0(\board_state[220] ),
    .A1(net46),
    .S(_2776_),
    .X(_0743_));
 sg13g2_nor2_1 _6592_ (.A(net159),
    .B(_2759_),
    .Y(_2777_));
 sg13g2_mux2_1 _6593_ (.A0(\board_state[221] ),
    .A1(net46),
    .S(_2777_),
    .X(_0744_));
 sg13g2_nor2_1 _6594_ (.A(net201),
    .B(_2759_),
    .Y(_2778_));
 sg13g2_mux2_1 _6595_ (.A0(\board_state[222] ),
    .A1(net46),
    .S(_2778_),
    .X(_0745_));
 sg13g2_nor2_1 _6596_ (.A(net158),
    .B(_2759_),
    .Y(_2779_));
 sg13g2_mux2_1 _6597_ (.A0(\board_state[223] ),
    .A1(net46),
    .S(_2779_),
    .X(_0746_));
 sg13g2_nand2_1 _6598_ (.Y(_2780_),
    .A(net316),
    .B(_2734_));
 sg13g2_buf_1 _6599_ (.A(_2780_),
    .X(_2781_));
 sg13g2_buf_1 _6600_ (.A(_2781_),
    .X(_2782_));
 sg13g2_nor2_1 _6601_ (.A(net207),
    .B(net242),
    .Y(_2783_));
 sg13g2_mux2_1 _6602_ (.A0(\board_state[224] ),
    .A1(_2771_),
    .S(_2783_),
    .X(_0747_));
 sg13g2_buf_1 _6603_ (.A(_2581_),
    .X(_2784_));
 sg13g2_nor2_1 _6604_ (.A(net200),
    .B(net242),
    .Y(_2785_));
 sg13g2_mux2_1 _6605_ (.A0(\board_state[225] ),
    .A1(_2771_),
    .S(_2785_),
    .X(_0748_));
 sg13g2_buf_1 _6606_ (.A(net66),
    .X(_2786_));
 sg13g2_buf_1 _6607_ (.A(_2585_),
    .X(_2787_));
 sg13g2_nor2_1 _6608_ (.A(net199),
    .B(net242),
    .Y(_2788_));
 sg13g2_mux2_1 _6609_ (.A0(\board_state[226] ),
    .A1(net45),
    .S(_2788_),
    .X(_0749_));
 sg13g2_buf_1 _6610_ (.A(_2589_),
    .X(_2789_));
 sg13g2_nor2_1 _6611_ (.A(net198),
    .B(net242),
    .Y(_2790_));
 sg13g2_mux2_1 _6612_ (.A0(\board_state[227] ),
    .A1(net45),
    .S(_2790_),
    .X(_0750_));
 sg13g2_nor2_1 _6613_ (.A(net166),
    .B(net242),
    .Y(_2791_));
 sg13g2_mux2_1 _6614_ (.A0(\board_state[228] ),
    .A1(net45),
    .S(_2791_),
    .X(_0751_));
 sg13g2_nor2_1 _6615_ (.A(net165),
    .B(net242),
    .Y(_2792_));
 sg13g2_mux2_1 _6616_ (.A0(\board_state[229] ),
    .A1(net45),
    .S(_2792_),
    .X(_0752_));
 sg13g2_nor2_1 _6617_ (.A(net164),
    .B(_2701_),
    .Y(_2793_));
 sg13g2_mux2_1 _6618_ (.A0(\board_state[22] ),
    .A1(_2786_),
    .S(_2793_),
    .X(_0753_));
 sg13g2_nor2_1 _6619_ (.A(net164),
    .B(net242),
    .Y(_2794_));
 sg13g2_mux2_1 _6620_ (.A0(\board_state[230] ),
    .A1(_2786_),
    .S(_2794_),
    .X(_0754_));
 sg13g2_nor2_1 _6621_ (.A(net163),
    .B(net242),
    .Y(_2795_));
 sg13g2_mux2_1 _6622_ (.A0(\board_state[231] ),
    .A1(net45),
    .S(_2795_),
    .X(_0755_));
 sg13g2_nor2_1 _6623_ (.A(net161),
    .B(_2782_),
    .Y(_2796_));
 sg13g2_mux2_1 _6624_ (.A0(\board_state[232] ),
    .A1(net45),
    .S(_2796_),
    .X(_0756_));
 sg13g2_nor2_1 _6625_ (.A(net160),
    .B(_2782_),
    .Y(_2797_));
 sg13g2_mux2_1 _6626_ (.A0(\board_state[233] ),
    .A1(net45),
    .S(_2797_),
    .X(_0757_));
 sg13g2_nor2_1 _6627_ (.A(net167),
    .B(_2781_),
    .Y(_2798_));
 sg13g2_mux2_1 _6628_ (.A0(\board_state[234] ),
    .A1(net45),
    .S(_2798_),
    .X(_0758_));
 sg13g2_buf_1 _6629_ (.A(net66),
    .X(_2799_));
 sg13g2_nor2_1 _6630_ (.A(net162),
    .B(_2781_),
    .Y(_2800_));
 sg13g2_mux2_1 _6631_ (.A0(\board_state[235] ),
    .A1(net44),
    .S(_2800_),
    .X(_0759_));
 sg13g2_nor2_1 _6632_ (.A(net202),
    .B(_2781_),
    .Y(_2801_));
 sg13g2_mux2_1 _6633_ (.A0(\board_state[236] ),
    .A1(net44),
    .S(_2801_),
    .X(_0760_));
 sg13g2_nor2_1 _6634_ (.A(net159),
    .B(_2781_),
    .Y(_2802_));
 sg13g2_mux2_1 _6635_ (.A0(\board_state[237] ),
    .A1(net44),
    .S(_2802_),
    .X(_0761_));
 sg13g2_nor2_1 _6636_ (.A(net201),
    .B(_2781_),
    .Y(_2803_));
 sg13g2_mux2_1 _6637_ (.A0(\board_state[238] ),
    .A1(_2799_),
    .S(_2803_),
    .X(_0762_));
 sg13g2_nor2_1 _6638_ (.A(net158),
    .B(_2781_),
    .Y(_2804_));
 sg13g2_mux2_1 _6639_ (.A0(\board_state[239] ),
    .A1(_2799_),
    .S(_2804_),
    .X(_0763_));
 sg13g2_nor2_1 _6640_ (.A(_2607_),
    .B(_2701_),
    .Y(_2805_));
 sg13g2_mux2_1 _6641_ (.A0(\board_state[23] ),
    .A1(net44),
    .S(_2805_),
    .X(_0764_));
 sg13g2_buf_1 _6642_ (.A(_2546_),
    .X(_2806_));
 sg13g2_nand2_1 _6643_ (.Y(_2807_),
    .A(net259),
    .B(_2734_));
 sg13g2_buf_1 _6644_ (.A(_2807_),
    .X(_2808_));
 sg13g2_buf_1 _6645_ (.A(_2808_),
    .X(_2809_));
 sg13g2_nor2_1 _6646_ (.A(net197),
    .B(net234),
    .Y(_2810_));
 sg13g2_mux2_1 _6647_ (.A0(\board_state[240] ),
    .A1(net44),
    .S(_2810_),
    .X(_0765_));
 sg13g2_nor2_1 _6648_ (.A(net200),
    .B(net234),
    .Y(_2811_));
 sg13g2_mux2_1 _6649_ (.A0(\board_state[241] ),
    .A1(net44),
    .S(_2811_),
    .X(_0766_));
 sg13g2_nor2_1 _6650_ (.A(net199),
    .B(net234),
    .Y(_2812_));
 sg13g2_mux2_1 _6651_ (.A0(\board_state[242] ),
    .A1(net44),
    .S(_2812_),
    .X(_0767_));
 sg13g2_nor2_1 _6652_ (.A(_2789_),
    .B(net234),
    .Y(_2813_));
 sg13g2_mux2_1 _6653_ (.A0(\board_state[243] ),
    .A1(net44),
    .S(_2813_),
    .X(_0768_));
 sg13g2_buf_1 _6654_ (.A(net66),
    .X(_2814_));
 sg13g2_buf_1 _6655_ (.A(_2593_),
    .X(_2815_));
 sg13g2_nor2_1 _6656_ (.A(net157),
    .B(net234),
    .Y(_2816_));
 sg13g2_mux2_1 _6657_ (.A0(\board_state[244] ),
    .A1(net43),
    .S(_2816_),
    .X(_0769_));
 sg13g2_buf_1 _6658_ (.A(_2597_),
    .X(_2817_));
 sg13g2_nor2_1 _6659_ (.A(net156),
    .B(net234),
    .Y(_2818_));
 sg13g2_mux2_1 _6660_ (.A0(\board_state[245] ),
    .A1(net43),
    .S(_2818_),
    .X(_0770_));
 sg13g2_buf_1 _6661_ (.A(_2602_),
    .X(_2819_));
 sg13g2_nor2_1 _6662_ (.A(_2819_),
    .B(_2809_),
    .Y(_2820_));
 sg13g2_mux2_1 _6663_ (.A0(\board_state[246] ),
    .A1(net43),
    .S(_2820_),
    .X(_0771_));
 sg13g2_buf_1 _6664_ (.A(_2606_),
    .X(_2821_));
 sg13g2_nor2_1 _6665_ (.A(_2821_),
    .B(_2809_),
    .Y(_2822_));
 sg13g2_mux2_1 _6666_ (.A0(\board_state[247] ),
    .A1(net43),
    .S(_2822_),
    .X(_0772_));
 sg13g2_nor2_1 _6667_ (.A(_2615_),
    .B(net234),
    .Y(_2823_));
 sg13g2_mux2_1 _6668_ (.A0(\board_state[248] ),
    .A1(net43),
    .S(_2823_),
    .X(_0773_));
 sg13g2_nor2_1 _6669_ (.A(_2619_),
    .B(net234),
    .Y(_2824_));
 sg13g2_mux2_1 _6670_ (.A0(\board_state[249] ),
    .A1(net43),
    .S(_2824_),
    .X(_0774_));
 sg13g2_buf_1 _6671_ (.A(_2614_),
    .X(_2825_));
 sg13g2_nor2_1 _6672_ (.A(net153),
    .B(net237),
    .Y(_2826_));
 sg13g2_mux2_1 _6673_ (.A0(\board_state[24] ),
    .A1(net43),
    .S(_2826_),
    .X(_0775_));
 sg13g2_nor2_1 _6674_ (.A(_2571_),
    .B(_2808_),
    .Y(_2827_));
 sg13g2_mux2_1 _6675_ (.A0(\board_state[250] ),
    .A1(_2814_),
    .S(_2827_),
    .X(_0776_));
 sg13g2_nor2_1 _6676_ (.A(_2611_),
    .B(_2808_),
    .Y(_2828_));
 sg13g2_mux2_1 _6677_ (.A0(\board_state[251] ),
    .A1(_2814_),
    .S(_2828_),
    .X(_0777_));
 sg13g2_nor2_1 _6678_ (.A(net202),
    .B(_2808_),
    .Y(_2829_));
 sg13g2_mux2_1 _6679_ (.A0(\board_state[252] ),
    .A1(net43),
    .S(_2829_),
    .X(_0778_));
 sg13g2_buf_1 _6680_ (.A(net66),
    .X(_2830_));
 sg13g2_nor2_1 _6681_ (.A(net159),
    .B(_2808_),
    .Y(_2831_));
 sg13g2_mux2_1 _6682_ (.A0(\board_state[253] ),
    .A1(net42),
    .S(_2831_),
    .X(_0779_));
 sg13g2_nor2_1 _6683_ (.A(net201),
    .B(_2808_),
    .Y(_2832_));
 sg13g2_mux2_1 _6684_ (.A0(\board_state[254] ),
    .A1(_2830_),
    .S(_2832_),
    .X(_0780_));
 sg13g2_nor2_1 _6685_ (.A(net158),
    .B(_2808_),
    .Y(_2833_));
 sg13g2_mux2_1 _6686_ (.A0(\board_state[255] ),
    .A1(_2830_),
    .S(_2833_),
    .X(_0781_));
 sg13g2_nand3_1 _6687_ (.B(net326),
    .C(_2032_),
    .A(net362),
    .Y(_2834_));
 sg13g2_buf_1 _6688_ (.A(_2834_),
    .X(_2835_));
 sg13g2_buf_1 _6689_ (.A(_2835_),
    .X(_2836_));
 sg13g2_nor2_1 _6690_ (.A(net197),
    .B(net256),
    .Y(_2837_));
 sg13g2_mux2_1 _6691_ (.A0(\board_state[256] ),
    .A1(net42),
    .S(_2837_),
    .X(_0782_));
 sg13g2_nor2_1 _6692_ (.A(net200),
    .B(net256),
    .Y(_2838_));
 sg13g2_mux2_1 _6693_ (.A0(\board_state[257] ),
    .A1(net42),
    .S(_2838_),
    .X(_0783_));
 sg13g2_nor2_1 _6694_ (.A(net199),
    .B(net256),
    .Y(_2839_));
 sg13g2_mux2_1 _6695_ (.A0(\board_state[258] ),
    .A1(net42),
    .S(_2839_),
    .X(_0784_));
 sg13g2_nor2_1 _6696_ (.A(net198),
    .B(_2836_),
    .Y(_2840_));
 sg13g2_mux2_1 _6697_ (.A0(\board_state[259] ),
    .A1(net42),
    .S(_2840_),
    .X(_0785_));
 sg13g2_buf_1 _6698_ (.A(_2618_),
    .X(_2841_));
 sg13g2_nor2_1 _6699_ (.A(net152),
    .B(net237),
    .Y(_2842_));
 sg13g2_mux2_1 _6700_ (.A0(\board_state[25] ),
    .A1(net42),
    .S(_2842_),
    .X(_0786_));
 sg13g2_nor2_1 _6701_ (.A(net157),
    .B(net256),
    .Y(_2843_));
 sg13g2_mux2_1 _6702_ (.A0(\board_state[260] ),
    .A1(net42),
    .S(_2843_),
    .X(_0787_));
 sg13g2_nor2_1 _6703_ (.A(net156),
    .B(net256),
    .Y(_2844_));
 sg13g2_mux2_1 _6704_ (.A0(\board_state[261] ),
    .A1(net42),
    .S(_2844_),
    .X(_0788_));
 sg13g2_buf_1 _6705_ (.A(_2533_),
    .X(_2845_));
 sg13g2_buf_1 _6706_ (.A(_2845_),
    .X(_2846_));
 sg13g2_nor2_1 _6707_ (.A(net155),
    .B(net256),
    .Y(_2847_));
 sg13g2_mux2_1 _6708_ (.A0(\board_state[262] ),
    .A1(_2846_),
    .S(_2847_),
    .X(_0789_));
 sg13g2_nor2_1 _6709_ (.A(net154),
    .B(_2836_),
    .Y(_2848_));
 sg13g2_mux2_1 _6710_ (.A0(\board_state[263] ),
    .A1(net41),
    .S(_2848_),
    .X(_0790_));
 sg13g2_nor2_1 _6711_ (.A(net153),
    .B(net256),
    .Y(_2849_));
 sg13g2_mux2_1 _6712_ (.A0(\board_state[264] ),
    .A1(net41),
    .S(_2849_),
    .X(_0791_));
 sg13g2_nor2_1 _6713_ (.A(net152),
    .B(net256),
    .Y(_2850_));
 sg13g2_mux2_1 _6714_ (.A0(\board_state[265] ),
    .A1(net41),
    .S(_2850_),
    .X(_0792_));
 sg13g2_buf_1 _6715_ (.A(_2570_),
    .X(_2851_));
 sg13g2_nor2_1 _6716_ (.A(net151),
    .B(_2835_),
    .Y(_2852_));
 sg13g2_mux2_1 _6717_ (.A0(\board_state[266] ),
    .A1(net41),
    .S(_2852_),
    .X(_0793_));
 sg13g2_buf_1 _6718_ (.A(_2610_),
    .X(_2853_));
 sg13g2_nor2_1 _6719_ (.A(net150),
    .B(_2835_),
    .Y(_2854_));
 sg13g2_mux2_1 _6720_ (.A0(\board_state[267] ),
    .A1(net41),
    .S(_2854_),
    .X(_0794_));
 sg13g2_buf_1 _6721_ (.A(_2624_),
    .X(_2855_));
 sg13g2_nor2_1 _6722_ (.A(net196),
    .B(_2835_),
    .Y(_2856_));
 sg13g2_mux2_1 _6723_ (.A0(\board_state[268] ),
    .A1(net41),
    .S(_2856_),
    .X(_0795_));
 sg13g2_buf_1 _6724_ (.A(_2628_),
    .X(_2857_));
 sg13g2_nor2_1 _6725_ (.A(net149),
    .B(_2835_),
    .Y(_2858_));
 sg13g2_mux2_1 _6726_ (.A0(\board_state[269] ),
    .A1(net41),
    .S(_2858_),
    .X(_0796_));
 sg13g2_nor2_1 _6727_ (.A(net151),
    .B(_2700_),
    .Y(_2859_));
 sg13g2_mux2_1 _6728_ (.A0(\board_state[26] ),
    .A1(_2846_),
    .S(_2859_),
    .X(_0797_));
 sg13g2_buf_1 _6729_ (.A(_2632_),
    .X(_2860_));
 sg13g2_nor2_1 _6730_ (.A(net195),
    .B(_2835_),
    .Y(_2861_));
 sg13g2_mux2_1 _6731_ (.A0(\board_state[270] ),
    .A1(net41),
    .S(_2861_),
    .X(_0798_));
 sg13g2_buf_1 _6732_ (.A(net65),
    .X(_2862_));
 sg13g2_buf_1 _6733_ (.A(_2637_),
    .X(_2863_));
 sg13g2_nor2_1 _6734_ (.A(net148),
    .B(_2835_),
    .Y(_2864_));
 sg13g2_mux2_1 _6735_ (.A0(\board_state[271] ),
    .A1(_2862_),
    .S(_2864_),
    .X(_0799_));
 sg13g2_nand3_1 _6736_ (.B(_2032_),
    .C(net258),
    .A(net362),
    .Y(_2865_));
 sg13g2_buf_1 _6737_ (.A(_2865_),
    .X(_2866_));
 sg13g2_buf_1 _6738_ (.A(_2866_),
    .X(_2867_));
 sg13g2_nor2_1 _6739_ (.A(net197),
    .B(net233),
    .Y(_2868_));
 sg13g2_mux2_1 _6740_ (.A0(\board_state[272] ),
    .A1(net40),
    .S(_2868_),
    .X(_0800_));
 sg13g2_nor2_1 _6741_ (.A(net200),
    .B(net233),
    .Y(_2869_));
 sg13g2_mux2_1 _6742_ (.A0(\board_state[273] ),
    .A1(net40),
    .S(_2869_),
    .X(_0801_));
 sg13g2_nor2_1 _6743_ (.A(net199),
    .B(net233),
    .Y(_2870_));
 sg13g2_mux2_1 _6744_ (.A0(\board_state[274] ),
    .A1(net40),
    .S(_2870_),
    .X(_0802_));
 sg13g2_nor2_1 _6745_ (.A(_2789_),
    .B(net233),
    .Y(_2871_));
 sg13g2_mux2_1 _6746_ (.A0(\board_state[275] ),
    .A1(net40),
    .S(_2871_),
    .X(_0803_));
 sg13g2_nor2_1 _6747_ (.A(_2815_),
    .B(net233),
    .Y(_2872_));
 sg13g2_mux2_1 _6748_ (.A0(\board_state[276] ),
    .A1(net40),
    .S(_2872_),
    .X(_0804_));
 sg13g2_nor2_1 _6749_ (.A(_2817_),
    .B(net233),
    .Y(_2873_));
 sg13g2_mux2_1 _6750_ (.A0(\board_state[277] ),
    .A1(net40),
    .S(_2873_),
    .X(_0805_));
 sg13g2_nor2_1 _6751_ (.A(net155),
    .B(_2867_),
    .Y(_2874_));
 sg13g2_mux2_1 _6752_ (.A0(\board_state[278] ),
    .A1(net40),
    .S(_2874_),
    .X(_0806_));
 sg13g2_nor2_1 _6753_ (.A(net154),
    .B(_2867_),
    .Y(_2875_));
 sg13g2_mux2_1 _6754_ (.A0(\board_state[279] ),
    .A1(net40),
    .S(_2875_),
    .X(_0807_));
 sg13g2_nor2_1 _6755_ (.A(net150),
    .B(_2700_),
    .Y(_2876_));
 sg13g2_mux2_1 _6756_ (.A0(\board_state[27] ),
    .A1(_2862_),
    .S(_2876_),
    .X(_0808_));
 sg13g2_buf_1 _6757_ (.A(net65),
    .X(_2877_));
 sg13g2_nor2_1 _6758_ (.A(net153),
    .B(net233),
    .Y(_2878_));
 sg13g2_mux2_1 _6759_ (.A0(\board_state[280] ),
    .A1(net39),
    .S(_2878_),
    .X(_0809_));
 sg13g2_nor2_1 _6760_ (.A(net152),
    .B(net233),
    .Y(_2879_));
 sg13g2_mux2_1 _6761_ (.A0(\board_state[281] ),
    .A1(net39),
    .S(_2879_),
    .X(_0810_));
 sg13g2_nor2_1 _6762_ (.A(net151),
    .B(_2866_),
    .Y(_2880_));
 sg13g2_mux2_1 _6763_ (.A0(\board_state[282] ),
    .A1(net39),
    .S(_2880_),
    .X(_0811_));
 sg13g2_nor2_1 _6764_ (.A(net150),
    .B(_2866_),
    .Y(_2881_));
 sg13g2_mux2_1 _6765_ (.A0(\board_state[283] ),
    .A1(net39),
    .S(_2881_),
    .X(_0812_));
 sg13g2_nor2_1 _6766_ (.A(net196),
    .B(_2866_),
    .Y(_2882_));
 sg13g2_mux2_1 _6767_ (.A0(\board_state[284] ),
    .A1(net39),
    .S(_2882_),
    .X(_0813_));
 sg13g2_nor2_1 _6768_ (.A(net149),
    .B(_2866_),
    .Y(_2883_));
 sg13g2_mux2_1 _6769_ (.A0(\board_state[285] ),
    .A1(net39),
    .S(_2883_),
    .X(_0814_));
 sg13g2_nor2_1 _6770_ (.A(net195),
    .B(_2866_),
    .Y(_2884_));
 sg13g2_mux2_1 _6771_ (.A0(\board_state[286] ),
    .A1(net39),
    .S(_2884_),
    .X(_0815_));
 sg13g2_nor2_1 _6772_ (.A(net148),
    .B(_2866_),
    .Y(_2885_));
 sg13g2_mux2_1 _6773_ (.A0(\board_state[287] ),
    .A1(_2877_),
    .S(_2885_),
    .X(_0816_));
 sg13g2_nand3_1 _6774_ (.B(_2032_),
    .C(net316),
    .A(net362),
    .Y(_2886_));
 sg13g2_buf_1 _6775_ (.A(_2886_),
    .X(_2887_));
 sg13g2_buf_1 _6776_ (.A(_2887_),
    .X(_2888_));
 sg13g2_nor2_1 _6777_ (.A(net197),
    .B(net255),
    .Y(_2889_));
 sg13g2_mux2_1 _6778_ (.A0(\board_state[288] ),
    .A1(net39),
    .S(_2889_),
    .X(_0817_));
 sg13g2_nor2_1 _6779_ (.A(net200),
    .B(net255),
    .Y(_2890_));
 sg13g2_mux2_1 _6780_ (.A0(\board_state[289] ),
    .A1(_2877_),
    .S(_2890_),
    .X(_0818_));
 sg13g2_buf_1 _6781_ (.A(net65),
    .X(_2891_));
 sg13g2_nor2_1 _6782_ (.A(net196),
    .B(_2700_),
    .Y(_2892_));
 sg13g2_mux2_1 _6783_ (.A0(\board_state[28] ),
    .A1(_2891_),
    .S(_2892_),
    .X(_0819_));
 sg13g2_nor2_1 _6784_ (.A(net199),
    .B(net255),
    .Y(_2893_));
 sg13g2_mux2_1 _6785_ (.A0(\board_state[290] ),
    .A1(net38),
    .S(_2893_),
    .X(_0820_));
 sg13g2_nor2_1 _6786_ (.A(net198),
    .B(net255),
    .Y(_2894_));
 sg13g2_mux2_1 _6787_ (.A0(\board_state[291] ),
    .A1(net38),
    .S(_2894_),
    .X(_0821_));
 sg13g2_nor2_1 _6788_ (.A(_2815_),
    .B(net255),
    .Y(_2895_));
 sg13g2_mux2_1 _6789_ (.A0(\board_state[292] ),
    .A1(net38),
    .S(_2895_),
    .X(_0822_));
 sg13g2_nor2_1 _6790_ (.A(_2817_),
    .B(net255),
    .Y(_2896_));
 sg13g2_mux2_1 _6791_ (.A0(\board_state[293] ),
    .A1(_2891_),
    .S(_2896_),
    .X(_0823_));
 sg13g2_nor2_1 _6792_ (.A(net155),
    .B(_2888_),
    .Y(_2897_));
 sg13g2_mux2_1 _6793_ (.A0(\board_state[294] ),
    .A1(net38),
    .S(_2897_),
    .X(_0824_));
 sg13g2_nor2_1 _6794_ (.A(net154),
    .B(_2888_),
    .Y(_2898_));
 sg13g2_mux2_1 _6795_ (.A0(\board_state[295] ),
    .A1(net38),
    .S(_2898_),
    .X(_0825_));
 sg13g2_nor2_1 _6796_ (.A(net153),
    .B(net255),
    .Y(_2899_));
 sg13g2_mux2_1 _6797_ (.A0(\board_state[296] ),
    .A1(net38),
    .S(_2899_),
    .X(_0826_));
 sg13g2_nor2_1 _6798_ (.A(net152),
    .B(net255),
    .Y(_2900_));
 sg13g2_mux2_1 _6799_ (.A0(\board_state[297] ),
    .A1(net38),
    .S(_2900_),
    .X(_0827_));
 sg13g2_nor2_1 _6800_ (.A(_2851_),
    .B(_2887_),
    .Y(_2901_));
 sg13g2_mux2_1 _6801_ (.A0(\board_state[298] ),
    .A1(net38),
    .S(_2901_),
    .X(_0828_));
 sg13g2_buf_1 _6802_ (.A(_2845_),
    .X(_2902_));
 sg13g2_nor2_1 _6803_ (.A(_2853_),
    .B(_2887_),
    .Y(_2903_));
 sg13g2_mux2_1 _6804_ (.A0(\board_state[299] ),
    .A1(net37),
    .S(_2903_),
    .X(_0829_));
 sg13g2_nor2_1 _6805_ (.A(net149),
    .B(_2700_),
    .Y(_2904_));
 sg13g2_mux2_1 _6806_ (.A0(\board_state[29] ),
    .A1(_2902_),
    .S(_2904_),
    .X(_0830_));
 sg13g2_nor2_1 _6807_ (.A(net247),
    .B(_2586_),
    .Y(_2905_));
 sg13g2_mux2_1 _6808_ (.A0(\board_state[2] ),
    .A1(_2902_),
    .S(_2905_),
    .X(_0831_));
 sg13g2_nor2_1 _6809_ (.A(_2855_),
    .B(_2887_),
    .Y(_2906_));
 sg13g2_mux2_1 _6810_ (.A0(\board_state[300] ),
    .A1(net37),
    .S(_2906_),
    .X(_0832_));
 sg13g2_nor2_1 _6811_ (.A(_2857_),
    .B(_2887_),
    .Y(_2907_));
 sg13g2_mux2_1 _6812_ (.A0(\board_state[301] ),
    .A1(net37),
    .S(_2907_),
    .X(_0833_));
 sg13g2_nor2_1 _6813_ (.A(_2860_),
    .B(_2887_),
    .Y(_2908_));
 sg13g2_mux2_1 _6814_ (.A0(\board_state[302] ),
    .A1(net37),
    .S(_2908_),
    .X(_0834_));
 sg13g2_nor2_1 _6815_ (.A(net148),
    .B(_2887_),
    .Y(_2909_));
 sg13g2_mux2_1 _6816_ (.A0(\board_state[303] ),
    .A1(net37),
    .S(_2909_),
    .X(_0835_));
 sg13g2_nand3_1 _6817_ (.B(_2032_),
    .C(net259),
    .A(net362),
    .Y(_2910_));
 sg13g2_buf_1 _6818_ (.A(_2910_),
    .X(_2911_));
 sg13g2_buf_1 _6819_ (.A(_2911_),
    .X(_2912_));
 sg13g2_nor2_1 _6820_ (.A(net197),
    .B(_2912_),
    .Y(_2913_));
 sg13g2_mux2_1 _6821_ (.A0(\board_state[304] ),
    .A1(net37),
    .S(_2913_),
    .X(_0836_));
 sg13g2_nor2_1 _6822_ (.A(_2784_),
    .B(net232),
    .Y(_2914_));
 sg13g2_mux2_1 _6823_ (.A0(\board_state[305] ),
    .A1(net37),
    .S(_2914_),
    .X(_0837_));
 sg13g2_nor2_1 _6824_ (.A(_2787_),
    .B(net232),
    .Y(_2915_));
 sg13g2_mux2_1 _6825_ (.A0(\board_state[306] ),
    .A1(net37),
    .S(_2915_),
    .X(_0838_));
 sg13g2_buf_1 _6826_ (.A(net65),
    .X(_2916_));
 sg13g2_nor2_1 _6827_ (.A(net198),
    .B(net232),
    .Y(_2917_));
 sg13g2_mux2_1 _6828_ (.A0(\board_state[307] ),
    .A1(net36),
    .S(_2917_),
    .X(_0839_));
 sg13g2_nor2_1 _6829_ (.A(net157),
    .B(net232),
    .Y(_2918_));
 sg13g2_mux2_1 _6830_ (.A0(\board_state[308] ),
    .A1(net36),
    .S(_2918_),
    .X(_0840_));
 sg13g2_nor2_1 _6831_ (.A(net156),
    .B(net232),
    .Y(_2919_));
 sg13g2_mux2_1 _6832_ (.A0(\board_state[309] ),
    .A1(net36),
    .S(_2919_),
    .X(_0841_));
 sg13g2_nor2_1 _6833_ (.A(net195),
    .B(_2700_),
    .Y(_2920_));
 sg13g2_mux2_1 _6834_ (.A0(\board_state[30] ),
    .A1(_2916_),
    .S(_2920_),
    .X(_0842_));
 sg13g2_nor2_1 _6835_ (.A(net155),
    .B(_2912_),
    .Y(_2921_));
 sg13g2_mux2_1 _6836_ (.A0(\board_state[310] ),
    .A1(_2916_),
    .S(_2921_),
    .X(_0843_));
 sg13g2_nor2_1 _6837_ (.A(net154),
    .B(net232),
    .Y(_2922_));
 sg13g2_mux2_1 _6838_ (.A0(\board_state[311] ),
    .A1(net36),
    .S(_2922_),
    .X(_0844_));
 sg13g2_nor2_1 _6839_ (.A(net153),
    .B(net232),
    .Y(_2923_));
 sg13g2_mux2_1 _6840_ (.A0(\board_state[312] ),
    .A1(net36),
    .S(_2923_),
    .X(_0845_));
 sg13g2_nor2_1 _6841_ (.A(net152),
    .B(net232),
    .Y(_2924_));
 sg13g2_mux2_1 _6842_ (.A0(\board_state[313] ),
    .A1(net36),
    .S(_2924_),
    .X(_0846_));
 sg13g2_nor2_1 _6843_ (.A(net151),
    .B(_2911_),
    .Y(_2925_));
 sg13g2_mux2_1 _6844_ (.A0(\board_state[314] ),
    .A1(net36),
    .S(_2925_),
    .X(_0847_));
 sg13g2_nor2_1 _6845_ (.A(net150),
    .B(_2911_),
    .Y(_2926_));
 sg13g2_mux2_1 _6846_ (.A0(\board_state[315] ),
    .A1(net36),
    .S(_2926_),
    .X(_0848_));
 sg13g2_buf_1 _6847_ (.A(net65),
    .X(_2927_));
 sg13g2_nor2_1 _6848_ (.A(net196),
    .B(_2911_),
    .Y(_2928_));
 sg13g2_mux2_1 _6849_ (.A0(\board_state[316] ),
    .A1(net35),
    .S(_2928_),
    .X(_0849_));
 sg13g2_nor2_1 _6850_ (.A(net149),
    .B(_2911_),
    .Y(_2929_));
 sg13g2_mux2_1 _6851_ (.A0(\board_state[317] ),
    .A1(_2927_),
    .S(_2929_),
    .X(_0850_));
 sg13g2_nor2_1 _6852_ (.A(net195),
    .B(_2911_),
    .Y(_2930_));
 sg13g2_mux2_1 _6853_ (.A0(\board_state[318] ),
    .A1(net35),
    .S(_2930_),
    .X(_0851_));
 sg13g2_nor2_1 _6854_ (.A(net148),
    .B(_2911_),
    .Y(_2931_));
 sg13g2_mux2_1 _6855_ (.A0(\board_state[319] ),
    .A1(net35),
    .S(_2931_),
    .X(_0852_));
 sg13g2_nor2_1 _6856_ (.A(_2863_),
    .B(_2700_),
    .Y(_2932_));
 sg13g2_mux2_1 _6857_ (.A0(\board_state[31] ),
    .A1(_2927_),
    .S(_2932_),
    .X(_0853_));
 sg13g2_nor3_2 _6858_ (.A(net394),
    .B(_2390_),
    .C(_2551_),
    .Y(_2933_));
 sg13g2_nand2_1 _6859_ (.Y(_2934_),
    .A(net326),
    .B(_2933_));
 sg13g2_buf_1 _6860_ (.A(_2934_),
    .X(_2935_));
 sg13g2_buf_1 _6861_ (.A(_2935_),
    .X(_2936_));
 sg13g2_nor2_1 _6862_ (.A(net197),
    .B(net254),
    .Y(_2937_));
 sg13g2_mux2_1 _6863_ (.A0(\board_state[320] ),
    .A1(net35),
    .S(_2937_),
    .X(_0854_));
 sg13g2_nor2_1 _6864_ (.A(net200),
    .B(net254),
    .Y(_2938_));
 sg13g2_mux2_1 _6865_ (.A0(\board_state[321] ),
    .A1(net35),
    .S(_2938_),
    .X(_0855_));
 sg13g2_nor2_1 _6866_ (.A(net199),
    .B(_2936_),
    .Y(_2939_));
 sg13g2_mux2_1 _6867_ (.A0(\board_state[322] ),
    .A1(net35),
    .S(_2939_),
    .X(_0856_));
 sg13g2_nor2_1 _6868_ (.A(net198),
    .B(_2936_),
    .Y(_2940_));
 sg13g2_mux2_1 _6869_ (.A0(\board_state[323] ),
    .A1(net35),
    .S(_2940_),
    .X(_0857_));
 sg13g2_nor2_1 _6870_ (.A(net157),
    .B(net254),
    .Y(_2941_));
 sg13g2_mux2_1 _6871_ (.A0(\board_state[324] ),
    .A1(net35),
    .S(_2941_),
    .X(_0858_));
 sg13g2_buf_1 _6872_ (.A(net65),
    .X(_2942_));
 sg13g2_nor2_1 _6873_ (.A(net156),
    .B(net254),
    .Y(_2943_));
 sg13g2_mux2_1 _6874_ (.A0(\board_state[325] ),
    .A1(net34),
    .S(_2943_),
    .X(_0859_));
 sg13g2_nor2_1 _6875_ (.A(net155),
    .B(net254),
    .Y(_2944_));
 sg13g2_mux2_1 _6876_ (.A0(\board_state[326] ),
    .A1(net34),
    .S(_2944_),
    .X(_0860_));
 sg13g2_nor2_1 _6877_ (.A(net154),
    .B(net254),
    .Y(_2945_));
 sg13g2_mux2_1 _6878_ (.A0(\board_state[327] ),
    .A1(_2942_),
    .S(_2945_),
    .X(_0861_));
 sg13g2_nor2_1 _6879_ (.A(net153),
    .B(net254),
    .Y(_2946_));
 sg13g2_mux2_1 _6880_ (.A0(\board_state[328] ),
    .A1(net34),
    .S(_2946_),
    .X(_0862_));
 sg13g2_nor2_1 _6881_ (.A(net152),
    .B(net254),
    .Y(_2947_));
 sg13g2_mux2_1 _6882_ (.A0(\board_state[329] ),
    .A1(net34),
    .S(_2947_),
    .X(_0863_));
 sg13g2_nand2_1 _6883_ (.Y(_2948_),
    .A(_2537_),
    .B(net316));
 sg13g2_buf_2 _6884_ (.A(_2948_),
    .X(_2949_));
 sg13g2_buf_1 _6885_ (.A(_2949_),
    .X(_2950_));
 sg13g2_nor2_1 _6886_ (.A(_2806_),
    .B(net241),
    .Y(_2951_));
 sg13g2_mux2_1 _6887_ (.A0(\board_state[32] ),
    .A1(_2942_),
    .S(_2951_),
    .X(_0864_));
 sg13g2_nor2_1 _6888_ (.A(net151),
    .B(_2935_),
    .Y(_2952_));
 sg13g2_mux2_1 _6889_ (.A0(\board_state[330] ),
    .A1(net34),
    .S(_2952_),
    .X(_0865_));
 sg13g2_nor2_1 _6890_ (.A(net150),
    .B(_2935_),
    .Y(_2953_));
 sg13g2_mux2_1 _6891_ (.A0(\board_state[331] ),
    .A1(net34),
    .S(_2953_),
    .X(_0866_));
 sg13g2_nor2_1 _6892_ (.A(net196),
    .B(_2935_),
    .Y(_2954_));
 sg13g2_mux2_1 _6893_ (.A0(\board_state[332] ),
    .A1(net34),
    .S(_2954_),
    .X(_0867_));
 sg13g2_nor2_1 _6894_ (.A(net149),
    .B(_2935_),
    .Y(_2955_));
 sg13g2_mux2_1 _6895_ (.A0(\board_state[333] ),
    .A1(net34),
    .S(_2955_),
    .X(_0868_));
 sg13g2_buf_1 _6896_ (.A(net65),
    .X(_2956_));
 sg13g2_nor2_1 _6897_ (.A(net195),
    .B(_2935_),
    .Y(_2957_));
 sg13g2_mux2_1 _6898_ (.A0(\board_state[334] ),
    .A1(net33),
    .S(_2957_),
    .X(_0869_));
 sg13g2_nor2_1 _6899_ (.A(net148),
    .B(_2935_),
    .Y(_2958_));
 sg13g2_mux2_1 _6900_ (.A0(\board_state[335] ),
    .A1(net33),
    .S(_2958_),
    .X(_0870_));
 sg13g2_nand2_1 _6901_ (.Y(_2959_),
    .A(net258),
    .B(_2933_));
 sg13g2_buf_2 _6902_ (.A(_2959_),
    .X(_2960_));
 sg13g2_buf_1 _6903_ (.A(_2960_),
    .X(_2961_));
 sg13g2_nor2_1 _6904_ (.A(net197),
    .B(net231),
    .Y(_2962_));
 sg13g2_mux2_1 _6905_ (.A0(\board_state[336] ),
    .A1(net33),
    .S(_2962_),
    .X(_0871_));
 sg13g2_nor2_1 _6906_ (.A(net200),
    .B(net231),
    .Y(_2963_));
 sg13g2_mux2_1 _6907_ (.A0(\board_state[337] ),
    .A1(_2956_),
    .S(_2963_),
    .X(_0872_));
 sg13g2_nor2_1 _6908_ (.A(net199),
    .B(net231),
    .Y(_2964_));
 sg13g2_mux2_1 _6909_ (.A0(\board_state[338] ),
    .A1(net33),
    .S(_2964_),
    .X(_0873_));
 sg13g2_nor2_1 _6910_ (.A(net198),
    .B(net231),
    .Y(_2965_));
 sg13g2_mux2_1 _6911_ (.A0(\board_state[339] ),
    .A1(net33),
    .S(_2965_),
    .X(_0874_));
 sg13g2_nor2_1 _6912_ (.A(_2784_),
    .B(net241),
    .Y(_2966_));
 sg13g2_mux2_1 _6913_ (.A0(\board_state[33] ),
    .A1(_2956_),
    .S(_2966_),
    .X(_0875_));
 sg13g2_nor2_1 _6914_ (.A(net157),
    .B(_2961_),
    .Y(_2967_));
 sg13g2_mux2_1 _6915_ (.A0(\board_state[340] ),
    .A1(net33),
    .S(_2967_),
    .X(_0876_));
 sg13g2_nor2_1 _6916_ (.A(net156),
    .B(net231),
    .Y(_2968_));
 sg13g2_mux2_1 _6917_ (.A0(\board_state[341] ),
    .A1(net33),
    .S(_2968_),
    .X(_0877_));
 sg13g2_nor2_1 _6918_ (.A(net155),
    .B(net231),
    .Y(_2969_));
 sg13g2_mux2_1 _6919_ (.A0(\board_state[342] ),
    .A1(net33),
    .S(_2969_),
    .X(_0878_));
 sg13g2_buf_1 _6920_ (.A(net65),
    .X(_2970_));
 sg13g2_nor2_1 _6921_ (.A(net154),
    .B(_2961_),
    .Y(_2971_));
 sg13g2_mux2_1 _6922_ (.A0(\board_state[343] ),
    .A1(net32),
    .S(_2971_),
    .X(_0879_));
 sg13g2_nor2_1 _6923_ (.A(net153),
    .B(net231),
    .Y(_2972_));
 sg13g2_mux2_1 _6924_ (.A0(\board_state[344] ),
    .A1(net32),
    .S(_2972_),
    .X(_0880_));
 sg13g2_nor2_1 _6925_ (.A(net152),
    .B(net231),
    .Y(_2973_));
 sg13g2_mux2_1 _6926_ (.A0(\board_state[345] ),
    .A1(_2970_),
    .S(_2973_),
    .X(_0881_));
 sg13g2_nor2_1 _6927_ (.A(net151),
    .B(_2960_),
    .Y(_2974_));
 sg13g2_mux2_1 _6928_ (.A0(\board_state[346] ),
    .A1(net32),
    .S(_2974_),
    .X(_0882_));
 sg13g2_nor2_1 _6929_ (.A(net150),
    .B(_2960_),
    .Y(_2975_));
 sg13g2_mux2_1 _6930_ (.A0(\board_state[347] ),
    .A1(net32),
    .S(_2975_),
    .X(_0883_));
 sg13g2_nor2_1 _6931_ (.A(net196),
    .B(_2960_),
    .Y(_2976_));
 sg13g2_mux2_1 _6932_ (.A0(\board_state[348] ),
    .A1(net32),
    .S(_2976_),
    .X(_0884_));
 sg13g2_nor2_1 _6933_ (.A(net149),
    .B(_2960_),
    .Y(_2977_));
 sg13g2_mux2_1 _6934_ (.A0(\board_state[349] ),
    .A1(net32),
    .S(_2977_),
    .X(_0885_));
 sg13g2_nor2_1 _6935_ (.A(_2787_),
    .B(net241),
    .Y(_2978_));
 sg13g2_mux2_1 _6936_ (.A0(\board_state[34] ),
    .A1(_2970_),
    .S(_2978_),
    .X(_0886_));
 sg13g2_nor2_1 _6937_ (.A(net195),
    .B(_2960_),
    .Y(_2979_));
 sg13g2_mux2_1 _6938_ (.A0(\board_state[350] ),
    .A1(net32),
    .S(_2979_),
    .X(_0887_));
 sg13g2_nor2_1 _6939_ (.A(net148),
    .B(_2960_),
    .Y(_2980_));
 sg13g2_mux2_1 _6940_ (.A0(\board_state[351] ),
    .A1(net32),
    .S(_2980_),
    .X(_0888_));
 sg13g2_buf_1 _6941_ (.A(_2533_),
    .X(_2981_));
 sg13g2_buf_1 _6942_ (.A(net64),
    .X(_2982_));
 sg13g2_nand2_1 _6943_ (.Y(_2983_),
    .A(net316),
    .B(_2933_));
 sg13g2_buf_1 _6944_ (.A(_2983_),
    .X(_2984_));
 sg13g2_buf_1 _6945_ (.A(_2984_),
    .X(_2985_));
 sg13g2_nor2_1 _6946_ (.A(net197),
    .B(net253),
    .Y(_2986_));
 sg13g2_mux2_1 _6947_ (.A0(\board_state[352] ),
    .A1(net31),
    .S(_2986_),
    .X(_0889_));
 sg13g2_nor2_1 _6948_ (.A(net200),
    .B(_2985_),
    .Y(_2987_));
 sg13g2_mux2_1 _6949_ (.A0(\board_state[353] ),
    .A1(net31),
    .S(_2987_),
    .X(_0890_));
 sg13g2_nor2_1 _6950_ (.A(net199),
    .B(_2985_),
    .Y(_2988_));
 sg13g2_mux2_1 _6951_ (.A0(\board_state[354] ),
    .A1(net31),
    .S(_2988_),
    .X(_0891_));
 sg13g2_nor2_1 _6952_ (.A(net198),
    .B(net253),
    .Y(_2989_));
 sg13g2_mux2_1 _6953_ (.A0(\board_state[355] ),
    .A1(net31),
    .S(_2989_),
    .X(_0892_));
 sg13g2_nor2_1 _6954_ (.A(net157),
    .B(net253),
    .Y(_2990_));
 sg13g2_mux2_1 _6955_ (.A0(\board_state[356] ),
    .A1(net31),
    .S(_2990_),
    .X(_0893_));
 sg13g2_nor2_1 _6956_ (.A(net156),
    .B(net253),
    .Y(_2991_));
 sg13g2_mux2_1 _6957_ (.A0(\board_state[357] ),
    .A1(net31),
    .S(_2991_),
    .X(_0894_));
 sg13g2_nor2_1 _6958_ (.A(net155),
    .B(net253),
    .Y(_2992_));
 sg13g2_mux2_1 _6959_ (.A0(\board_state[358] ),
    .A1(net31),
    .S(_2992_),
    .X(_0895_));
 sg13g2_nor2_1 _6960_ (.A(net154),
    .B(net253),
    .Y(_2993_));
 sg13g2_mux2_1 _6961_ (.A0(\board_state[359] ),
    .A1(net31),
    .S(_2993_),
    .X(_0896_));
 sg13g2_nor2_1 _6962_ (.A(net198),
    .B(net241),
    .Y(_2994_));
 sg13g2_mux2_1 _6963_ (.A0(\board_state[35] ),
    .A1(_2982_),
    .S(_2994_),
    .X(_0897_));
 sg13g2_nor2_1 _6964_ (.A(_2825_),
    .B(net253),
    .Y(_2995_));
 sg13g2_mux2_1 _6965_ (.A0(\board_state[360] ),
    .A1(_2982_),
    .S(_2995_),
    .X(_0898_));
 sg13g2_buf_1 _6966_ (.A(net64),
    .X(_2996_));
 sg13g2_nor2_1 _6967_ (.A(net152),
    .B(net253),
    .Y(_2997_));
 sg13g2_mux2_1 _6968_ (.A0(\board_state[361] ),
    .A1(net30),
    .S(_2997_),
    .X(_0899_));
 sg13g2_nor2_1 _6969_ (.A(_2851_),
    .B(_2984_),
    .Y(_2998_));
 sg13g2_mux2_1 _6970_ (.A0(\board_state[362] ),
    .A1(net30),
    .S(_2998_),
    .X(_0900_));
 sg13g2_nor2_1 _6971_ (.A(_2853_),
    .B(_2984_),
    .Y(_2999_));
 sg13g2_mux2_1 _6972_ (.A0(\board_state[363] ),
    .A1(net30),
    .S(_2999_),
    .X(_0901_));
 sg13g2_nor2_1 _6973_ (.A(net196),
    .B(_2984_),
    .Y(_3000_));
 sg13g2_mux2_1 _6974_ (.A0(\board_state[364] ),
    .A1(net30),
    .S(_3000_),
    .X(_0902_));
 sg13g2_nor2_1 _6975_ (.A(net149),
    .B(_2984_),
    .Y(_3001_));
 sg13g2_mux2_1 _6976_ (.A0(\board_state[365] ),
    .A1(net30),
    .S(_3001_),
    .X(_0903_));
 sg13g2_nor2_1 _6977_ (.A(net195),
    .B(_2984_),
    .Y(_3002_));
 sg13g2_mux2_1 _6978_ (.A0(\board_state[366] ),
    .A1(net30),
    .S(_3002_),
    .X(_0904_));
 sg13g2_nor2_1 _6979_ (.A(net148),
    .B(_2984_),
    .Y(_3003_));
 sg13g2_mux2_1 _6980_ (.A0(\board_state[367] ),
    .A1(net30),
    .S(_3003_),
    .X(_0905_));
 sg13g2_nand2_1 _6981_ (.Y(_3004_),
    .A(net259),
    .B(_2933_));
 sg13g2_buf_1 _6982_ (.A(_3004_),
    .X(_3005_));
 sg13g2_buf_1 _6983_ (.A(_3005_),
    .X(_3006_));
 sg13g2_nor2_1 _6984_ (.A(_2806_),
    .B(net230),
    .Y(_3007_));
 sg13g2_mux2_1 _6985_ (.A0(\board_state[368] ),
    .A1(_2996_),
    .S(_3007_),
    .X(_0906_));
 sg13g2_buf_1 _6986_ (.A(_2581_),
    .X(_3008_));
 sg13g2_nor2_1 _6987_ (.A(net194),
    .B(_3006_),
    .Y(_3009_));
 sg13g2_mux2_1 _6988_ (.A0(\board_state[369] ),
    .A1(net30),
    .S(_3009_),
    .X(_0907_));
 sg13g2_nor2_1 _6989_ (.A(net157),
    .B(net241),
    .Y(_3010_));
 sg13g2_mux2_1 _6990_ (.A0(\board_state[36] ),
    .A1(_2996_),
    .S(_3010_),
    .X(_0908_));
 sg13g2_buf_1 _6991_ (.A(net64),
    .X(_3011_));
 sg13g2_buf_1 _6992_ (.A(_2585_),
    .X(_3012_));
 sg13g2_nor2_1 _6993_ (.A(net193),
    .B(net230),
    .Y(_3013_));
 sg13g2_mux2_1 _6994_ (.A0(\board_state[370] ),
    .A1(net29),
    .S(_3013_),
    .X(_0909_));
 sg13g2_buf_1 _6995_ (.A(_2589_),
    .X(_3014_));
 sg13g2_nor2_1 _6996_ (.A(net192),
    .B(net230),
    .Y(_3015_));
 sg13g2_mux2_1 _6997_ (.A0(\board_state[371] ),
    .A1(net29),
    .S(_3015_),
    .X(_0910_));
 sg13g2_nor2_1 _6998_ (.A(net157),
    .B(net230),
    .Y(_3016_));
 sg13g2_mux2_1 _6999_ (.A0(\board_state[372] ),
    .A1(net29),
    .S(_3016_),
    .X(_0911_));
 sg13g2_nor2_1 _7000_ (.A(net156),
    .B(net230),
    .Y(_3017_));
 sg13g2_mux2_1 _7001_ (.A0(\board_state[373] ),
    .A1(net29),
    .S(_3017_),
    .X(_0912_));
 sg13g2_nor2_1 _7002_ (.A(_2819_),
    .B(net230),
    .Y(_3018_));
 sg13g2_mux2_1 _7003_ (.A0(\board_state[374] ),
    .A1(net29),
    .S(_3018_),
    .X(_0913_));
 sg13g2_nor2_1 _7004_ (.A(net154),
    .B(net230),
    .Y(_3019_));
 sg13g2_mux2_1 _7005_ (.A0(\board_state[375] ),
    .A1(net29),
    .S(_3019_),
    .X(_0914_));
 sg13g2_nor2_1 _7006_ (.A(net153),
    .B(net230),
    .Y(_3020_));
 sg13g2_mux2_1 _7007_ (.A0(\board_state[376] ),
    .A1(net29),
    .S(_3020_),
    .X(_0915_));
 sg13g2_nor2_1 _7008_ (.A(_2841_),
    .B(_3006_),
    .Y(_3021_));
 sg13g2_mux2_1 _7009_ (.A0(\board_state[377] ),
    .A1(_3011_),
    .S(_3021_),
    .X(_0916_));
 sg13g2_nor2_1 _7010_ (.A(net151),
    .B(_3005_),
    .Y(_3022_));
 sg13g2_mux2_1 _7011_ (.A0(\board_state[378] ),
    .A1(_3011_),
    .S(_3022_),
    .X(_0917_));
 sg13g2_nor2_1 _7012_ (.A(net150),
    .B(_3005_),
    .Y(_3023_));
 sg13g2_mux2_1 _7013_ (.A0(\board_state[379] ),
    .A1(net29),
    .S(_3023_),
    .X(_0918_));
 sg13g2_buf_1 _7014_ (.A(net64),
    .X(_3024_));
 sg13g2_nor2_1 _7015_ (.A(net156),
    .B(net241),
    .Y(_3025_));
 sg13g2_mux2_1 _7016_ (.A0(\board_state[37] ),
    .A1(_3024_),
    .S(_3025_),
    .X(_0919_));
 sg13g2_nor2_1 _7017_ (.A(net196),
    .B(_3005_),
    .Y(_3026_));
 sg13g2_mux2_1 _7018_ (.A0(\board_state[380] ),
    .A1(net28),
    .S(_3026_),
    .X(_0920_));
 sg13g2_nor2_1 _7019_ (.A(net149),
    .B(_3005_),
    .Y(_3027_));
 sg13g2_mux2_1 _7020_ (.A0(\board_state[381] ),
    .A1(net28),
    .S(_3027_),
    .X(_0921_));
 sg13g2_nor2_1 _7021_ (.A(net195),
    .B(_3005_),
    .Y(_3028_));
 sg13g2_mux2_1 _7022_ (.A0(\board_state[382] ),
    .A1(net28),
    .S(_3028_),
    .X(_0922_));
 sg13g2_nor2_1 _7023_ (.A(net148),
    .B(_3005_),
    .Y(_3029_));
 sg13g2_mux2_1 _7024_ (.A0(\board_state[383] ),
    .A1(_3024_),
    .S(_3029_),
    .X(_0923_));
 sg13g2_buf_1 _7025_ (.A(_2546_),
    .X(_3030_));
 sg13g2_nand2_1 _7026_ (.Y(_3031_),
    .A(net326),
    .B(_2456_));
 sg13g2_buf_1 _7027_ (.A(_3031_),
    .X(_3032_));
 sg13g2_buf_1 _7028_ (.A(_3032_),
    .X(_3033_));
 sg13g2_nor2_1 _7029_ (.A(net191),
    .B(net252),
    .Y(_3034_));
 sg13g2_mux2_1 _7030_ (.A0(\board_state[384] ),
    .A1(net28),
    .S(_3034_),
    .X(_0924_));
 sg13g2_nor2_1 _7031_ (.A(net194),
    .B(net252),
    .Y(_3035_));
 sg13g2_mux2_1 _7032_ (.A0(\board_state[385] ),
    .A1(net28),
    .S(_3035_),
    .X(_0925_));
 sg13g2_nor2_1 _7033_ (.A(net193),
    .B(net252),
    .Y(_3036_));
 sg13g2_mux2_1 _7034_ (.A0(\board_state[386] ),
    .A1(net28),
    .S(_3036_),
    .X(_0926_));
 sg13g2_nor2_1 _7035_ (.A(net192),
    .B(_3033_),
    .Y(_3037_));
 sg13g2_mux2_1 _7036_ (.A0(\board_state[387] ),
    .A1(net28),
    .S(_3037_),
    .X(_0927_));
 sg13g2_buf_1 _7037_ (.A(_2593_),
    .X(_3038_));
 sg13g2_nor2_1 _7038_ (.A(net147),
    .B(net252),
    .Y(_3039_));
 sg13g2_mux2_1 _7039_ (.A0(\board_state[388] ),
    .A1(net28),
    .S(_3039_),
    .X(_0928_));
 sg13g2_buf_1 _7040_ (.A(net64),
    .X(_3040_));
 sg13g2_buf_1 _7041_ (.A(_2597_),
    .X(_3041_));
 sg13g2_nor2_1 _7042_ (.A(net146),
    .B(net252),
    .Y(_3042_));
 sg13g2_mux2_1 _7043_ (.A0(\board_state[389] ),
    .A1(net27),
    .S(_3042_),
    .X(_0929_));
 sg13g2_nor2_1 _7044_ (.A(net155),
    .B(net241),
    .Y(_3043_));
 sg13g2_mux2_1 _7045_ (.A0(\board_state[38] ),
    .A1(_3040_),
    .S(_3043_),
    .X(_0930_));
 sg13g2_buf_1 _7046_ (.A(_2602_),
    .X(_3044_));
 sg13g2_nor2_1 _7047_ (.A(net145),
    .B(net252),
    .Y(_3045_));
 sg13g2_mux2_1 _7048_ (.A0(\board_state[390] ),
    .A1(net27),
    .S(_3045_),
    .X(_0931_));
 sg13g2_nor2_1 _7049_ (.A(_2821_),
    .B(net252),
    .Y(_3046_));
 sg13g2_mux2_1 _7050_ (.A0(\board_state[391] ),
    .A1(net27),
    .S(_3046_),
    .X(_0932_));
 sg13g2_nor2_1 _7051_ (.A(_2825_),
    .B(_3033_),
    .Y(_3047_));
 sg13g2_mux2_1 _7052_ (.A0(\board_state[392] ),
    .A1(net27),
    .S(_3047_),
    .X(_0933_));
 sg13g2_nor2_1 _7053_ (.A(_2841_),
    .B(net252),
    .Y(_3048_));
 sg13g2_mux2_1 _7054_ (.A0(\board_state[393] ),
    .A1(net27),
    .S(_3048_),
    .X(_0934_));
 sg13g2_nor2_1 _7055_ (.A(net151),
    .B(_3032_),
    .Y(_3049_));
 sg13g2_mux2_1 _7056_ (.A0(\board_state[394] ),
    .A1(net27),
    .S(_3049_),
    .X(_0935_));
 sg13g2_nor2_1 _7057_ (.A(net150),
    .B(_3032_),
    .Y(_3050_));
 sg13g2_mux2_1 _7058_ (.A0(\board_state[395] ),
    .A1(net27),
    .S(_3050_),
    .X(_0936_));
 sg13g2_nor2_1 _7059_ (.A(_2855_),
    .B(_3032_),
    .Y(_3051_));
 sg13g2_mux2_1 _7060_ (.A0(\board_state[396] ),
    .A1(net27),
    .S(_3051_),
    .X(_0937_));
 sg13g2_nor2_1 _7061_ (.A(_2857_),
    .B(_3032_),
    .Y(_3052_));
 sg13g2_mux2_1 _7062_ (.A0(\board_state[397] ),
    .A1(_3040_),
    .S(_3052_),
    .X(_0938_));
 sg13g2_buf_1 _7063_ (.A(net64),
    .X(_3053_));
 sg13g2_nor2_1 _7064_ (.A(_2860_),
    .B(_3032_),
    .Y(_3054_));
 sg13g2_mux2_1 _7065_ (.A0(\board_state[398] ),
    .A1(net26),
    .S(_3054_),
    .X(_0939_));
 sg13g2_nor2_1 _7066_ (.A(_2863_),
    .B(_3032_),
    .Y(_3055_));
 sg13g2_mux2_1 _7067_ (.A0(\board_state[399] ),
    .A1(net26),
    .S(_3055_),
    .X(_0940_));
 sg13g2_buf_1 _7068_ (.A(_2606_),
    .X(_3056_));
 sg13g2_nor2_1 _7069_ (.A(net144),
    .B(net241),
    .Y(_3057_));
 sg13g2_mux2_1 _7070_ (.A0(\board_state[39] ),
    .A1(_3053_),
    .S(_3057_),
    .X(_0941_));
 sg13g2_nor2_1 _7071_ (.A(net247),
    .B(net203),
    .Y(_3058_));
 sg13g2_mux2_1 _7072_ (.A0(\board_state[3] ),
    .A1(_3053_),
    .S(_3058_),
    .X(_0942_));
 sg13g2_nand2_1 _7073_ (.Y(_3059_),
    .A(net258),
    .B(_2456_));
 sg13g2_buf_1 _7074_ (.A(_3059_),
    .X(_3060_));
 sg13g2_buf_1 _7075_ (.A(_3060_),
    .X(_3061_));
 sg13g2_nor2_1 _7076_ (.A(net191),
    .B(net229),
    .Y(_3062_));
 sg13g2_mux2_1 _7077_ (.A0(\board_state[400] ),
    .A1(net26),
    .S(_3062_),
    .X(_0943_));
 sg13g2_nor2_1 _7078_ (.A(net194),
    .B(net229),
    .Y(_3063_));
 sg13g2_mux2_1 _7079_ (.A0(\board_state[401] ),
    .A1(net26),
    .S(_3063_),
    .X(_0944_));
 sg13g2_nor2_1 _7080_ (.A(net193),
    .B(net229),
    .Y(_3064_));
 sg13g2_mux2_1 _7081_ (.A0(\board_state[402] ),
    .A1(net26),
    .S(_3064_),
    .X(_0945_));
 sg13g2_nor2_1 _7082_ (.A(net192),
    .B(net229),
    .Y(_3065_));
 sg13g2_mux2_1 _7083_ (.A0(\board_state[403] ),
    .A1(net26),
    .S(_3065_),
    .X(_0946_));
 sg13g2_nor2_1 _7084_ (.A(net147),
    .B(net229),
    .Y(_3066_));
 sg13g2_mux2_1 _7085_ (.A0(\board_state[404] ),
    .A1(net26),
    .S(_3066_),
    .X(_0947_));
 sg13g2_nor2_1 _7086_ (.A(net146),
    .B(net229),
    .Y(_3067_));
 sg13g2_mux2_1 _7087_ (.A0(\board_state[405] ),
    .A1(net26),
    .S(_3067_),
    .X(_0948_));
 sg13g2_buf_1 _7088_ (.A(net64),
    .X(_3068_));
 sg13g2_nor2_1 _7089_ (.A(net145),
    .B(_3061_),
    .Y(_3069_));
 sg13g2_mux2_1 _7090_ (.A0(\board_state[406] ),
    .A1(net25),
    .S(_3069_),
    .X(_0949_));
 sg13g2_nor2_1 _7091_ (.A(net144),
    .B(_3061_),
    .Y(_3070_));
 sg13g2_mux2_1 _7092_ (.A0(\board_state[407] ),
    .A1(net25),
    .S(_3070_),
    .X(_0950_));
 sg13g2_buf_1 _7093_ (.A(_2614_),
    .X(_3071_));
 sg13g2_nor2_1 _7094_ (.A(net143),
    .B(net229),
    .Y(_3072_));
 sg13g2_mux2_1 _7095_ (.A0(\board_state[408] ),
    .A1(net25),
    .S(_3072_),
    .X(_0951_));
 sg13g2_buf_1 _7096_ (.A(_2618_),
    .X(_3073_));
 sg13g2_nor2_1 _7097_ (.A(net142),
    .B(net229),
    .Y(_3074_));
 sg13g2_mux2_1 _7098_ (.A0(\board_state[409] ),
    .A1(net25),
    .S(_3074_),
    .X(_0952_));
 sg13g2_nor2_1 _7099_ (.A(net143),
    .B(_2950_),
    .Y(_3075_));
 sg13g2_mux2_1 _7100_ (.A0(\board_state[40] ),
    .A1(_3068_),
    .S(_3075_),
    .X(_0953_));
 sg13g2_buf_1 _7101_ (.A(_2570_),
    .X(_3076_));
 sg13g2_nor2_1 _7102_ (.A(net141),
    .B(_3060_),
    .Y(_3077_));
 sg13g2_mux2_1 _7103_ (.A0(\board_state[410] ),
    .A1(net25),
    .S(_3077_),
    .X(_0954_));
 sg13g2_buf_1 _7104_ (.A(_2610_),
    .X(_3078_));
 sg13g2_nor2_1 _7105_ (.A(net140),
    .B(_3060_),
    .Y(_3079_));
 sg13g2_mux2_1 _7106_ (.A0(\board_state[411] ),
    .A1(net25),
    .S(_3079_),
    .X(_0955_));
 sg13g2_buf_1 _7107_ (.A(_2624_),
    .X(_3080_));
 sg13g2_nor2_1 _7108_ (.A(net190),
    .B(_3060_),
    .Y(_3081_));
 sg13g2_mux2_1 _7109_ (.A0(\board_state[412] ),
    .A1(_3068_),
    .S(_3081_),
    .X(_0956_));
 sg13g2_buf_1 _7110_ (.A(_2628_),
    .X(_3082_));
 sg13g2_nor2_1 _7111_ (.A(net139),
    .B(_3060_),
    .Y(_3083_));
 sg13g2_mux2_1 _7112_ (.A0(\board_state[413] ),
    .A1(net25),
    .S(_3083_),
    .X(_0957_));
 sg13g2_buf_1 _7113_ (.A(_2632_),
    .X(_3084_));
 sg13g2_nor2_1 _7114_ (.A(net189),
    .B(_3060_),
    .Y(_3085_));
 sg13g2_mux2_1 _7115_ (.A0(\board_state[414] ),
    .A1(net25),
    .S(_3085_),
    .X(_0958_));
 sg13g2_buf_1 _7116_ (.A(_2981_),
    .X(_3086_));
 sg13g2_buf_1 _7117_ (.A(_2637_),
    .X(_3087_));
 sg13g2_nor2_1 _7118_ (.A(net138),
    .B(_3060_),
    .Y(_3088_));
 sg13g2_mux2_1 _7119_ (.A0(\board_state[415] ),
    .A1(net24),
    .S(_3088_),
    .X(_0959_));
 sg13g2_nand2_1 _7120_ (.Y(_3089_),
    .A(_2456_),
    .B(net316));
 sg13g2_buf_1 _7121_ (.A(_3089_),
    .X(_3090_));
 sg13g2_buf_1 _7122_ (.A(_3090_),
    .X(_3091_));
 sg13g2_nor2_1 _7123_ (.A(net191),
    .B(net251),
    .Y(_3092_));
 sg13g2_mux2_1 _7124_ (.A0(\board_state[416] ),
    .A1(net24),
    .S(_3092_),
    .X(_0960_));
 sg13g2_nor2_1 _7125_ (.A(net194),
    .B(net251),
    .Y(_3093_));
 sg13g2_mux2_1 _7126_ (.A0(\board_state[417] ),
    .A1(net24),
    .S(_3093_),
    .X(_0961_));
 sg13g2_nor2_1 _7127_ (.A(net193),
    .B(net251),
    .Y(_3094_));
 sg13g2_mux2_1 _7128_ (.A0(\board_state[418] ),
    .A1(net24),
    .S(_3094_),
    .X(_0962_));
 sg13g2_nor2_1 _7129_ (.A(net192),
    .B(net251),
    .Y(_3095_));
 sg13g2_mux2_1 _7130_ (.A0(\board_state[419] ),
    .A1(net24),
    .S(_3095_),
    .X(_0963_));
 sg13g2_nor2_1 _7131_ (.A(net142),
    .B(_2950_),
    .Y(_3096_));
 sg13g2_mux2_1 _7132_ (.A0(\board_state[41] ),
    .A1(_3086_),
    .S(_3096_),
    .X(_0964_));
 sg13g2_nor2_1 _7133_ (.A(net147),
    .B(_3091_),
    .Y(_3097_));
 sg13g2_mux2_1 _7134_ (.A0(\board_state[420] ),
    .A1(_3086_),
    .S(_3097_),
    .X(_0965_));
 sg13g2_nor2_1 _7135_ (.A(_3041_),
    .B(net251),
    .Y(_3098_));
 sg13g2_mux2_1 _7136_ (.A0(\board_state[421] ),
    .A1(net24),
    .S(_3098_),
    .X(_0966_));
 sg13g2_nor2_1 _7137_ (.A(net145),
    .B(net251),
    .Y(_3099_));
 sg13g2_mux2_1 _7138_ (.A0(\board_state[422] ),
    .A1(net24),
    .S(_3099_),
    .X(_0967_));
 sg13g2_nor2_1 _7139_ (.A(net144),
    .B(net251),
    .Y(_3100_));
 sg13g2_mux2_1 _7140_ (.A0(\board_state[423] ),
    .A1(net24),
    .S(_3100_),
    .X(_0968_));
 sg13g2_buf_1 _7141_ (.A(_2981_),
    .X(_3101_));
 sg13g2_nor2_1 _7142_ (.A(_3071_),
    .B(net251),
    .Y(_3102_));
 sg13g2_mux2_1 _7143_ (.A0(\board_state[424] ),
    .A1(net23),
    .S(_3102_),
    .X(_0969_));
 sg13g2_nor2_1 _7144_ (.A(net142),
    .B(_3091_),
    .Y(_3103_));
 sg13g2_mux2_1 _7145_ (.A0(\board_state[425] ),
    .A1(_3101_),
    .S(_3103_),
    .X(_0970_));
 sg13g2_nor2_1 _7146_ (.A(_3076_),
    .B(_3090_),
    .Y(_3104_));
 sg13g2_mux2_1 _7147_ (.A0(\board_state[426] ),
    .A1(net23),
    .S(_3104_),
    .X(_0971_));
 sg13g2_nor2_1 _7148_ (.A(_3078_),
    .B(_3090_),
    .Y(_3105_));
 sg13g2_mux2_1 _7149_ (.A0(\board_state[427] ),
    .A1(net23),
    .S(_3105_),
    .X(_0972_));
 sg13g2_nor2_1 _7150_ (.A(net190),
    .B(_3090_),
    .Y(_3106_));
 sg13g2_mux2_1 _7151_ (.A0(\board_state[428] ),
    .A1(net23),
    .S(_3106_),
    .X(_0973_));
 sg13g2_nor2_1 _7152_ (.A(net139),
    .B(_3090_),
    .Y(_3107_));
 sg13g2_mux2_1 _7153_ (.A0(\board_state[429] ),
    .A1(net23),
    .S(_3107_),
    .X(_0974_));
 sg13g2_nor2_1 _7154_ (.A(net141),
    .B(_2949_),
    .Y(_3108_));
 sg13g2_mux2_1 _7155_ (.A0(\board_state[42] ),
    .A1(_3101_),
    .S(_3108_),
    .X(_0975_));
 sg13g2_nor2_1 _7156_ (.A(net189),
    .B(_3090_),
    .Y(_3109_));
 sg13g2_mux2_1 _7157_ (.A0(\board_state[430] ),
    .A1(net23),
    .S(_3109_),
    .X(_0976_));
 sg13g2_nor2_1 _7158_ (.A(net138),
    .B(_3090_),
    .Y(_3110_));
 sg13g2_mux2_1 _7159_ (.A0(\board_state[431] ),
    .A1(net23),
    .S(_3110_),
    .X(_0977_));
 sg13g2_nand2_1 _7160_ (.Y(_3111_),
    .A(net259),
    .B(_2456_));
 sg13g2_buf_1 _7161_ (.A(_3111_),
    .X(_3112_));
 sg13g2_buf_1 _7162_ (.A(_3112_),
    .X(_3113_));
 sg13g2_nor2_1 _7163_ (.A(net191),
    .B(net228),
    .Y(_3114_));
 sg13g2_mux2_1 _7164_ (.A0(\board_state[432] ),
    .A1(net23),
    .S(_3114_),
    .X(_0978_));
 sg13g2_buf_1 _7165_ (.A(net64),
    .X(_3115_));
 sg13g2_nor2_1 _7166_ (.A(net194),
    .B(net228),
    .Y(_3116_));
 sg13g2_mux2_1 _7167_ (.A0(\board_state[433] ),
    .A1(net22),
    .S(_3116_),
    .X(_0979_));
 sg13g2_nor2_1 _7168_ (.A(net193),
    .B(net228),
    .Y(_3117_));
 sg13g2_mux2_1 _7169_ (.A0(\board_state[434] ),
    .A1(net22),
    .S(_3117_),
    .X(_0980_));
 sg13g2_nor2_1 _7170_ (.A(net192),
    .B(net228),
    .Y(_3118_));
 sg13g2_mux2_1 _7171_ (.A0(\board_state[435] ),
    .A1(net22),
    .S(_3118_),
    .X(_0981_));
 sg13g2_nor2_1 _7172_ (.A(net147),
    .B(net228),
    .Y(_3119_));
 sg13g2_mux2_1 _7173_ (.A0(\board_state[436] ),
    .A1(net22),
    .S(_3119_),
    .X(_0982_));
 sg13g2_nor2_1 _7174_ (.A(net146),
    .B(_3113_),
    .Y(_3120_));
 sg13g2_mux2_1 _7175_ (.A0(\board_state[437] ),
    .A1(net22),
    .S(_3120_),
    .X(_0983_));
 sg13g2_nor2_1 _7176_ (.A(net145),
    .B(net228),
    .Y(_3121_));
 sg13g2_mux2_1 _7177_ (.A0(\board_state[438] ),
    .A1(net22),
    .S(_3121_),
    .X(_0984_));
 sg13g2_nor2_1 _7178_ (.A(net144),
    .B(net228),
    .Y(_3122_));
 sg13g2_mux2_1 _7179_ (.A0(\board_state[439] ),
    .A1(net22),
    .S(_3122_),
    .X(_0985_));
 sg13g2_nor2_1 _7180_ (.A(net140),
    .B(_2949_),
    .Y(_3123_));
 sg13g2_mux2_1 _7181_ (.A0(\board_state[43] ),
    .A1(net22),
    .S(_3123_),
    .X(_0986_));
 sg13g2_nor2_1 _7182_ (.A(net143),
    .B(net228),
    .Y(_3124_));
 sg13g2_mux2_1 _7183_ (.A0(\board_state[440] ),
    .A1(_3115_),
    .S(_3124_),
    .X(_0987_));
 sg13g2_nor2_1 _7184_ (.A(net142),
    .B(_3113_),
    .Y(_3125_));
 sg13g2_mux2_1 _7185_ (.A0(\board_state[441] ),
    .A1(_3115_),
    .S(_3125_),
    .X(_0988_));
 sg13g2_buf_1 _7186_ (.A(_2533_),
    .X(_3126_));
 sg13g2_buf_1 _7187_ (.A(net63),
    .X(_3127_));
 sg13g2_nor2_1 _7188_ (.A(_3076_),
    .B(_3112_),
    .Y(_3128_));
 sg13g2_mux2_1 _7189_ (.A0(\board_state[442] ),
    .A1(net21),
    .S(_3128_),
    .X(_0989_));
 sg13g2_nor2_1 _7190_ (.A(net140),
    .B(_3112_),
    .Y(_3129_));
 sg13g2_mux2_1 _7191_ (.A0(\board_state[443] ),
    .A1(net21),
    .S(_3129_),
    .X(_0990_));
 sg13g2_nor2_1 _7192_ (.A(net190),
    .B(_3112_),
    .Y(_3130_));
 sg13g2_mux2_1 _7193_ (.A0(\board_state[444] ),
    .A1(net21),
    .S(_3130_),
    .X(_0991_));
 sg13g2_nor2_1 _7194_ (.A(net139),
    .B(_3112_),
    .Y(_3131_));
 sg13g2_mux2_1 _7195_ (.A0(\board_state[445] ),
    .A1(net21),
    .S(_3131_),
    .X(_0992_));
 sg13g2_nor2_1 _7196_ (.A(net189),
    .B(_3112_),
    .Y(_3132_));
 sg13g2_mux2_1 _7197_ (.A0(\board_state[446] ),
    .A1(net21),
    .S(_3132_),
    .X(_0993_));
 sg13g2_nor2_1 _7198_ (.A(net138),
    .B(_3112_),
    .Y(_3133_));
 sg13g2_mux2_1 _7199_ (.A0(\board_state[447] ),
    .A1(_3127_),
    .S(_3133_),
    .X(_0994_));
 sg13g2_nor2_2 _7200_ (.A(_2551_),
    .B(_2455_),
    .Y(_3134_));
 sg13g2_nand2_1 _7201_ (.Y(_3135_),
    .A(net326),
    .B(_3134_));
 sg13g2_buf_1 _7202_ (.A(_3135_),
    .X(_3136_));
 sg13g2_buf_1 _7203_ (.A(_3136_),
    .X(_3137_));
 sg13g2_nor2_1 _7204_ (.A(net191),
    .B(net250),
    .Y(_3138_));
 sg13g2_mux2_1 _7205_ (.A0(\board_state[448] ),
    .A1(net21),
    .S(_3138_),
    .X(_0995_));
 sg13g2_nor2_1 _7206_ (.A(_3008_),
    .B(net250),
    .Y(_3139_));
 sg13g2_mux2_1 _7207_ (.A0(\board_state[449] ),
    .A1(net21),
    .S(_3139_),
    .X(_0996_));
 sg13g2_nor2_1 _7208_ (.A(net190),
    .B(_2949_),
    .Y(_3140_));
 sg13g2_mux2_1 _7209_ (.A0(\board_state[44] ),
    .A1(_3127_),
    .S(_3140_),
    .X(_0997_));
 sg13g2_nor2_1 _7210_ (.A(_3012_),
    .B(net250),
    .Y(_3141_));
 sg13g2_mux2_1 _7211_ (.A0(\board_state[450] ),
    .A1(net21),
    .S(_3141_),
    .X(_0998_));
 sg13g2_buf_1 _7212_ (.A(_3126_),
    .X(_3142_));
 sg13g2_nor2_1 _7213_ (.A(_3014_),
    .B(net250),
    .Y(_3143_));
 sg13g2_mux2_1 _7214_ (.A0(\board_state[451] ),
    .A1(net20),
    .S(_3143_),
    .X(_0999_));
 sg13g2_nor2_1 _7215_ (.A(net147),
    .B(net250),
    .Y(_3144_));
 sg13g2_mux2_1 _7216_ (.A0(\board_state[452] ),
    .A1(net20),
    .S(_3144_),
    .X(_1000_));
 sg13g2_nor2_1 _7217_ (.A(net146),
    .B(net250),
    .Y(_3145_));
 sg13g2_mux2_1 _7218_ (.A0(\board_state[453] ),
    .A1(net20),
    .S(_3145_),
    .X(_1001_));
 sg13g2_nor2_1 _7219_ (.A(net145),
    .B(_3137_),
    .Y(_3146_));
 sg13g2_mux2_1 _7220_ (.A0(\board_state[454] ),
    .A1(net20),
    .S(_3146_),
    .X(_1002_));
 sg13g2_nor2_1 _7221_ (.A(net144),
    .B(_3137_),
    .Y(_3147_));
 sg13g2_mux2_1 _7222_ (.A0(\board_state[455] ),
    .A1(net20),
    .S(_3147_),
    .X(_1003_));
 sg13g2_nor2_1 _7223_ (.A(net143),
    .B(net250),
    .Y(_3148_));
 sg13g2_mux2_1 _7224_ (.A0(\board_state[456] ),
    .A1(net20),
    .S(_3148_),
    .X(_1004_));
 sg13g2_nor2_1 _7225_ (.A(net142),
    .B(net250),
    .Y(_3149_));
 sg13g2_mux2_1 _7226_ (.A0(\board_state[457] ),
    .A1(net20),
    .S(_3149_),
    .X(_1005_));
 sg13g2_nor2_1 _7227_ (.A(net141),
    .B(_3136_),
    .Y(_3150_));
 sg13g2_mux2_1 _7228_ (.A0(\board_state[458] ),
    .A1(net20),
    .S(_3150_),
    .X(_1006_));
 sg13g2_nor2_1 _7229_ (.A(net140),
    .B(_3136_),
    .Y(_3151_));
 sg13g2_mux2_1 _7230_ (.A0(\board_state[459] ),
    .A1(_3142_),
    .S(_3151_),
    .X(_1007_));
 sg13g2_nor2_1 _7231_ (.A(net139),
    .B(_2949_),
    .Y(_3152_));
 sg13g2_mux2_1 _7232_ (.A0(\board_state[45] ),
    .A1(_3142_),
    .S(_3152_),
    .X(_1008_));
 sg13g2_buf_1 _7233_ (.A(net63),
    .X(_3153_));
 sg13g2_nor2_1 _7234_ (.A(net190),
    .B(_3136_),
    .Y(_3154_));
 sg13g2_mux2_1 _7235_ (.A0(\board_state[460] ),
    .A1(net19),
    .S(_3154_),
    .X(_1009_));
 sg13g2_nor2_1 _7236_ (.A(net139),
    .B(_3136_),
    .Y(_3155_));
 sg13g2_mux2_1 _7237_ (.A0(\board_state[461] ),
    .A1(net19),
    .S(_3155_),
    .X(_1010_));
 sg13g2_nor2_1 _7238_ (.A(net189),
    .B(_3136_),
    .Y(_3156_));
 sg13g2_mux2_1 _7239_ (.A0(\board_state[462] ),
    .A1(_3153_),
    .S(_3156_),
    .X(_1011_));
 sg13g2_nor2_1 _7240_ (.A(net138),
    .B(_3136_),
    .Y(_3157_));
 sg13g2_mux2_1 _7241_ (.A0(\board_state[463] ),
    .A1(_3153_),
    .S(_3157_),
    .X(_1012_));
 sg13g2_nand2_1 _7242_ (.Y(_3158_),
    .A(net258),
    .B(_3134_));
 sg13g2_buf_1 _7243_ (.A(_3158_),
    .X(_3159_));
 sg13g2_buf_1 _7244_ (.A(_3159_),
    .X(_3160_));
 sg13g2_nor2_1 _7245_ (.A(net191),
    .B(net227),
    .Y(_3161_));
 sg13g2_mux2_1 _7246_ (.A0(\board_state[464] ),
    .A1(net19),
    .S(_3161_),
    .X(_1013_));
 sg13g2_nor2_1 _7247_ (.A(_3008_),
    .B(net227),
    .Y(_3162_));
 sg13g2_mux2_1 _7248_ (.A0(\board_state[465] ),
    .A1(net19),
    .S(_3162_),
    .X(_1014_));
 sg13g2_nor2_1 _7249_ (.A(_3012_),
    .B(net227),
    .Y(_3163_));
 sg13g2_mux2_1 _7250_ (.A0(\board_state[466] ),
    .A1(net19),
    .S(_3163_),
    .X(_1015_));
 sg13g2_nor2_1 _7251_ (.A(_3014_),
    .B(net227),
    .Y(_3164_));
 sg13g2_mux2_1 _7252_ (.A0(\board_state[467] ),
    .A1(net19),
    .S(_3164_),
    .X(_1016_));
 sg13g2_nor2_1 _7253_ (.A(net147),
    .B(net227),
    .Y(_3165_));
 sg13g2_mux2_1 _7254_ (.A0(\board_state[468] ),
    .A1(net19),
    .S(_3165_),
    .X(_1017_));
 sg13g2_nor2_1 _7255_ (.A(net146),
    .B(net227),
    .Y(_3166_));
 sg13g2_mux2_1 _7256_ (.A0(\board_state[469] ),
    .A1(net19),
    .S(_3166_),
    .X(_1018_));
 sg13g2_buf_1 _7257_ (.A(_3126_),
    .X(_3167_));
 sg13g2_nor2_1 _7258_ (.A(net189),
    .B(_2949_),
    .Y(_3168_));
 sg13g2_mux2_1 _7259_ (.A0(\board_state[46] ),
    .A1(_3167_),
    .S(_3168_),
    .X(_1019_));
 sg13g2_nor2_1 _7260_ (.A(net145),
    .B(net227),
    .Y(_3169_));
 sg13g2_mux2_1 _7261_ (.A0(\board_state[470] ),
    .A1(net18),
    .S(_3169_),
    .X(_1020_));
 sg13g2_nor2_1 _7262_ (.A(net144),
    .B(net227),
    .Y(_3170_));
 sg13g2_mux2_1 _7263_ (.A0(\board_state[471] ),
    .A1(net18),
    .S(_3170_),
    .X(_1021_));
 sg13g2_nor2_1 _7264_ (.A(net143),
    .B(_3160_),
    .Y(_3171_));
 sg13g2_mux2_1 _7265_ (.A0(\board_state[472] ),
    .A1(net18),
    .S(_3171_),
    .X(_1022_));
 sg13g2_nor2_1 _7266_ (.A(net142),
    .B(_3160_),
    .Y(_3172_));
 sg13g2_mux2_1 _7267_ (.A0(\board_state[473] ),
    .A1(net18),
    .S(_3172_),
    .X(_1023_));
 sg13g2_nor2_1 _7268_ (.A(net141),
    .B(_3159_),
    .Y(_3173_));
 sg13g2_mux2_1 _7269_ (.A0(\board_state[474] ),
    .A1(net18),
    .S(_3173_),
    .X(_1024_));
 sg13g2_nor2_1 _7270_ (.A(net140),
    .B(_3159_),
    .Y(_3174_));
 sg13g2_mux2_1 _7271_ (.A0(\board_state[475] ),
    .A1(net18),
    .S(_3174_),
    .X(_1025_));
 sg13g2_nor2_1 _7272_ (.A(net190),
    .B(_3159_),
    .Y(_3175_));
 sg13g2_mux2_1 _7273_ (.A0(\board_state[476] ),
    .A1(net18),
    .S(_3175_),
    .X(_1026_));
 sg13g2_nor2_1 _7274_ (.A(net139),
    .B(_3159_),
    .Y(_3176_));
 sg13g2_mux2_1 _7275_ (.A0(\board_state[477] ),
    .A1(net18),
    .S(_3176_),
    .X(_1027_));
 sg13g2_nor2_1 _7276_ (.A(net189),
    .B(_3159_),
    .Y(_3177_));
 sg13g2_mux2_1 _7277_ (.A0(\board_state[478] ),
    .A1(_3167_),
    .S(_3177_),
    .X(_1028_));
 sg13g2_buf_1 _7278_ (.A(net63),
    .X(_3178_));
 sg13g2_nor2_1 _7279_ (.A(net138),
    .B(_3159_),
    .Y(_3179_));
 sg13g2_mux2_1 _7280_ (.A0(\board_state[479] ),
    .A1(net17),
    .S(_3179_),
    .X(_1029_));
 sg13g2_nor2_1 _7281_ (.A(_3087_),
    .B(_2949_),
    .Y(_3180_));
 sg13g2_mux2_1 _7282_ (.A0(\board_state[47] ),
    .A1(_3178_),
    .S(_3180_),
    .X(_1030_));
 sg13g2_nand2_1 _7283_ (.Y(_3181_),
    .A(net316),
    .B(_3134_));
 sg13g2_buf_1 _7284_ (.A(_3181_),
    .X(_3182_));
 sg13g2_buf_1 _7285_ (.A(_3182_),
    .X(_3183_));
 sg13g2_nor2_1 _7286_ (.A(net191),
    .B(net249),
    .Y(_3184_));
 sg13g2_mux2_1 _7287_ (.A0(\board_state[480] ),
    .A1(net17),
    .S(_3184_),
    .X(_1031_));
 sg13g2_nor2_1 _7288_ (.A(net194),
    .B(net249),
    .Y(_3185_));
 sg13g2_mux2_1 _7289_ (.A0(\board_state[481] ),
    .A1(net17),
    .S(_3185_),
    .X(_1032_));
 sg13g2_nor2_1 _7290_ (.A(net193),
    .B(_3183_),
    .Y(_3186_));
 sg13g2_mux2_1 _7291_ (.A0(\board_state[482] ),
    .A1(net17),
    .S(_3186_),
    .X(_1033_));
 sg13g2_nor2_1 _7292_ (.A(net192),
    .B(_3183_),
    .Y(_3187_));
 sg13g2_mux2_1 _7293_ (.A0(\board_state[483] ),
    .A1(_3178_),
    .S(_3187_),
    .X(_1034_));
 sg13g2_nor2_1 _7294_ (.A(net147),
    .B(net249),
    .Y(_3188_));
 sg13g2_mux2_1 _7295_ (.A0(\board_state[484] ),
    .A1(net17),
    .S(_3188_),
    .X(_1035_));
 sg13g2_nor2_1 _7296_ (.A(net146),
    .B(net249),
    .Y(_3189_));
 sg13g2_mux2_1 _7297_ (.A0(\board_state[485] ),
    .A1(net17),
    .S(_3189_),
    .X(_1036_));
 sg13g2_nor2_1 _7298_ (.A(net145),
    .B(net249),
    .Y(_3190_));
 sg13g2_mux2_1 _7299_ (.A0(\board_state[486] ),
    .A1(net17),
    .S(_3190_),
    .X(_1037_));
 sg13g2_nor2_1 _7300_ (.A(net144),
    .B(net249),
    .Y(_3191_));
 sg13g2_mux2_1 _7301_ (.A0(\board_state[487] ),
    .A1(net17),
    .S(_3191_),
    .X(_1038_));
 sg13g2_buf_1 _7302_ (.A(net63),
    .X(_3192_));
 sg13g2_nor2_1 _7303_ (.A(net143),
    .B(net249),
    .Y(_3193_));
 sg13g2_mux2_1 _7304_ (.A0(\board_state[488] ),
    .A1(net16),
    .S(_3193_),
    .X(_1039_));
 sg13g2_nor2_1 _7305_ (.A(net142),
    .B(net249),
    .Y(_3194_));
 sg13g2_mux2_1 _7306_ (.A0(\board_state[489] ),
    .A1(net16),
    .S(_3194_),
    .X(_1040_));
 sg13g2_nand2_1 _7307_ (.Y(_3195_),
    .A(_2537_),
    .B(net259));
 sg13g2_buf_1 _7308_ (.A(_3195_),
    .X(_3196_));
 sg13g2_buf_1 _7309_ (.A(_3196_),
    .X(_3197_));
 sg13g2_nor2_1 _7310_ (.A(_3030_),
    .B(net226),
    .Y(_3198_));
 sg13g2_mux2_1 _7311_ (.A0(\board_state[48] ),
    .A1(_3192_),
    .S(_3198_),
    .X(_1041_));
 sg13g2_nor2_1 _7312_ (.A(net141),
    .B(_3182_),
    .Y(_3199_));
 sg13g2_mux2_1 _7313_ (.A0(\board_state[490] ),
    .A1(net16),
    .S(_3199_),
    .X(_1042_));
 sg13g2_nor2_1 _7314_ (.A(net140),
    .B(_3182_),
    .Y(_3200_));
 sg13g2_mux2_1 _7315_ (.A0(\board_state[491] ),
    .A1(net16),
    .S(_3200_),
    .X(_1043_));
 sg13g2_nor2_1 _7316_ (.A(_3080_),
    .B(_3182_),
    .Y(_3201_));
 sg13g2_mux2_1 _7317_ (.A0(\board_state[492] ),
    .A1(net16),
    .S(_3201_),
    .X(_1044_));
 sg13g2_nor2_1 _7318_ (.A(_3082_),
    .B(_3182_),
    .Y(_3202_));
 sg13g2_mux2_1 _7319_ (.A0(\board_state[493] ),
    .A1(net16),
    .S(_3202_),
    .X(_1045_));
 sg13g2_nor2_1 _7320_ (.A(net189),
    .B(_3182_),
    .Y(_3203_));
 sg13g2_mux2_1 _7321_ (.A0(\board_state[494] ),
    .A1(net16),
    .S(_3203_),
    .X(_1046_));
 sg13g2_nor2_1 _7322_ (.A(_3087_),
    .B(_3182_),
    .Y(_3204_));
 sg13g2_mux2_1 _7323_ (.A0(\board_state[495] ),
    .A1(net16),
    .S(_3204_),
    .X(_1047_));
 sg13g2_nand2_1 _7324_ (.Y(_3205_),
    .A(net259),
    .B(_3134_));
 sg13g2_buf_1 _7325_ (.A(_3205_),
    .X(_3206_));
 sg13g2_buf_1 _7326_ (.A(_3206_),
    .X(_3207_));
 sg13g2_nor2_1 _7327_ (.A(net191),
    .B(net225),
    .Y(_3208_));
 sg13g2_mux2_1 _7328_ (.A0(\board_state[496] ),
    .A1(_3192_),
    .S(_3208_),
    .X(_1048_));
 sg13g2_buf_1 _7329_ (.A(net63),
    .X(_3209_));
 sg13g2_nor2_1 _7330_ (.A(net194),
    .B(net225),
    .Y(_3210_));
 sg13g2_mux2_1 _7331_ (.A0(\board_state[497] ),
    .A1(net15),
    .S(_3210_),
    .X(_1049_));
 sg13g2_nor2_1 _7332_ (.A(net193),
    .B(_3207_),
    .Y(_3211_));
 sg13g2_mux2_1 _7333_ (.A0(\board_state[498] ),
    .A1(net15),
    .S(_3211_),
    .X(_1050_));
 sg13g2_nor2_1 _7334_ (.A(net192),
    .B(net225),
    .Y(_3212_));
 sg13g2_mux2_1 _7335_ (.A0(\board_state[499] ),
    .A1(net15),
    .S(_3212_),
    .X(_1051_));
 sg13g2_nor2_1 _7336_ (.A(net194),
    .B(net226),
    .Y(_3213_));
 sg13g2_mux2_1 _7337_ (.A0(\board_state[49] ),
    .A1(net15),
    .S(_3213_),
    .X(_1052_));
 sg13g2_nor2_1 _7338_ (.A(_2539_),
    .B(_2594_),
    .Y(_3214_));
 sg13g2_mux2_1 _7339_ (.A0(\board_state[4] ),
    .A1(net15),
    .S(_3214_),
    .X(_1053_));
 sg13g2_nor2_1 _7340_ (.A(_3038_),
    .B(net225),
    .Y(_3215_));
 sg13g2_mux2_1 _7341_ (.A0(\board_state[500] ),
    .A1(net15),
    .S(_3215_),
    .X(_1054_));
 sg13g2_nor2_1 _7342_ (.A(_3041_),
    .B(net225),
    .Y(_3216_));
 sg13g2_mux2_1 _7343_ (.A0(\board_state[501] ),
    .A1(net15),
    .S(_3216_),
    .X(_1055_));
 sg13g2_nor2_1 _7344_ (.A(net145),
    .B(net225),
    .Y(_3217_));
 sg13g2_mux2_1 _7345_ (.A0(\board_state[502] ),
    .A1(net15),
    .S(_3217_),
    .X(_1056_));
 sg13g2_nor2_1 _7346_ (.A(_3056_),
    .B(_3207_),
    .Y(_3218_));
 sg13g2_mux2_1 _7347_ (.A0(\board_state[503] ),
    .A1(_3209_),
    .S(_3218_),
    .X(_1057_));
 sg13g2_nor2_1 _7348_ (.A(net143),
    .B(net225),
    .Y(_3219_));
 sg13g2_mux2_1 _7349_ (.A0(\board_state[504] ),
    .A1(_3209_),
    .S(_3219_),
    .X(_1058_));
 sg13g2_buf_1 _7350_ (.A(net63),
    .X(_3220_));
 sg13g2_nor2_1 _7351_ (.A(net142),
    .B(net225),
    .Y(_3221_));
 sg13g2_mux2_1 _7352_ (.A0(\board_state[505] ),
    .A1(net14),
    .S(_3221_),
    .X(_1059_));
 sg13g2_nor2_1 _7353_ (.A(net141),
    .B(_3206_),
    .Y(_3222_));
 sg13g2_mux2_1 _7354_ (.A0(\board_state[506] ),
    .A1(net14),
    .S(_3222_),
    .X(_1060_));
 sg13g2_nor2_1 _7355_ (.A(net140),
    .B(_3206_),
    .Y(_3223_));
 sg13g2_mux2_1 _7356_ (.A0(\board_state[507] ),
    .A1(net14),
    .S(_3223_),
    .X(_1061_));
 sg13g2_nor2_1 _7357_ (.A(net190),
    .B(_3206_),
    .Y(_3224_));
 sg13g2_mux2_1 _7358_ (.A0(\board_state[508] ),
    .A1(net14),
    .S(_3224_),
    .X(_1062_));
 sg13g2_nor2_1 _7359_ (.A(net139),
    .B(_3206_),
    .Y(_3225_));
 sg13g2_mux2_1 _7360_ (.A0(\board_state[509] ),
    .A1(net14),
    .S(_3225_),
    .X(_1063_));
 sg13g2_nor2_1 _7361_ (.A(net193),
    .B(net226),
    .Y(_3226_));
 sg13g2_mux2_1 _7362_ (.A0(\board_state[50] ),
    .A1(net14),
    .S(_3226_),
    .X(_1064_));
 sg13g2_nor2_1 _7363_ (.A(net189),
    .B(_3206_),
    .Y(_3227_));
 sg13g2_mux2_1 _7364_ (.A0(\board_state[510] ),
    .A1(_3220_),
    .S(_3227_),
    .X(_1065_));
 sg13g2_nor2_1 _7365_ (.A(net138),
    .B(_3206_),
    .Y(_3228_));
 sg13g2_mux2_1 _7366_ (.A0(\board_state[511] ),
    .A1(_3220_),
    .S(_3228_),
    .X(_1066_));
 sg13g2_nor2_1 _7367_ (.A(net192),
    .B(net226),
    .Y(_3229_));
 sg13g2_mux2_1 _7368_ (.A0(\board_state[51] ),
    .A1(net14),
    .S(_3229_),
    .X(_1067_));
 sg13g2_nor2_1 _7369_ (.A(_3038_),
    .B(net226),
    .Y(_3230_));
 sg13g2_mux2_1 _7370_ (.A0(\board_state[52] ),
    .A1(net14),
    .S(_3230_),
    .X(_1068_));
 sg13g2_buf_1 _7371_ (.A(net63),
    .X(_3231_));
 sg13g2_nor2_1 _7372_ (.A(net146),
    .B(net226),
    .Y(_3232_));
 sg13g2_mux2_1 _7373_ (.A0(\board_state[53] ),
    .A1(net13),
    .S(_3232_),
    .X(_1069_));
 sg13g2_nor2_1 _7374_ (.A(_3044_),
    .B(net226),
    .Y(_3233_));
 sg13g2_mux2_1 _7375_ (.A0(\board_state[54] ),
    .A1(net13),
    .S(_3233_),
    .X(_1070_));
 sg13g2_nor2_1 _7376_ (.A(_3056_),
    .B(_3197_),
    .Y(_3234_));
 sg13g2_mux2_1 _7377_ (.A0(\board_state[55] ),
    .A1(net13),
    .S(_3234_),
    .X(_1071_));
 sg13g2_nor2_1 _7378_ (.A(_3071_),
    .B(net226),
    .Y(_3235_));
 sg13g2_mux2_1 _7379_ (.A0(\board_state[56] ),
    .A1(_3231_),
    .S(_3235_),
    .X(_1072_));
 sg13g2_nor2_1 _7380_ (.A(_3073_),
    .B(_3197_),
    .Y(_3236_));
 sg13g2_mux2_1 _7381_ (.A0(\board_state[57] ),
    .A1(net13),
    .S(_3236_),
    .X(_1073_));
 sg13g2_nor2_1 _7382_ (.A(net141),
    .B(_3196_),
    .Y(_3237_));
 sg13g2_mux2_1 _7383_ (.A0(\board_state[58] ),
    .A1(net13),
    .S(_3237_),
    .X(_1074_));
 sg13g2_nor2_1 _7384_ (.A(_3078_),
    .B(_3196_),
    .Y(_3238_));
 sg13g2_mux2_1 _7385_ (.A0(\board_state[59] ),
    .A1(net13),
    .S(_3238_),
    .X(_1075_));
 sg13g2_nor2_1 _7386_ (.A(_2539_),
    .B(_2598_),
    .Y(_3239_));
 sg13g2_mux2_1 _7387_ (.A0(\board_state[5] ),
    .A1(net13),
    .S(_3239_),
    .X(_1076_));
 sg13g2_nor2_1 _7388_ (.A(_3080_),
    .B(_3196_),
    .Y(_3240_));
 sg13g2_mux2_1 _7389_ (.A0(\board_state[60] ),
    .A1(net13),
    .S(_3240_),
    .X(_1077_));
 sg13g2_nor2_1 _7390_ (.A(_3082_),
    .B(_3196_),
    .Y(_3241_));
 sg13g2_mux2_1 _7391_ (.A0(\board_state[61] ),
    .A1(_3231_),
    .S(_3241_),
    .X(_1078_));
 sg13g2_buf_1 _7392_ (.A(net63),
    .X(_3242_));
 sg13g2_nor2_1 _7393_ (.A(_3084_),
    .B(_3196_),
    .Y(_3243_));
 sg13g2_mux2_1 _7394_ (.A0(\board_state[62] ),
    .A1(net12),
    .S(_3243_),
    .X(_1079_));
 sg13g2_nor2_1 _7395_ (.A(net138),
    .B(_3196_),
    .Y(_3244_));
 sg13g2_mux2_1 _7396_ (.A0(\board_state[63] ),
    .A1(_3242_),
    .S(_3244_),
    .X(_1080_));
 sg13g2_nand2_1 _7397_ (.Y(_3245_),
    .A(_2031_),
    .B(_2552_));
 sg13g2_buf_2 _7398_ (.A(_3245_),
    .X(_3246_));
 sg13g2_buf_1 _7399_ (.A(_3246_),
    .X(_3247_));
 sg13g2_nor2_1 _7400_ (.A(_3030_),
    .B(net248),
    .Y(_3248_));
 sg13g2_mux2_1 _7401_ (.A0(\board_state[64] ),
    .A1(net12),
    .S(_3248_),
    .X(_1081_));
 sg13g2_nor2_1 _7402_ (.A(_2581_),
    .B(net248),
    .Y(_3249_));
 sg13g2_mux2_1 _7403_ (.A0(\board_state[65] ),
    .A1(net12),
    .S(_3249_),
    .X(_1082_));
 sg13g2_nor2_1 _7404_ (.A(_2585_),
    .B(net248),
    .Y(_3250_));
 sg13g2_mux2_1 _7405_ (.A0(\board_state[66] ),
    .A1(net12),
    .S(_3250_),
    .X(_1083_));
 sg13g2_nor2_1 _7406_ (.A(_2589_),
    .B(net248),
    .Y(_3251_));
 sg13g2_mux2_1 _7407_ (.A0(\board_state[67] ),
    .A1(_3242_),
    .S(_3251_),
    .X(_1084_));
 sg13g2_nor2_1 _7408_ (.A(net147),
    .B(net248),
    .Y(_3252_));
 sg13g2_mux2_1 _7409_ (.A0(\board_state[68] ),
    .A1(net12),
    .S(_3252_),
    .X(_1085_));
 sg13g2_nor2_1 _7410_ (.A(net146),
    .B(net248),
    .Y(_3253_));
 sg13g2_mux2_1 _7411_ (.A0(\board_state[69] ),
    .A1(net12),
    .S(_3253_),
    .X(_1086_));
 sg13g2_nor2_1 _7412_ (.A(_2539_),
    .B(_2603_),
    .Y(_3254_));
 sg13g2_mux2_1 _7413_ (.A0(\board_state[6] ),
    .A1(net12),
    .S(_3254_),
    .X(_1087_));
 sg13g2_nor2_1 _7414_ (.A(_3044_),
    .B(net248),
    .Y(_3255_));
 sg13g2_mux2_1 _7415_ (.A0(\board_state[70] ),
    .A1(net12),
    .S(_3255_),
    .X(_1088_));
 sg13g2_buf_1 _7416_ (.A(_2533_),
    .X(_3256_));
 sg13g2_nor2_1 _7417_ (.A(net144),
    .B(_3247_),
    .Y(_3257_));
 sg13g2_mux2_1 _7418_ (.A0(\board_state[71] ),
    .A1(net62),
    .S(_3257_),
    .X(_1089_));
 sg13g2_nor2_1 _7419_ (.A(net143),
    .B(_3247_),
    .Y(_3258_));
 sg13g2_mux2_1 _7420_ (.A0(\board_state[72] ),
    .A1(_3256_),
    .S(_3258_),
    .X(_1090_));
 sg13g2_nor2_1 _7421_ (.A(_3073_),
    .B(net248),
    .Y(_3259_));
 sg13g2_mux2_1 _7422_ (.A0(\board_state[73] ),
    .A1(net62),
    .S(_3259_),
    .X(_1091_));
 sg13g2_nor2_1 _7423_ (.A(net141),
    .B(_3246_),
    .Y(_3260_));
 sg13g2_mux2_1 _7424_ (.A0(\board_state[74] ),
    .A1(net62),
    .S(_3260_),
    .X(_1092_));
 sg13g2_nor2_1 _7425_ (.A(net140),
    .B(_3246_),
    .Y(_3261_));
 sg13g2_mux2_1 _7426_ (.A0(\board_state[75] ),
    .A1(net62),
    .S(_3261_),
    .X(_1093_));
 sg13g2_nor2_1 _7427_ (.A(net190),
    .B(_3246_),
    .Y(_3262_));
 sg13g2_mux2_1 _7428_ (.A0(\board_state[76] ),
    .A1(net62),
    .S(_3262_),
    .X(_1094_));
 sg13g2_nor2_1 _7429_ (.A(net139),
    .B(_3246_),
    .Y(_3263_));
 sg13g2_mux2_1 _7430_ (.A0(\board_state[77] ),
    .A1(net62),
    .S(_3263_),
    .X(_1095_));
 sg13g2_nor2_1 _7431_ (.A(_3084_),
    .B(_3246_),
    .Y(_3264_));
 sg13g2_mux2_1 _7432_ (.A0(\board_state[78] ),
    .A1(net62),
    .S(_3264_),
    .X(_1096_));
 sg13g2_nor2_1 _7433_ (.A(net138),
    .B(_3246_),
    .Y(_3265_));
 sg13g2_mux2_1 _7434_ (.A0(\board_state[79] ),
    .A1(net62),
    .S(_3265_),
    .X(_1097_));
 sg13g2_nor2_1 _7435_ (.A(_2539_),
    .B(_2607_),
    .Y(_3266_));
 sg13g2_mux2_1 _7436_ (.A0(\board_state[7] ),
    .A1(_3256_),
    .S(_3266_),
    .X(_1098_));
 sg13g2_buf_1 _7437_ (.A(_2533_),
    .X(_3267_));
 sg13g2_nand2_1 _7438_ (.Y(_3268_),
    .A(net258),
    .B(_2552_));
 sg13g2_buf_1 _7439_ (.A(_3268_),
    .X(_3269_));
 sg13g2_buf_1 _7440_ (.A(_3269_),
    .X(_3270_));
 sg13g2_nor2_1 _7441_ (.A(_2546_),
    .B(net224),
    .Y(_3271_));
 sg13g2_mux2_1 _7442_ (.A0(\board_state[80] ),
    .A1(net61),
    .S(_3271_),
    .X(_1099_));
 sg13g2_nor2_1 _7443_ (.A(_2581_),
    .B(net224),
    .Y(_3272_));
 sg13g2_mux2_1 _7444_ (.A0(\board_state[81] ),
    .A1(net61),
    .S(_3272_),
    .X(_1100_));
 sg13g2_nor2_1 _7445_ (.A(_2585_),
    .B(net224),
    .Y(_3273_));
 sg13g2_mux2_1 _7446_ (.A0(\board_state[82] ),
    .A1(net61),
    .S(_3273_),
    .X(_1101_));
 sg13g2_nor2_1 _7447_ (.A(_2589_),
    .B(_3270_),
    .Y(_3274_));
 sg13g2_mux2_1 _7448_ (.A0(\board_state[83] ),
    .A1(_3267_),
    .S(_3274_),
    .X(_1102_));
 sg13g2_nor2_1 _7449_ (.A(_2593_),
    .B(net224),
    .Y(_3275_));
 sg13g2_mux2_1 _7450_ (.A0(\board_state[84] ),
    .A1(net61),
    .S(_3275_),
    .X(_1103_));
 sg13g2_nor2_1 _7451_ (.A(_2597_),
    .B(net224),
    .Y(_3276_));
 sg13g2_mux2_1 _7452_ (.A0(\board_state[85] ),
    .A1(net61),
    .S(_3276_),
    .X(_1104_));
 sg13g2_nor2_1 _7453_ (.A(_2602_),
    .B(net224),
    .Y(_3277_));
 sg13g2_mux2_1 _7454_ (.A0(\board_state[86] ),
    .A1(net61),
    .S(_3277_),
    .X(_1105_));
 sg13g2_nor2_1 _7455_ (.A(_2606_),
    .B(net224),
    .Y(_3278_));
 sg13g2_mux2_1 _7456_ (.A0(\board_state[87] ),
    .A1(net61),
    .S(_3278_),
    .X(_1106_));
 sg13g2_nor2_1 _7457_ (.A(_2614_),
    .B(net224),
    .Y(_3279_));
 sg13g2_mux2_1 _7458_ (.A0(\board_state[88] ),
    .A1(_3267_),
    .S(_3279_),
    .X(_1107_));
 sg13g2_nor2_1 _7459_ (.A(_2618_),
    .B(_3270_),
    .Y(_3280_));
 sg13g2_mux2_1 _7460_ (.A0(\board_state[89] ),
    .A1(net61),
    .S(_3280_),
    .X(_1108_));
 sg13g2_buf_1 _7461_ (.A(_2533_),
    .X(_3281_));
 sg13g2_nor2_1 _7462_ (.A(_2539_),
    .B(net161),
    .Y(_3282_));
 sg13g2_mux2_1 _7463_ (.A0(\board_state[8] ),
    .A1(net60),
    .S(_3282_),
    .X(_1109_));
 sg13g2_nor2_1 _7464_ (.A(_2570_),
    .B(_3269_),
    .Y(_3283_));
 sg13g2_mux2_1 _7465_ (.A0(\board_state[90] ),
    .A1(net60),
    .S(_3283_),
    .X(_1110_));
 sg13g2_nor2_1 _7466_ (.A(_2610_),
    .B(_3269_),
    .Y(_3284_));
 sg13g2_mux2_1 _7467_ (.A0(\board_state[91] ),
    .A1(net60),
    .S(_3284_),
    .X(_1111_));
 sg13g2_nor2_1 _7468_ (.A(_2624_),
    .B(_3269_),
    .Y(_3285_));
 sg13g2_mux2_1 _7469_ (.A0(\board_state[92] ),
    .A1(net60),
    .S(_3285_),
    .X(_1112_));
 sg13g2_nor2_1 _7470_ (.A(_2628_),
    .B(_3269_),
    .Y(_3286_));
 sg13g2_mux2_1 _7471_ (.A0(\board_state[93] ),
    .A1(net60),
    .S(_3286_),
    .X(_1113_));
 sg13g2_nor2_1 _7472_ (.A(_2632_),
    .B(_3269_),
    .Y(_3287_));
 sg13g2_mux2_1 _7473_ (.A0(\board_state[94] ),
    .A1(_3281_),
    .S(_3287_),
    .X(_1114_));
 sg13g2_nor2_1 _7474_ (.A(_2637_),
    .B(_3269_),
    .Y(_3288_));
 sg13g2_mux2_1 _7475_ (.A0(\board_state[95] ),
    .A1(_3281_),
    .S(_3288_),
    .X(_1115_));
 sg13g2_nor2_1 _7476_ (.A(_2546_),
    .B(_2554_),
    .Y(_3289_));
 sg13g2_mux2_1 _7477_ (.A0(\board_state[96] ),
    .A1(net60),
    .S(_3289_),
    .X(_1116_));
 sg13g2_nor2_1 _7478_ (.A(_2554_),
    .B(net205),
    .Y(_3290_));
 sg13g2_mux2_1 _7479_ (.A0(\board_state[97] ),
    .A1(net60),
    .S(_3290_),
    .X(_1117_));
 sg13g2_nor2_1 _7480_ (.A(_2554_),
    .B(net204),
    .Y(_3291_));
 sg13g2_mux2_1 _7481_ (.A0(\board_state[98] ),
    .A1(net60),
    .S(_3291_),
    .X(_1118_));
 sg13g2_nor2_1 _7482_ (.A(_2554_),
    .B(_2590_),
    .Y(_3292_));
 sg13g2_mux2_1 _7483_ (.A0(\board_state[99] ),
    .A1(net67),
    .S(_3292_),
    .X(_1119_));
 sg13g2_nor2_1 _7484_ (.A(_2539_),
    .B(_2619_),
    .Y(_3293_));
 sg13g2_mux2_1 _7485_ (.A0(\board_state[9] ),
    .A1(net67),
    .S(_3293_),
    .X(_1120_));
 sg13g2_inv_1 _7486_ (.Y(_3294_),
    .A(\num_neighbors[0] ));
 sg13g2_buf_1 _7487_ (.A(_0002_),
    .X(_3295_));
 sg13g2_buf_2 _7488_ (.A(_3295_),
    .X(_3296_));
 sg13g2_buf_2 _7489_ (.A(net361),
    .X(_3297_));
 sg13g2_buf_1 _7490_ (.A(_0000_),
    .X(_3298_));
 sg13g2_buf_1 _7491_ (.A(_3298_),
    .X(_3299_));
 sg13g2_buf_1 _7492_ (.A(net360),
    .X(_3300_));
 sg13g2_mux4_1 _7493_ (.S0(net315),
    .A0(_0082_),
    .A1(_0087_),
    .A2(_0083_),
    .A3(_0088_),
    .S1(net314),
    .X(_3301_));
 sg13g2_mux4_1 _7494_ (.S0(net315),
    .A0(_0085_),
    .A1(_0089_),
    .A2(_0086_),
    .A3(_0090_),
    .S1(net314),
    .X(_3302_));
 sg13g2_buf_1 _7495_ (.A(_3295_),
    .X(_3303_));
 sg13g2_buf_2 _7496_ (.A(_3303_),
    .X(_3304_));
 sg13g2_buf_1 _7497_ (.A(_3298_),
    .X(_3305_));
 sg13g2_buf_1 _7498_ (.A(_3305_),
    .X(_3306_));
 sg13g2_mux4_1 _7499_ (.S0(net313),
    .A0(_0099_),
    .A1(_0103_),
    .A2(_0100_),
    .A3(_0104_),
    .S1(net312),
    .X(_3307_));
 sg13g2_mux4_1 _7500_ (.S0(net313),
    .A0(_0101_),
    .A1(_0105_),
    .A2(_0102_),
    .A3(_0106_),
    .S1(net312),
    .X(_3308_));
 sg13g2_buf_2 _7501_ (.A(_0001_),
    .X(_3309_));
 sg13g2_buf_2 _7502_ (.A(_3309_),
    .X(_3310_));
 sg13g2_buf_2 _7503_ (.A(_0004_),
    .X(_3311_));
 sg13g2_buf_1 _7504_ (.A(_3311_),
    .X(_3312_));
 sg13g2_mux4_1 _7505_ (.S0(_3310_),
    .A0(_3301_),
    .A1(_3302_),
    .A2(_3307_),
    .A3(_3308_),
    .S1(_3312_),
    .X(_3313_));
 sg13g2_mux4_1 _7506_ (.S0(net315),
    .A0(_0091_),
    .A1(_0095_),
    .A2(_0092_),
    .A3(_0096_),
    .S1(net314),
    .X(_3314_));
 sg13g2_mux4_1 _7507_ (.S0(net315),
    .A0(_0093_),
    .A1(_0097_),
    .A2(_0094_),
    .A3(_0098_),
    .S1(net314),
    .X(_3315_));
 sg13g2_mux4_1 _7508_ (.S0(net313),
    .A0(_0107_),
    .A1(_0111_),
    .A2(_0108_),
    .A3(_0112_),
    .S1(net312),
    .X(_3316_));
 sg13g2_buf_2 _7509_ (.A(_3303_),
    .X(_3317_));
 sg13g2_buf_1 _7510_ (.A(_3305_),
    .X(_3318_));
 sg13g2_mux4_1 _7511_ (.S0(net311),
    .A0(_0109_),
    .A1(_0113_),
    .A2(_0110_),
    .A3(_0114_),
    .S1(net310),
    .X(_3319_));
 sg13g2_mux4_1 _7512_ (.S0(net359),
    .A0(_3314_),
    .A1(_3315_),
    .A2(_3316_),
    .A3(_3319_),
    .S1(net358),
    .X(_3320_));
 sg13g2_mux4_1 _7513_ (.S0(net313),
    .A0(_0147_),
    .A1(_0151_),
    .A2(_0148_),
    .A3(_0152_),
    .S1(net312),
    .X(_3321_));
 sg13g2_mux4_1 _7514_ (.S0(net313),
    .A0(_0149_),
    .A1(_0153_),
    .A2(_0150_),
    .A3(_0154_),
    .S1(net312),
    .X(_3322_));
 sg13g2_buf_2 _7515_ (.A(_3303_),
    .X(_3323_));
 sg13g2_buf_1 _7516_ (.A(_3305_),
    .X(_3324_));
 sg13g2_mux4_1 _7517_ (.S0(_3323_),
    .A0(_0163_),
    .A1(_0167_),
    .A2(_0164_),
    .A3(_0168_),
    .S1(_3324_),
    .X(_3325_));
 sg13g2_mux4_1 _7518_ (.S0(_3323_),
    .A0(_0165_),
    .A1(_0169_),
    .A2(_0166_),
    .A3(_0170_),
    .S1(_3324_),
    .X(_3326_));
 sg13g2_buf_2 _7519_ (.A(_3309_),
    .X(_3327_));
 sg13g2_buf_1 _7520_ (.A(_3311_),
    .X(_3328_));
 sg13g2_mux4_1 _7521_ (.S0(net357),
    .A0(_3321_),
    .A1(_3322_),
    .A2(_3325_),
    .A3(_3326_),
    .S1(net356),
    .X(_3329_));
 sg13g2_mux4_1 _7522_ (.S0(net313),
    .A0(_0155_),
    .A1(_0159_),
    .A2(_0156_),
    .A3(_0160_),
    .S1(net312),
    .X(_3330_));
 sg13g2_mux4_1 _7523_ (.S0(net311),
    .A0(_0157_),
    .A1(_0161_),
    .A2(_0158_),
    .A3(_0162_),
    .S1(net310),
    .X(_3331_));
 sg13g2_mux4_1 _7524_ (.S0(net309),
    .A0(_0171_),
    .A1(_0175_),
    .A2(_0172_),
    .A3(_0176_),
    .S1(net308),
    .X(_3332_));
 sg13g2_buf_2 _7525_ (.A(_3303_),
    .X(_3333_));
 sg13g2_buf_1 _7526_ (.A(_3305_),
    .X(_3334_));
 sg13g2_mux4_1 _7527_ (.S0(net307),
    .A0(_0173_),
    .A1(_0177_),
    .A2(_0174_),
    .A3(_0178_),
    .S1(net306),
    .X(_3335_));
 sg13g2_mux4_1 _7528_ (.S0(net357),
    .A0(_3330_),
    .A1(_3331_),
    .A2(_3332_),
    .A3(_3335_),
    .S1(net356),
    .X(_3336_));
 sg13g2_buf_8 _7529_ (.A(_0003_),
    .X(_3337_));
 sg13g2_buf_4 _7530_ (.X(_3338_),
    .A(_0006_));
 sg13g2_mux4_1 _7531_ (.S0(_3337_),
    .A0(_3313_),
    .A1(_3320_),
    .A2(_3329_),
    .A3(_3336_),
    .S1(_3338_),
    .X(_3339_));
 sg13g2_mux4_1 _7532_ (.S0(net315),
    .A0(_0115_),
    .A1(_0119_),
    .A2(_0116_),
    .A3(_0120_),
    .S1(net314),
    .X(_3340_));
 sg13g2_mux4_1 _7533_ (.S0(net315),
    .A0(_0117_),
    .A1(_0121_),
    .A2(_0118_),
    .A3(_0122_),
    .S1(net314),
    .X(_3341_));
 sg13g2_mux4_1 _7534_ (.S0(_3304_),
    .A0(_0131_),
    .A1(_0135_),
    .A2(_0132_),
    .A3(_0136_),
    .S1(_3306_),
    .X(_3342_));
 sg13g2_mux4_1 _7535_ (.S0(_3317_),
    .A0(_0133_),
    .A1(_0137_),
    .A2(_0134_),
    .A3(_0138_),
    .S1(_3318_),
    .X(_3343_));
 sg13g2_mux4_1 _7536_ (.S0(net359),
    .A0(_3340_),
    .A1(_3341_),
    .A2(_3342_),
    .A3(_3343_),
    .S1(net358),
    .X(_3344_));
 sg13g2_mux4_1 _7537_ (.S0(net315),
    .A0(_0123_),
    .A1(_0127_),
    .A2(_0124_),
    .A3(_0128_),
    .S1(net314),
    .X(_3345_));
 sg13g2_mux4_1 _7538_ (.S0(net315),
    .A0(_0125_),
    .A1(_0129_),
    .A2(_0126_),
    .A3(_0130_),
    .S1(net314),
    .X(_3346_));
 sg13g2_mux4_1 _7539_ (.S0(net311),
    .A0(_0139_),
    .A1(_0143_),
    .A2(_0140_),
    .A3(_0144_),
    .S1(net310),
    .X(_3347_));
 sg13g2_buf_2 _7540_ (.A(net361),
    .X(_3348_));
 sg13g2_buf_1 _7541_ (.A(net360),
    .X(_3349_));
 sg13g2_mux4_1 _7542_ (.S0(net305),
    .A0(_0141_),
    .A1(_0145_),
    .A2(_0142_),
    .A3(_0146_),
    .S1(net304),
    .X(_3350_));
 sg13g2_mux4_1 _7543_ (.S0(net359),
    .A0(_3345_),
    .A1(_3346_),
    .A2(_3347_),
    .A3(_3350_),
    .S1(net358),
    .X(_3351_));
 sg13g2_mux4_1 _7544_ (.S0(_3304_),
    .A0(_0179_),
    .A1(_0183_),
    .A2(_0180_),
    .A3(_0184_),
    .S1(_3306_),
    .X(_3352_));
 sg13g2_mux4_1 _7545_ (.S0(_3317_),
    .A0(_0181_),
    .A1(_0185_),
    .A2(_0182_),
    .A3(_0186_),
    .S1(_3318_),
    .X(_3353_));
 sg13g2_mux4_1 _7546_ (.S0(net307),
    .A0(_0195_),
    .A1(_0199_),
    .A2(_0196_),
    .A3(_0200_),
    .S1(net306),
    .X(_3354_));
 sg13g2_mux4_1 _7547_ (.S0(_3333_),
    .A0(_0197_),
    .A1(_0201_),
    .A2(_0198_),
    .A3(_0202_),
    .S1(_3334_),
    .X(_3355_));
 sg13g2_mux4_1 _7548_ (.S0(net357),
    .A0(_3352_),
    .A1(_3353_),
    .A2(_3354_),
    .A3(_3355_),
    .S1(net356),
    .X(_3356_));
 sg13g2_mux4_1 _7549_ (.S0(net311),
    .A0(_0187_),
    .A1(_0191_),
    .A2(_0188_),
    .A3(_0192_),
    .S1(net310),
    .X(_3357_));
 sg13g2_mux4_1 _7550_ (.S0(net305),
    .A0(_0189_),
    .A1(_0193_),
    .A2(_0190_),
    .A3(_0194_),
    .S1(net304),
    .X(_3358_));
 sg13g2_mux4_1 _7551_ (.S0(_3333_),
    .A0(_0203_),
    .A1(_0207_),
    .A2(_0204_),
    .A3(_0208_),
    .S1(_3334_),
    .X(_3359_));
 sg13g2_buf_2 _7552_ (.A(_3303_),
    .X(_3360_));
 sg13g2_buf_1 _7553_ (.A(_3305_),
    .X(_3361_));
 sg13g2_mux4_1 _7554_ (.S0(net303),
    .A0(_0205_),
    .A1(_0209_),
    .A2(_0206_),
    .A3(_0210_),
    .S1(net302),
    .X(_3362_));
 sg13g2_mux4_1 _7555_ (.S0(_3310_),
    .A0(_3357_),
    .A1(_3358_),
    .A2(_3359_),
    .A3(_3362_),
    .S1(_3312_),
    .X(_3363_));
 sg13g2_mux4_1 _7556_ (.S0(_3337_),
    .A0(_3344_),
    .A1(_3351_),
    .A2(_3356_),
    .A3(_3363_),
    .S1(_3338_),
    .X(_3364_));
 sg13g2_mux4_1 _7557_ (.S0(net313),
    .A0(_0339_),
    .A1(_0343_),
    .A2(_0340_),
    .A3(_0344_),
    .S1(net312),
    .X(_3365_));
 sg13g2_mux4_1 _7558_ (.S0(net311),
    .A0(_0341_),
    .A1(_0345_),
    .A2(_0342_),
    .A3(_0346_),
    .S1(net310),
    .X(_3366_));
 sg13g2_mux4_1 _7559_ (.S0(net309),
    .A0(_0355_),
    .A1(_0359_),
    .A2(_0356_),
    .A3(_0360_),
    .S1(net308),
    .X(_3367_));
 sg13g2_mux4_1 _7560_ (.S0(net309),
    .A0(_0357_),
    .A1(_0361_),
    .A2(_0358_),
    .A3(_0362_),
    .S1(net306),
    .X(_3368_));
 sg13g2_mux4_1 _7561_ (.S0(net357),
    .A0(_3365_),
    .A1(_3366_),
    .A2(_3367_),
    .A3(_3368_),
    .S1(net356),
    .X(_3369_));
 sg13g2_mux4_1 _7562_ (.S0(net311),
    .A0(_0347_),
    .A1(_0351_),
    .A2(_0348_),
    .A3(_0352_),
    .S1(net310),
    .X(_3370_));
 sg13g2_mux4_1 _7563_ (.S0(net305),
    .A0(_0349_),
    .A1(_0353_),
    .A2(_0350_),
    .A3(_0354_),
    .S1(net304),
    .X(_3371_));
 sg13g2_mux4_1 _7564_ (.S0(net307),
    .A0(_0363_),
    .A1(_0367_),
    .A2(_0364_),
    .A3(_0368_),
    .S1(net306),
    .X(_3372_));
 sg13g2_mux4_1 _7565_ (.S0(net303),
    .A0(_0365_),
    .A1(_0369_),
    .A2(_0366_),
    .A3(_0370_),
    .S1(net302),
    .X(_3373_));
 sg13g2_mux4_1 _7566_ (.S0(net357),
    .A0(_3370_),
    .A1(_3371_),
    .A2(_3372_),
    .A3(_3373_),
    .S1(net356),
    .X(_3374_));
 sg13g2_mux4_1 _7567_ (.S0(net309),
    .A0(_0403_),
    .A1(_0407_),
    .A2(_0404_),
    .A3(_0408_),
    .S1(net308),
    .X(_3375_));
 sg13g2_mux4_1 _7568_ (.S0(net307),
    .A0(_0405_),
    .A1(_0409_),
    .A2(_0406_),
    .A3(_0410_),
    .S1(net306),
    .X(_3376_));
 sg13g2_buf_2 _7569_ (.A(_3295_),
    .X(_3377_));
 sg13g2_buf_1 _7570_ (.A(_3298_),
    .X(_3378_));
 sg13g2_mux4_1 _7571_ (.S0(net355),
    .A0(_0419_),
    .A1(_0423_),
    .A2(_0420_),
    .A3(_0424_),
    .S1(net354),
    .X(_3379_));
 sg13g2_mux4_1 _7572_ (.S0(net355),
    .A0(_0421_),
    .A1(_0425_),
    .A2(_0422_),
    .A3(_0426_),
    .S1(net354),
    .X(_3380_));
 sg13g2_buf_2 _7573_ (.A(_3309_),
    .X(_3381_));
 sg13g2_buf_1 _7574_ (.A(_3311_),
    .X(_3382_));
 sg13g2_mux4_1 _7575_ (.S0(net353),
    .A0(_3375_),
    .A1(_3376_),
    .A2(_3379_),
    .A3(_3380_),
    .S1(net352),
    .X(_3383_));
 sg13g2_mux4_1 _7576_ (.S0(net307),
    .A0(_0411_),
    .A1(_0415_),
    .A2(_0412_),
    .A3(_0416_),
    .S1(net308),
    .X(_3384_));
 sg13g2_mux4_1 _7577_ (.S0(net303),
    .A0(_0413_),
    .A1(_0417_),
    .A2(_0414_),
    .A3(_0418_),
    .S1(net302),
    .X(_3385_));
 sg13g2_mux4_1 _7578_ (.S0(net355),
    .A0(_0427_),
    .A1(_0431_),
    .A2(_0428_),
    .A3(_0432_),
    .S1(net354),
    .X(_3386_));
 sg13g2_mux4_1 _7579_ (.S0(net355),
    .A0(_0429_),
    .A1(_0433_),
    .A2(_0430_),
    .A3(_0434_),
    .S1(net354),
    .X(_3387_));
 sg13g2_mux4_1 _7580_ (.S0(net353),
    .A0(_3384_),
    .A1(_3385_),
    .A2(_3386_),
    .A3(_3387_),
    .S1(net352),
    .X(_3388_));
 sg13g2_mux4_1 _7581_ (.S0(_3337_),
    .A0(_3369_),
    .A1(_3374_),
    .A2(_3383_),
    .A3(_3388_),
    .S1(_3338_),
    .X(_3389_));
 sg13g2_mux4_1 _7582_ (.S0(net313),
    .A0(_0371_),
    .A1(_0375_),
    .A2(_0372_),
    .A3(_0376_),
    .S1(net312),
    .X(_3390_));
 sg13g2_mux4_1 _7583_ (.S0(net311),
    .A0(_0373_),
    .A1(_0377_),
    .A2(_0374_),
    .A3(_0378_),
    .S1(net310),
    .X(_3391_));
 sg13g2_mux4_1 _7584_ (.S0(net309),
    .A0(_0387_),
    .A1(_0391_),
    .A2(_0388_),
    .A3(_0392_),
    .S1(net308),
    .X(_3392_));
 sg13g2_mux4_1 _7585_ (.S0(net307),
    .A0(_0389_),
    .A1(_0393_),
    .A2(_0390_),
    .A3(_0394_),
    .S1(net306),
    .X(_3393_));
 sg13g2_mux4_1 _7586_ (.S0(net357),
    .A0(_3390_),
    .A1(_3391_),
    .A2(_3392_),
    .A3(_3393_),
    .S1(net356),
    .X(_3394_));
 sg13g2_mux4_1 _7587_ (.S0(net311),
    .A0(_0379_),
    .A1(_0383_),
    .A2(_0380_),
    .A3(_0384_),
    .S1(net310),
    .X(_3395_));
 sg13g2_mux4_1 _7588_ (.S0(net305),
    .A0(_0381_),
    .A1(_0385_),
    .A2(_0382_),
    .A3(_0386_),
    .S1(net304),
    .X(_3396_));
 sg13g2_mux4_1 _7589_ (.S0(net303),
    .A0(_0395_),
    .A1(_0399_),
    .A2(_0396_),
    .A3(_0400_),
    .S1(net302),
    .X(_3397_));
 sg13g2_mux4_1 _7590_ (.S0(net303),
    .A0(_0397_),
    .A1(_0401_),
    .A2(_0398_),
    .A3(_0402_),
    .S1(net302),
    .X(_3398_));
 sg13g2_mux4_1 _7591_ (.S0(net359),
    .A0(_3395_),
    .A1(_3396_),
    .A2(_3397_),
    .A3(_3398_),
    .S1(net358),
    .X(_3399_));
 sg13g2_mux4_1 _7592_ (.S0(net309),
    .A0(_0435_),
    .A1(_0439_),
    .A2(_0436_),
    .A3(_0440_),
    .S1(net308),
    .X(_3400_));
 sg13g2_mux4_1 _7593_ (.S0(net307),
    .A0(_0437_),
    .A1(_0441_),
    .A2(_0438_),
    .A3(_0442_),
    .S1(net306),
    .X(_3401_));
 sg13g2_mux4_1 _7594_ (.S0(net355),
    .A0(_0451_),
    .A1(_0455_),
    .A2(_0452_),
    .A3(_0456_),
    .S1(net354),
    .X(_3402_));
 sg13g2_mux4_1 _7595_ (.S0(net355),
    .A0(_0453_),
    .A1(_0457_),
    .A2(_0454_),
    .A3(_0458_),
    .S1(net354),
    .X(_3403_));
 sg13g2_mux4_1 _7596_ (.S0(net353),
    .A0(_3400_),
    .A1(_3401_),
    .A2(_3402_),
    .A3(_3403_),
    .S1(net352),
    .X(_3404_));
 sg13g2_mux4_1 _7597_ (.S0(net307),
    .A0(_0443_),
    .A1(_0447_),
    .A2(_0444_),
    .A3(_0448_),
    .S1(net306),
    .X(_3405_));
 sg13g2_mux4_1 _7598_ (.S0(net303),
    .A0(_0445_),
    .A1(_0449_),
    .A2(_0446_),
    .A3(_0450_),
    .S1(net302),
    .X(_3406_));
 sg13g2_mux4_1 _7599_ (.S0(net355),
    .A0(_0459_),
    .A1(_0463_),
    .A2(_0460_),
    .A3(_0464_),
    .S1(net354),
    .X(_3407_));
 sg13g2_mux4_1 _7600_ (.S0(_3377_),
    .A0(_0461_),
    .A1(_0465_),
    .A2(_0462_),
    .A3(_0466_),
    .S1(_3378_),
    .X(_3408_));
 sg13g2_mux4_1 _7601_ (.S0(net353),
    .A0(_3405_),
    .A1(_3406_),
    .A2(_3407_),
    .A3(_3408_),
    .S1(net352),
    .X(_3409_));
 sg13g2_mux4_1 _7602_ (.S0(_3337_),
    .A0(_3394_),
    .A1(_3399_),
    .A2(_3404_),
    .A3(_3409_),
    .S1(_3338_),
    .X(_3410_));
 sg13g2_mux4_1 _7603_ (.S0(_0005_),
    .A0(_3339_),
    .A1(_3364_),
    .A2(_3389_),
    .A3(_3410_),
    .S1(_0008_),
    .X(_3411_));
 sg13g2_mux4_1 _7604_ (.S0(net305),
    .A0(_0211_),
    .A1(_0215_),
    .A2(_0212_),
    .A3(_0216_),
    .S1(net304),
    .X(_3412_));
 sg13g2_mux4_1 _7605_ (.S0(net305),
    .A0(_0213_),
    .A1(_0217_),
    .A2(_0214_),
    .A3(_0218_),
    .S1(net304),
    .X(_3413_));
 sg13g2_mux4_1 _7606_ (.S0(net303),
    .A0(_0227_),
    .A1(_0231_),
    .A2(_0228_),
    .A3(_0232_),
    .S1(net302),
    .X(_3414_));
 sg13g2_buf_1 _7607_ (.A(_3305_),
    .X(_3415_));
 sg13g2_mux4_1 _7608_ (.S0(_3360_),
    .A0(_0229_),
    .A1(_0233_),
    .A2(_0230_),
    .A3(_0234_),
    .S1(net301),
    .X(_3416_));
 sg13g2_mux4_1 _7609_ (.S0(net359),
    .A0(_3412_),
    .A1(_3413_),
    .A2(_3414_),
    .A3(_3416_),
    .S1(net358),
    .X(_3417_));
 sg13g2_mux4_1 _7610_ (.S0(net305),
    .A0(_0219_),
    .A1(_0223_),
    .A2(_0220_),
    .A3(_0224_),
    .S1(net304),
    .X(_3418_));
 sg13g2_mux4_1 _7611_ (.S0(net305),
    .A0(_0221_),
    .A1(_0225_),
    .A2(_0222_),
    .A3(_0226_),
    .S1(net304),
    .X(_3419_));
 sg13g2_buf_2 _7612_ (.A(_3303_),
    .X(_3420_));
 sg13g2_mux4_1 _7613_ (.S0(net300),
    .A0(_0235_),
    .A1(_0239_),
    .A2(_0236_),
    .A3(_0240_),
    .S1(net301),
    .X(_3421_));
 sg13g2_buf_2 _7614_ (.A(_3303_),
    .X(_3422_));
 sg13g2_buf_1 _7615_ (.A(_3305_),
    .X(_3423_));
 sg13g2_mux4_1 _7616_ (.S0(net299),
    .A0(_0237_),
    .A1(_0241_),
    .A2(_0238_),
    .A3(_0242_),
    .S1(net298),
    .X(_3424_));
 sg13g2_mux4_1 _7617_ (.S0(net359),
    .A0(_3418_),
    .A1(_3419_),
    .A2(_3421_),
    .A3(_3424_),
    .S1(net358),
    .X(_3425_));
 sg13g2_mux4_1 _7618_ (.S0(_3360_),
    .A0(_0275_),
    .A1(_0279_),
    .A2(_0276_),
    .A3(_0280_),
    .S1(_3361_),
    .X(_3426_));
 sg13g2_mux4_1 _7619_ (.S0(net300),
    .A0(_0277_),
    .A1(_0281_),
    .A2(_0278_),
    .A3(_0282_),
    .S1(net301),
    .X(_3427_));
 sg13g2_mux4_1 _7620_ (.S0(net355),
    .A0(_0291_),
    .A1(_0295_),
    .A2(_0292_),
    .A3(_0296_),
    .S1(net354),
    .X(_3428_));
 sg13g2_buf_2 _7621_ (.A(_3295_),
    .X(_3429_));
 sg13g2_buf_1 _7622_ (.A(_3298_),
    .X(_3430_));
 sg13g2_mux4_1 _7623_ (.S0(net351),
    .A0(_0293_),
    .A1(_0297_),
    .A2(_0294_),
    .A3(_0298_),
    .S1(net350),
    .X(_3431_));
 sg13g2_mux4_1 _7624_ (.S0(net353),
    .A0(_3426_),
    .A1(_3427_),
    .A2(_3428_),
    .A3(_3431_),
    .S1(net352),
    .X(_3432_));
 sg13g2_mux4_1 _7625_ (.S0(net300),
    .A0(_0283_),
    .A1(_0287_),
    .A2(_0284_),
    .A3(_0288_),
    .S1(_3361_),
    .X(_3433_));
 sg13g2_mux4_1 _7626_ (.S0(net300),
    .A0(_0285_),
    .A1(_0289_),
    .A2(_0286_),
    .A3(_0290_),
    .S1(net301),
    .X(_3434_));
 sg13g2_mux4_1 _7627_ (.S0(net351),
    .A0(_0299_),
    .A1(_0303_),
    .A2(_0300_),
    .A3(_0304_),
    .S1(net350),
    .X(_3435_));
 sg13g2_buf_2 _7628_ (.A(_3295_),
    .X(_3436_));
 sg13g2_buf_1 _7629_ (.A(_3298_),
    .X(_3437_));
 sg13g2_mux4_1 _7630_ (.S0(net349),
    .A0(_0301_),
    .A1(_0305_),
    .A2(_0302_),
    .A3(_0306_),
    .S1(net348),
    .X(_3438_));
 sg13g2_mux4_1 _7631_ (.S0(net353),
    .A0(_3433_),
    .A1(_3434_),
    .A2(_3435_),
    .A3(_3438_),
    .S1(net352),
    .X(_3439_));
 sg13g2_mux4_1 _7632_ (.S0(_3337_),
    .A0(_3417_),
    .A1(_3425_),
    .A2(_3432_),
    .A3(_3439_),
    .S1(_3338_),
    .X(_3440_));
 sg13g2_mux4_1 _7633_ (.S0(_3348_),
    .A0(_0243_),
    .A1(_0247_),
    .A2(_0244_),
    .A3(_0248_),
    .S1(_3349_),
    .X(_3441_));
 sg13g2_mux4_1 _7634_ (.S0(_3297_),
    .A0(_0245_),
    .A1(_0249_),
    .A2(_0246_),
    .A3(_0250_),
    .S1(_3349_),
    .X(_3442_));
 sg13g2_mux4_1 _7635_ (.S0(net300),
    .A0(_0259_),
    .A1(_0263_),
    .A2(_0260_),
    .A3(_0264_),
    .S1(net301),
    .X(_3443_));
 sg13g2_mux4_1 _7636_ (.S0(_3420_),
    .A0(_0261_),
    .A1(_0265_),
    .A2(_0262_),
    .A3(_0266_),
    .S1(net298),
    .X(_3444_));
 sg13g2_mux4_1 _7637_ (.S0(net359),
    .A0(_3441_),
    .A1(_3442_),
    .A2(_3443_),
    .A3(_3444_),
    .S1(net358),
    .X(_3445_));
 sg13g2_mux4_1 _7638_ (.S0(_3348_),
    .A0(_0251_),
    .A1(_0255_),
    .A2(_0252_),
    .A3(_0256_),
    .S1(_3300_),
    .X(_3446_));
 sg13g2_mux4_1 _7639_ (.S0(_3297_),
    .A0(_0253_),
    .A1(_0257_),
    .A2(_0254_),
    .A3(_0258_),
    .S1(_3300_),
    .X(_3447_));
 sg13g2_mux4_1 _7640_ (.S0(net299),
    .A0(_0267_),
    .A1(_0271_),
    .A2(_0268_),
    .A3(_0272_),
    .S1(net298),
    .X(_3448_));
 sg13g2_mux4_1 _7641_ (.S0(net299),
    .A0(_0269_),
    .A1(_0273_),
    .A2(_0270_),
    .A3(_0274_),
    .S1(net298),
    .X(_3449_));
 sg13g2_mux4_1 _7642_ (.S0(net359),
    .A0(_3446_),
    .A1(_3447_),
    .A2(_3448_),
    .A3(_3449_),
    .S1(net358),
    .X(_3450_));
 sg13g2_mux4_1 _7643_ (.S0(_3420_),
    .A0(_0307_),
    .A1(_0311_),
    .A2(_0308_),
    .A3(_0312_),
    .S1(_3415_),
    .X(_3451_));
 sg13g2_mux4_1 _7644_ (.S0(net299),
    .A0(_0309_),
    .A1(_0313_),
    .A2(_0310_),
    .A3(_0314_),
    .S1(_3423_),
    .X(_3452_));
 sg13g2_mux4_1 _7645_ (.S0(net351),
    .A0(_0323_),
    .A1(_0327_),
    .A2(_0324_),
    .A3(_0328_),
    .S1(net350),
    .X(_3453_));
 sg13g2_mux4_1 _7646_ (.S0(net349),
    .A0(_0325_),
    .A1(_0329_),
    .A2(_0326_),
    .A3(_0330_),
    .S1(net348),
    .X(_3454_));
 sg13g2_mux4_1 _7647_ (.S0(net357),
    .A0(_3451_),
    .A1(_3452_),
    .A2(_3453_),
    .A3(_3454_),
    .S1(net356),
    .X(_3455_));
 sg13g2_mux4_1 _7648_ (.S0(_3422_),
    .A0(_0315_),
    .A1(_0319_),
    .A2(_0316_),
    .A3(_0320_),
    .S1(_3415_),
    .X(_3456_));
 sg13g2_mux4_1 _7649_ (.S0(_3422_),
    .A0(_0317_),
    .A1(_0321_),
    .A2(_0318_),
    .A3(_0322_),
    .S1(_3423_),
    .X(_3457_));
 sg13g2_mux4_1 _7650_ (.S0(net349),
    .A0(_0331_),
    .A1(_0335_),
    .A2(_0332_),
    .A3(_0336_),
    .S1(net348),
    .X(_3458_));
 sg13g2_mux4_1 _7651_ (.S0(net349),
    .A0(_0333_),
    .A1(_0337_),
    .A2(_0334_),
    .A3(_0338_),
    .S1(net348),
    .X(_3459_));
 sg13g2_mux4_1 _7652_ (.S0(net357),
    .A0(_3456_),
    .A1(_3457_),
    .A2(_3458_),
    .A3(_3459_),
    .S1(net356),
    .X(_3460_));
 sg13g2_mux4_1 _7653_ (.S0(_3337_),
    .A0(_3445_),
    .A1(_3450_),
    .A2(_3455_),
    .A3(_3460_),
    .S1(_3338_),
    .X(_3461_));
 sg13g2_mux4_1 _7654_ (.S0(net303),
    .A0(_0467_),
    .A1(_0471_),
    .A2(_0468_),
    .A3(_0472_),
    .S1(net302),
    .X(_3462_));
 sg13g2_mux4_1 _7655_ (.S0(net300),
    .A0(_0469_),
    .A1(_0473_),
    .A2(_0470_),
    .A3(_0474_),
    .S1(net301),
    .X(_3463_));
 sg13g2_mux4_1 _7656_ (.S0(_3377_),
    .A0(_0483_),
    .A1(_0487_),
    .A2(_0484_),
    .A3(_0488_),
    .S1(_3378_),
    .X(_3464_));
 sg13g2_mux4_1 _7657_ (.S0(net351),
    .A0(_0485_),
    .A1(_0489_),
    .A2(_0486_),
    .A3(_0490_),
    .S1(net350),
    .X(_3465_));
 sg13g2_mux4_1 _7658_ (.S0(net353),
    .A0(_3462_),
    .A1(_3463_),
    .A2(_3464_),
    .A3(_3465_),
    .S1(net352),
    .X(_3466_));
 sg13g2_mux4_1 _7659_ (.S0(net300),
    .A0(_0475_),
    .A1(_0479_),
    .A2(_0476_),
    .A3(_0480_),
    .S1(net301),
    .X(_3467_));
 sg13g2_mux4_1 _7660_ (.S0(net299),
    .A0(_0477_),
    .A1(_0481_),
    .A2(_0478_),
    .A3(_0482_),
    .S1(net298),
    .X(_3468_));
 sg13g2_mux4_1 _7661_ (.S0(net351),
    .A0(_0491_),
    .A1(_0495_),
    .A2(_0492_),
    .A3(_0496_),
    .S1(net350),
    .X(_3469_));
 sg13g2_mux4_1 _7662_ (.S0(net349),
    .A0(_0493_),
    .A1(_0497_),
    .A2(_0494_),
    .A3(_0498_),
    .S1(net348),
    .X(_3470_));
 sg13g2_mux4_1 _7663_ (.S0(_3327_),
    .A0(_3467_),
    .A1(_3468_),
    .A2(_3469_),
    .A3(_3470_),
    .S1(_3328_),
    .X(_3471_));
 sg13g2_mux4_1 _7664_ (.S0(net351),
    .A0(_0531_),
    .A1(_0535_),
    .A2(_0532_),
    .A3(_0536_),
    .S1(net350),
    .X(_3472_));
 sg13g2_mux4_1 _7665_ (.S0(net351),
    .A0(_0533_),
    .A1(_0537_),
    .A2(_0534_),
    .A3(_0538_),
    .S1(net350),
    .X(_3473_));
 sg13g2_mux4_1 _7666_ (.S0(net361),
    .A0(_0547_),
    .A1(_0551_),
    .A2(_0548_),
    .A3(_0552_),
    .S1(net360),
    .X(_3474_));
 sg13g2_mux4_1 _7667_ (.S0(net361),
    .A0(_0549_),
    .A1(_0553_),
    .A2(_0550_),
    .A3(_0554_),
    .S1(net360),
    .X(_3475_));
 sg13g2_mux4_1 _7668_ (.S0(_3309_),
    .A0(_3472_),
    .A1(_3473_),
    .A2(_3474_),
    .A3(_3475_),
    .S1(_3311_),
    .X(_3476_));
 sg13g2_mux4_1 _7669_ (.S0(net351),
    .A0(_0539_),
    .A1(_0543_),
    .A2(_0540_),
    .A3(_0544_),
    .S1(net350),
    .X(_3477_));
 sg13g2_mux4_1 _7670_ (.S0(net349),
    .A0(_0541_),
    .A1(_0545_),
    .A2(_0542_),
    .A3(_0546_),
    .S1(net348),
    .X(_3478_));
 sg13g2_mux4_1 _7671_ (.S0(net361),
    .A0(_0555_),
    .A1(_0559_),
    .A2(_0556_),
    .A3(_0560_),
    .S1(net360),
    .X(_3479_));
 sg13g2_mux4_1 _7672_ (.S0(net361),
    .A0(_0557_),
    .A1(_0561_),
    .A2(_0558_),
    .A3(_0562_),
    .S1(net360),
    .X(_3480_));
 sg13g2_mux4_1 _7673_ (.S0(net353),
    .A0(_3477_),
    .A1(_3478_),
    .A2(_3479_),
    .A3(_3480_),
    .S1(net352),
    .X(_3481_));
 sg13g2_mux4_1 _7674_ (.S0(_3337_),
    .A0(_3466_),
    .A1(_3471_),
    .A2(_3476_),
    .A3(_3481_),
    .S1(_3338_),
    .X(_3482_));
 sg13g2_mux4_1 _7675_ (.S0(net300),
    .A0(_0499_),
    .A1(_0503_),
    .A2(_0500_),
    .A3(_0504_),
    .S1(net301),
    .X(_3483_));
 sg13g2_mux4_1 _7676_ (.S0(net299),
    .A0(_0501_),
    .A1(_0505_),
    .A2(_0502_),
    .A3(_0506_),
    .S1(net298),
    .X(_3484_));
 sg13g2_mux4_1 _7677_ (.S0(_3429_),
    .A0(_0515_),
    .A1(_0519_),
    .A2(_0516_),
    .A3(_0520_),
    .S1(_3430_),
    .X(_3485_));
 sg13g2_mux4_1 _7678_ (.S0(net349),
    .A0(_0517_),
    .A1(_0521_),
    .A2(_0518_),
    .A3(_0522_),
    .S1(net348),
    .X(_3486_));
 sg13g2_mux4_1 _7679_ (.S0(_3381_),
    .A0(_3483_),
    .A1(_3484_),
    .A2(_3485_),
    .A3(_3486_),
    .S1(_3382_),
    .X(_3487_));
 sg13g2_mux4_1 _7680_ (.S0(net299),
    .A0(_0507_),
    .A1(_0511_),
    .A2(_0508_),
    .A3(_0512_),
    .S1(net298),
    .X(_3488_));
 sg13g2_mux4_1 _7681_ (.S0(net299),
    .A0(_0509_),
    .A1(_0513_),
    .A2(_0510_),
    .A3(_0514_),
    .S1(net298),
    .X(_3489_));
 sg13g2_mux4_1 _7682_ (.S0(net349),
    .A0(_0523_),
    .A1(_0527_),
    .A2(_0524_),
    .A3(_0528_),
    .S1(net348),
    .X(_3490_));
 sg13g2_mux4_1 _7683_ (.S0(net309),
    .A0(_0525_),
    .A1(_0529_),
    .A2(_0526_),
    .A3(_0530_),
    .S1(net308),
    .X(_3491_));
 sg13g2_mux4_1 _7684_ (.S0(_3327_),
    .A0(_3488_),
    .A1(_3489_),
    .A2(_3490_),
    .A3(_3491_),
    .S1(_3328_),
    .X(_3492_));
 sg13g2_mux4_1 _7685_ (.S0(_3429_),
    .A0(_0563_),
    .A1(_0567_),
    .A2(_0564_),
    .A3(_0568_),
    .S1(_3430_),
    .X(_3493_));
 sg13g2_mux4_1 _7686_ (.S0(_3436_),
    .A0(_0565_),
    .A1(_0569_),
    .A2(_0566_),
    .A3(_0570_),
    .S1(_3437_),
    .X(_3494_));
 sg13g2_mux4_1 _7687_ (.S0(net361),
    .A0(_0579_),
    .A1(_0583_),
    .A2(_0580_),
    .A3(_0584_),
    .S1(net360),
    .X(_3495_));
 sg13g2_mux4_1 _7688_ (.S0(net361),
    .A0(_0581_),
    .A1(_0585_),
    .A2(_0582_),
    .A3(_0586_),
    .S1(net360),
    .X(_3496_));
 sg13g2_mux4_1 _7689_ (.S0(_3309_),
    .A0(_3493_),
    .A1(_3494_),
    .A2(_3495_),
    .A3(_3496_),
    .S1(_3311_),
    .X(_3497_));
 sg13g2_mux4_1 _7690_ (.S0(_3436_),
    .A0(_0571_),
    .A1(_0575_),
    .A2(_0572_),
    .A3(_0576_),
    .S1(_3437_),
    .X(_3498_));
 sg13g2_mux4_1 _7691_ (.S0(net309),
    .A0(_0573_),
    .A1(_0577_),
    .A2(_0574_),
    .A3(_0578_),
    .S1(net308),
    .X(_3499_));
 sg13g2_mux4_1 _7692_ (.S0(_3296_),
    .A0(_0587_),
    .A1(_0591_),
    .A2(_0588_),
    .A3(_0592_),
    .S1(_3299_),
    .X(_3500_));
 sg13g2_mux4_1 _7693_ (.S0(_3296_),
    .A0(_0589_),
    .A1(_0593_),
    .A2(_0590_),
    .A3(_0594_),
    .S1(_3299_),
    .X(_3501_));
 sg13g2_mux4_1 _7694_ (.S0(_3381_),
    .A0(_3498_),
    .A1(_3499_),
    .A2(_3500_),
    .A3(_3501_),
    .S1(_3382_),
    .X(_3502_));
 sg13g2_mux4_1 _7695_ (.S0(_3337_),
    .A0(_3487_),
    .A1(_3492_),
    .A2(_3497_),
    .A3(_3502_),
    .S1(_3338_),
    .X(_3503_));
 sg13g2_mux4_1 _7696_ (.S0(_0005_),
    .A0(_3440_),
    .A1(_3461_),
    .A2(_3482_),
    .A3(_3503_),
    .S1(_0008_),
    .X(_3504_));
 sg13g2_mux2_1 _7697_ (.A0(_3411_),
    .A1(_3504_),
    .S(_0007_),
    .X(_3505_));
 sg13g2_inv_1 _7698_ (.Y(_3506_),
    .A(\num_neighbors[1] ));
 sg13g2_buf_1 _7699_ (.A(\num_neighbors[2] ),
    .X(_3507_));
 sg13g2_or4_1 _7700_ (.A(_1785_),
    .B(_3506_),
    .C(_3507_),
    .D(\num_neighbors[3] ),
    .X(_3508_));
 sg13g2_a21oi_1 _7701_ (.A1(_3294_),
    .A2(_3505_),
    .Y(_3509_),
    .B1(_3508_));
 sg13g2_a22oi_1 _7702_ (.Y(_3510_),
    .B1(_2011_),
    .B2(_2086_),
    .A2(_2007_),
    .A1(_1785_));
 sg13g2_or2_1 _7703_ (.X(_3511_),
    .B(_2011_),
    .A(_1785_));
 sg13g2_and3_1 _7704_ (.X(_3512_),
    .A(_1793_),
    .B(_3510_),
    .C(_3511_));
 sg13g2_buf_1 _7705_ (.A(_3512_),
    .X(_3513_));
 sg13g2_buf_1 _7706_ (.A(_3513_),
    .X(_3514_));
 sg13g2_buf_2 _7707_ (.A(_3514_),
    .X(_3515_));
 sg13g2_buf_1 _7708_ (.A(_3515_),
    .X(_3516_));
 sg13g2_mux2_1 _7709_ (.A0(\board_state_next[0] ),
    .A1(_3509_),
    .S(net102),
    .X(_1121_));
 sg13g2_mux2_1 _7710_ (.A0(\board_state_next[100] ),
    .A1(\board_state_next[99] ),
    .S(net102),
    .X(_1122_));
 sg13g2_mux2_1 _7711_ (.A0(\board_state_next[101] ),
    .A1(\board_state_next[100] ),
    .S(_3516_),
    .X(_1123_));
 sg13g2_mux2_1 _7712_ (.A0(\board_state_next[102] ),
    .A1(\board_state_next[101] ),
    .S(_3516_),
    .X(_1124_));
 sg13g2_mux2_1 _7713_ (.A0(\board_state_next[103] ),
    .A1(\board_state_next[102] ),
    .S(net102),
    .X(_1125_));
 sg13g2_mux2_1 _7714_ (.A0(\board_state_next[104] ),
    .A1(\board_state_next[103] ),
    .S(net102),
    .X(_1126_));
 sg13g2_mux2_1 _7715_ (.A0(\board_state_next[105] ),
    .A1(\board_state_next[104] ),
    .S(net102),
    .X(_1127_));
 sg13g2_mux2_1 _7716_ (.A0(\board_state_next[106] ),
    .A1(\board_state_next[105] ),
    .S(net102),
    .X(_1128_));
 sg13g2_mux2_1 _7717_ (.A0(\board_state_next[107] ),
    .A1(\board_state_next[106] ),
    .S(net102),
    .X(_1129_));
 sg13g2_mux2_1 _7718_ (.A0(\board_state_next[108] ),
    .A1(\board_state_next[107] ),
    .S(net102),
    .X(_1130_));
 sg13g2_buf_1 _7719_ (.A(_3515_),
    .X(_3517_));
 sg13g2_mux2_1 _7720_ (.A0(\board_state_next[109] ),
    .A1(\board_state_next[108] ),
    .S(_3517_),
    .X(_1131_));
 sg13g2_mux2_1 _7721_ (.A0(\board_state_next[10] ),
    .A1(\board_state_next[9] ),
    .S(net101),
    .X(_1132_));
 sg13g2_mux2_1 _7722_ (.A0(\board_state_next[110] ),
    .A1(\board_state_next[109] ),
    .S(net101),
    .X(_1133_));
 sg13g2_mux2_1 _7723_ (.A0(\board_state_next[111] ),
    .A1(\board_state_next[110] ),
    .S(net101),
    .X(_1134_));
 sg13g2_mux2_1 _7724_ (.A0(\board_state_next[112] ),
    .A1(\board_state_next[111] ),
    .S(net101),
    .X(_1135_));
 sg13g2_mux2_1 _7725_ (.A0(\board_state_next[113] ),
    .A1(\board_state_next[112] ),
    .S(net101),
    .X(_1136_));
 sg13g2_mux2_1 _7726_ (.A0(\board_state_next[114] ),
    .A1(\board_state_next[113] ),
    .S(net101),
    .X(_1137_));
 sg13g2_mux2_1 _7727_ (.A0(\board_state_next[115] ),
    .A1(\board_state_next[114] ),
    .S(_3517_),
    .X(_1138_));
 sg13g2_mux2_1 _7728_ (.A0(\board_state_next[116] ),
    .A1(\board_state_next[115] ),
    .S(net101),
    .X(_1139_));
 sg13g2_mux2_1 _7729_ (.A0(\board_state_next[117] ),
    .A1(\board_state_next[116] ),
    .S(net101),
    .X(_1140_));
 sg13g2_buf_1 _7730_ (.A(_3515_),
    .X(_3518_));
 sg13g2_mux2_1 _7731_ (.A0(\board_state_next[118] ),
    .A1(\board_state_next[117] ),
    .S(_3518_),
    .X(_1141_));
 sg13g2_mux2_1 _7732_ (.A0(\board_state_next[119] ),
    .A1(\board_state_next[118] ),
    .S(net100),
    .X(_1142_));
 sg13g2_mux2_1 _7733_ (.A0(\board_state_next[11] ),
    .A1(\board_state_next[10] ),
    .S(_3518_),
    .X(_1143_));
 sg13g2_mux2_1 _7734_ (.A0(\board_state_next[120] ),
    .A1(\board_state_next[119] ),
    .S(net100),
    .X(_1144_));
 sg13g2_mux2_1 _7735_ (.A0(\board_state_next[121] ),
    .A1(\board_state_next[120] ),
    .S(net100),
    .X(_1145_));
 sg13g2_mux2_1 _7736_ (.A0(\board_state_next[122] ),
    .A1(\board_state_next[121] ),
    .S(net100),
    .X(_1146_));
 sg13g2_mux2_1 _7737_ (.A0(\board_state_next[123] ),
    .A1(\board_state_next[122] ),
    .S(net100),
    .X(_1147_));
 sg13g2_mux2_1 _7738_ (.A0(\board_state_next[124] ),
    .A1(\board_state_next[123] ),
    .S(net100),
    .X(_1148_));
 sg13g2_mux2_1 _7739_ (.A0(\board_state_next[125] ),
    .A1(\board_state_next[124] ),
    .S(net100),
    .X(_1149_));
 sg13g2_mux2_1 _7740_ (.A0(\board_state_next[126] ),
    .A1(\board_state_next[125] ),
    .S(net100),
    .X(_1150_));
 sg13g2_buf_1 _7741_ (.A(_3515_),
    .X(_3519_));
 sg13g2_mux2_1 _7742_ (.A0(\board_state_next[127] ),
    .A1(\board_state_next[126] ),
    .S(net99),
    .X(_1151_));
 sg13g2_mux2_1 _7743_ (.A0(\board_state_next[128] ),
    .A1(\board_state_next[127] ),
    .S(_3519_),
    .X(_1152_));
 sg13g2_mux2_1 _7744_ (.A0(\board_state_next[129] ),
    .A1(\board_state_next[128] ),
    .S(_3519_),
    .X(_1153_));
 sg13g2_mux2_1 _7745_ (.A0(\board_state_next[12] ),
    .A1(\board_state_next[11] ),
    .S(net99),
    .X(_1154_));
 sg13g2_mux2_1 _7746_ (.A0(\board_state_next[130] ),
    .A1(\board_state_next[129] ),
    .S(net99),
    .X(_1155_));
 sg13g2_mux2_1 _7747_ (.A0(\board_state_next[131] ),
    .A1(\board_state_next[130] ),
    .S(net99),
    .X(_1156_));
 sg13g2_mux2_1 _7748_ (.A0(\board_state_next[132] ),
    .A1(\board_state_next[131] ),
    .S(net99),
    .X(_1157_));
 sg13g2_mux2_1 _7749_ (.A0(\board_state_next[133] ),
    .A1(\board_state_next[132] ),
    .S(net99),
    .X(_1158_));
 sg13g2_mux2_1 _7750_ (.A0(\board_state_next[134] ),
    .A1(\board_state_next[133] ),
    .S(net99),
    .X(_1159_));
 sg13g2_mux2_1 _7751_ (.A0(\board_state_next[135] ),
    .A1(\board_state_next[134] ),
    .S(net99),
    .X(_1160_));
 sg13g2_buf_1 _7752_ (.A(_3515_),
    .X(_3520_));
 sg13g2_mux2_1 _7753_ (.A0(\board_state_next[136] ),
    .A1(\board_state_next[135] ),
    .S(net98),
    .X(_1161_));
 sg13g2_mux2_1 _7754_ (.A0(\board_state_next[137] ),
    .A1(\board_state_next[136] ),
    .S(net98),
    .X(_1162_));
 sg13g2_mux2_1 _7755_ (.A0(\board_state_next[138] ),
    .A1(\board_state_next[137] ),
    .S(net98),
    .X(_1163_));
 sg13g2_mux2_1 _7756_ (.A0(\board_state_next[139] ),
    .A1(\board_state_next[138] ),
    .S(net98),
    .X(_1164_));
 sg13g2_mux2_1 _7757_ (.A0(\board_state_next[13] ),
    .A1(\board_state_next[12] ),
    .S(_3520_),
    .X(_1165_));
 sg13g2_mux2_1 _7758_ (.A0(\board_state_next[140] ),
    .A1(\board_state_next[139] ),
    .S(net98),
    .X(_1166_));
 sg13g2_mux2_1 _7759_ (.A0(\board_state_next[141] ),
    .A1(\board_state_next[140] ),
    .S(net98),
    .X(_1167_));
 sg13g2_mux2_1 _7760_ (.A0(\board_state_next[142] ),
    .A1(\board_state_next[141] ),
    .S(net98),
    .X(_1168_));
 sg13g2_mux2_1 _7761_ (.A0(\board_state_next[143] ),
    .A1(\board_state_next[142] ),
    .S(net98),
    .X(_1169_));
 sg13g2_mux2_1 _7762_ (.A0(\board_state_next[144] ),
    .A1(\board_state_next[143] ),
    .S(_3520_),
    .X(_1170_));
 sg13g2_buf_1 _7763_ (.A(_3515_),
    .X(_3521_));
 sg13g2_mux2_1 _7764_ (.A0(\board_state_next[145] ),
    .A1(\board_state_next[144] ),
    .S(net97),
    .X(_1171_));
 sg13g2_mux2_1 _7765_ (.A0(\board_state_next[146] ),
    .A1(\board_state_next[145] ),
    .S(net97),
    .X(_1172_));
 sg13g2_mux2_1 _7766_ (.A0(\board_state_next[147] ),
    .A1(\board_state_next[146] ),
    .S(_3521_),
    .X(_1173_));
 sg13g2_mux2_1 _7767_ (.A0(\board_state_next[148] ),
    .A1(\board_state_next[147] ),
    .S(net97),
    .X(_1174_));
 sg13g2_mux2_1 _7768_ (.A0(\board_state_next[149] ),
    .A1(\board_state_next[148] ),
    .S(net97),
    .X(_1175_));
 sg13g2_mux2_1 _7769_ (.A0(\board_state_next[14] ),
    .A1(\board_state_next[13] ),
    .S(_3521_),
    .X(_1176_));
 sg13g2_mux2_1 _7770_ (.A0(\board_state_next[150] ),
    .A1(\board_state_next[149] ),
    .S(net97),
    .X(_1177_));
 sg13g2_mux2_1 _7771_ (.A0(\board_state_next[151] ),
    .A1(\board_state_next[150] ),
    .S(net97),
    .X(_1178_));
 sg13g2_mux2_1 _7772_ (.A0(\board_state_next[152] ),
    .A1(\board_state_next[151] ),
    .S(net97),
    .X(_1179_));
 sg13g2_mux2_1 _7773_ (.A0(\board_state_next[153] ),
    .A1(\board_state_next[152] ),
    .S(net97),
    .X(_1180_));
 sg13g2_buf_1 _7774_ (.A(_3514_),
    .X(_3522_));
 sg13g2_buf_1 _7775_ (.A(_3522_),
    .X(_3523_));
 sg13g2_mux2_1 _7776_ (.A0(\board_state_next[154] ),
    .A1(\board_state_next[153] ),
    .S(net96),
    .X(_1181_));
 sg13g2_mux2_1 _7777_ (.A0(\board_state_next[155] ),
    .A1(\board_state_next[154] ),
    .S(net96),
    .X(_1182_));
 sg13g2_mux2_1 _7778_ (.A0(\board_state_next[156] ),
    .A1(\board_state_next[155] ),
    .S(net96),
    .X(_1183_));
 sg13g2_mux2_1 _7779_ (.A0(\board_state_next[157] ),
    .A1(\board_state_next[156] ),
    .S(net96),
    .X(_1184_));
 sg13g2_mux2_1 _7780_ (.A0(\board_state_next[158] ),
    .A1(\board_state_next[157] ),
    .S(net96),
    .X(_1185_));
 sg13g2_mux2_1 _7781_ (.A0(\board_state_next[159] ),
    .A1(\board_state_next[158] ),
    .S(net96),
    .X(_1186_));
 sg13g2_mux2_1 _7782_ (.A0(\board_state_next[15] ),
    .A1(\board_state_next[14] ),
    .S(net96),
    .X(_1187_));
 sg13g2_mux2_1 _7783_ (.A0(\board_state_next[160] ),
    .A1(\board_state_next[159] ),
    .S(net96),
    .X(_1188_));
 sg13g2_mux2_1 _7784_ (.A0(\board_state_next[161] ),
    .A1(\board_state_next[160] ),
    .S(_3523_),
    .X(_1189_));
 sg13g2_mux2_1 _7785_ (.A0(\board_state_next[162] ),
    .A1(\board_state_next[161] ),
    .S(_3523_),
    .X(_1190_));
 sg13g2_buf_1 _7786_ (.A(_3522_),
    .X(_3524_));
 sg13g2_mux2_1 _7787_ (.A0(\board_state_next[163] ),
    .A1(\board_state_next[162] ),
    .S(net95),
    .X(_1191_));
 sg13g2_mux2_1 _7788_ (.A0(\board_state_next[164] ),
    .A1(\board_state_next[163] ),
    .S(net95),
    .X(_1192_));
 sg13g2_mux2_1 _7789_ (.A0(\board_state_next[165] ),
    .A1(\board_state_next[164] ),
    .S(net95),
    .X(_1193_));
 sg13g2_mux2_1 _7790_ (.A0(\board_state_next[166] ),
    .A1(\board_state_next[165] ),
    .S(net95),
    .X(_1194_));
 sg13g2_mux2_1 _7791_ (.A0(\board_state_next[167] ),
    .A1(\board_state_next[166] ),
    .S(net95),
    .X(_1195_));
 sg13g2_mux2_1 _7792_ (.A0(\board_state_next[168] ),
    .A1(\board_state_next[167] ),
    .S(net95),
    .X(_1196_));
 sg13g2_mux2_1 _7793_ (.A0(\board_state_next[169] ),
    .A1(\board_state_next[168] ),
    .S(net95),
    .X(_1197_));
 sg13g2_mux2_1 _7794_ (.A0(\board_state_next[16] ),
    .A1(\board_state_next[15] ),
    .S(_3524_),
    .X(_1198_));
 sg13g2_mux2_1 _7795_ (.A0(\board_state_next[170] ),
    .A1(\board_state_next[169] ),
    .S(net95),
    .X(_1199_));
 sg13g2_mux2_1 _7796_ (.A0(\board_state_next[171] ),
    .A1(\board_state_next[170] ),
    .S(_3524_),
    .X(_1200_));
 sg13g2_buf_1 _7797_ (.A(_3522_),
    .X(_3525_));
 sg13g2_mux2_1 _7798_ (.A0(\board_state_next[172] ),
    .A1(\board_state_next[171] ),
    .S(net94),
    .X(_1201_));
 sg13g2_mux2_1 _7799_ (.A0(\board_state_next[173] ),
    .A1(\board_state_next[172] ),
    .S(net94),
    .X(_1202_));
 sg13g2_mux2_1 _7800_ (.A0(\board_state_next[174] ),
    .A1(\board_state_next[173] ),
    .S(net94),
    .X(_1203_));
 sg13g2_mux2_1 _7801_ (.A0(\board_state_next[175] ),
    .A1(\board_state_next[174] ),
    .S(net94),
    .X(_1204_));
 sg13g2_mux2_1 _7802_ (.A0(\board_state_next[176] ),
    .A1(\board_state_next[175] ),
    .S(_3525_),
    .X(_1205_));
 sg13g2_mux2_1 _7803_ (.A0(\board_state_next[177] ),
    .A1(\board_state_next[176] ),
    .S(_3525_),
    .X(_1206_));
 sg13g2_mux2_1 _7804_ (.A0(\board_state_next[178] ),
    .A1(\board_state_next[177] ),
    .S(net94),
    .X(_1207_));
 sg13g2_mux2_1 _7805_ (.A0(\board_state_next[179] ),
    .A1(\board_state_next[178] ),
    .S(net94),
    .X(_1208_));
 sg13g2_mux2_1 _7806_ (.A0(\board_state_next[17] ),
    .A1(\board_state_next[16] ),
    .S(net94),
    .X(_1209_));
 sg13g2_mux2_1 _7807_ (.A0(\board_state_next[180] ),
    .A1(\board_state_next[179] ),
    .S(net94),
    .X(_1210_));
 sg13g2_buf_1 _7808_ (.A(_3522_),
    .X(_3526_));
 sg13g2_mux2_1 _7809_ (.A0(\board_state_next[181] ),
    .A1(\board_state_next[180] ),
    .S(_3526_),
    .X(_1211_));
 sg13g2_mux2_1 _7810_ (.A0(\board_state_next[182] ),
    .A1(\board_state_next[181] ),
    .S(net93),
    .X(_1212_));
 sg13g2_mux2_1 _7811_ (.A0(\board_state_next[183] ),
    .A1(\board_state_next[182] ),
    .S(net93),
    .X(_1213_));
 sg13g2_mux2_1 _7812_ (.A0(\board_state_next[184] ),
    .A1(\board_state_next[183] ),
    .S(net93),
    .X(_1214_));
 sg13g2_mux2_1 _7813_ (.A0(\board_state_next[185] ),
    .A1(\board_state_next[184] ),
    .S(net93),
    .X(_1215_));
 sg13g2_mux2_1 _7814_ (.A0(\board_state_next[186] ),
    .A1(\board_state_next[185] ),
    .S(net93),
    .X(_1216_));
 sg13g2_mux2_1 _7815_ (.A0(\board_state_next[187] ),
    .A1(\board_state_next[186] ),
    .S(net93),
    .X(_1217_));
 sg13g2_mux2_1 _7816_ (.A0(\board_state_next[188] ),
    .A1(\board_state_next[187] ),
    .S(net93),
    .X(_1218_));
 sg13g2_mux2_1 _7817_ (.A0(\board_state_next[189] ),
    .A1(\board_state_next[188] ),
    .S(net93),
    .X(_1219_));
 sg13g2_mux2_1 _7818_ (.A0(\board_state_next[18] ),
    .A1(\board_state_next[17] ),
    .S(_3526_),
    .X(_1220_));
 sg13g2_buf_1 _7819_ (.A(_3522_),
    .X(_3527_));
 sg13g2_mux2_1 _7820_ (.A0(\board_state_next[190] ),
    .A1(\board_state_next[189] ),
    .S(net92),
    .X(_1221_));
 sg13g2_mux2_1 _7821_ (.A0(\board_state_next[191] ),
    .A1(\board_state_next[190] ),
    .S(net92),
    .X(_1222_));
 sg13g2_mux2_1 _7822_ (.A0(\board_state_next[192] ),
    .A1(\board_state_next[191] ),
    .S(net92),
    .X(_1223_));
 sg13g2_mux2_1 _7823_ (.A0(\board_state_next[193] ),
    .A1(\board_state_next[192] ),
    .S(net92),
    .X(_1224_));
 sg13g2_mux2_1 _7824_ (.A0(\board_state_next[194] ),
    .A1(\board_state_next[193] ),
    .S(net92),
    .X(_1225_));
 sg13g2_mux2_1 _7825_ (.A0(\board_state_next[195] ),
    .A1(\board_state_next[194] ),
    .S(net92),
    .X(_1226_));
 sg13g2_mux2_1 _7826_ (.A0(\board_state_next[196] ),
    .A1(\board_state_next[195] ),
    .S(net92),
    .X(_1227_));
 sg13g2_mux2_1 _7827_ (.A0(\board_state_next[197] ),
    .A1(\board_state_next[196] ),
    .S(net92),
    .X(_1228_));
 sg13g2_mux2_1 _7828_ (.A0(\board_state_next[198] ),
    .A1(\board_state_next[197] ),
    .S(_3527_),
    .X(_1229_));
 sg13g2_mux2_1 _7829_ (.A0(\board_state_next[199] ),
    .A1(\board_state_next[198] ),
    .S(_3527_),
    .X(_1230_));
 sg13g2_buf_1 _7830_ (.A(_3522_),
    .X(_3528_));
 sg13g2_mux2_1 _7831_ (.A0(\board_state_next[19] ),
    .A1(\board_state_next[18] ),
    .S(net91),
    .X(_1231_));
 sg13g2_mux2_1 _7832_ (.A0(\board_state_next[1] ),
    .A1(\board_state_next[0] ),
    .S(net91),
    .X(_1232_));
 sg13g2_mux2_1 _7833_ (.A0(\board_state_next[200] ),
    .A1(\board_state_next[199] ),
    .S(net91),
    .X(_1233_));
 sg13g2_mux2_1 _7834_ (.A0(\board_state_next[201] ),
    .A1(\board_state_next[200] ),
    .S(net91),
    .X(_1234_));
 sg13g2_mux2_1 _7835_ (.A0(\board_state_next[202] ),
    .A1(\board_state_next[201] ),
    .S(net91),
    .X(_1235_));
 sg13g2_mux2_1 _7836_ (.A0(\board_state_next[203] ),
    .A1(\board_state_next[202] ),
    .S(net91),
    .X(_1236_));
 sg13g2_mux2_1 _7837_ (.A0(\board_state_next[204] ),
    .A1(\board_state_next[203] ),
    .S(net91),
    .X(_1237_));
 sg13g2_mux2_1 _7838_ (.A0(\board_state_next[205] ),
    .A1(\board_state_next[204] ),
    .S(_3528_),
    .X(_1238_));
 sg13g2_mux2_1 _7839_ (.A0(\board_state_next[206] ),
    .A1(\board_state_next[205] ),
    .S(_3528_),
    .X(_1239_));
 sg13g2_mux2_1 _7840_ (.A0(\board_state_next[207] ),
    .A1(\board_state_next[206] ),
    .S(net91),
    .X(_1240_));
 sg13g2_buf_1 _7841_ (.A(_3522_),
    .X(_3529_));
 sg13g2_mux2_1 _7842_ (.A0(\board_state_next[208] ),
    .A1(\board_state_next[207] ),
    .S(net90),
    .X(_1241_));
 sg13g2_mux2_1 _7843_ (.A0(\board_state_next[209] ),
    .A1(\board_state_next[208] ),
    .S(net90),
    .X(_1242_));
 sg13g2_mux2_1 _7844_ (.A0(\board_state_next[20] ),
    .A1(\board_state_next[19] ),
    .S(net90),
    .X(_1243_));
 sg13g2_mux2_1 _7845_ (.A0(\board_state_next[210] ),
    .A1(\board_state_next[209] ),
    .S(net90),
    .X(_1244_));
 sg13g2_mux2_1 _7846_ (.A0(\board_state_next[211] ),
    .A1(\board_state_next[210] ),
    .S(_3529_),
    .X(_1245_));
 sg13g2_mux2_1 _7847_ (.A0(\board_state_next[212] ),
    .A1(\board_state_next[211] ),
    .S(_3529_),
    .X(_1246_));
 sg13g2_mux2_1 _7848_ (.A0(\board_state_next[213] ),
    .A1(\board_state_next[212] ),
    .S(net90),
    .X(_1247_));
 sg13g2_mux2_1 _7849_ (.A0(\board_state_next[214] ),
    .A1(\board_state_next[213] ),
    .S(net90),
    .X(_1248_));
 sg13g2_mux2_1 _7850_ (.A0(\board_state_next[215] ),
    .A1(\board_state_next[214] ),
    .S(net90),
    .X(_1249_));
 sg13g2_mux2_1 _7851_ (.A0(\board_state_next[216] ),
    .A1(\board_state_next[215] ),
    .S(net90),
    .X(_1250_));
 sg13g2_buf_1 _7852_ (.A(_3514_),
    .X(_3530_));
 sg13g2_buf_1 _7853_ (.A(_3530_),
    .X(_3531_));
 sg13g2_mux2_1 _7854_ (.A0(\board_state_next[217] ),
    .A1(\board_state_next[216] ),
    .S(net89),
    .X(_1251_));
 sg13g2_mux2_1 _7855_ (.A0(\board_state_next[218] ),
    .A1(\board_state_next[217] ),
    .S(_3531_),
    .X(_1252_));
 sg13g2_mux2_1 _7856_ (.A0(\board_state_next[219] ),
    .A1(\board_state_next[218] ),
    .S(net89),
    .X(_1253_));
 sg13g2_mux2_1 _7857_ (.A0(\board_state_next[21] ),
    .A1(\board_state_next[20] ),
    .S(_3531_),
    .X(_1254_));
 sg13g2_mux2_1 _7858_ (.A0(\board_state_next[220] ),
    .A1(\board_state_next[219] ),
    .S(net89),
    .X(_1255_));
 sg13g2_mux2_1 _7859_ (.A0(\board_state_next[221] ),
    .A1(\board_state_next[220] ),
    .S(net89),
    .X(_1256_));
 sg13g2_mux2_1 _7860_ (.A0(\board_state_next[222] ),
    .A1(\board_state_next[221] ),
    .S(net89),
    .X(_1257_));
 sg13g2_mux2_1 _7861_ (.A0(\board_state_next[223] ),
    .A1(\board_state_next[222] ),
    .S(net89),
    .X(_1258_));
 sg13g2_mux2_1 _7862_ (.A0(\board_state_next[224] ),
    .A1(\board_state_next[223] ),
    .S(net89),
    .X(_1259_));
 sg13g2_mux2_1 _7863_ (.A0(\board_state_next[225] ),
    .A1(\board_state_next[224] ),
    .S(net89),
    .X(_1260_));
 sg13g2_buf_1 _7864_ (.A(_3530_),
    .X(_3532_));
 sg13g2_mux2_1 _7865_ (.A0(\board_state_next[226] ),
    .A1(\board_state_next[225] ),
    .S(net88),
    .X(_1261_));
 sg13g2_mux2_1 _7866_ (.A0(\board_state_next[227] ),
    .A1(\board_state_next[226] ),
    .S(net88),
    .X(_1262_));
 sg13g2_mux2_1 _7867_ (.A0(\board_state_next[228] ),
    .A1(\board_state_next[227] ),
    .S(net88),
    .X(_1263_));
 sg13g2_mux2_1 _7868_ (.A0(\board_state_next[229] ),
    .A1(\board_state_next[228] ),
    .S(net88),
    .X(_1264_));
 sg13g2_mux2_1 _7869_ (.A0(\board_state_next[22] ),
    .A1(\board_state_next[21] ),
    .S(net88),
    .X(_1265_));
 sg13g2_mux2_1 _7870_ (.A0(\board_state_next[230] ),
    .A1(\board_state_next[229] ),
    .S(_3532_),
    .X(_1266_));
 sg13g2_mux2_1 _7871_ (.A0(\board_state_next[231] ),
    .A1(\board_state_next[230] ),
    .S(net88),
    .X(_1267_));
 sg13g2_mux2_1 _7872_ (.A0(\board_state_next[232] ),
    .A1(\board_state_next[231] ),
    .S(_3532_),
    .X(_1268_));
 sg13g2_mux2_1 _7873_ (.A0(\board_state_next[233] ),
    .A1(\board_state_next[232] ),
    .S(net88),
    .X(_1269_));
 sg13g2_mux2_1 _7874_ (.A0(\board_state_next[234] ),
    .A1(\board_state_next[233] ),
    .S(net88),
    .X(_1270_));
 sg13g2_buf_1 _7875_ (.A(_3530_),
    .X(_3533_));
 sg13g2_mux2_1 _7876_ (.A0(\board_state_next[235] ),
    .A1(\board_state_next[234] ),
    .S(net87),
    .X(_1271_));
 sg13g2_mux2_1 _7877_ (.A0(\board_state_next[236] ),
    .A1(\board_state_next[235] ),
    .S(net87),
    .X(_1272_));
 sg13g2_mux2_1 _7878_ (.A0(\board_state_next[237] ),
    .A1(\board_state_next[236] ),
    .S(net87),
    .X(_1273_));
 sg13g2_mux2_1 _7879_ (.A0(\board_state_next[238] ),
    .A1(\board_state_next[237] ),
    .S(_3533_),
    .X(_1274_));
 sg13g2_mux2_1 _7880_ (.A0(\board_state_next[239] ),
    .A1(\board_state_next[238] ),
    .S(net87),
    .X(_1275_));
 sg13g2_mux2_1 _7881_ (.A0(\board_state_next[23] ),
    .A1(\board_state_next[22] ),
    .S(net87),
    .X(_1276_));
 sg13g2_mux2_1 _7882_ (.A0(\board_state_next[240] ),
    .A1(\board_state_next[239] ),
    .S(net87),
    .X(_1277_));
 sg13g2_mux2_1 _7883_ (.A0(\board_state_next[241] ),
    .A1(\board_state_next[240] ),
    .S(net87),
    .X(_1278_));
 sg13g2_mux2_1 _7884_ (.A0(\board_state_next[242] ),
    .A1(\board_state_next[241] ),
    .S(_3533_),
    .X(_1279_));
 sg13g2_mux2_1 _7885_ (.A0(\board_state_next[243] ),
    .A1(\board_state_next[242] ),
    .S(net87),
    .X(_1280_));
 sg13g2_buf_1 _7886_ (.A(_3530_),
    .X(_3534_));
 sg13g2_mux2_1 _7887_ (.A0(\board_state_next[244] ),
    .A1(\board_state_next[243] ),
    .S(net86),
    .X(_1281_));
 sg13g2_mux2_1 _7888_ (.A0(\board_state_next[245] ),
    .A1(\board_state_next[244] ),
    .S(net86),
    .X(_1282_));
 sg13g2_mux2_1 _7889_ (.A0(\board_state_next[246] ),
    .A1(\board_state_next[245] ),
    .S(_3534_),
    .X(_1283_));
 sg13g2_mux2_1 _7890_ (.A0(\board_state_next[247] ),
    .A1(\board_state_next[246] ),
    .S(_3534_),
    .X(_1284_));
 sg13g2_mux2_1 _7891_ (.A0(\board_state_next[248] ),
    .A1(\board_state_next[247] ),
    .S(net86),
    .X(_1285_));
 sg13g2_mux2_1 _7892_ (.A0(\board_state_next[249] ),
    .A1(\board_state_next[248] ),
    .S(net86),
    .X(_1286_));
 sg13g2_mux2_1 _7893_ (.A0(\board_state_next[24] ),
    .A1(\board_state_next[23] ),
    .S(net86),
    .X(_1287_));
 sg13g2_mux2_1 _7894_ (.A0(\board_state_next[250] ),
    .A1(\board_state_next[249] ),
    .S(net86),
    .X(_1288_));
 sg13g2_mux2_1 _7895_ (.A0(\board_state_next[251] ),
    .A1(\board_state_next[250] ),
    .S(net86),
    .X(_1289_));
 sg13g2_mux2_1 _7896_ (.A0(\board_state_next[252] ),
    .A1(\board_state_next[251] ),
    .S(net86),
    .X(_1290_));
 sg13g2_buf_1 _7897_ (.A(_3530_),
    .X(_3535_));
 sg13g2_mux2_1 _7898_ (.A0(\board_state_next[253] ),
    .A1(\board_state_next[252] ),
    .S(net85),
    .X(_1291_));
 sg13g2_mux2_1 _7899_ (.A0(\board_state_next[254] ),
    .A1(\board_state_next[253] ),
    .S(net85),
    .X(_1292_));
 sg13g2_mux2_1 _7900_ (.A0(\board_state_next[255] ),
    .A1(\board_state_next[254] ),
    .S(net85),
    .X(_1293_));
 sg13g2_mux2_1 _7901_ (.A0(\board_state_next[256] ),
    .A1(\board_state_next[255] ),
    .S(net85),
    .X(_1294_));
 sg13g2_mux2_1 _7902_ (.A0(\board_state_next[257] ),
    .A1(\board_state_next[256] ),
    .S(net85),
    .X(_1295_));
 sg13g2_mux2_1 _7903_ (.A0(\board_state_next[258] ),
    .A1(\board_state_next[257] ),
    .S(_3535_),
    .X(_1296_));
 sg13g2_mux2_1 _7904_ (.A0(\board_state_next[259] ),
    .A1(\board_state_next[258] ),
    .S(_3535_),
    .X(_1297_));
 sg13g2_mux2_1 _7905_ (.A0(\board_state_next[25] ),
    .A1(\board_state_next[24] ),
    .S(net85),
    .X(_1298_));
 sg13g2_mux2_1 _7906_ (.A0(\board_state_next[260] ),
    .A1(\board_state_next[259] ),
    .S(net85),
    .X(_1299_));
 sg13g2_mux2_1 _7907_ (.A0(\board_state_next[261] ),
    .A1(\board_state_next[260] ),
    .S(net85),
    .X(_1300_));
 sg13g2_buf_1 _7908_ (.A(_3530_),
    .X(_3536_));
 sg13g2_mux2_1 _7909_ (.A0(\board_state_next[262] ),
    .A1(\board_state_next[261] ),
    .S(net84),
    .X(_1301_));
 sg13g2_mux2_1 _7910_ (.A0(\board_state_next[263] ),
    .A1(\board_state_next[262] ),
    .S(net84),
    .X(_1302_));
 sg13g2_mux2_1 _7911_ (.A0(\board_state_next[264] ),
    .A1(\board_state_next[263] ),
    .S(net84),
    .X(_1303_));
 sg13g2_mux2_1 _7912_ (.A0(\board_state_next[265] ),
    .A1(\board_state_next[264] ),
    .S(_3536_),
    .X(_1304_));
 sg13g2_mux2_1 _7913_ (.A0(\board_state_next[266] ),
    .A1(\board_state_next[265] ),
    .S(_3536_),
    .X(_1305_));
 sg13g2_mux2_1 _7914_ (.A0(\board_state_next[267] ),
    .A1(\board_state_next[266] ),
    .S(net84),
    .X(_1306_));
 sg13g2_mux2_1 _7915_ (.A0(\board_state_next[268] ),
    .A1(\board_state_next[267] ),
    .S(net84),
    .X(_1307_));
 sg13g2_mux2_1 _7916_ (.A0(\board_state_next[269] ),
    .A1(\board_state_next[268] ),
    .S(net84),
    .X(_1308_));
 sg13g2_mux2_1 _7917_ (.A0(\board_state_next[26] ),
    .A1(\board_state_next[25] ),
    .S(net84),
    .X(_1309_));
 sg13g2_mux2_1 _7918_ (.A0(\board_state_next[270] ),
    .A1(\board_state_next[269] ),
    .S(net84),
    .X(_1310_));
 sg13g2_buf_1 _7919_ (.A(_3530_),
    .X(_3537_));
 sg13g2_mux2_1 _7920_ (.A0(\board_state_next[271] ),
    .A1(\board_state_next[270] ),
    .S(net83),
    .X(_1311_));
 sg13g2_mux2_1 _7921_ (.A0(\board_state_next[272] ),
    .A1(\board_state_next[271] ),
    .S(_3537_),
    .X(_1312_));
 sg13g2_mux2_1 _7922_ (.A0(\board_state_next[273] ),
    .A1(\board_state_next[272] ),
    .S(net83),
    .X(_1313_));
 sg13g2_mux2_1 _7923_ (.A0(\board_state_next[274] ),
    .A1(\board_state_next[273] ),
    .S(net83),
    .X(_1314_));
 sg13g2_mux2_1 _7924_ (.A0(\board_state_next[275] ),
    .A1(\board_state_next[274] ),
    .S(net83),
    .X(_1315_));
 sg13g2_mux2_1 _7925_ (.A0(\board_state_next[276] ),
    .A1(\board_state_next[275] ),
    .S(net83),
    .X(_1316_));
 sg13g2_mux2_1 _7926_ (.A0(\board_state_next[277] ),
    .A1(\board_state_next[276] ),
    .S(net83),
    .X(_1317_));
 sg13g2_mux2_1 _7927_ (.A0(\board_state_next[278] ),
    .A1(\board_state_next[277] ),
    .S(net83),
    .X(_1318_));
 sg13g2_mux2_1 _7928_ (.A0(\board_state_next[279] ),
    .A1(\board_state_next[278] ),
    .S(_3537_),
    .X(_1319_));
 sg13g2_mux2_1 _7929_ (.A0(\board_state_next[27] ),
    .A1(\board_state_next[26] ),
    .S(net83),
    .X(_1320_));
 sg13g2_buf_1 _7930_ (.A(_3514_),
    .X(_3538_));
 sg13g2_buf_1 _7931_ (.A(_3538_),
    .X(_3539_));
 sg13g2_mux2_1 _7932_ (.A0(\board_state_next[280] ),
    .A1(\board_state_next[279] ),
    .S(net82),
    .X(_1321_));
 sg13g2_mux2_1 _7933_ (.A0(\board_state_next[281] ),
    .A1(\board_state_next[280] ),
    .S(net82),
    .X(_1322_));
 sg13g2_mux2_1 _7934_ (.A0(\board_state_next[282] ),
    .A1(\board_state_next[281] ),
    .S(net82),
    .X(_1323_));
 sg13g2_mux2_1 _7935_ (.A0(\board_state_next[283] ),
    .A1(\board_state_next[282] ),
    .S(net82),
    .X(_1324_));
 sg13g2_mux2_1 _7936_ (.A0(\board_state_next[284] ),
    .A1(\board_state_next[283] ),
    .S(net82),
    .X(_1325_));
 sg13g2_mux2_1 _7937_ (.A0(\board_state_next[285] ),
    .A1(\board_state_next[284] ),
    .S(net82),
    .X(_1326_));
 sg13g2_mux2_1 _7938_ (.A0(\board_state_next[286] ),
    .A1(\board_state_next[285] ),
    .S(net82),
    .X(_1327_));
 sg13g2_mux2_1 _7939_ (.A0(\board_state_next[287] ),
    .A1(\board_state_next[286] ),
    .S(_3539_),
    .X(_1328_));
 sg13g2_mux2_1 _7940_ (.A0(\board_state_next[288] ),
    .A1(\board_state_next[287] ),
    .S(net82),
    .X(_1329_));
 sg13g2_mux2_1 _7941_ (.A0(\board_state_next[289] ),
    .A1(\board_state_next[288] ),
    .S(_3539_),
    .X(_1330_));
 sg13g2_buf_1 _7942_ (.A(_3538_),
    .X(_3540_));
 sg13g2_mux2_1 _7943_ (.A0(\board_state_next[28] ),
    .A1(\board_state_next[27] ),
    .S(net81),
    .X(_1331_));
 sg13g2_mux2_1 _7944_ (.A0(\board_state_next[290] ),
    .A1(\board_state_next[289] ),
    .S(net81),
    .X(_1332_));
 sg13g2_mux2_1 _7945_ (.A0(\board_state_next[291] ),
    .A1(\board_state_next[290] ),
    .S(net81),
    .X(_1333_));
 sg13g2_mux2_1 _7946_ (.A0(\board_state_next[292] ),
    .A1(\board_state_next[291] ),
    .S(_3540_),
    .X(_1334_));
 sg13g2_mux2_1 _7947_ (.A0(\board_state_next[293] ),
    .A1(\board_state_next[292] ),
    .S(_3540_),
    .X(_1335_));
 sg13g2_mux2_1 _7948_ (.A0(\board_state_next[294] ),
    .A1(\board_state_next[293] ),
    .S(net81),
    .X(_1336_));
 sg13g2_mux2_1 _7949_ (.A0(\board_state_next[295] ),
    .A1(\board_state_next[294] ),
    .S(net81),
    .X(_1337_));
 sg13g2_mux2_1 _7950_ (.A0(\board_state_next[296] ),
    .A1(\board_state_next[295] ),
    .S(net81),
    .X(_1338_));
 sg13g2_mux2_1 _7951_ (.A0(\board_state_next[297] ),
    .A1(\board_state_next[296] ),
    .S(net81),
    .X(_1339_));
 sg13g2_mux2_1 _7952_ (.A0(\board_state_next[298] ),
    .A1(\board_state_next[297] ),
    .S(net81),
    .X(_1340_));
 sg13g2_buf_1 _7953_ (.A(_3538_),
    .X(_3541_));
 sg13g2_mux2_1 _7954_ (.A0(\board_state_next[299] ),
    .A1(\board_state_next[298] ),
    .S(net80),
    .X(_1341_));
 sg13g2_mux2_1 _7955_ (.A0(\board_state_next[29] ),
    .A1(\board_state_next[28] ),
    .S(_3541_),
    .X(_1342_));
 sg13g2_mux2_1 _7956_ (.A0(\board_state_next[2] ),
    .A1(\board_state_next[1] ),
    .S(net80),
    .X(_1343_));
 sg13g2_mux2_1 _7957_ (.A0(\board_state_next[300] ),
    .A1(\board_state_next[299] ),
    .S(net80),
    .X(_1344_));
 sg13g2_mux2_1 _7958_ (.A0(\board_state_next[301] ),
    .A1(\board_state_next[300] ),
    .S(_3541_),
    .X(_1345_));
 sg13g2_mux2_1 _7959_ (.A0(\board_state_next[302] ),
    .A1(\board_state_next[301] ),
    .S(net80),
    .X(_1346_));
 sg13g2_mux2_1 _7960_ (.A0(\board_state_next[303] ),
    .A1(\board_state_next[302] ),
    .S(net80),
    .X(_1347_));
 sg13g2_mux2_1 _7961_ (.A0(\board_state_next[304] ),
    .A1(\board_state_next[303] ),
    .S(net80),
    .X(_1348_));
 sg13g2_mux2_1 _7962_ (.A0(\board_state_next[305] ),
    .A1(\board_state_next[304] ),
    .S(net80),
    .X(_1349_));
 sg13g2_mux2_1 _7963_ (.A0(\board_state_next[306] ),
    .A1(\board_state_next[305] ),
    .S(net80),
    .X(_1350_));
 sg13g2_buf_1 _7964_ (.A(_3538_),
    .X(_3542_));
 sg13g2_mux2_1 _7965_ (.A0(\board_state_next[307] ),
    .A1(\board_state_next[306] ),
    .S(net79),
    .X(_1351_));
 sg13g2_mux2_1 _7966_ (.A0(\board_state_next[308] ),
    .A1(\board_state_next[307] ),
    .S(net79),
    .X(_1352_));
 sg13g2_mux2_1 _7967_ (.A0(\board_state_next[309] ),
    .A1(\board_state_next[308] ),
    .S(net79),
    .X(_1353_));
 sg13g2_mux2_1 _7968_ (.A0(\board_state_next[30] ),
    .A1(\board_state_next[29] ),
    .S(net79),
    .X(_1354_));
 sg13g2_mux2_1 _7969_ (.A0(\board_state_next[310] ),
    .A1(\board_state_next[309] ),
    .S(net79),
    .X(_1355_));
 sg13g2_mux2_1 _7970_ (.A0(\board_state_next[311] ),
    .A1(\board_state_next[310] ),
    .S(net79),
    .X(_1356_));
 sg13g2_mux2_1 _7971_ (.A0(\board_state_next[312] ),
    .A1(\board_state_next[311] ),
    .S(net79),
    .X(_1357_));
 sg13g2_mux2_1 _7972_ (.A0(\board_state_next[313] ),
    .A1(\board_state_next[312] ),
    .S(net79),
    .X(_1358_));
 sg13g2_mux2_1 _7973_ (.A0(\board_state_next[314] ),
    .A1(\board_state_next[313] ),
    .S(_3542_),
    .X(_1359_));
 sg13g2_mux2_1 _7974_ (.A0(\board_state_next[315] ),
    .A1(\board_state_next[314] ),
    .S(_3542_),
    .X(_1360_));
 sg13g2_buf_1 _7975_ (.A(_3538_),
    .X(_3543_));
 sg13g2_mux2_1 _7976_ (.A0(\board_state_next[316] ),
    .A1(\board_state_next[315] ),
    .S(net78),
    .X(_1361_));
 sg13g2_mux2_1 _7977_ (.A0(\board_state_next[317] ),
    .A1(\board_state_next[316] ),
    .S(net78),
    .X(_1362_));
 sg13g2_mux2_1 _7978_ (.A0(\board_state_next[318] ),
    .A1(\board_state_next[317] ),
    .S(_3543_),
    .X(_1363_));
 sg13g2_mux2_1 _7979_ (.A0(\board_state_next[319] ),
    .A1(\board_state_next[318] ),
    .S(_3543_),
    .X(_1364_));
 sg13g2_mux2_1 _7980_ (.A0(\board_state_next[31] ),
    .A1(\board_state_next[30] ),
    .S(net78),
    .X(_1365_));
 sg13g2_mux2_1 _7981_ (.A0(\board_state_next[320] ),
    .A1(\board_state_next[319] ),
    .S(net78),
    .X(_1366_));
 sg13g2_mux2_1 _7982_ (.A0(\board_state_next[321] ),
    .A1(\board_state_next[320] ),
    .S(net78),
    .X(_1367_));
 sg13g2_mux2_1 _7983_ (.A0(\board_state_next[322] ),
    .A1(\board_state_next[321] ),
    .S(net78),
    .X(_1368_));
 sg13g2_mux2_1 _7984_ (.A0(\board_state_next[323] ),
    .A1(\board_state_next[322] ),
    .S(net78),
    .X(_1369_));
 sg13g2_mux2_1 _7985_ (.A0(\board_state_next[324] ),
    .A1(\board_state_next[323] ),
    .S(net78),
    .X(_1370_));
 sg13g2_buf_1 _7986_ (.A(_3538_),
    .X(_3544_));
 sg13g2_mux2_1 _7987_ (.A0(\board_state_next[325] ),
    .A1(\board_state_next[324] ),
    .S(net77),
    .X(_1371_));
 sg13g2_mux2_1 _7988_ (.A0(\board_state_next[326] ),
    .A1(\board_state_next[325] ),
    .S(net77),
    .X(_1372_));
 sg13g2_mux2_1 _7989_ (.A0(\board_state_next[327] ),
    .A1(\board_state_next[326] ),
    .S(net77),
    .X(_1373_));
 sg13g2_mux2_1 _7990_ (.A0(\board_state_next[328] ),
    .A1(\board_state_next[327] ),
    .S(_3544_),
    .X(_1374_));
 sg13g2_mux2_1 _7991_ (.A0(\board_state_next[329] ),
    .A1(\board_state_next[328] ),
    .S(net77),
    .X(_1375_));
 sg13g2_mux2_1 _7992_ (.A0(\board_state_next[32] ),
    .A1(\board_state_next[31] ),
    .S(net77),
    .X(_1376_));
 sg13g2_mux2_1 _7993_ (.A0(\board_state_next[330] ),
    .A1(\board_state_next[329] ),
    .S(net77),
    .X(_1377_));
 sg13g2_mux2_1 _7994_ (.A0(\board_state_next[331] ),
    .A1(\board_state_next[330] ),
    .S(net77),
    .X(_1378_));
 sg13g2_mux2_1 _7995_ (.A0(\board_state_next[332] ),
    .A1(\board_state_next[331] ),
    .S(net77),
    .X(_1379_));
 sg13g2_mux2_1 _7996_ (.A0(\board_state_next[333] ),
    .A1(\board_state_next[332] ),
    .S(_3544_),
    .X(_1380_));
 sg13g2_buf_1 _7997_ (.A(_3538_),
    .X(_3545_));
 sg13g2_mux2_1 _7998_ (.A0(\board_state_next[334] ),
    .A1(\board_state_next[333] ),
    .S(net76),
    .X(_1381_));
 sg13g2_mux2_1 _7999_ (.A0(\board_state_next[335] ),
    .A1(\board_state_next[334] ),
    .S(net76),
    .X(_1382_));
 sg13g2_mux2_1 _8000_ (.A0(\board_state_next[336] ),
    .A1(\board_state_next[335] ),
    .S(_3545_),
    .X(_1383_));
 sg13g2_mux2_1 _8001_ (.A0(\board_state_next[337] ),
    .A1(\board_state_next[336] ),
    .S(_3545_),
    .X(_1384_));
 sg13g2_mux2_1 _8002_ (.A0(\board_state_next[338] ),
    .A1(\board_state_next[337] ),
    .S(net76),
    .X(_1385_));
 sg13g2_mux2_1 _8003_ (.A0(\board_state_next[339] ),
    .A1(\board_state_next[338] ),
    .S(net76),
    .X(_1386_));
 sg13g2_mux2_1 _8004_ (.A0(\board_state_next[33] ),
    .A1(\board_state_next[32] ),
    .S(net76),
    .X(_1387_));
 sg13g2_mux2_1 _8005_ (.A0(\board_state_next[340] ),
    .A1(\board_state_next[339] ),
    .S(net76),
    .X(_1388_));
 sg13g2_mux2_1 _8006_ (.A0(\board_state_next[341] ),
    .A1(\board_state_next[340] ),
    .S(net76),
    .X(_1389_));
 sg13g2_mux2_1 _8007_ (.A0(\board_state_next[342] ),
    .A1(\board_state_next[341] ),
    .S(net76),
    .X(_1390_));
 sg13g2_buf_1 _8008_ (.A(_3513_),
    .X(_3546_));
 sg13g2_buf_1 _8009_ (.A(_3546_),
    .X(_3547_));
 sg13g2_mux2_1 _8010_ (.A0(\board_state_next[343] ),
    .A1(\board_state_next[342] ),
    .S(net137),
    .X(_1391_));
 sg13g2_mux2_1 _8011_ (.A0(\board_state_next[344] ),
    .A1(\board_state_next[343] ),
    .S(net137),
    .X(_1392_));
 sg13g2_mux2_1 _8012_ (.A0(\board_state_next[345] ),
    .A1(\board_state_next[344] ),
    .S(net137),
    .X(_1393_));
 sg13g2_mux2_1 _8013_ (.A0(\board_state_next[346] ),
    .A1(\board_state_next[345] ),
    .S(net137),
    .X(_1394_));
 sg13g2_mux2_1 _8014_ (.A0(\board_state_next[347] ),
    .A1(\board_state_next[346] ),
    .S(net137),
    .X(_1395_));
 sg13g2_mux2_1 _8015_ (.A0(\board_state_next[348] ),
    .A1(\board_state_next[347] ),
    .S(net137),
    .X(_1396_));
 sg13g2_mux2_1 _8016_ (.A0(\board_state_next[349] ),
    .A1(\board_state_next[348] ),
    .S(net137),
    .X(_1397_));
 sg13g2_mux2_1 _8017_ (.A0(\board_state_next[34] ),
    .A1(\board_state_next[33] ),
    .S(net137),
    .X(_1398_));
 sg13g2_mux2_1 _8018_ (.A0(\board_state_next[350] ),
    .A1(\board_state_next[349] ),
    .S(_3547_),
    .X(_1399_));
 sg13g2_mux2_1 _8019_ (.A0(\board_state_next[351] ),
    .A1(\board_state_next[350] ),
    .S(_3547_),
    .X(_1400_));
 sg13g2_buf_1 _8020_ (.A(_3546_),
    .X(_3548_));
 sg13g2_mux2_1 _8021_ (.A0(\board_state_next[352] ),
    .A1(\board_state_next[351] ),
    .S(net136),
    .X(_1401_));
 sg13g2_mux2_1 _8022_ (.A0(\board_state_next[353] ),
    .A1(\board_state_next[352] ),
    .S(net136),
    .X(_1402_));
 sg13g2_mux2_1 _8023_ (.A0(\board_state_next[354] ),
    .A1(\board_state_next[353] ),
    .S(net136),
    .X(_1403_));
 sg13g2_mux2_1 _8024_ (.A0(\board_state_next[355] ),
    .A1(\board_state_next[354] ),
    .S(net136),
    .X(_1404_));
 sg13g2_mux2_1 _8025_ (.A0(\board_state_next[356] ),
    .A1(\board_state_next[355] ),
    .S(_3548_),
    .X(_1405_));
 sg13g2_mux2_1 _8026_ (.A0(\board_state_next[357] ),
    .A1(\board_state_next[356] ),
    .S(net136),
    .X(_1406_));
 sg13g2_mux2_1 _8027_ (.A0(\board_state_next[358] ),
    .A1(\board_state_next[357] ),
    .S(net136),
    .X(_1407_));
 sg13g2_mux2_1 _8028_ (.A0(\board_state_next[359] ),
    .A1(\board_state_next[358] ),
    .S(_3548_),
    .X(_1408_));
 sg13g2_mux2_1 _8029_ (.A0(\board_state_next[35] ),
    .A1(\board_state_next[34] ),
    .S(net136),
    .X(_1409_));
 sg13g2_mux2_1 _8030_ (.A0(\board_state_next[360] ),
    .A1(\board_state_next[359] ),
    .S(net136),
    .X(_1410_));
 sg13g2_buf_1 _8031_ (.A(_3546_),
    .X(_3549_));
 sg13g2_mux2_1 _8032_ (.A0(\board_state_next[361] ),
    .A1(\board_state_next[360] ),
    .S(net135),
    .X(_1411_));
 sg13g2_mux2_1 _8033_ (.A0(\board_state_next[362] ),
    .A1(\board_state_next[361] ),
    .S(_3549_),
    .X(_1412_));
 sg13g2_mux2_1 _8034_ (.A0(\board_state_next[363] ),
    .A1(\board_state_next[362] ),
    .S(net135),
    .X(_1413_));
 sg13g2_mux2_1 _8035_ (.A0(\board_state_next[364] ),
    .A1(\board_state_next[363] ),
    .S(net135),
    .X(_1414_));
 sg13g2_mux2_1 _8036_ (.A0(\board_state_next[365] ),
    .A1(\board_state_next[364] ),
    .S(net135),
    .X(_1415_));
 sg13g2_mux2_1 _8037_ (.A0(\board_state_next[366] ),
    .A1(\board_state_next[365] ),
    .S(net135),
    .X(_1416_));
 sg13g2_mux2_1 _8038_ (.A0(\board_state_next[367] ),
    .A1(\board_state_next[366] ),
    .S(net135),
    .X(_1417_));
 sg13g2_mux2_1 _8039_ (.A0(\board_state_next[368] ),
    .A1(\board_state_next[367] ),
    .S(net135),
    .X(_1418_));
 sg13g2_mux2_1 _8040_ (.A0(\board_state_next[369] ),
    .A1(\board_state_next[368] ),
    .S(_3549_),
    .X(_1419_));
 sg13g2_mux2_1 _8041_ (.A0(\board_state_next[36] ),
    .A1(\board_state_next[35] ),
    .S(net135),
    .X(_1420_));
 sg13g2_buf_1 _8042_ (.A(_3546_),
    .X(_3550_));
 sg13g2_mux2_1 _8043_ (.A0(\board_state_next[370] ),
    .A1(\board_state_next[369] ),
    .S(_3550_),
    .X(_1421_));
 sg13g2_mux2_1 _8044_ (.A0(\board_state_next[371] ),
    .A1(\board_state_next[370] ),
    .S(net134),
    .X(_1422_));
 sg13g2_mux2_1 _8045_ (.A0(\board_state_next[372] ),
    .A1(\board_state_next[371] ),
    .S(_3550_),
    .X(_1423_));
 sg13g2_mux2_1 _8046_ (.A0(\board_state_next[373] ),
    .A1(\board_state_next[372] ),
    .S(net134),
    .X(_1424_));
 sg13g2_mux2_1 _8047_ (.A0(\board_state_next[374] ),
    .A1(\board_state_next[373] ),
    .S(net134),
    .X(_1425_));
 sg13g2_mux2_1 _8048_ (.A0(\board_state_next[375] ),
    .A1(\board_state_next[374] ),
    .S(net134),
    .X(_1426_));
 sg13g2_mux2_1 _8049_ (.A0(\board_state_next[376] ),
    .A1(\board_state_next[375] ),
    .S(net134),
    .X(_1427_));
 sg13g2_mux2_1 _8050_ (.A0(\board_state_next[377] ),
    .A1(\board_state_next[376] ),
    .S(net134),
    .X(_1428_));
 sg13g2_mux2_1 _8051_ (.A0(\board_state_next[378] ),
    .A1(\board_state_next[377] ),
    .S(net134),
    .X(_1429_));
 sg13g2_mux2_1 _8052_ (.A0(\board_state_next[379] ),
    .A1(\board_state_next[378] ),
    .S(net134),
    .X(_1430_));
 sg13g2_buf_1 _8053_ (.A(_3546_),
    .X(_3551_));
 sg13g2_mux2_1 _8054_ (.A0(\board_state_next[37] ),
    .A1(\board_state_next[36] ),
    .S(net133),
    .X(_1431_));
 sg13g2_mux2_1 _8055_ (.A0(\board_state_next[380] ),
    .A1(\board_state_next[379] ),
    .S(net133),
    .X(_1432_));
 sg13g2_mux2_1 _8056_ (.A0(\board_state_next[381] ),
    .A1(\board_state_next[380] ),
    .S(net133),
    .X(_1433_));
 sg13g2_mux2_1 _8057_ (.A0(\board_state_next[382] ),
    .A1(\board_state_next[381] ),
    .S(net133),
    .X(_1434_));
 sg13g2_mux2_1 _8058_ (.A0(\board_state_next[383] ),
    .A1(\board_state_next[382] ),
    .S(_3551_),
    .X(_1435_));
 sg13g2_mux2_1 _8059_ (.A0(\board_state_next[384] ),
    .A1(\board_state_next[383] ),
    .S(net133),
    .X(_1436_));
 sg13g2_mux2_1 _8060_ (.A0(\board_state_next[385] ),
    .A1(\board_state_next[384] ),
    .S(_3551_),
    .X(_1437_));
 sg13g2_mux2_1 _8061_ (.A0(\board_state_next[386] ),
    .A1(\board_state_next[385] ),
    .S(net133),
    .X(_1438_));
 sg13g2_mux2_1 _8062_ (.A0(\board_state_next[387] ),
    .A1(\board_state_next[386] ),
    .S(net133),
    .X(_1439_));
 sg13g2_mux2_1 _8063_ (.A0(\board_state_next[388] ),
    .A1(\board_state_next[387] ),
    .S(net133),
    .X(_1440_));
 sg13g2_buf_1 _8064_ (.A(_3546_),
    .X(_3552_));
 sg13g2_mux2_1 _8065_ (.A0(\board_state_next[389] ),
    .A1(\board_state_next[388] ),
    .S(net132),
    .X(_1441_));
 sg13g2_mux2_1 _8066_ (.A0(\board_state_next[38] ),
    .A1(\board_state_next[37] ),
    .S(net132),
    .X(_1442_));
 sg13g2_mux2_1 _8067_ (.A0(\board_state_next[390] ),
    .A1(\board_state_next[389] ),
    .S(_3552_),
    .X(_1443_));
 sg13g2_mux2_1 _8068_ (.A0(\board_state_next[391] ),
    .A1(\board_state_next[390] ),
    .S(_3552_),
    .X(_1444_));
 sg13g2_mux2_1 _8069_ (.A0(\board_state_next[392] ),
    .A1(\board_state_next[391] ),
    .S(net132),
    .X(_1445_));
 sg13g2_mux2_1 _8070_ (.A0(\board_state_next[393] ),
    .A1(\board_state_next[392] ),
    .S(net132),
    .X(_1446_));
 sg13g2_mux2_1 _8071_ (.A0(\board_state_next[394] ),
    .A1(\board_state_next[393] ),
    .S(net132),
    .X(_1447_));
 sg13g2_mux2_1 _8072_ (.A0(\board_state_next[395] ),
    .A1(\board_state_next[394] ),
    .S(net132),
    .X(_1448_));
 sg13g2_mux2_1 _8073_ (.A0(\board_state_next[396] ),
    .A1(\board_state_next[395] ),
    .S(net132),
    .X(_1449_));
 sg13g2_mux2_1 _8074_ (.A0(\board_state_next[397] ),
    .A1(\board_state_next[396] ),
    .S(net132),
    .X(_1450_));
 sg13g2_buf_1 _8075_ (.A(_3546_),
    .X(_3553_));
 sg13g2_mux2_1 _8076_ (.A0(\board_state_next[398] ),
    .A1(\board_state_next[397] ),
    .S(net131),
    .X(_1451_));
 sg13g2_mux2_1 _8077_ (.A0(\board_state_next[399] ),
    .A1(\board_state_next[398] ),
    .S(net131),
    .X(_1452_));
 sg13g2_mux2_1 _8078_ (.A0(\board_state_next[39] ),
    .A1(\board_state_next[38] ),
    .S(_3553_),
    .X(_1453_));
 sg13g2_mux2_1 _8079_ (.A0(\board_state_next[3] ),
    .A1(\board_state_next[2] ),
    .S(net131),
    .X(_1454_));
 sg13g2_mux2_1 _8080_ (.A0(\board_state_next[400] ),
    .A1(\board_state_next[399] ),
    .S(net131),
    .X(_1455_));
 sg13g2_mux2_1 _8081_ (.A0(\board_state_next[401] ),
    .A1(\board_state_next[400] ),
    .S(net131),
    .X(_1456_));
 sg13g2_mux2_1 _8082_ (.A0(\board_state_next[402] ),
    .A1(\board_state_next[401] ),
    .S(net131),
    .X(_1457_));
 sg13g2_mux2_1 _8083_ (.A0(\board_state_next[403] ),
    .A1(\board_state_next[402] ),
    .S(net131),
    .X(_1458_));
 sg13g2_mux2_1 _8084_ (.A0(\board_state_next[404] ),
    .A1(\board_state_next[403] ),
    .S(net131),
    .X(_1459_));
 sg13g2_mux2_1 _8085_ (.A0(\board_state_next[405] ),
    .A1(\board_state_next[404] ),
    .S(_3553_),
    .X(_1460_));
 sg13g2_buf_1 _8086_ (.A(_3513_),
    .X(_3554_));
 sg13g2_buf_1 _8087_ (.A(_3554_),
    .X(_3555_));
 sg13g2_mux2_1 _8088_ (.A0(\board_state_next[406] ),
    .A1(\board_state_next[405] ),
    .S(net130),
    .X(_1461_));
 sg13g2_mux2_1 _8089_ (.A0(\board_state_next[407] ),
    .A1(\board_state_next[406] ),
    .S(net130),
    .X(_1462_));
 sg13g2_mux2_1 _8090_ (.A0(\board_state_next[408] ),
    .A1(\board_state_next[407] ),
    .S(net130),
    .X(_1463_));
 sg13g2_mux2_1 _8091_ (.A0(\board_state_next[409] ),
    .A1(\board_state_next[408] ),
    .S(net130),
    .X(_1464_));
 sg13g2_mux2_1 _8092_ (.A0(\board_state_next[40] ),
    .A1(\board_state_next[39] ),
    .S(net130),
    .X(_1465_));
 sg13g2_mux2_1 _8093_ (.A0(\board_state_next[410] ),
    .A1(\board_state_next[409] ),
    .S(net130),
    .X(_1466_));
 sg13g2_mux2_1 _8094_ (.A0(\board_state_next[411] ),
    .A1(\board_state_next[410] ),
    .S(net130),
    .X(_1467_));
 sg13g2_mux2_1 _8095_ (.A0(\board_state_next[412] ),
    .A1(\board_state_next[411] ),
    .S(net130),
    .X(_1468_));
 sg13g2_mux2_1 _8096_ (.A0(\board_state_next[413] ),
    .A1(\board_state_next[412] ),
    .S(_3555_),
    .X(_1469_));
 sg13g2_mux2_1 _8097_ (.A0(\board_state_next[414] ),
    .A1(\board_state_next[413] ),
    .S(_3555_),
    .X(_1470_));
 sg13g2_buf_1 _8098_ (.A(_3554_),
    .X(_3556_));
 sg13g2_mux2_1 _8099_ (.A0(\board_state_next[415] ),
    .A1(\board_state_next[414] ),
    .S(net129),
    .X(_1471_));
 sg13g2_mux2_1 _8100_ (.A0(\board_state_next[416] ),
    .A1(\board_state_next[415] ),
    .S(net129),
    .X(_1472_));
 sg13g2_mux2_1 _8101_ (.A0(\board_state_next[417] ),
    .A1(\board_state_next[416] ),
    .S(net129),
    .X(_1473_));
 sg13g2_mux2_1 _8102_ (.A0(\board_state_next[418] ),
    .A1(\board_state_next[417] ),
    .S(net129),
    .X(_1474_));
 sg13g2_mux2_1 _8103_ (.A0(\board_state_next[419] ),
    .A1(\board_state_next[418] ),
    .S(net129),
    .X(_1475_));
 sg13g2_mux2_1 _8104_ (.A0(\board_state_next[41] ),
    .A1(\board_state_next[40] ),
    .S(net129),
    .X(_1476_));
 sg13g2_mux2_1 _8105_ (.A0(\board_state_next[420] ),
    .A1(\board_state_next[419] ),
    .S(net129),
    .X(_1477_));
 sg13g2_mux2_1 _8106_ (.A0(\board_state_next[421] ),
    .A1(\board_state_next[420] ),
    .S(net129),
    .X(_1478_));
 sg13g2_mux2_1 _8107_ (.A0(\board_state_next[422] ),
    .A1(\board_state_next[421] ),
    .S(_3556_),
    .X(_1479_));
 sg13g2_mux2_1 _8108_ (.A0(\board_state_next[423] ),
    .A1(\board_state_next[422] ),
    .S(_3556_),
    .X(_1480_));
 sg13g2_buf_1 _8109_ (.A(_3554_),
    .X(_3557_));
 sg13g2_mux2_1 _8110_ (.A0(\board_state_next[424] ),
    .A1(\board_state_next[423] ),
    .S(net128),
    .X(_1481_));
 sg13g2_mux2_1 _8111_ (.A0(\board_state_next[425] ),
    .A1(\board_state_next[424] ),
    .S(_3557_),
    .X(_1482_));
 sg13g2_mux2_1 _8112_ (.A0(\board_state_next[426] ),
    .A1(\board_state_next[425] ),
    .S(net128),
    .X(_1483_));
 sg13g2_mux2_1 _8113_ (.A0(\board_state_next[427] ),
    .A1(\board_state_next[426] ),
    .S(net128),
    .X(_1484_));
 sg13g2_mux2_1 _8114_ (.A0(\board_state_next[428] ),
    .A1(\board_state_next[427] ),
    .S(net128),
    .X(_1485_));
 sg13g2_mux2_1 _8115_ (.A0(\board_state_next[429] ),
    .A1(\board_state_next[428] ),
    .S(net128),
    .X(_1486_));
 sg13g2_mux2_1 _8116_ (.A0(\board_state_next[42] ),
    .A1(\board_state_next[41] ),
    .S(_3557_),
    .X(_1487_));
 sg13g2_mux2_1 _8117_ (.A0(\board_state_next[430] ),
    .A1(\board_state_next[429] ),
    .S(net128),
    .X(_1488_));
 sg13g2_mux2_1 _8118_ (.A0(\board_state_next[431] ),
    .A1(\board_state_next[430] ),
    .S(net128),
    .X(_1489_));
 sg13g2_mux2_1 _8119_ (.A0(\board_state_next[432] ),
    .A1(\board_state_next[431] ),
    .S(net128),
    .X(_1490_));
 sg13g2_buf_1 _8120_ (.A(_3554_),
    .X(_3558_));
 sg13g2_mux2_1 _8121_ (.A0(\board_state_next[433] ),
    .A1(\board_state_next[432] ),
    .S(net127),
    .X(_1491_));
 sg13g2_mux2_1 _8122_ (.A0(\board_state_next[434] ),
    .A1(\board_state_next[433] ),
    .S(net127),
    .X(_1492_));
 sg13g2_mux2_1 _8123_ (.A0(\board_state_next[435] ),
    .A1(\board_state_next[434] ),
    .S(_3558_),
    .X(_1493_));
 sg13g2_mux2_1 _8124_ (.A0(\board_state_next[436] ),
    .A1(\board_state_next[435] ),
    .S(net127),
    .X(_1494_));
 sg13g2_mux2_1 _8125_ (.A0(\board_state_next[437] ),
    .A1(\board_state_next[436] ),
    .S(net127),
    .X(_1495_));
 sg13g2_mux2_1 _8126_ (.A0(\board_state_next[438] ),
    .A1(\board_state_next[437] ),
    .S(net127),
    .X(_1496_));
 sg13g2_mux2_1 _8127_ (.A0(\board_state_next[439] ),
    .A1(\board_state_next[438] ),
    .S(net127),
    .X(_1497_));
 sg13g2_mux2_1 _8128_ (.A0(\board_state_next[43] ),
    .A1(\board_state_next[42] ),
    .S(_3558_),
    .X(_1498_));
 sg13g2_mux2_1 _8129_ (.A0(\board_state_next[440] ),
    .A1(\board_state_next[439] ),
    .S(net127),
    .X(_1499_));
 sg13g2_mux2_1 _8130_ (.A0(\board_state_next[441] ),
    .A1(\board_state_next[440] ),
    .S(net127),
    .X(_1500_));
 sg13g2_buf_1 _8131_ (.A(_3554_),
    .X(_3559_));
 sg13g2_mux2_1 _8132_ (.A0(\board_state_next[442] ),
    .A1(\board_state_next[441] ),
    .S(_3559_),
    .X(_1501_));
 sg13g2_mux2_1 _8133_ (.A0(\board_state_next[443] ),
    .A1(\board_state_next[442] ),
    .S(net126),
    .X(_1502_));
 sg13g2_mux2_1 _8134_ (.A0(\board_state_next[444] ),
    .A1(\board_state_next[443] ),
    .S(net126),
    .X(_1503_));
 sg13g2_mux2_1 _8135_ (.A0(\board_state_next[445] ),
    .A1(\board_state_next[444] ),
    .S(net126),
    .X(_1504_));
 sg13g2_mux2_1 _8136_ (.A0(\board_state_next[446] ),
    .A1(\board_state_next[445] ),
    .S(net126),
    .X(_1505_));
 sg13g2_mux2_1 _8137_ (.A0(\board_state_next[447] ),
    .A1(\board_state_next[446] ),
    .S(net126),
    .X(_1506_));
 sg13g2_mux2_1 _8138_ (.A0(\board_state_next[448] ),
    .A1(\board_state_next[447] ),
    .S(net126),
    .X(_1507_));
 sg13g2_mux2_1 _8139_ (.A0(\board_state_next[449] ),
    .A1(\board_state_next[448] ),
    .S(net126),
    .X(_1508_));
 sg13g2_mux2_1 _8140_ (.A0(\board_state_next[44] ),
    .A1(\board_state_next[43] ),
    .S(_3559_),
    .X(_1509_));
 sg13g2_mux2_1 _8141_ (.A0(\board_state_next[450] ),
    .A1(\board_state_next[449] ),
    .S(net126),
    .X(_1510_));
 sg13g2_buf_1 _8142_ (.A(_3554_),
    .X(_3560_));
 sg13g2_mux2_1 _8143_ (.A0(\board_state_next[451] ),
    .A1(\board_state_next[450] ),
    .S(net125),
    .X(_1511_));
 sg13g2_mux2_1 _8144_ (.A0(\board_state_next[452] ),
    .A1(\board_state_next[451] ),
    .S(net125),
    .X(_1512_));
 sg13g2_mux2_1 _8145_ (.A0(\board_state_next[453] ),
    .A1(\board_state_next[452] ),
    .S(net125),
    .X(_1513_));
 sg13g2_mux2_1 _8146_ (.A0(\board_state_next[454] ),
    .A1(\board_state_next[453] ),
    .S(net125),
    .X(_1514_));
 sg13g2_mux2_1 _8147_ (.A0(\board_state_next[455] ),
    .A1(\board_state_next[454] ),
    .S(_3560_),
    .X(_1515_));
 sg13g2_mux2_1 _8148_ (.A0(\board_state_next[456] ),
    .A1(\board_state_next[455] ),
    .S(_3560_),
    .X(_1516_));
 sg13g2_mux2_1 _8149_ (.A0(\board_state_next[457] ),
    .A1(\board_state_next[456] ),
    .S(net125),
    .X(_1517_));
 sg13g2_mux2_1 _8150_ (.A0(\board_state_next[458] ),
    .A1(\board_state_next[457] ),
    .S(net125),
    .X(_1518_));
 sg13g2_mux2_1 _8151_ (.A0(\board_state_next[459] ),
    .A1(\board_state_next[458] ),
    .S(net125),
    .X(_1519_));
 sg13g2_mux2_1 _8152_ (.A0(\board_state_next[45] ),
    .A1(\board_state_next[44] ),
    .S(net125),
    .X(_1520_));
 sg13g2_buf_1 _8153_ (.A(_3554_),
    .X(_3561_));
 sg13g2_mux2_1 _8154_ (.A0(\board_state_next[460] ),
    .A1(\board_state_next[459] ),
    .S(net124),
    .X(_1521_));
 sg13g2_mux2_1 _8155_ (.A0(\board_state_next[461] ),
    .A1(\board_state_next[460] ),
    .S(net124),
    .X(_1522_));
 sg13g2_mux2_1 _8156_ (.A0(\board_state_next[462] ),
    .A1(\board_state_next[461] ),
    .S(_3561_),
    .X(_1523_));
 sg13g2_mux2_1 _8157_ (.A0(\board_state_next[463] ),
    .A1(\board_state_next[462] ),
    .S(net124),
    .X(_1524_));
 sg13g2_mux2_1 _8158_ (.A0(\board_state_next[464] ),
    .A1(\board_state_next[463] ),
    .S(_3561_),
    .X(_1525_));
 sg13g2_mux2_1 _8159_ (.A0(\board_state_next[465] ),
    .A1(\board_state_next[464] ),
    .S(net124),
    .X(_1526_));
 sg13g2_mux2_1 _8160_ (.A0(\board_state_next[466] ),
    .A1(\board_state_next[465] ),
    .S(net124),
    .X(_1527_));
 sg13g2_mux2_1 _8161_ (.A0(\board_state_next[467] ),
    .A1(\board_state_next[466] ),
    .S(net124),
    .X(_1528_));
 sg13g2_mux2_1 _8162_ (.A0(\board_state_next[468] ),
    .A1(\board_state_next[467] ),
    .S(net124),
    .X(_1529_));
 sg13g2_mux2_1 _8163_ (.A0(\board_state_next[469] ),
    .A1(\board_state_next[468] ),
    .S(net124),
    .X(_1530_));
 sg13g2_buf_1 _8164_ (.A(_3513_),
    .X(_3562_));
 sg13g2_buf_1 _8165_ (.A(_3562_),
    .X(_3563_));
 sg13g2_mux2_1 _8166_ (.A0(\board_state_next[46] ),
    .A1(\board_state_next[45] ),
    .S(net123),
    .X(_1531_));
 sg13g2_mux2_1 _8167_ (.A0(\board_state_next[470] ),
    .A1(\board_state_next[469] ),
    .S(net123),
    .X(_1532_));
 sg13g2_mux2_1 _8168_ (.A0(\board_state_next[471] ),
    .A1(\board_state_next[470] ),
    .S(net123),
    .X(_1533_));
 sg13g2_mux2_1 _8169_ (.A0(\board_state_next[472] ),
    .A1(\board_state_next[471] ),
    .S(net123),
    .X(_1534_));
 sg13g2_mux2_1 _8170_ (.A0(\board_state_next[473] ),
    .A1(\board_state_next[472] ),
    .S(_3563_),
    .X(_1535_));
 sg13g2_mux2_1 _8171_ (.A0(\board_state_next[474] ),
    .A1(\board_state_next[473] ),
    .S(net123),
    .X(_1536_));
 sg13g2_mux2_1 _8172_ (.A0(\board_state_next[475] ),
    .A1(\board_state_next[474] ),
    .S(_3563_),
    .X(_1537_));
 sg13g2_mux2_1 _8173_ (.A0(\board_state_next[476] ),
    .A1(\board_state_next[475] ),
    .S(net123),
    .X(_1538_));
 sg13g2_mux2_1 _8174_ (.A0(\board_state_next[477] ),
    .A1(\board_state_next[476] ),
    .S(net123),
    .X(_1539_));
 sg13g2_mux2_1 _8175_ (.A0(\board_state_next[478] ),
    .A1(\board_state_next[477] ),
    .S(net123),
    .X(_1540_));
 sg13g2_buf_1 _8176_ (.A(_3562_),
    .X(_3564_));
 sg13g2_mux2_1 _8177_ (.A0(\board_state_next[479] ),
    .A1(\board_state_next[478] ),
    .S(net122),
    .X(_1541_));
 sg13g2_mux2_1 _8178_ (.A0(\board_state_next[47] ),
    .A1(\board_state_next[46] ),
    .S(_3564_),
    .X(_1542_));
 sg13g2_mux2_1 _8179_ (.A0(\board_state_next[480] ),
    .A1(\board_state_next[479] ),
    .S(_3564_),
    .X(_1543_));
 sg13g2_mux2_1 _8180_ (.A0(\board_state_next[481] ),
    .A1(\board_state_next[480] ),
    .S(net122),
    .X(_1544_));
 sg13g2_mux2_1 _8181_ (.A0(\board_state_next[482] ),
    .A1(\board_state_next[481] ),
    .S(net122),
    .X(_1545_));
 sg13g2_mux2_1 _8182_ (.A0(\board_state_next[483] ),
    .A1(\board_state_next[482] ),
    .S(net122),
    .X(_1546_));
 sg13g2_mux2_1 _8183_ (.A0(\board_state_next[484] ),
    .A1(\board_state_next[483] ),
    .S(net122),
    .X(_1547_));
 sg13g2_mux2_1 _8184_ (.A0(\board_state_next[485] ),
    .A1(\board_state_next[484] ),
    .S(net122),
    .X(_1548_));
 sg13g2_mux2_1 _8185_ (.A0(\board_state_next[486] ),
    .A1(\board_state_next[485] ),
    .S(net122),
    .X(_1549_));
 sg13g2_mux2_1 _8186_ (.A0(\board_state_next[487] ),
    .A1(\board_state_next[486] ),
    .S(net122),
    .X(_1550_));
 sg13g2_buf_1 _8187_ (.A(_3562_),
    .X(_3565_));
 sg13g2_mux2_1 _8188_ (.A0(\board_state_next[488] ),
    .A1(\board_state_next[487] ),
    .S(net121),
    .X(_1551_));
 sg13g2_mux2_1 _8189_ (.A0(\board_state_next[489] ),
    .A1(\board_state_next[488] ),
    .S(net121),
    .X(_1552_));
 sg13g2_mux2_1 _8190_ (.A0(\board_state_next[48] ),
    .A1(\board_state_next[47] ),
    .S(net121),
    .X(_1553_));
 sg13g2_mux2_1 _8191_ (.A0(\board_state_next[490] ),
    .A1(\board_state_next[489] ),
    .S(net121),
    .X(_1554_));
 sg13g2_mux2_1 _8192_ (.A0(\board_state_next[491] ),
    .A1(\board_state_next[490] ),
    .S(net121),
    .X(_1555_));
 sg13g2_mux2_1 _8193_ (.A0(\board_state_next[492] ),
    .A1(\board_state_next[491] ),
    .S(_3565_),
    .X(_1556_));
 sg13g2_mux2_1 _8194_ (.A0(\board_state_next[493] ),
    .A1(\board_state_next[492] ),
    .S(_3565_),
    .X(_1557_));
 sg13g2_mux2_1 _8195_ (.A0(\board_state_next[494] ),
    .A1(\board_state_next[493] ),
    .S(net121),
    .X(_1558_));
 sg13g2_mux2_1 _8196_ (.A0(\board_state_next[495] ),
    .A1(\board_state_next[494] ),
    .S(net121),
    .X(_1559_));
 sg13g2_mux2_1 _8197_ (.A0(\board_state_next[496] ),
    .A1(\board_state_next[495] ),
    .S(net121),
    .X(_1560_));
 sg13g2_buf_1 _8198_ (.A(_3562_),
    .X(_3566_));
 sg13g2_mux2_1 _8199_ (.A0(\board_state_next[497] ),
    .A1(\board_state_next[496] ),
    .S(net120),
    .X(_1561_));
 sg13g2_mux2_1 _8200_ (.A0(\board_state_next[498] ),
    .A1(\board_state_next[497] ),
    .S(net120),
    .X(_1562_));
 sg13g2_mux2_1 _8201_ (.A0(\board_state_next[499] ),
    .A1(\board_state_next[498] ),
    .S(net120),
    .X(_1563_));
 sg13g2_mux2_1 _8202_ (.A0(\board_state_next[49] ),
    .A1(\board_state_next[48] ),
    .S(net120),
    .X(_1564_));
 sg13g2_mux2_1 _8203_ (.A0(\board_state_next[4] ),
    .A1(\board_state_next[3] ),
    .S(net120),
    .X(_1565_));
 sg13g2_mux2_1 _8204_ (.A0(\board_state_next[500] ),
    .A1(\board_state_next[499] ),
    .S(net120),
    .X(_1566_));
 sg13g2_mux2_1 _8205_ (.A0(\board_state_next[501] ),
    .A1(\board_state_next[500] ),
    .S(net120),
    .X(_1567_));
 sg13g2_mux2_1 _8206_ (.A0(\board_state_next[502] ),
    .A1(\board_state_next[501] ),
    .S(_3566_),
    .X(_1568_));
 sg13g2_mux2_1 _8207_ (.A0(\board_state_next[503] ),
    .A1(\board_state_next[502] ),
    .S(net120),
    .X(_1569_));
 sg13g2_mux2_1 _8208_ (.A0(\board_state_next[504] ),
    .A1(\board_state_next[503] ),
    .S(_3566_),
    .X(_1570_));
 sg13g2_buf_1 _8209_ (.A(_3562_),
    .X(_3567_));
 sg13g2_mux2_1 _8210_ (.A0(\board_state_next[505] ),
    .A1(\board_state_next[504] ),
    .S(net119),
    .X(_1571_));
 sg13g2_mux2_1 _8211_ (.A0(\board_state_next[506] ),
    .A1(\board_state_next[505] ),
    .S(net119),
    .X(_1572_));
 sg13g2_mux2_1 _8212_ (.A0(\board_state_next[507] ),
    .A1(\board_state_next[506] ),
    .S(net119),
    .X(_1573_));
 sg13g2_mux2_1 _8213_ (.A0(\board_state_next[508] ),
    .A1(\board_state_next[507] ),
    .S(net119),
    .X(_1574_));
 sg13g2_mux2_1 _8214_ (.A0(\board_state_next[509] ),
    .A1(\board_state_next[508] ),
    .S(net119),
    .X(_1575_));
 sg13g2_mux2_1 _8215_ (.A0(\board_state_next[50] ),
    .A1(\board_state_next[49] ),
    .S(_3567_),
    .X(_1576_));
 sg13g2_mux2_1 _8216_ (.A0(\board_state_next[510] ),
    .A1(\board_state_next[509] ),
    .S(net119),
    .X(_1577_));
 sg13g2_mux2_1 _8217_ (.A0(\board_state_next[511] ),
    .A1(\board_state_next[510] ),
    .S(net119),
    .X(_1578_));
 sg13g2_mux2_1 _8218_ (.A0(\board_state_next[51] ),
    .A1(\board_state_next[50] ),
    .S(_3567_),
    .X(_1579_));
 sg13g2_mux2_1 _8219_ (.A0(\board_state_next[52] ),
    .A1(\board_state_next[51] ),
    .S(net119),
    .X(_1580_));
 sg13g2_buf_1 _8220_ (.A(_3562_),
    .X(_3568_));
 sg13g2_mux2_1 _8221_ (.A0(\board_state_next[53] ),
    .A1(\board_state_next[52] ),
    .S(net118),
    .X(_1581_));
 sg13g2_mux2_1 _8222_ (.A0(\board_state_next[54] ),
    .A1(\board_state_next[53] ),
    .S(net118),
    .X(_1582_));
 sg13g2_mux2_1 _8223_ (.A0(\board_state_next[55] ),
    .A1(\board_state_next[54] ),
    .S(net118),
    .X(_1583_));
 sg13g2_mux2_1 _8224_ (.A0(\board_state_next[56] ),
    .A1(\board_state_next[55] ),
    .S(net118),
    .X(_1584_));
 sg13g2_mux2_1 _8225_ (.A0(\board_state_next[57] ),
    .A1(\board_state_next[56] ),
    .S(net118),
    .X(_1585_));
 sg13g2_mux2_1 _8226_ (.A0(\board_state_next[58] ),
    .A1(\board_state_next[57] ),
    .S(net118),
    .X(_1586_));
 sg13g2_mux2_1 _8227_ (.A0(\board_state_next[59] ),
    .A1(\board_state_next[58] ),
    .S(_3568_),
    .X(_1587_));
 sg13g2_mux2_1 _8228_ (.A0(\board_state_next[5] ),
    .A1(\board_state_next[4] ),
    .S(_3568_),
    .X(_1588_));
 sg13g2_mux2_1 _8229_ (.A0(\board_state_next[60] ),
    .A1(\board_state_next[59] ),
    .S(net118),
    .X(_1589_));
 sg13g2_mux2_1 _8230_ (.A0(\board_state_next[61] ),
    .A1(\board_state_next[60] ),
    .S(net118),
    .X(_1590_));
 sg13g2_buf_1 _8231_ (.A(_3562_),
    .X(_3569_));
 sg13g2_mux2_1 _8232_ (.A0(\board_state_next[62] ),
    .A1(\board_state_next[61] ),
    .S(net117),
    .X(_1591_));
 sg13g2_mux2_1 _8233_ (.A0(\board_state_next[63] ),
    .A1(\board_state_next[62] ),
    .S(net117),
    .X(_1592_));
 sg13g2_mux2_1 _8234_ (.A0(\board_state_next[64] ),
    .A1(\board_state_next[63] ),
    .S(net117),
    .X(_1593_));
 sg13g2_mux2_1 _8235_ (.A0(\board_state_next[65] ),
    .A1(\board_state_next[64] ),
    .S(_3569_),
    .X(_1594_));
 sg13g2_mux2_1 _8236_ (.A0(\board_state_next[66] ),
    .A1(\board_state_next[65] ),
    .S(_3569_),
    .X(_1595_));
 sg13g2_mux2_1 _8237_ (.A0(\board_state_next[67] ),
    .A1(\board_state_next[66] ),
    .S(net117),
    .X(_1596_));
 sg13g2_mux2_1 _8238_ (.A0(\board_state_next[68] ),
    .A1(\board_state_next[67] ),
    .S(net117),
    .X(_1597_));
 sg13g2_mux2_1 _8239_ (.A0(\board_state_next[69] ),
    .A1(\board_state_next[68] ),
    .S(net117),
    .X(_1598_));
 sg13g2_mux2_1 _8240_ (.A0(\board_state_next[6] ),
    .A1(\board_state_next[5] ),
    .S(net117),
    .X(_1599_));
 sg13g2_mux2_1 _8241_ (.A0(\board_state_next[70] ),
    .A1(\board_state_next[69] ),
    .S(net117),
    .X(_1600_));
 sg13g2_buf_1 _8242_ (.A(_3514_),
    .X(_3570_));
 sg13g2_mux2_1 _8243_ (.A0(\board_state_next[71] ),
    .A1(\board_state_next[70] ),
    .S(net116),
    .X(_1601_));
 sg13g2_mux2_1 _8244_ (.A0(\board_state_next[72] ),
    .A1(\board_state_next[71] ),
    .S(net116),
    .X(_1602_));
 sg13g2_mux2_1 _8245_ (.A0(\board_state_next[73] ),
    .A1(\board_state_next[72] ),
    .S(net116),
    .X(_1603_));
 sg13g2_mux2_1 _8246_ (.A0(\board_state_next[74] ),
    .A1(\board_state_next[73] ),
    .S(_3570_),
    .X(_1604_));
 sg13g2_mux2_1 _8247_ (.A0(\board_state_next[75] ),
    .A1(\board_state_next[74] ),
    .S(_3570_),
    .X(_1605_));
 sg13g2_mux2_1 _8248_ (.A0(\board_state_next[76] ),
    .A1(\board_state_next[75] ),
    .S(net116),
    .X(_1606_));
 sg13g2_mux2_1 _8249_ (.A0(\board_state_next[77] ),
    .A1(\board_state_next[76] ),
    .S(net116),
    .X(_1607_));
 sg13g2_mux2_1 _8250_ (.A0(\board_state_next[78] ),
    .A1(\board_state_next[77] ),
    .S(net116),
    .X(_1608_));
 sg13g2_mux2_1 _8251_ (.A0(\board_state_next[79] ),
    .A1(\board_state_next[78] ),
    .S(net116),
    .X(_1609_));
 sg13g2_mux2_1 _8252_ (.A0(\board_state_next[7] ),
    .A1(\board_state_next[6] ),
    .S(net116),
    .X(_1610_));
 sg13g2_buf_1 _8253_ (.A(_3514_),
    .X(_3571_));
 sg13g2_mux2_1 _8254_ (.A0(\board_state_next[80] ),
    .A1(\board_state_next[79] ),
    .S(_3571_),
    .X(_1611_));
 sg13g2_mux2_1 _8255_ (.A0(\board_state_next[81] ),
    .A1(\board_state_next[80] ),
    .S(net115),
    .X(_1612_));
 sg13g2_mux2_1 _8256_ (.A0(\board_state_next[82] ),
    .A1(\board_state_next[81] ),
    .S(_3571_),
    .X(_1613_));
 sg13g2_mux2_1 _8257_ (.A0(\board_state_next[83] ),
    .A1(\board_state_next[82] ),
    .S(net115),
    .X(_1614_));
 sg13g2_mux2_1 _8258_ (.A0(\board_state_next[84] ),
    .A1(\board_state_next[83] ),
    .S(net115),
    .X(_1615_));
 sg13g2_mux2_1 _8259_ (.A0(\board_state_next[85] ),
    .A1(\board_state_next[84] ),
    .S(net115),
    .X(_1616_));
 sg13g2_mux2_1 _8260_ (.A0(\board_state_next[86] ),
    .A1(\board_state_next[85] ),
    .S(net115),
    .X(_1617_));
 sg13g2_mux2_1 _8261_ (.A0(\board_state_next[87] ),
    .A1(\board_state_next[86] ),
    .S(net115),
    .X(_1618_));
 sg13g2_mux2_1 _8262_ (.A0(\board_state_next[88] ),
    .A1(\board_state_next[87] ),
    .S(net115),
    .X(_1619_));
 sg13g2_mux2_1 _8263_ (.A0(\board_state_next[89] ),
    .A1(\board_state_next[88] ),
    .S(net115),
    .X(_1620_));
 sg13g2_buf_1 _8264_ (.A(_3514_),
    .X(_3572_));
 sg13g2_mux2_1 _8265_ (.A0(\board_state_next[8] ),
    .A1(\board_state_next[7] ),
    .S(net114),
    .X(_1621_));
 sg13g2_mux2_1 _8266_ (.A0(\board_state_next[90] ),
    .A1(\board_state_next[89] ),
    .S(net114),
    .X(_1622_));
 sg13g2_mux2_1 _8267_ (.A0(\board_state_next[91] ),
    .A1(\board_state_next[90] ),
    .S(net114),
    .X(_1623_));
 sg13g2_mux2_1 _8268_ (.A0(\board_state_next[92] ),
    .A1(\board_state_next[91] ),
    .S(net114),
    .X(_1624_));
 sg13g2_mux2_1 _8269_ (.A0(\board_state_next[93] ),
    .A1(\board_state_next[92] ),
    .S(_3572_),
    .X(_1625_));
 sg13g2_mux2_1 _8270_ (.A0(\board_state_next[94] ),
    .A1(\board_state_next[93] ),
    .S(net114),
    .X(_1626_));
 sg13g2_mux2_1 _8271_ (.A0(\board_state_next[95] ),
    .A1(\board_state_next[94] ),
    .S(_3572_),
    .X(_1627_));
 sg13g2_mux2_1 _8272_ (.A0(\board_state_next[96] ),
    .A1(\board_state_next[95] ),
    .S(net114),
    .X(_1628_));
 sg13g2_mux2_1 _8273_ (.A0(\board_state_next[97] ),
    .A1(\board_state_next[96] ),
    .S(net114),
    .X(_1629_));
 sg13g2_mux2_1 _8274_ (.A0(\board_state_next[98] ),
    .A1(\board_state_next[97] ),
    .S(net114),
    .X(_1630_));
 sg13g2_mux2_1 _8275_ (.A0(\board_state_next[99] ),
    .A1(\board_state_next[98] ),
    .S(_3515_),
    .X(_1631_));
 sg13g2_mux2_1 _8276_ (.A0(\board_state_next[9] ),
    .A1(\board_state_next[8] ),
    .S(_3515_),
    .X(_1632_));
 sg13g2_o21ai_1 _8277_ (.B1(_2153_),
    .Y(_1651_),
    .A1(_2098_),
    .A2(_2150_));
 sg13g2_xor2_1 _8278_ (.B(_2138_),
    .A(_0070_),
    .X(_3573_));
 sg13g2_a22oi_1 _8279_ (.Y(_3574_),
    .B1(_2136_),
    .B2(_3573_),
    .A2(_2140_),
    .A1(\hvsync_inst.vpos[3] ));
 sg13g2_inv_1 _8280_ (.Y(_1652_),
    .A(_3574_));
 sg13g2_buf_1 _8281_ (.A(_2095_),
    .X(_3575_));
 sg13g2_inv_1 _8282_ (.Y(_3576_),
    .A(\hvsync_inst.vpos[3] ));
 sg13g2_nor2_1 _8283_ (.A(_3576_),
    .B(_2138_),
    .Y(_3577_));
 sg13g2_nand2_1 _8284_ (.Y(_3578_),
    .A(_2136_),
    .B(_3577_));
 sg13g2_nor2b_1 _8285_ (.A(_3577_),
    .B_N(_2134_),
    .Y(_3579_));
 sg13g2_o21ai_1 _8286_ (.B1(net347),
    .Y(_3580_),
    .A1(net213),
    .A2(_3579_));
 sg13g2_o21ai_1 _8287_ (.B1(_3580_),
    .Y(_1653_),
    .A1(net347),
    .A2(_3578_));
 sg13g2_nand2_1 _8288_ (.Y(_3581_),
    .A(_2095_),
    .B(_3577_));
 sg13g2_a21o_1 _8289_ (.A2(_3581_),
    .A1(_2134_),
    .B1(net213),
    .X(_3582_));
 sg13g2_nor3_1 _8290_ (.A(_2092_),
    .B(_2142_),
    .C(_3581_),
    .Y(_3583_));
 sg13g2_a21o_1 _8291_ (.A2(_3582_),
    .A1(_2092_),
    .B1(_3583_),
    .X(_1654_));
 sg13g2_nand3_1 _8292_ (.B(net347),
    .C(_3577_),
    .A(_2092_),
    .Y(_3584_));
 sg13g2_a21o_1 _8293_ (.A2(_3584_),
    .A1(_2134_),
    .B1(net213),
    .X(_3585_));
 sg13g2_nor2_1 _8294_ (.A(_2093_),
    .B(_3584_),
    .Y(_3586_));
 sg13g2_a22oi_1 _8295_ (.Y(_3587_),
    .B1(_3586_),
    .B2(_2136_),
    .A2(_3585_),
    .A1(_2093_));
 sg13g2_inv_1 _8296_ (.Y(_1655_),
    .A(_3587_));
 sg13g2_nor2_1 _8297_ (.A(_2094_),
    .B(_3581_),
    .Y(_3588_));
 sg13g2_nand2_1 _8298_ (.Y(_3589_),
    .A(_2136_),
    .B(_3588_));
 sg13g2_nor2b_1 _8299_ (.A(_3588_),
    .B_N(_2134_),
    .Y(_3590_));
 sg13g2_o21ai_1 _8300_ (.B1(_2099_),
    .Y(_3591_),
    .A1(net213),
    .A2(_3590_));
 sg13g2_o21ai_1 _8301_ (.B1(_3591_),
    .Y(_1656_),
    .A1(_2099_),
    .A2(_3589_));
 sg13g2_and2_1 _8302_ (.A(_2099_),
    .B(_3588_),
    .X(_3592_));
 sg13g2_buf_1 _8303_ (.A(_3592_),
    .X(_3593_));
 sg13g2_nand2_1 _8304_ (.Y(_3594_),
    .A(_2136_),
    .B(_3593_));
 sg13g2_nor2b_1 _8305_ (.A(_3593_),
    .B_N(_2134_),
    .Y(_3595_));
 sg13g2_o21ai_1 _8306_ (.B1(_2090_),
    .Y(_3596_),
    .A1(net213),
    .A2(_3595_));
 sg13g2_o21ai_1 _8307_ (.B1(_3596_),
    .Y(_1657_),
    .A1(_2090_),
    .A2(_3594_));
 sg13g2_a21oi_1 _8308_ (.A1(_2090_),
    .A2(_3593_),
    .Y(_3597_),
    .B1(_2142_));
 sg13g2_o21ai_1 _8309_ (.B1(\hvsync_inst.vpos[9] ),
    .Y(_3598_),
    .A1(net213),
    .A2(_3597_));
 sg13g2_o21ai_1 _8310_ (.B1(_3598_),
    .Y(_1658_),
    .A1(_2091_),
    .A2(_3594_));
 sg13g2_buf_1 _8311_ (.A(_2065_),
    .X(_3599_));
 sg13g2_nor2_1 _8312_ (.A(_1888_),
    .B(_1886_),
    .Y(_3600_));
 sg13g2_nor3_1 _8313_ (.A(_1887_),
    .B(net388),
    .C(_2064_),
    .Y(_3601_));
 sg13g2_nor2_1 _8314_ (.A(_3600_),
    .B(_3601_),
    .Y(_3602_));
 sg13g2_and2_1 _8315_ (.A(net297),
    .B(_3602_),
    .X(_3603_));
 sg13g2_nor3_1 _8316_ (.A(_1935_),
    .B(_1877_),
    .C(_1922_),
    .Y(_3604_));
 sg13g2_a21oi_1 _8317_ (.A1(_3602_),
    .A2(_3604_),
    .Y(_3605_),
    .B1(\uart_rx_inst.out_latched ));
 sg13g2_nor4_1 _8318_ (.A(net271),
    .B(net274),
    .C(_3603_),
    .D(_3605_),
    .Y(_1744_));
 sg13g2_nand3b_1 _8319_ (.B(_2070_),
    .C(net262),
    .Y(_3606_),
    .A_N(_1800_));
 sg13g2_a21oi_1 _8320_ (.A1(_1801_),
    .A2(_3606_),
    .Y(_1773_),
    .B1(net272));
 sg13g2_nand2_1 _8321_ (.Y(_3607_),
    .A(_1998_),
    .B(_1997_));
 sg13g2_nor4_1 _8322_ (.A(net381),
    .B(net400),
    .C(_2008_),
    .D(_1990_),
    .Y(_3608_));
 sg13g2_a22oi_1 _8323_ (.Y(_3609_),
    .B1(_3608_),
    .B2(_2085_),
    .A2(_3607_),
    .A1(net381));
 sg13g2_a21oi_1 _8324_ (.A1(_3510_),
    .A2(_3609_),
    .Y(_3610_),
    .B1(_2346_));
 sg13g2_nor2_1 _8325_ (.A(net381),
    .B(_2346_),
    .Y(_3611_));
 sg13g2_nand2_1 _8326_ (.Y(_3612_),
    .A(_3510_),
    .B(_3609_));
 sg13g2_buf_1 _8327_ (.A(_3612_),
    .X(_3613_));
 sg13g2_a221oi_1 _8328_ (.B2(_3611_),
    .C1(_3613_),
    .B1(_1827_),
    .A1(net381),
    .Y(_3614_),
    .A2(net396));
 sg13g2_nor3_1 _8329_ (.A(net271),
    .B(_3610_),
    .C(_3614_),
    .Y(_0600_));
 sg13g2_a21oi_1 _8330_ (.A1(_1892_),
    .A2(_1991_),
    .Y(_3615_),
    .B1(net223));
 sg13g2_buf_2 _8331_ (.A(_3615_),
    .X(_3616_));
 sg13g2_xor2_1 _8332_ (.B(_2027_),
    .A(_1814_),
    .X(_3617_));
 sg13g2_a22oi_1 _8333_ (.Y(_3618_),
    .B1(_3616_),
    .B2(_3617_),
    .A2(_3613_),
    .A1(_1817_));
 sg13g2_nor2_1 _8334_ (.A(net275),
    .B(_3618_),
    .Y(_0601_));
 sg13g2_xnor2_1 _8335_ (.Y(_3619_),
    .A(_2378_),
    .B(_2484_));
 sg13g2_a22oi_1 _8336_ (.Y(_3620_),
    .B1(_3616_),
    .B2(_3619_),
    .A2(net223),
    .A1(_2336_));
 sg13g2_nor2_1 _8337_ (.A(net275),
    .B(_3620_),
    .Y(_0602_));
 sg13g2_buf_2 _8338_ (.A(_0074_),
    .X(_3621_));
 sg13g2_xnor2_1 _8339_ (.Y(_3622_),
    .A(_3621_),
    .B(_2352_));
 sg13g2_a22oi_1 _8340_ (.Y(_3623_),
    .B1(_3616_),
    .B2(_3622_),
    .A2(net223),
    .A1(net318));
 sg13g2_nor2_1 _8341_ (.A(net275),
    .B(_3623_),
    .Y(_0603_));
 sg13g2_buf_1 _8342_ (.A(_0075_),
    .X(_3624_));
 sg13g2_xnor2_1 _8343_ (.Y(_3625_),
    .A(_3624_),
    .B(_2503_));
 sg13g2_a22oi_1 _8344_ (.Y(_3626_),
    .B1(_3616_),
    .B2(_3625_),
    .A2(net223),
    .A1(net363));
 sg13g2_nor2_1 _8345_ (.A(net275),
    .B(_3626_),
    .Y(_0604_));
 sg13g2_xnor2_1 _8346_ (.Y(_3627_),
    .A(_0076_),
    .B(_2353_));
 sg13g2_a22oi_1 _8347_ (.Y(_3628_),
    .B1(_3616_),
    .B2(_3627_),
    .A2(net223),
    .A1(net375));
 sg13g2_nor2_1 _8348_ (.A(net275),
    .B(_3628_),
    .Y(_0605_));
 sg13g2_nor2_1 _8349_ (.A(_2423_),
    .B(_2574_),
    .Y(_3629_));
 sg13g2_xnor2_1 _8350_ (.Y(_3630_),
    .A(_2551_),
    .B(_3629_));
 sg13g2_a22oi_1 _8351_ (.Y(_3631_),
    .B1(_3616_),
    .B2(_3630_),
    .A2(net223),
    .A1(net376));
 sg13g2_nor2_1 _8352_ (.A(net275),
    .B(_3631_),
    .Y(_0606_));
 sg13g2_buf_1 _8353_ (.A(net330),
    .X(_3632_));
 sg13g2_nand2_1 _8354_ (.Y(_3633_),
    .A(net376),
    .B(_3629_));
 sg13g2_xor2_1 _8355_ (.B(_3633_),
    .A(_0078_),
    .X(_3634_));
 sg13g2_a22oi_1 _8356_ (.Y(_3635_),
    .B1(_3616_),
    .B2(_3634_),
    .A2(net223),
    .A1(net394));
 sg13g2_nor2_1 _8357_ (.A(net265),
    .B(_3635_),
    .Y(_0607_));
 sg13g2_nand3_1 _8358_ (.B(net376),
    .C(_3629_),
    .A(net394),
    .Y(_3636_));
 sg13g2_xor2_1 _8359_ (.B(_3636_),
    .A(_0065_),
    .X(_3637_));
 sg13g2_a22oi_1 _8360_ (.Y(_3638_),
    .B1(_3616_),
    .B2(_3637_),
    .A2(net223),
    .A1(net362));
 sg13g2_nor2_1 _8361_ (.A(net265),
    .B(_3638_),
    .Y(_0608_));
 sg13g2_o21ai_1 _8362_ (.B1(_1795_),
    .Y(_3639_),
    .A1(_2040_),
    .A2(_1998_));
 sg13g2_nor2_2 _8363_ (.A(_2043_),
    .B(_3639_),
    .Y(_3640_));
 sg13g2_buf_1 _8364_ (.A(\colindex[0] ),
    .X(_3641_));
 sg13g2_inv_1 _8365_ (.Y(_3642_),
    .A(_0079_));
 sg13g2_nor3_1 _8366_ (.A(_1996_),
    .B(_3641_),
    .C(_3642_),
    .Y(_3643_));
 sg13g2_nor2b_1 _8367_ (.A(_3640_),
    .B_N(_3641_),
    .Y(_3644_));
 sg13g2_a21oi_1 _8368_ (.A1(_3640_),
    .A2(_3643_),
    .Y(_3645_),
    .B1(_3644_));
 sg13g2_nor2_1 _8369_ (.A(_3632_),
    .B(_3645_),
    .Y(_1633_));
 sg13g2_o21ai_1 _8370_ (.B1(_3640_),
    .Y(_3646_),
    .A1(_1996_),
    .A2(_3642_));
 sg13g2_nand2_1 _8371_ (.Y(_3647_),
    .A(net372),
    .B(_3646_));
 sg13g2_nand2_1 _8372_ (.Y(_3648_),
    .A(_3641_),
    .B(_3640_));
 sg13g2_xor2_1 _8373_ (.B(_3648_),
    .A(\colindex[1] ),
    .X(_3649_));
 sg13g2_nor2_1 _8374_ (.A(_3647_),
    .B(_3649_),
    .Y(_1634_));
 sg13g2_nand3_1 _8375_ (.B(_3641_),
    .C(_3640_),
    .A(\colindex[1] ),
    .Y(_3650_));
 sg13g2_xor2_1 _8376_ (.B(_3650_),
    .A(\colindex[2] ),
    .X(_3651_));
 sg13g2_nor2_1 _8377_ (.A(_3647_),
    .B(_3651_),
    .Y(_1635_));
 sg13g2_inv_1 _8378_ (.Y(_3652_),
    .A(\colindex[3] ));
 sg13g2_nand4_1 _8379_ (.B(\colindex[1] ),
    .C(_3641_),
    .A(\colindex[2] ),
    .Y(_3653_),
    .D(_3640_));
 sg13g2_xnor2_1 _8380_ (.Y(_3654_),
    .A(_3652_),
    .B(_3653_));
 sg13g2_nor2_1 _8381_ (.A(_3647_),
    .B(_3654_),
    .Y(_1636_));
 sg13g2_nor2_1 _8382_ (.A(_3652_),
    .B(_3653_),
    .Y(_3655_));
 sg13g2_xnor2_1 _8383_ (.Y(_3656_),
    .A(\colindex[4] ),
    .B(_3655_));
 sg13g2_nor2_1 _8384_ (.A(_3647_),
    .B(_3656_),
    .Y(_1637_));
 sg13g2_o21ai_1 _8385_ (.B1(_1996_),
    .Y(_3657_),
    .A1(_2043_),
    .A2(_3639_));
 sg13g2_nand4_1 _8386_ (.B(\colindex[4] ),
    .C(_0079_),
    .A(_1997_),
    .Y(_3658_),
    .D(_3655_));
 sg13g2_a21oi_1 _8387_ (.A1(_3657_),
    .A2(_3658_),
    .Y(_1638_),
    .B1(net272));
 sg13g2_and2_1 _8388_ (.A(_0598_),
    .B(_2140_),
    .X(_1639_));
 sg13g2_xnor2_1 _8389_ (.Y(_3659_),
    .A(_2119_),
    .B(_2120_));
 sg13g2_nor2_1 _8390_ (.A(_2150_),
    .B(_3659_),
    .Y(_1640_));
 sg13g2_xnor2_1 _8391_ (.Y(_3660_),
    .A(_2117_),
    .B(_2122_));
 sg13g2_nor2_1 _8392_ (.A(net265),
    .B(_3660_),
    .Y(_1641_));
 sg13g2_nand2_1 _8393_ (.Y(_3661_),
    .A(_2117_),
    .B(_2122_));
 sg13g2_xor2_1 _8394_ (.B(_3661_),
    .A(_2118_),
    .X(_3662_));
 sg13g2_nor2_1 _8395_ (.A(net265),
    .B(_3662_),
    .Y(_1642_));
 sg13g2_xnor2_1 _8396_ (.Y(_3663_),
    .A(_2116_),
    .B(_2123_));
 sg13g2_nor2_1 _8397_ (.A(_2150_),
    .B(_3663_),
    .Y(_1643_));
 sg13g2_xnor2_1 _8398_ (.Y(_3664_),
    .A(net324),
    .B(_2124_));
 sg13g2_nor2_1 _8399_ (.A(_2150_),
    .B(_3664_),
    .Y(_1644_));
 sg13g2_nand2_1 _8400_ (.Y(_3665_),
    .A(net324),
    .B(_2124_));
 sg13g2_xor2_1 _8401_ (.B(_3665_),
    .A(net323),
    .X(_3666_));
 sg13g2_nor2_1 _8402_ (.A(_2150_),
    .B(_3666_),
    .Y(_1645_));
 sg13g2_nand3_1 _8403_ (.B(net323),
    .C(_2124_),
    .A(net324),
    .Y(_3667_));
 sg13g2_xor2_1 _8404_ (.B(_3667_),
    .A(net366),
    .X(_3668_));
 sg13g2_nor2_1 _8405_ (.A(net265),
    .B(_3668_),
    .Y(_1646_));
 sg13g2_buf_2 _8406_ (.A(_2125_),
    .X(_3669_));
 sg13g2_nand4_1 _8407_ (.B(net366),
    .C(net323),
    .A(net324),
    .Y(_3670_),
    .D(_2124_));
 sg13g2_xnor2_1 _8408_ (.Y(_3671_),
    .A(net346),
    .B(_3670_));
 sg13g2_nor2_1 _8409_ (.A(_2150_),
    .B(_3671_),
    .Y(_1647_));
 sg13g2_or2_1 _8410_ (.X(_3672_),
    .B(_3670_),
    .A(net346));
 sg13g2_xor2_1 _8411_ (.B(_3672_),
    .A(_2114_),
    .X(_3673_));
 sg13g2_nor2_1 _8412_ (.A(_2150_),
    .B(_3673_),
    .Y(_1648_));
 sg13g2_xor2_1 _8413_ (.B(\lfsr.lfsr_reg[12] ),
    .A(\lfsr.lfsr_reg[15] ),
    .X(_3674_));
 sg13g2_xor2_1 _8414_ (.B(\lfsr.lfsr_reg[10] ),
    .A(\lfsr.lfsr_reg[13] ),
    .X(_3675_));
 sg13g2_xnor2_1 _8415_ (.Y(_3676_),
    .A(_3674_),
    .B(_3675_));
 sg13g2_nand2_1 _8416_ (.Y(_1659_),
    .A(net329),
    .B(_3676_));
 sg13g2_and2_1 _8417_ (.A(net329),
    .B(\lfsr.lfsr_reg[9] ),
    .X(_1660_));
 sg13g2_and2_1 _8418_ (.A(net329),
    .B(\lfsr.lfsr_reg[10] ),
    .X(_1661_));
 sg13g2_buf_1 _8419_ (.A(net372),
    .X(_3677_));
 sg13g2_and2_1 _8420_ (.A(net296),
    .B(\lfsr.lfsr_reg[11] ),
    .X(_1662_));
 sg13g2_and2_1 _8421_ (.A(net296),
    .B(\lfsr.lfsr_reg[12] ),
    .X(_1663_));
 sg13g2_and2_1 _8422_ (.A(net296),
    .B(\lfsr.lfsr_reg[13] ),
    .X(_1664_));
 sg13g2_and2_1 _8423_ (.A(net296),
    .B(\lfsr.lfsr_reg[14] ),
    .X(_1665_));
 sg13g2_and2_1 _8424_ (.A(net296),
    .B(\lfsr.lfsr_reg[0] ),
    .X(_1666_));
 sg13g2_and2_1 _8425_ (.A(net296),
    .B(\lfsr.lfsr_reg[1] ),
    .X(_1667_));
 sg13g2_and2_1 _8426_ (.A(net296),
    .B(\lfsr.lfsr_reg[2] ),
    .X(_1668_));
 sg13g2_and2_1 _8427_ (.A(_3677_),
    .B(\lfsr.lfsr_reg[3] ),
    .X(_1669_));
 sg13g2_and2_1 _8428_ (.A(net296),
    .B(\lfsr.lfsr_reg[4] ),
    .X(_1670_));
 sg13g2_and2_1 _8429_ (.A(_3677_),
    .B(\lfsr.lfsr_reg[5] ),
    .X(_1671_));
 sg13g2_and2_1 _8430_ (.A(net322),
    .B(\lfsr.lfsr_reg[6] ),
    .X(_1672_));
 sg13g2_and2_1 _8431_ (.A(net322),
    .B(\lfsr.lfsr_reg[7] ),
    .X(_1673_));
 sg13g2_and2_1 _8432_ (.A(net322),
    .B(\lfsr.lfsr_reg[8] ),
    .X(_1674_));
 sg13g2_inv_2 _8433_ (.Y(_3678_),
    .A(_2017_));
 sg13g2_nor2_1 _8434_ (.A(_2085_),
    .B(net371),
    .Y(_3679_));
 sg13g2_nor2_1 _8435_ (.A(net387),
    .B(net345),
    .Y(_3680_));
 sg13g2_a21oi_1 _8436_ (.A1(net345),
    .A2(_3679_),
    .Y(_3681_),
    .B1(_3680_));
 sg13g2_nor2_1 _8437_ (.A(net265),
    .B(_3681_),
    .Y(_1675_));
 sg13g2_buf_1 _8438_ (.A(net386),
    .X(_3682_));
 sg13g2_inv_2 _8439_ (.Y(_3683_),
    .A(_2012_));
 sg13g2_nor2b_1 _8440_ (.A(net386),
    .B_N(_2017_),
    .Y(_3684_));
 sg13g2_buf_2 _8441_ (.A(_3684_),
    .X(_3685_));
 sg13g2_buf_1 _8442_ (.A(_2017_),
    .X(_3686_));
 sg13g2_buf_1 _8443_ (.A(net343),
    .X(_3687_));
 sg13g2_inv_1 _8444_ (.Y(_3688_),
    .A(net386));
 sg13g2_nor2_1 _8445_ (.A(net295),
    .B(_3688_),
    .Y(_3689_));
 sg13g2_a21o_1 _8446_ (.A2(_3685_),
    .A1(net387),
    .B1(_3689_),
    .X(_3690_));
 sg13g2_a22oi_1 _8447_ (.Y(_3691_),
    .B1(_3683_),
    .B2(_3690_),
    .A2(_3682_),
    .A1(_2085_));
 sg13g2_nor2_1 _8448_ (.A(net265),
    .B(_3691_),
    .Y(_1676_));
 sg13g2_nand2_1 _8449_ (.Y(_3692_),
    .A(net343),
    .B(net344));
 sg13g2_or2_1 _8450_ (.X(_3693_),
    .B(_2012_),
    .A(net370));
 sg13g2_buf_1 _8451_ (.A(_3693_),
    .X(_3694_));
 sg13g2_nor2_1 _8452_ (.A(_3692_),
    .B(_3694_),
    .Y(_3695_));
 sg13g2_and2_1 _8453_ (.A(net343),
    .B(net386),
    .X(_3696_));
 sg13g2_buf_1 _8454_ (.A(_3696_),
    .X(_3697_));
 sg13g2_o21ai_1 _8455_ (.B1(net387),
    .Y(_3698_),
    .A1(net371),
    .A2(_3697_));
 sg13g2_a22oi_1 _8456_ (.Y(_3699_),
    .B1(_3698_),
    .B2(net327),
    .A2(_3695_),
    .A1(net387));
 sg13g2_nor2_1 _8457_ (.A(net265),
    .B(_3699_),
    .Y(_1677_));
 sg13g2_nand2_1 _8458_ (.Y(_3700_),
    .A(_2085_),
    .B(_2013_));
 sg13g2_nand3_1 _8459_ (.B(_3679_),
    .C(_3697_),
    .A(_2016_),
    .Y(_3701_));
 sg13g2_a21oi_1 _8460_ (.A1(_3700_),
    .A2(_3701_),
    .Y(_1678_),
    .B1(net272));
 sg13g2_nor3_1 _8461_ (.A(net374),
    .B(_2085_),
    .C(_2013_),
    .Y(_3702_));
 sg13g2_nor2_2 _8462_ (.A(net327),
    .B(net371),
    .Y(_3703_));
 sg13g2_mux2_1 _8463_ (.A0(_2029_),
    .A1(_2503_),
    .S(net344),
    .X(_3704_));
 sg13g2_a22oi_1 _8464_ (.Y(_3705_),
    .B1(_3704_),
    .B2(net345),
    .A2(_3697_),
    .A1(_2029_));
 sg13g2_xnor2_1 _8465_ (.Y(_3706_),
    .A(_3624_),
    .B(_3705_));
 sg13g2_inv_1 _8466_ (.Y(_3707_),
    .A(_3624_));
 sg13g2_nor2b_1 _8467_ (.A(_2012_),
    .B_N(net370),
    .Y(_3708_));
 sg13g2_o21ai_1 _8468_ (.B1(_3708_),
    .Y(_3709_),
    .A1(_3688_),
    .A2(_2503_));
 sg13g2_a21oi_1 _8469_ (.A1(_3688_),
    .A2(_2503_),
    .Y(_3710_),
    .B1(net295));
 sg13g2_or2_1 _8470_ (.X(_3711_),
    .B(_3710_),
    .A(_3709_));
 sg13g2_nand2_1 _8471_ (.Y(_3712_),
    .A(net370),
    .B(_3624_));
 sg13g2_mux2_1 _8472_ (.A0(_3624_),
    .A1(_3712_),
    .S(_2029_),
    .X(_3713_));
 sg13g2_inv_1 _8473_ (.Y(_3714_),
    .A(net370));
 sg13g2_nor2_1 _8474_ (.A(_3714_),
    .B(_3685_),
    .Y(_3715_));
 sg13g2_a21oi_1 _8475_ (.A1(_3685_),
    .A2(_3713_),
    .Y(_3716_),
    .B1(_3715_));
 sg13g2_nor2_1 _8476_ (.A(net343),
    .B(net386),
    .Y(_3717_));
 sg13g2_a21oi_1 _8477_ (.A1(net327),
    .A2(_3717_),
    .Y(_3718_),
    .B1(_3697_));
 sg13g2_nor4_1 _8478_ (.A(_2012_),
    .B(_3707_),
    .C(_2574_),
    .D(_3718_),
    .Y(_3719_));
 sg13g2_a221oi_1 _8479_ (.B2(_3683_),
    .C1(_3719_),
    .B1(_3716_),
    .A1(_3707_),
    .Y(_3720_),
    .A2(_3711_));
 sg13g2_a21o_1 _8480_ (.A2(_3706_),
    .A1(_3703_),
    .B1(_3720_),
    .X(_3721_));
 sg13g2_buf_1 _8481_ (.A(_3721_),
    .X(_3722_));
 sg13g2_nand2_1 _8482_ (.Y(_3723_),
    .A(_3621_),
    .B(_2352_));
 sg13g2_a21oi_1 _8483_ (.A1(_2020_),
    .A2(_3692_),
    .Y(_3724_),
    .B1(_3723_));
 sg13g2_nor3_1 _8484_ (.A(net295),
    .B(_3621_),
    .C(_2352_),
    .Y(_3725_));
 sg13g2_o21ai_1 _8485_ (.B1(_3683_),
    .Y(_3726_),
    .A1(_3724_),
    .A2(_3725_));
 sg13g2_nand2b_1 _8486_ (.Y(_3727_),
    .B(net344),
    .A_N(_3621_));
 sg13g2_a21oi_1 _8487_ (.A1(net295),
    .A2(_2352_),
    .Y(_3728_),
    .B1(_3727_));
 sg13g2_o21ai_1 _8488_ (.B1(_3685_),
    .Y(_3729_),
    .A1(_3621_),
    .A2(_2433_));
 sg13g2_or2_1 _8489_ (.X(_3730_),
    .B(_2014_),
    .A(net386));
 sg13g2_buf_1 _8490_ (.A(_3730_),
    .X(_3731_));
 sg13g2_o21ai_1 _8491_ (.B1(_3683_),
    .Y(_3732_),
    .A1(_3678_),
    .A2(_3731_));
 sg13g2_and3_1 _8492_ (.X(_3733_),
    .A(net327),
    .B(_3621_),
    .C(_2433_));
 sg13g2_a221oi_1 _8493_ (.B2(_3621_),
    .C1(_3733_),
    .B1(_3732_),
    .A1(_3708_),
    .Y(_3734_),
    .A2(_3729_));
 sg13g2_nor2_1 _8494_ (.A(_3728_),
    .B(_3734_),
    .Y(_3735_));
 sg13g2_a21oi_1 _8495_ (.A1(_2020_),
    .A2(_3692_),
    .Y(_3736_),
    .B1(_2433_));
 sg13g2_a21oi_1 _8496_ (.A1(_2352_),
    .A2(_3689_),
    .Y(_3737_),
    .B1(_3736_));
 sg13g2_xnor2_1 _8497_ (.Y(_3738_),
    .A(_3621_),
    .B(_3737_));
 sg13g2_a22oi_1 _8498_ (.Y(_3739_),
    .B1(_3738_),
    .B2(_3703_),
    .A2(_3735_),
    .A1(_3726_));
 sg13g2_buf_4 _8499_ (.X(_3740_),
    .A(_3739_));
 sg13g2_nand2_1 _8500_ (.Y(_3741_),
    .A(_3722_),
    .B(_3740_));
 sg13g2_buf_2 _8501_ (.A(_3741_),
    .X(_3742_));
 sg13g2_buf_8 _8502_ (.A(_3742_),
    .X(_3743_));
 sg13g2_nor2_1 _8503_ (.A(_3678_),
    .B(_3731_),
    .Y(_3744_));
 sg13g2_nand2_1 _8504_ (.Y(_3745_),
    .A(_2018_),
    .B(_2014_));
 sg13g2_o21ai_1 _8505_ (.B1(_3683_),
    .Y(_3746_),
    .A1(net343),
    .A2(_3745_));
 sg13g2_a21oi_1 _8506_ (.A1(_3682_),
    .A2(_2015_),
    .Y(_3747_),
    .B1(net369));
 sg13g2_nor3_1 _8507_ (.A(_3744_),
    .B(_3746_),
    .C(_3747_),
    .Y(_3748_));
 sg13g2_nand4_1 _8508_ (.B(_3686_),
    .C(net320),
    .A(net396),
    .Y(_3749_),
    .D(_3731_));
 sg13g2_nor2_1 _8509_ (.A(net343),
    .B(net369),
    .Y(_3750_));
 sg13g2_and4_1 _8510_ (.A(_1806_),
    .B(_3686_),
    .C(net386),
    .D(_2014_),
    .X(_3751_));
 sg13g2_a21oi_1 _8511_ (.A1(_3745_),
    .A2(_3750_),
    .Y(_3752_),
    .B1(_3751_));
 sg13g2_a21o_1 _8512_ (.A2(_3752_),
    .A1(_3749_),
    .B1(_2012_),
    .X(_3753_));
 sg13g2_o21ai_1 _8513_ (.B1(_3753_),
    .Y(_3754_),
    .A1(_1806_),
    .A2(_3748_));
 sg13g2_buf_1 _8514_ (.A(_3754_),
    .X(_3755_));
 sg13g2_buf_4 _8515_ (.X(_3756_),
    .A(_3755_));
 sg13g2_buf_8 _8516_ (.A(_3756_),
    .X(_3757_));
 sg13g2_buf_2 _8517_ (.A(net188),
    .X(_3758_));
 sg13g2_and2_1 _8518_ (.A(net370),
    .B(_3685_),
    .X(_3759_));
 sg13g2_xor2_1 _8519_ (.B(_3617_),
    .A(net370),
    .X(_3760_));
 sg13g2_xnor2_1 _8520_ (.Y(_3761_),
    .A(net343),
    .B(net344));
 sg13g2_nor4_1 _8521_ (.A(net343),
    .B(_3688_),
    .C(net370),
    .D(_3617_),
    .Y(_3762_));
 sg13g2_a221oi_1 _8522_ (.B2(_3761_),
    .C1(_3762_),
    .B1(_3760_),
    .A1(_3617_),
    .Y(_3763_),
    .A2(_3759_));
 sg13g2_o21ai_1 _8523_ (.B1(_0084_),
    .Y(_3764_),
    .A1(_3744_),
    .A2(_3746_));
 sg13g2_o21ai_1 _8524_ (.B1(_3764_),
    .Y(_3765_),
    .A1(_2012_),
    .A2(_3763_));
 sg13g2_buf_1 _8525_ (.A(_3765_),
    .X(_3766_));
 sg13g2_buf_1 _8526_ (.A(_3766_),
    .X(_3767_));
 sg13g2_buf_8 _8527_ (.A(net222),
    .X(_3768_));
 sg13g2_buf_2 _8528_ (.A(net187),
    .X(_3769_));
 sg13g2_mux4_1 _8529_ (.S0(net113),
    .A0(_0225_),
    .A1(_0226_),
    .A2(_0223_),
    .A3(_0224_),
    .S1(net112),
    .X(_3770_));
 sg13g2_mux4_1 _8530_ (.S0(net113),
    .A0(_0221_),
    .A1(_0222_),
    .A2(_0219_),
    .A3(_0220_),
    .S1(net112),
    .X(_3771_));
 sg13g2_xnor2_1 _8531_ (.Y(_3772_),
    .A(_1811_),
    .B(_2356_));
 sg13g2_nand2b_1 _8532_ (.Y(_3773_),
    .B(net295),
    .A_N(net384));
 sg13g2_o21ai_1 _8533_ (.B1(_3773_),
    .Y(_3774_),
    .A1(net295),
    .A2(_3772_));
 sg13g2_nor2_1 _8534_ (.A(net344),
    .B(_3694_),
    .Y(_3775_));
 sg13g2_nand3_1 _8535_ (.B(net384),
    .C(_2360_),
    .A(net345),
    .Y(_3776_));
 sg13g2_a21oi_1 _8536_ (.A1(net344),
    .A2(_3776_),
    .Y(_3777_),
    .B1(net327));
 sg13g2_nor4_1 _8537_ (.A(_3714_),
    .B(net384),
    .C(_2360_),
    .D(_3692_),
    .Y(_3778_));
 sg13g2_o21ai_1 _8538_ (.B1(_3683_),
    .Y(_3779_),
    .A1(_3777_),
    .A2(_3778_));
 sg13g2_and2_1 _8539_ (.A(net344),
    .B(_2015_),
    .X(_3780_));
 sg13g2_a21oi_1 _8540_ (.A1(net345),
    .A2(_2360_),
    .Y(_3781_),
    .B1(_3780_));
 sg13g2_nor2_1 _8541_ (.A(net345),
    .B(_2360_),
    .Y(_3782_));
 sg13g2_o21ai_1 _8542_ (.B1(_3683_),
    .Y(_3783_),
    .A1(_3781_),
    .A2(_3782_));
 sg13g2_nor3_1 _8543_ (.A(_3687_),
    .B(net384),
    .C(_2360_),
    .Y(_3784_));
 sg13g2_a21o_1 _8544_ (.A2(_3772_),
    .A1(_3687_),
    .B1(_3784_),
    .X(_3785_));
 sg13g2_nor2_1 _8545_ (.A(net371),
    .B(_3780_),
    .Y(_3786_));
 sg13g2_a22oi_1 _8546_ (.Y(_3787_),
    .B1(_3785_),
    .B2(_3786_),
    .A2(_3783_),
    .A1(net384));
 sg13g2_a22oi_1 _8547_ (.Y(_3788_),
    .B1(_3779_),
    .B2(_3787_),
    .A2(_3775_),
    .A1(_3774_));
 sg13g2_buf_2 _8548_ (.A(_3788_),
    .X(_3789_));
 sg13g2_buf_2 _8549_ (.A(_3789_),
    .X(_3790_));
 sg13g2_buf_2 _8550_ (.A(net111),
    .X(_3791_));
 sg13g2_mux2_1 _8551_ (.A0(_3770_),
    .A1(_3771_),
    .S(_3791_),
    .X(_3792_));
 sg13g2_nand2b_1 _8552_ (.Y(_3793_),
    .B(_3722_),
    .A_N(_3740_));
 sg13g2_buf_2 _8553_ (.A(_3793_),
    .X(_3794_));
 sg13g2_buf_8 _8554_ (.A(_3794_),
    .X(_3795_));
 sg13g2_buf_2 _8555_ (.A(_3756_),
    .X(_3796_));
 sg13g2_buf_1 _8556_ (.A(_3766_),
    .X(_3797_));
 sg13g2_buf_2 _8557_ (.A(net221),
    .X(_3798_));
 sg13g2_mux4_1 _8558_ (.S0(net186),
    .A0(_0217_),
    .A1(_0218_),
    .A2(_0215_),
    .A3(_0216_),
    .S1(net185),
    .X(_3799_));
 sg13g2_buf_2 _8559_ (.A(_3756_),
    .X(_3800_));
 sg13g2_mux4_1 _8560_ (.S0(net184),
    .A0(_0213_),
    .A1(_0214_),
    .A2(_0211_),
    .A3(_0212_),
    .S1(net185),
    .X(_3801_));
 sg13g2_buf_1 _8561_ (.A(_3789_),
    .X(_3802_));
 sg13g2_mux2_1 _8562_ (.A0(_3799_),
    .A1(_3801_),
    .S(net110),
    .X(_3803_));
 sg13g2_nand2_1 _8563_ (.Y(_3804_),
    .A(_3717_),
    .B(_3708_));
 sg13g2_nand3_1 _8564_ (.B(_3694_),
    .C(_3804_),
    .A(_2366_),
    .Y(_3805_));
 sg13g2_nor2_1 _8565_ (.A(_3697_),
    .B(_3694_),
    .Y(_3806_));
 sg13g2_nand3_1 _8566_ (.B(net393),
    .C(_3806_),
    .A(_1821_),
    .Y(_3807_));
 sg13g2_o21ai_1 _8567_ (.B1(_3807_),
    .Y(_3808_),
    .A1(_1821_),
    .A2(_3805_));
 sg13g2_xor2_1 _8568_ (.B(_3808_),
    .A(_0078_),
    .X(_3809_));
 sg13g2_nor2_1 _8569_ (.A(net345),
    .B(_0076_),
    .Y(_3810_));
 sg13g2_a22oi_1 _8570_ (.Y(_3811_),
    .B1(_3703_),
    .B2(_3810_),
    .A2(net345),
    .A1(_2367_));
 sg13g2_nand3b_1 _8571_ (.B(net344),
    .C(net295),
    .Y(_3812_),
    .A_N(net327));
 sg13g2_nand2b_1 _8572_ (.Y(_3813_),
    .B(net327),
    .A_N(net295));
 sg13g2_a21oi_1 _8573_ (.A1(_3812_),
    .A2(_3813_),
    .Y(_3814_),
    .B1(net371));
 sg13g2_mux2_1 _8574_ (.A0(_3804_),
    .A1(_3814_),
    .S(_2366_),
    .X(_3815_));
 sg13g2_o21ai_1 _8575_ (.B1(_3815_),
    .Y(_3816_),
    .A1(_3688_),
    .A2(_3811_));
 sg13g2_buf_1 _8576_ (.A(_3816_),
    .X(_3817_));
 sg13g2_xnor2_1 _8577_ (.Y(_3818_),
    .A(_1821_),
    .B(net393));
 sg13g2_nor2_1 _8578_ (.A(_3806_),
    .B(_3818_),
    .Y(_3819_));
 sg13g2_nand2b_1 _8579_ (.Y(_3820_),
    .B(_3804_),
    .A_N(_3695_));
 sg13g2_mux2_1 _8580_ (.A0(_3819_),
    .A1(_2551_),
    .S(_3820_),
    .X(_3821_));
 sg13g2_a21oi_1 _8581_ (.A1(_3806_),
    .A2(_3818_),
    .Y(_3822_),
    .B1(_3821_));
 sg13g2_buf_2 _8582_ (.A(_3822_),
    .X(_3823_));
 sg13g2_nor3_2 _8583_ (.A(_3809_),
    .B(_3817_),
    .C(_3823_),
    .Y(_3824_));
 sg13g2_o21ai_1 _8584_ (.B1(_3824_),
    .Y(_3825_),
    .A1(net71),
    .A2(_3803_));
 sg13g2_a21oi_2 _8585_ (.B1(_3720_),
    .Y(_3826_),
    .A2(_3706_),
    .A1(_3703_));
 sg13g2_nand2_1 _8586_ (.Y(_3827_),
    .A(_3826_),
    .B(_3740_));
 sg13g2_buf_2 _8587_ (.A(_3827_),
    .X(_3828_));
 sg13g2_buf_1 _8588_ (.A(_3828_),
    .X(_3829_));
 sg13g2_buf_2 _8589_ (.A(_3755_),
    .X(_3830_));
 sg13g2_buf_2 _8590_ (.A(net220),
    .X(_3831_));
 sg13g2_buf_1 _8591_ (.A(_3766_),
    .X(_3832_));
 sg13g2_buf_1 _8592_ (.A(net219),
    .X(_3833_));
 sg13g2_buf_1 _8593_ (.A(net182),
    .X(_3834_));
 sg13g2_mux4_1 _8594_ (.S0(net183),
    .A0(_0241_),
    .A1(_0242_),
    .A2(_0239_),
    .A3(_0240_),
    .S1(net109),
    .X(_3835_));
 sg13g2_buf_8 _8595_ (.A(net219),
    .X(_3836_));
 sg13g2_buf_2 _8596_ (.A(net181),
    .X(_3837_));
 sg13g2_mux4_1 _8597_ (.S0(net186),
    .A0(_0237_),
    .A1(_0238_),
    .A2(_0235_),
    .A3(_0236_),
    .S1(net108),
    .X(_3838_));
 sg13g2_buf_1 _8598_ (.A(_3789_),
    .X(_3839_));
 sg13g2_mux2_1 _8599_ (.A0(_3835_),
    .A1(_3838_),
    .S(net107),
    .X(_3840_));
 sg13g2_nor2_1 _8600_ (.A(net70),
    .B(_3840_),
    .Y(_3841_));
 sg13g2_or2_1 _8601_ (.X(_3842_),
    .B(_3740_),
    .A(_3722_));
 sg13g2_buf_2 _8602_ (.A(_3842_),
    .X(_3843_));
 sg13g2_buf_8 _8603_ (.A(_3843_),
    .X(_3844_));
 sg13g2_mux2_1 _8604_ (.A0(_0233_),
    .A1(_0231_),
    .S(net187),
    .X(_3845_));
 sg13g2_mux2_1 _8605_ (.A0(_0234_),
    .A1(_0232_),
    .S(net187),
    .X(_3846_));
 sg13g2_buf_2 _8606_ (.A(net219),
    .X(_3847_));
 sg13g2_mux2_1 _8607_ (.A0(_0229_),
    .A1(_0227_),
    .S(_3847_),
    .X(_3848_));
 sg13g2_mux2_1 _8608_ (.A0(_0230_),
    .A1(_0228_),
    .S(_3847_),
    .X(_3849_));
 sg13g2_mux4_1 _8609_ (.S0(_3758_),
    .A0(_3845_),
    .A1(_3846_),
    .A2(_3848_),
    .A3(_3849_),
    .S1(net107),
    .X(_3850_));
 sg13g2_nor2_1 _8610_ (.A(net69),
    .B(_3850_),
    .Y(_3851_));
 sg13g2_nor3_1 _8611_ (.A(_3825_),
    .B(_3841_),
    .C(_3851_),
    .Y(_3852_));
 sg13g2_o21ai_1 _8612_ (.B1(_3852_),
    .Y(_3853_),
    .A1(net72),
    .A2(_3792_));
 sg13g2_mux4_1 _8613_ (.S0(net113),
    .A0(_0137_),
    .A1(_0138_),
    .A2(_0135_),
    .A3(_0136_),
    .S1(net112),
    .X(_3854_));
 sg13g2_mux4_1 _8614_ (.S0(net113),
    .A0(_0145_),
    .A1(_0146_),
    .A2(_0143_),
    .A3(_0144_),
    .S1(net112),
    .X(_3855_));
 sg13g2_mux4_1 _8615_ (.S0(net113),
    .A0(_0133_),
    .A1(_0134_),
    .A2(_0131_),
    .A3(_0132_),
    .S1(_3769_),
    .X(_3856_));
 sg13g2_mux4_1 _8616_ (.S0(net113),
    .A0(_0141_),
    .A1(_0142_),
    .A2(_0139_),
    .A3(_0140_),
    .S1(_3769_),
    .X(_3857_));
 sg13g2_mux4_1 _8617_ (.S0(_3740_),
    .A0(_3854_),
    .A1(_3855_),
    .A2(_3856_),
    .A3(_3857_),
    .S1(net75),
    .X(_3858_));
 sg13g2_buf_1 _8618_ (.A(net219),
    .X(_3859_));
 sg13g2_mux2_1 _8619_ (.A0(_0121_),
    .A1(_0119_),
    .S(net179),
    .X(_3860_));
 sg13g2_mux2_1 _8620_ (.A0(_0122_),
    .A1(_0120_),
    .S(net179),
    .X(_3861_));
 sg13g2_buf_2 _8621_ (.A(net219),
    .X(_3862_));
 sg13g2_mux2_1 _8622_ (.A0(_0117_),
    .A1(_0115_),
    .S(net178),
    .X(_3863_));
 sg13g2_mux2_1 _8623_ (.A0(_0118_),
    .A1(_0116_),
    .S(net178),
    .X(_3864_));
 sg13g2_mux4_1 _8624_ (.S0(net113),
    .A0(_3860_),
    .A1(_3861_),
    .A2(_3863_),
    .A3(_3864_),
    .S1(_3839_),
    .X(_3865_));
 sg13g2_xnor2_1 _8625_ (.Y(_3866_),
    .A(_0078_),
    .B(_3808_));
 sg13g2_inv_1 _8626_ (.Y(_3867_),
    .A(_3817_));
 sg13g2_nor3_1 _8627_ (.A(_3866_),
    .B(_3867_),
    .C(_3823_),
    .Y(_3868_));
 sg13g2_o21ai_1 _8628_ (.B1(_3868_),
    .Y(_3869_),
    .A1(net71),
    .A2(_3865_));
 sg13g2_buf_2 _8629_ (.A(_3830_),
    .X(_3870_));
 sg13g2_mux4_1 _8630_ (.S0(net177),
    .A0(_0129_),
    .A1(_0130_),
    .A2(_0127_),
    .A3(_0128_),
    .S1(_3834_),
    .X(_3871_));
 sg13g2_mux4_1 _8631_ (.S0(net183),
    .A0(_0125_),
    .A1(_0126_),
    .A2(_0123_),
    .A3(_0124_),
    .S1(_3834_),
    .X(_3872_));
 sg13g2_mux2_1 _8632_ (.A0(_3871_),
    .A1(_3872_),
    .S(_3839_),
    .X(_3873_));
 sg13g2_nor2_1 _8633_ (.A(net72),
    .B(_3873_),
    .Y(_3874_));
 sg13g2_nor2_1 _8634_ (.A(_3869_),
    .B(_3874_),
    .Y(_3875_));
 sg13g2_o21ai_1 _8635_ (.B1(_3875_),
    .Y(_3876_),
    .A1(_3722_),
    .A2(_3858_));
 sg13g2_mux4_1 _8636_ (.S0(net183),
    .A0(_0193_),
    .A1(_0194_),
    .A2(_0191_),
    .A3(_0192_),
    .S1(net109),
    .X(_3877_));
 sg13g2_mux4_1 _8637_ (.S0(net183),
    .A0(_0189_),
    .A1(_0190_),
    .A2(_0187_),
    .A3(_0188_),
    .S1(net109),
    .X(_3878_));
 sg13g2_mux2_1 _8638_ (.A0(_3877_),
    .A1(_3878_),
    .S(net107),
    .X(_3879_));
 sg13g2_nor2_1 _8639_ (.A(net72),
    .B(_3879_),
    .Y(_3880_));
 sg13g2_mux4_1 _8640_ (.S0(net183),
    .A0(_0209_),
    .A1(_0210_),
    .A2(_0207_),
    .A3(_0208_),
    .S1(net109),
    .X(_3881_));
 sg13g2_mux4_1 _8641_ (.S0(_3831_),
    .A0(_0205_),
    .A1(_0206_),
    .A2(_0203_),
    .A3(_0204_),
    .S1(net109),
    .X(_3882_));
 sg13g2_mux2_1 _8642_ (.A0(_3881_),
    .A1(_3882_),
    .S(net107),
    .X(_3883_));
 sg13g2_nor2_1 _8643_ (.A(net70),
    .B(_3883_),
    .Y(_3884_));
 sg13g2_mux4_1 _8644_ (.S0(net183),
    .A0(_0185_),
    .A1(_0186_),
    .A2(_0183_),
    .A3(_0184_),
    .S1(net109),
    .X(_3885_));
 sg13g2_mux4_1 _8645_ (.S0(net183),
    .A0(_0181_),
    .A1(_0182_),
    .A2(_0179_),
    .A3(_0180_),
    .S1(net109),
    .X(_3886_));
 sg13g2_mux2_1 _8646_ (.A0(_3885_),
    .A1(_3886_),
    .S(net107),
    .X(_3887_));
 sg13g2_nor2_1 _8647_ (.A(net71),
    .B(_3887_),
    .Y(_3888_));
 sg13g2_mux4_1 _8648_ (.S0(_3831_),
    .A0(_0201_),
    .A1(_0202_),
    .A2(_0199_),
    .A3(_0200_),
    .S1(net108),
    .X(_3889_));
 sg13g2_mux4_1 _8649_ (.S0(net186),
    .A0(_0197_),
    .A1(_0198_),
    .A2(_0195_),
    .A3(_0196_),
    .S1(net108),
    .X(_3890_));
 sg13g2_mux2_1 _8650_ (.A0(_3889_),
    .A1(_3890_),
    .S(net107),
    .X(_3891_));
 sg13g2_and3_1 _8651_ (.X(_3892_),
    .A(_3809_),
    .B(_3817_),
    .C(_3823_));
 sg13g2_o21ai_1 _8652_ (.B1(_3892_),
    .Y(_3893_),
    .A1(net69),
    .A2(_3891_));
 sg13g2_or4_1 _8653_ (.A(_3880_),
    .B(_3884_),
    .C(_3888_),
    .D(_3893_),
    .X(_3894_));
 sg13g2_and3_1 _8654_ (.X(_3895_),
    .A(_3853_),
    .B(_3876_),
    .C(_3894_));
 sg13g2_buf_1 _8655_ (.A(net179),
    .X(_3896_));
 sg13g2_mux4_1 _8656_ (.S0(net177),
    .A0(_0089_),
    .A1(_0090_),
    .A2(_0087_),
    .A3(_0088_),
    .S1(net106),
    .X(_3897_));
 sg13g2_mux4_1 _8657_ (.S0(net177),
    .A0(_0085_),
    .A1(_0086_),
    .A2(_0082_),
    .A3(_0083_),
    .S1(net106),
    .X(_3898_));
 sg13g2_mux2_1 _8658_ (.A0(_3897_),
    .A1(_3898_),
    .S(net75),
    .X(_3899_));
 sg13g2_nor2_1 _8659_ (.A(net71),
    .B(_3899_),
    .Y(_3900_));
 sg13g2_mux4_1 _8660_ (.S0(net177),
    .A0(_0097_),
    .A1(_0098_),
    .A2(_0095_),
    .A3(_0096_),
    .S1(net106),
    .X(_3901_));
 sg13g2_mux4_1 _8661_ (.S0(net177),
    .A0(_0093_),
    .A1(_0094_),
    .A2(_0091_),
    .A3(_0092_),
    .S1(net106),
    .X(_3902_));
 sg13g2_mux2_1 _8662_ (.A0(_3901_),
    .A1(_3902_),
    .S(net75),
    .X(_3903_));
 sg13g2_nor2_1 _8663_ (.A(_3743_),
    .B(_3903_),
    .Y(_3904_));
 sg13g2_buf_2 _8664_ (.A(_3755_),
    .X(_3905_));
 sg13g2_buf_2 _8665_ (.A(net218),
    .X(_3906_));
 sg13g2_mux4_1 _8666_ (.S0(_3906_),
    .A0(_0113_),
    .A1(_0114_),
    .A2(_0111_),
    .A3(_0112_),
    .S1(net106),
    .X(_3907_));
 sg13g2_mux4_1 _8667_ (.S0(_3906_),
    .A0(_0109_),
    .A1(_0110_),
    .A2(_0107_),
    .A3(_0108_),
    .S1(net106),
    .X(_3908_));
 sg13g2_mux2_1 _8668_ (.A0(_3907_),
    .A1(_3908_),
    .S(net75),
    .X(_3909_));
 sg13g2_nor2_1 _8669_ (.A(_3829_),
    .B(_3909_),
    .Y(_3910_));
 sg13g2_mux4_1 _8670_ (.S0(net177),
    .A0(_0105_),
    .A1(_0106_),
    .A2(_0103_),
    .A3(_0104_),
    .S1(net106),
    .X(_3911_));
 sg13g2_mux4_1 _8671_ (.S0(net177),
    .A0(_0101_),
    .A1(_0102_),
    .A2(_0099_),
    .A3(_0100_),
    .S1(net106),
    .X(_3912_));
 sg13g2_mux2_1 _8672_ (.A0(_3911_),
    .A1(_3912_),
    .S(net107),
    .X(_3913_));
 sg13g2_nor3_1 _8673_ (.A(_3866_),
    .B(_3817_),
    .C(_3823_),
    .Y(_3914_));
 sg13g2_o21ai_1 _8674_ (.B1(_3914_),
    .Y(_3915_),
    .A1(_3844_),
    .A2(_3913_));
 sg13g2_nor4_1 _8675_ (.A(_3900_),
    .B(_3904_),
    .C(_3910_),
    .D(_3915_),
    .Y(_3916_));
 sg13g2_mux4_1 _8676_ (.S0(net176),
    .A0(_0273_),
    .A1(_0274_),
    .A2(_0271_),
    .A3(_0272_),
    .S1(_3896_),
    .X(_3917_));
 sg13g2_mux4_1 _8677_ (.S0(_3870_),
    .A0(_0269_),
    .A1(_0270_),
    .A2(_0267_),
    .A3(_0268_),
    .S1(_3896_),
    .X(_3918_));
 sg13g2_mux2_1 _8678_ (.A0(_3917_),
    .A1(_3918_),
    .S(_3791_),
    .X(_3919_));
 sg13g2_nor2_1 _8679_ (.A(_3829_),
    .B(_3919_),
    .Y(_3920_));
 sg13g2_mux4_1 _8680_ (.S0(net186),
    .A0(_0261_),
    .A1(_0262_),
    .A2(_0259_),
    .A3(_0260_),
    .S1(net108),
    .X(_3921_));
 sg13g2_a21o_1 _8681_ (.A2(_3921_),
    .A1(net75),
    .B1(_3843_),
    .X(_3922_));
 sg13g2_mux4_1 _8682_ (.S0(_3870_),
    .A0(_0265_),
    .A1(_0266_),
    .A2(_0263_),
    .A3(_0264_),
    .S1(net109),
    .X(_3923_));
 sg13g2_nor2b_1 _8683_ (.A(net75),
    .B_N(_3923_),
    .Y(_3924_));
 sg13g2_nor3_1 _8684_ (.A(_3809_),
    .B(_3867_),
    .C(_3823_),
    .Y(_3925_));
 sg13g2_o21ai_1 _8685_ (.B1(_3925_),
    .Y(_3926_),
    .A1(_3922_),
    .A2(_3924_));
 sg13g2_mux4_1 _8686_ (.S0(net176),
    .A0(_0257_),
    .A1(_0258_),
    .A2(_0255_),
    .A3(_0256_),
    .S1(net112),
    .X(_3927_));
 sg13g2_mux4_1 _8687_ (.S0(net176),
    .A0(_0253_),
    .A1(_0254_),
    .A2(_0251_),
    .A3(_0252_),
    .S1(net112),
    .X(_3928_));
 sg13g2_mux2_1 _8688_ (.A0(_3927_),
    .A1(_3928_),
    .S(net75),
    .X(_3929_));
 sg13g2_nor2_1 _8689_ (.A(_3743_),
    .B(_3929_),
    .Y(_3930_));
 sg13g2_mux4_1 _8690_ (.S0(_3758_),
    .A0(_0249_),
    .A1(_0250_),
    .A2(_0247_),
    .A3(_0248_),
    .S1(net112),
    .X(_3931_));
 sg13g2_mux4_1 _8691_ (.S0(net176),
    .A0(_0245_),
    .A1(_0246_),
    .A2(_0243_),
    .A3(_0244_),
    .S1(net112),
    .X(_3932_));
 sg13g2_mux2_1 _8692_ (.A0(_3931_),
    .A1(_3932_),
    .S(net75),
    .X(_3933_));
 sg13g2_nor2_1 _8693_ (.A(net71),
    .B(_3933_),
    .Y(_3934_));
 sg13g2_nor4_1 _8694_ (.A(_3920_),
    .B(_3926_),
    .C(_3930_),
    .D(_3934_),
    .Y(_3935_));
 sg13g2_nand4_1 _8695_ (.B(net376),
    .C(net375),
    .A(net394),
    .Y(_3936_),
    .D(_3806_));
 sg13g2_o21ai_1 _8696_ (.B1(_3936_),
    .Y(_3937_),
    .A1(_2536_),
    .A2(_3805_));
 sg13g2_xnor2_1 _8697_ (.Y(_3938_),
    .A(_0065_),
    .B(_3937_));
 sg13g2_buf_2 _8698_ (.A(_3755_),
    .X(_3939_));
 sg13g2_mux4_1 _8699_ (.S0(net217),
    .A0(_0329_),
    .A1(_0330_),
    .A2(_0327_),
    .A3(_0328_),
    .S1(net178),
    .X(_3940_));
 sg13g2_mux4_1 _8700_ (.S0(net217),
    .A0(_0325_),
    .A1(_0326_),
    .A2(_0323_),
    .A3(_0324_),
    .S1(net178),
    .X(_3941_));
 sg13g2_buf_2 _8701_ (.A(_3789_),
    .X(_3942_));
 sg13g2_mux2_1 _8702_ (.A0(_3940_),
    .A1(_3941_),
    .S(net105),
    .X(_3943_));
 sg13g2_nor2_1 _8703_ (.A(_3843_),
    .B(_3943_),
    .Y(_3944_));
 sg13g2_mux4_1 _8704_ (.S0(_3756_),
    .A0(_0313_),
    .A1(_0314_),
    .A2(_0311_),
    .A3(_0312_),
    .S1(net182),
    .X(_3945_));
 sg13g2_mux4_1 _8705_ (.S0(_3756_),
    .A0(_0309_),
    .A1(_0310_),
    .A2(_0307_),
    .A3(_0308_),
    .S1(net181),
    .X(_3946_));
 sg13g2_mux2_1 _8706_ (.A0(_3945_),
    .A1(_3946_),
    .S(_3789_),
    .X(_3947_));
 sg13g2_and3_1 _8707_ (.X(_3948_),
    .A(_3866_),
    .B(_3817_),
    .C(_3823_));
 sg13g2_o21ai_1 _8708_ (.B1(_3948_),
    .Y(_3949_),
    .A1(_3794_),
    .A2(_3947_));
 sg13g2_buf_2 _8709_ (.A(_3832_),
    .X(_3950_));
 sg13g2_mux4_1 _8710_ (.S0(net218),
    .A0(_0321_),
    .A1(_0322_),
    .A2(_0319_),
    .A3(_0320_),
    .S1(net175),
    .X(_3951_));
 sg13g2_mux4_1 _8711_ (.S0(net218),
    .A0(_0317_),
    .A1(_0318_),
    .A2(_0315_),
    .A3(_0316_),
    .S1(net175),
    .X(_3952_));
 sg13g2_mux2_1 _8712_ (.A0(_3951_),
    .A1(_3952_),
    .S(net111),
    .X(_3953_));
 sg13g2_nor2_1 _8713_ (.A(net72),
    .B(_3953_),
    .Y(_3954_));
 sg13g2_mux2_1 _8714_ (.A0(_0337_),
    .A1(_0335_),
    .S(net181),
    .X(_3955_));
 sg13g2_mux2_1 _8715_ (.A0(_0338_),
    .A1(_0336_),
    .S(net181),
    .X(_3956_));
 sg13g2_mux2_1 _8716_ (.A0(_0333_),
    .A1(_0331_),
    .S(net221),
    .X(_3957_));
 sg13g2_mux2_1 _8717_ (.A0(_0334_),
    .A1(_0332_),
    .S(net221),
    .X(_3958_));
 sg13g2_buf_2 _8718_ (.A(_3789_),
    .X(_3959_));
 sg13g2_mux4_1 _8719_ (.S0(net176),
    .A0(_3955_),
    .A1(_3956_),
    .A2(_3957_),
    .A3(_3958_),
    .S1(net104),
    .X(_3960_));
 sg13g2_nor2_1 _8720_ (.A(net70),
    .B(_3960_),
    .Y(_3961_));
 sg13g2_nor4_1 _8721_ (.A(_3944_),
    .B(_3949_),
    .C(_3954_),
    .D(_3961_),
    .Y(_3962_));
 sg13g2_mux4_1 _8722_ (.S0(_3905_),
    .A0(_0161_),
    .A1(_0162_),
    .A2(_0159_),
    .A3(_0160_),
    .S1(net179),
    .X(_3963_));
 sg13g2_mux4_1 _8723_ (.S0(_3905_),
    .A0(_0157_),
    .A1(_0158_),
    .A2(_0155_),
    .A3(_0156_),
    .S1(_3859_),
    .X(_3964_));
 sg13g2_mux2_1 _8724_ (.A0(_3963_),
    .A1(_3964_),
    .S(_3942_),
    .X(_3965_));
 sg13g2_nor2_1 _8725_ (.A(_3742_),
    .B(_3965_),
    .Y(_3966_));
 sg13g2_mux4_1 _8726_ (.S0(net220),
    .A0(_0153_),
    .A1(_0154_),
    .A2(_0151_),
    .A3(_0152_),
    .S1(net182),
    .X(_3967_));
 sg13g2_mux4_1 _8727_ (.S0(_3756_),
    .A0(_0149_),
    .A1(_0150_),
    .A2(_0147_),
    .A3(_0148_),
    .S1(net182),
    .X(_3968_));
 sg13g2_mux2_1 _8728_ (.A0(_3967_),
    .A1(_3968_),
    .S(_3789_),
    .X(_3969_));
 sg13g2_and3_1 _8729_ (.X(_3970_),
    .A(_3809_),
    .B(_3867_),
    .C(_3823_));
 sg13g2_o21ai_1 _8730_ (.B1(_3970_),
    .Y(_3971_),
    .A1(_3794_),
    .A2(_3969_));
 sg13g2_buf_2 _8731_ (.A(_3756_),
    .X(_3972_));
 sg13g2_mux4_1 _8732_ (.S0(net174),
    .A0(_0177_),
    .A1(_0178_),
    .A2(_0175_),
    .A3(_0176_),
    .S1(net175),
    .X(_3973_));
 sg13g2_mux4_1 _8733_ (.S0(net218),
    .A0(_0173_),
    .A1(_0174_),
    .A2(_0171_),
    .A3(_0172_),
    .S1(net175),
    .X(_3974_));
 sg13g2_mux2_1 _8734_ (.A0(_3973_),
    .A1(_3974_),
    .S(net111),
    .X(_3975_));
 sg13g2_nor2_1 _8735_ (.A(_3828_),
    .B(_3975_),
    .Y(_3976_));
 sg13g2_mux2_1 _8736_ (.A0(_0169_),
    .A1(_0167_),
    .S(_3836_),
    .X(_3977_));
 sg13g2_mux2_1 _8737_ (.A0(_0170_),
    .A1(_0168_),
    .S(_3836_),
    .X(_3978_));
 sg13g2_mux2_1 _8738_ (.A0(_0165_),
    .A1(_0163_),
    .S(_3797_),
    .X(_3979_));
 sg13g2_mux2_1 _8739_ (.A0(_0166_),
    .A1(_0164_),
    .S(_3797_),
    .X(_3980_));
 sg13g2_mux4_1 _8740_ (.S0(net176),
    .A0(_3977_),
    .A1(_3978_),
    .A2(_3979_),
    .A3(_3980_),
    .S1(net110),
    .X(_3981_));
 sg13g2_nor2_1 _8741_ (.A(net69),
    .B(_3981_),
    .Y(_3982_));
 sg13g2_nor4_1 _8742_ (.A(_3966_),
    .B(_3971_),
    .C(_3976_),
    .D(_3982_),
    .Y(_3983_));
 sg13g2_mux4_1 _8743_ (.S0(net218),
    .A0(_0297_),
    .A1(_0298_),
    .A2(_0295_),
    .A3(_0296_),
    .S1(net175),
    .X(_3984_));
 sg13g2_mux4_1 _8744_ (.S0(net218),
    .A0(_0293_),
    .A1(_0294_),
    .A2(_0291_),
    .A3(_0292_),
    .S1(net179),
    .X(_3985_));
 sg13g2_mux2_1 _8745_ (.A0(_3984_),
    .A1(_3985_),
    .S(net111),
    .X(_3986_));
 sg13g2_and3_1 _8746_ (.X(_3987_),
    .A(_3866_),
    .B(_3867_),
    .C(_3823_));
 sg13g2_o21ai_1 _8747_ (.B1(_3987_),
    .Y(_3988_),
    .A1(_3844_),
    .A2(_3986_));
 sg13g2_buf_2 _8748_ (.A(net222),
    .X(_3989_));
 sg13g2_mux4_1 _8749_ (.S0(net188),
    .A0(_0305_),
    .A1(_0306_),
    .A2(_0303_),
    .A3(_0304_),
    .S1(net173),
    .X(_3990_));
 sg13g2_mux4_1 _8750_ (.S0(net188),
    .A0(_0301_),
    .A1(_0302_),
    .A2(_0299_),
    .A3(_0300_),
    .S1(net173),
    .X(_3991_));
 sg13g2_mux2_1 _8751_ (.A0(_3990_),
    .A1(_3991_),
    .S(net104),
    .X(_3992_));
 sg13g2_nor2_1 _8752_ (.A(net70),
    .B(_3992_),
    .Y(_3993_));
 sg13g2_mux4_1 _8753_ (.S0(net220),
    .A0(_0281_),
    .A1(_0282_),
    .A2(_0279_),
    .A3(_0280_),
    .S1(net182),
    .X(_3994_));
 sg13g2_mux4_1 _8754_ (.S0(net220),
    .A0(_0277_),
    .A1(_0278_),
    .A2(_0275_),
    .A3(_0276_),
    .S1(net182),
    .X(_3995_));
 sg13g2_mux4_1 _8755_ (.S0(net220),
    .A0(_0289_),
    .A1(_0290_),
    .A2(_0287_),
    .A3(_0288_),
    .S1(net182),
    .X(_3996_));
 sg13g2_mux4_1 _8756_ (.S0(net220),
    .A0(_0285_),
    .A1(_0286_),
    .A2(_0283_),
    .A3(_0284_),
    .S1(net182),
    .X(_3997_));
 sg13g2_mux4_1 _8757_ (.S0(net105),
    .A0(_3994_),
    .A1(_3995_),
    .A2(_3996_),
    .A3(_3997_),
    .S1(_3740_),
    .X(_3998_));
 sg13g2_nor2_1 _8758_ (.A(_3826_),
    .B(_3998_),
    .Y(_3999_));
 sg13g2_nor3_1 _8759_ (.A(_3988_),
    .B(_3993_),
    .C(_3999_),
    .Y(_4000_));
 sg13g2_or3_1 _8760_ (.A(_3962_),
    .B(_3983_),
    .C(_4000_),
    .X(_4001_));
 sg13g2_nor4_1 _8761_ (.A(_3916_),
    .B(_3935_),
    .C(_3938_),
    .D(_4001_),
    .Y(_4002_));
 sg13g2_mux4_1 _8762_ (.S0(net217),
    .A0(_0505_),
    .A1(_0506_),
    .A2(_0503_),
    .A3(_0504_),
    .S1(net178),
    .X(_4003_));
 sg13g2_mux4_1 _8763_ (.S0(net217),
    .A0(_0501_),
    .A1(_0502_),
    .A2(_0499_),
    .A3(_0500_),
    .S1(_3862_),
    .X(_4004_));
 sg13g2_mux2_1 _8764_ (.A0(_4003_),
    .A1(_4004_),
    .S(net105),
    .X(_4005_));
 sg13g2_nor2_1 _8765_ (.A(_3794_),
    .B(_4005_),
    .Y(_4006_));
 sg13g2_mux4_1 _8766_ (.S0(_3939_),
    .A0(_0521_),
    .A1(_0522_),
    .A2(_0519_),
    .A3(_0520_),
    .S1(_3859_),
    .X(_4007_));
 sg13g2_mux4_1 _8767_ (.S0(_3939_),
    .A0(_0517_),
    .A1(_0518_),
    .A2(_0515_),
    .A3(_0516_),
    .S1(_3862_),
    .X(_4008_));
 sg13g2_mux2_1 _8768_ (.A0(_4007_),
    .A1(_4008_),
    .S(net105),
    .X(_4009_));
 sg13g2_nor2_1 _8769_ (.A(_3843_),
    .B(_4009_),
    .Y(_4010_));
 sg13g2_mux2_1 _8770_ (.A0(_0513_),
    .A1(_0511_),
    .S(net221),
    .X(_4011_));
 sg13g2_mux2_1 _8771_ (.A0(_0514_),
    .A1(_0512_),
    .S(net221),
    .X(_4012_));
 sg13g2_mux2_1 _8772_ (.A0(_0509_),
    .A1(_0507_),
    .S(_3767_),
    .X(_4013_));
 sg13g2_mux2_1 _8773_ (.A0(_0510_),
    .A1(_0508_),
    .S(_3767_),
    .X(_4014_));
 sg13g2_mux4_1 _8774_ (.S0(net176),
    .A0(_4011_),
    .A1(_4012_),
    .A2(_4013_),
    .A3(_4014_),
    .S1(_3959_),
    .X(_4015_));
 sg13g2_nor2_1 _8775_ (.A(_3742_),
    .B(_4015_),
    .Y(_4016_));
 sg13g2_mux4_1 _8776_ (.S0(net220),
    .A0(_0529_),
    .A1(_0530_),
    .A2(_0527_),
    .A3(_0528_),
    .S1(_3833_),
    .X(_4017_));
 sg13g2_mux4_1 _8777_ (.S0(_3830_),
    .A0(_0525_),
    .A1(_0526_),
    .A2(_0523_),
    .A3(_0524_),
    .S1(_3833_),
    .X(_4018_));
 sg13g2_mux2_1 _8778_ (.A0(_4017_),
    .A1(_4018_),
    .S(_3942_),
    .X(_4019_));
 sg13g2_o21ai_1 _8779_ (.B1(_3925_),
    .Y(_4020_),
    .A1(_3828_),
    .A2(_4019_));
 sg13g2_nor4_1 _8780_ (.A(_4006_),
    .B(_4010_),
    .C(_4016_),
    .D(_4020_),
    .Y(_4021_));
 sg13g2_mux4_1 _8781_ (.S0(net217),
    .A0(_0449_),
    .A1(_0450_),
    .A2(_0447_),
    .A3(_0448_),
    .S1(net179),
    .X(_4022_));
 sg13g2_mux4_1 _8782_ (.S0(net217),
    .A0(_0445_),
    .A1(_0446_),
    .A2(_0443_),
    .A3(_0444_),
    .S1(net178),
    .X(_4023_));
 sg13g2_mux2_1 _8783_ (.A0(_4022_),
    .A1(_4023_),
    .S(net105),
    .X(_4024_));
 sg13g2_nor2_1 _8784_ (.A(_3742_),
    .B(_4024_),
    .Y(_4025_));
 sg13g2_mux4_1 _8785_ (.S0(net218),
    .A0(_0465_),
    .A1(_0466_),
    .A2(_0463_),
    .A3(_0464_),
    .S1(net179),
    .X(_4026_));
 sg13g2_mux4_1 _8786_ (.S0(net217),
    .A0(_0461_),
    .A1(_0462_),
    .A2(_0459_),
    .A3(_0460_),
    .S1(net179),
    .X(_4027_));
 sg13g2_mux2_1 _8787_ (.A0(_4026_),
    .A1(_4027_),
    .S(net105),
    .X(_4028_));
 sg13g2_nor2_1 _8788_ (.A(_3828_),
    .B(_4028_),
    .Y(_4029_));
 sg13g2_mux2_1 _8789_ (.A0(_0457_),
    .A1(_0455_),
    .S(net221),
    .X(_4030_));
 sg13g2_mux2_1 _8790_ (.A0(_0458_),
    .A1(_0456_),
    .S(net221),
    .X(_4031_));
 sg13g2_mux2_1 _8791_ (.A0(_0453_),
    .A1(_0451_),
    .S(net222),
    .X(_4032_));
 sg13g2_mux2_1 _8792_ (.A0(_0454_),
    .A1(_0452_),
    .S(net221),
    .X(_4033_));
 sg13g2_mux4_1 _8793_ (.S0(net176),
    .A0(_4030_),
    .A1(_4031_),
    .A2(_4032_),
    .A3(_4033_),
    .S1(net104),
    .X(_4034_));
 sg13g2_nor2_1 _8794_ (.A(net69),
    .B(_4034_),
    .Y(_4035_));
 sg13g2_mux4_1 _8795_ (.S0(net217),
    .A0(_0441_),
    .A1(_0442_),
    .A2(_0439_),
    .A3(_0440_),
    .S1(net178),
    .X(_4036_));
 sg13g2_mux4_1 _8796_ (.S0(net220),
    .A0(_0437_),
    .A1(_0438_),
    .A2(_0435_),
    .A3(_0436_),
    .S1(net178),
    .X(_4037_));
 sg13g2_mux2_1 _8797_ (.A0(_4036_),
    .A1(_4037_),
    .S(net105),
    .X(_4038_));
 sg13g2_o21ai_1 _8798_ (.B1(_3892_),
    .Y(_4039_),
    .A1(_3794_),
    .A2(_4038_));
 sg13g2_nor4_1 _8799_ (.A(_4025_),
    .B(_4029_),
    .C(_4035_),
    .D(_4039_),
    .Y(_4040_));
 sg13g2_mux2_1 _8800_ (.A0(_0393_),
    .A1(_0391_),
    .S(net219),
    .X(_4041_));
 sg13g2_mux2_1 _8801_ (.A0(_0394_),
    .A1(_0392_),
    .S(net222),
    .X(_4042_));
 sg13g2_mux2_1 _8802_ (.A0(_0389_),
    .A1(_0387_),
    .S(net219),
    .X(_4043_));
 sg13g2_mux2_1 _8803_ (.A0(_0390_),
    .A1(_0388_),
    .S(net219),
    .X(_4044_));
 sg13g2_mux4_1 _8804_ (.S0(net183),
    .A0(_4041_),
    .A1(_4042_),
    .A2(_4043_),
    .A3(_4044_),
    .S1(net105),
    .X(_4045_));
 sg13g2_o21ai_1 _8805_ (.B1(_3868_),
    .Y(_4046_),
    .A1(_3843_),
    .A2(_4045_));
 sg13g2_mux4_1 _8806_ (.S0(net174),
    .A0(_0401_),
    .A1(_0402_),
    .A2(_0399_),
    .A3(_0400_),
    .S1(net175),
    .X(_4047_));
 sg13g2_mux4_1 _8807_ (.S0(net218),
    .A0(_0397_),
    .A1(_0398_),
    .A2(_0395_),
    .A3(_0396_),
    .S1(net175),
    .X(_4048_));
 sg13g2_mux2_1 _8808_ (.A0(_4047_),
    .A1(_4048_),
    .S(net111),
    .X(_4049_));
 sg13g2_nor2_1 _8809_ (.A(_3828_),
    .B(_4049_),
    .Y(_4050_));
 sg13g2_mux4_1 _8810_ (.S0(net174),
    .A0(_0385_),
    .A1(_0386_),
    .A2(_0383_),
    .A3(_0384_),
    .S1(net180),
    .X(_4051_));
 sg13g2_mux4_1 _8811_ (.S0(net174),
    .A0(_0381_),
    .A1(_0382_),
    .A2(_0379_),
    .A3(_0380_),
    .S1(net180),
    .X(_4052_));
 sg13g2_mux2_1 _8812_ (.A0(_4051_),
    .A1(_4052_),
    .S(net111),
    .X(_4053_));
 sg13g2_nor2_1 _8813_ (.A(net72),
    .B(_4053_),
    .Y(_4054_));
 sg13g2_buf_2 _8814_ (.A(_3756_),
    .X(_4055_));
 sg13g2_mux4_1 _8815_ (.S0(net172),
    .A0(_0377_),
    .A1(_0378_),
    .A2(_0375_),
    .A3(_0376_),
    .S1(net187),
    .X(_4056_));
 sg13g2_mux4_1 _8816_ (.S0(net172),
    .A0(_0373_),
    .A1(_0374_),
    .A2(_0371_),
    .A3(_0372_),
    .S1(net187),
    .X(_4057_));
 sg13g2_mux2_1 _8817_ (.A0(_4056_),
    .A1(_4057_),
    .S(net104),
    .X(_4058_));
 sg13g2_nor2_1 _8818_ (.A(net71),
    .B(_4058_),
    .Y(_4059_));
 sg13g2_nor4_1 _8819_ (.A(_4046_),
    .B(_4050_),
    .C(_4054_),
    .D(_4059_),
    .Y(_4060_));
 sg13g2_mux2_1 _8820_ (.A0(_0545_),
    .A1(_0543_),
    .S(net222),
    .X(_4061_));
 sg13g2_mux2_1 _8821_ (.A0(_0546_),
    .A1(_0544_),
    .S(net222),
    .X(_4062_));
 sg13g2_mux2_1 _8822_ (.A0(_0541_),
    .A1(_0539_),
    .S(net222),
    .X(_4063_));
 sg13g2_mux2_1 _8823_ (.A0(_0542_),
    .A1(_0540_),
    .S(net222),
    .X(_4064_));
 sg13g2_mux4_1 _8824_ (.S0(net177),
    .A0(_4061_),
    .A1(_4062_),
    .A2(_4063_),
    .A3(_4064_),
    .S1(net111),
    .X(_4065_));
 sg13g2_o21ai_1 _8825_ (.B1(_3987_),
    .Y(_4066_),
    .A1(_3742_),
    .A2(_4065_));
 sg13g2_mux4_1 _8826_ (.S0(net172),
    .A0(_0537_),
    .A1(_0538_),
    .A2(_0535_),
    .A3(_0536_),
    .S1(net187),
    .X(_4067_));
 sg13g2_mux4_1 _8827_ (.S0(net172),
    .A0(_0533_),
    .A1(_0534_),
    .A2(_0531_),
    .A3(_0532_),
    .S1(net180),
    .X(_4068_));
 sg13g2_mux2_1 _8828_ (.A0(_4067_),
    .A1(_4068_),
    .S(_3790_),
    .X(_4069_));
 sg13g2_nor2_1 _8829_ (.A(_3795_),
    .B(_4069_),
    .Y(_4070_));
 sg13g2_mux4_1 _8830_ (.S0(_4055_),
    .A0(_0561_),
    .A1(_0562_),
    .A2(_0559_),
    .A3(_0560_),
    .S1(_3768_),
    .X(_4071_));
 sg13g2_mux4_1 _8831_ (.S0(_4055_),
    .A0(_0557_),
    .A1(_0558_),
    .A2(_0555_),
    .A3(_0556_),
    .S1(_3768_),
    .X(_4072_));
 sg13g2_mux2_1 _8832_ (.A0(_4071_),
    .A1(_4072_),
    .S(_3959_),
    .X(_4073_));
 sg13g2_nor2_1 _8833_ (.A(net70),
    .B(_4073_),
    .Y(_4074_));
 sg13g2_mux4_1 _8834_ (.S0(net184),
    .A0(_0553_),
    .A1(_0554_),
    .A2(_0551_),
    .A3(_0552_),
    .S1(net185),
    .X(_4075_));
 sg13g2_mux4_1 _8835_ (.S0(net184),
    .A0(_0549_),
    .A1(_0550_),
    .A2(_0547_),
    .A3(_0548_),
    .S1(net185),
    .X(_4076_));
 sg13g2_mux2_1 _8836_ (.A0(_4075_),
    .A1(_4076_),
    .S(net110),
    .X(_4077_));
 sg13g2_nor2_1 _8837_ (.A(net69),
    .B(_4077_),
    .Y(_4078_));
 sg13g2_nor4_1 _8838_ (.A(_4066_),
    .B(_4070_),
    .C(_4074_),
    .D(_4078_),
    .Y(_4079_));
 sg13g2_nor4_1 _8839_ (.A(_4021_),
    .B(_4040_),
    .C(_4060_),
    .D(_4079_),
    .Y(_4080_));
 sg13g2_mux4_1 _8840_ (.S0(net188),
    .A0(_0409_),
    .A1(_0410_),
    .A2(_0407_),
    .A3(_0408_),
    .S1(net173),
    .X(_4081_));
 sg13g2_mux4_1 _8841_ (.S0(net188),
    .A0(_0405_),
    .A1(_0406_),
    .A2(_0403_),
    .A3(_0404_),
    .S1(net173),
    .X(_4082_));
 sg13g2_mux2_1 _8842_ (.A0(_4081_),
    .A1(_4082_),
    .S(net104),
    .X(_4083_));
 sg13g2_nor2_1 _8843_ (.A(net71),
    .B(_4083_),
    .Y(_4084_));
 sg13g2_mux4_1 _8844_ (.S0(net184),
    .A0(_0417_),
    .A1(_0418_),
    .A2(_0415_),
    .A3(_0416_),
    .S1(net185),
    .X(_4085_));
 sg13g2_mux4_1 _8845_ (.S0(net184),
    .A0(_0413_),
    .A1(_0414_),
    .A2(_0411_),
    .A3(_0412_),
    .S1(net173),
    .X(_4086_));
 sg13g2_mux2_1 _8846_ (.A0(_4085_),
    .A1(_4086_),
    .S(net110),
    .X(_4087_));
 sg13g2_nor2_1 _8847_ (.A(net72),
    .B(_4087_),
    .Y(_4088_));
 sg13g2_mux4_1 _8848_ (.S0(net184),
    .A0(_0433_),
    .A1(_0434_),
    .A2(_0431_),
    .A3(_0432_),
    .S1(net185),
    .X(_4089_));
 sg13g2_mux4_1 _8849_ (.S0(net184),
    .A0(_0429_),
    .A1(_0430_),
    .A2(_0427_),
    .A3(_0428_),
    .S1(net185),
    .X(_4090_));
 sg13g2_mux2_1 _8850_ (.A0(_4089_),
    .A1(_4090_),
    .S(net110),
    .X(_4091_));
 sg13g2_nor2_1 _8851_ (.A(net70),
    .B(_4091_),
    .Y(_4092_));
 sg13g2_mux4_1 _8852_ (.S0(net188),
    .A0(_0425_),
    .A1(_0426_),
    .A2(_0423_),
    .A3(_0424_),
    .S1(net173),
    .X(_4093_));
 sg13g2_mux4_1 _8853_ (.S0(net188),
    .A0(_0421_),
    .A1(_0422_),
    .A2(_0419_),
    .A3(_0420_),
    .S1(net173),
    .X(_4094_));
 sg13g2_mux2_1 _8854_ (.A0(_4093_),
    .A1(_4094_),
    .S(net104),
    .X(_4095_));
 sg13g2_o21ai_1 _8855_ (.B1(_3970_),
    .Y(_4096_),
    .A1(net69),
    .A2(_4095_));
 sg13g2_nor4_1 _8856_ (.A(_4084_),
    .B(_4088_),
    .C(_4092_),
    .D(_4096_),
    .Y(_4097_));
 sg13g2_mux2_1 _8857_ (.A0(_0497_),
    .A1(_0495_),
    .S(net181),
    .X(_4098_));
 sg13g2_mux2_1 _8858_ (.A0(_0498_),
    .A1(_0496_),
    .S(net181),
    .X(_4099_));
 sg13g2_mux2_1 _8859_ (.A0(_0493_),
    .A1(_0491_),
    .S(net181),
    .X(_4100_));
 sg13g2_mux2_1 _8860_ (.A0(_0494_),
    .A1(_0492_),
    .S(net181),
    .X(_4101_));
 sg13g2_mux4_1 _8861_ (.S0(net113),
    .A0(_4098_),
    .A1(_4099_),
    .A2(_4100_),
    .A3(_4101_),
    .S1(net110),
    .X(_4102_));
 sg13g2_o21ai_1 _8862_ (.B1(_3824_),
    .Y(_4103_),
    .A1(net70),
    .A2(_4102_));
 sg13g2_mux4_1 _8863_ (.S0(net174),
    .A0(_0473_),
    .A1(_0474_),
    .A2(_0471_),
    .A3(_0472_),
    .S1(net180),
    .X(_4104_));
 sg13g2_mux4_1 _8864_ (.S0(net172),
    .A0(_0469_),
    .A1(_0470_),
    .A2(_0467_),
    .A3(_0468_),
    .S1(net180),
    .X(_4105_));
 sg13g2_mux4_1 _8865_ (.S0(net174),
    .A0(_0481_),
    .A1(_0482_),
    .A2(_0479_),
    .A3(_0480_),
    .S1(net175),
    .X(_4106_));
 sg13g2_mux4_1 _8866_ (.S0(net174),
    .A0(_0477_),
    .A1(_0478_),
    .A2(_0475_),
    .A3(_0476_),
    .S1(net180),
    .X(_4107_));
 sg13g2_mux4_1 _8867_ (.S0(net111),
    .A0(_4104_),
    .A1(_4105_),
    .A2(_4106_),
    .A3(_4107_),
    .S1(_3740_),
    .X(_4108_));
 sg13g2_nor2_1 _8868_ (.A(_3826_),
    .B(_4108_),
    .Y(_4109_));
 sg13g2_mux4_1 _8869_ (.S0(net186),
    .A0(_0489_),
    .A1(_0490_),
    .A2(_0487_),
    .A3(_0488_),
    .S1(net108),
    .X(_4110_));
 sg13g2_mux4_1 _8870_ (.S0(net186),
    .A0(_0485_),
    .A1(_0486_),
    .A2(_0483_),
    .A3(_0484_),
    .S1(net108),
    .X(_4111_));
 sg13g2_mux2_1 _8871_ (.A0(_4110_),
    .A1(_4111_),
    .S(net110),
    .X(_4112_));
 sg13g2_nor2_1 _8872_ (.A(net69),
    .B(_4112_),
    .Y(_4113_));
 sg13g2_nor3_1 _8873_ (.A(_4103_),
    .B(_4109_),
    .C(_4113_),
    .Y(_4114_));
 sg13g2_nor2_1 _8874_ (.A(_4097_),
    .B(_4114_),
    .Y(_4115_));
 sg13g2_mux4_1 _8875_ (.S0(_3757_),
    .A0(_0585_),
    .A1(_0586_),
    .A2(_0583_),
    .A3(_0584_),
    .S1(_3989_),
    .X(_4116_));
 sg13g2_mux4_1 _8876_ (.S0(_3757_),
    .A0(_0581_),
    .A1(_0582_),
    .A2(_0579_),
    .A3(_0580_),
    .S1(_3989_),
    .X(_4117_));
 sg13g2_mux2_1 _8877_ (.A0(_4116_),
    .A1(_4117_),
    .S(net104),
    .X(_4118_));
 sg13g2_nor2_1 _8878_ (.A(net69),
    .B(_4118_),
    .Y(_4119_));
 sg13g2_mux4_1 _8879_ (.S0(_3972_),
    .A0(_0577_),
    .A1(_0578_),
    .A2(_0575_),
    .A3(_0576_),
    .S1(_3950_),
    .X(_4120_));
 sg13g2_mux4_1 _8880_ (.S0(_3972_),
    .A0(_0573_),
    .A1(_0574_),
    .A2(_0571_),
    .A3(_0572_),
    .S1(_3950_),
    .X(_4121_));
 sg13g2_mux2_1 _8881_ (.A0(_4120_),
    .A1(_4121_),
    .S(_3790_),
    .X(_4122_));
 sg13g2_o21ai_1 _8882_ (.B1(_3948_),
    .Y(_4123_),
    .A1(net72),
    .A2(_4122_));
 sg13g2_mux4_1 _8883_ (.S0(_3800_),
    .A0(_0593_),
    .A1(_0594_),
    .A2(_0591_),
    .A3(_0592_),
    .S1(_3798_),
    .X(_4124_));
 sg13g2_mux4_1 _8884_ (.S0(_3800_),
    .A0(_0589_),
    .A1(_0590_),
    .A2(_0587_),
    .A3(_0588_),
    .S1(_3798_),
    .X(_4125_));
 sg13g2_mux2_1 _8885_ (.A0(_4124_),
    .A1(_4125_),
    .S(_3802_),
    .X(_4126_));
 sg13g2_nor2_1 _8886_ (.A(net70),
    .B(_4126_),
    .Y(_4127_));
 sg13g2_mux4_1 _8887_ (.S0(_3796_),
    .A0(_0569_),
    .A1(_0570_),
    .A2(_0567_),
    .A3(_0568_),
    .S1(_3837_),
    .X(_4128_));
 sg13g2_mux4_1 _8888_ (.S0(_3796_),
    .A0(_0565_),
    .A1(_0566_),
    .A2(_0563_),
    .A3(_0564_),
    .S1(_3837_),
    .X(_4129_));
 sg13g2_mux2_1 _8889_ (.A0(_4128_),
    .A1(_4129_),
    .S(_3802_),
    .X(_4130_));
 sg13g2_nor2_1 _8890_ (.A(_3795_),
    .B(_4130_),
    .Y(_4131_));
 sg13g2_nor4_1 _8891_ (.A(_4119_),
    .B(_4123_),
    .C(_4127_),
    .D(_4131_),
    .Y(_4132_));
 sg13g2_mux4_1 _8892_ (.S0(net184),
    .A0(_0353_),
    .A1(_0354_),
    .A2(_0351_),
    .A3(_0352_),
    .S1(net185),
    .X(_4133_));
 sg13g2_mux4_1 _8893_ (.S0(net188),
    .A0(_0349_),
    .A1(_0350_),
    .A2(_0347_),
    .A3(_0348_),
    .S1(net173),
    .X(_4134_));
 sg13g2_mux2_1 _8894_ (.A0(_4133_),
    .A1(_4134_),
    .S(net104),
    .X(_4135_));
 sg13g2_o21ai_1 _8895_ (.B1(_3914_),
    .Y(_4136_),
    .A1(net72),
    .A2(_4135_));
 sg13g2_mux4_1 _8896_ (.S0(net186),
    .A0(_0345_),
    .A1(_0346_),
    .A2(_0343_),
    .A3(_0344_),
    .S1(net108),
    .X(_4137_));
 sg13g2_mux4_1 _8897_ (.S0(net186),
    .A0(_0341_),
    .A1(_0342_),
    .A2(_0339_),
    .A3(_0340_),
    .S1(net108),
    .X(_4138_));
 sg13g2_mux2_1 _8898_ (.A0(_4137_),
    .A1(_4138_),
    .S(net110),
    .X(_4139_));
 sg13g2_nor2_1 _8899_ (.A(net71),
    .B(_4139_),
    .Y(_4140_));
 sg13g2_mux4_1 _8900_ (.S0(net172),
    .A0(_0361_),
    .A1(_0362_),
    .A2(_0359_),
    .A3(_0360_),
    .S1(net187),
    .X(_4141_));
 sg13g2_mux4_1 _8901_ (.S0(net172),
    .A0(_0369_),
    .A1(_0370_),
    .A2(_0367_),
    .A3(_0368_),
    .S1(net187),
    .X(_4142_));
 sg13g2_mux4_1 _8902_ (.S0(net174),
    .A0(_0357_),
    .A1(_0358_),
    .A2(_0355_),
    .A3(_0356_),
    .S1(net180),
    .X(_4143_));
 sg13g2_mux4_1 _8903_ (.S0(net172),
    .A0(_0365_),
    .A1(_0366_),
    .A2(_0363_),
    .A3(_0364_),
    .S1(net180),
    .X(_4144_));
 sg13g2_mux4_1 _8904_ (.S0(_3740_),
    .A0(_4141_),
    .A1(_4142_),
    .A2(_4143_),
    .A3(_4144_),
    .S1(net107),
    .X(_4145_));
 sg13g2_nor2_1 _8905_ (.A(_3722_),
    .B(_4145_),
    .Y(_4146_));
 sg13g2_nor3_1 _8906_ (.A(_4136_),
    .B(_4140_),
    .C(_4146_),
    .Y(_4147_));
 sg13g2_nor2_1 _8907_ (.A(_4132_),
    .B(_4147_),
    .Y(_4148_));
 sg13g2_and4_1 _8908_ (.A(_3938_),
    .B(_4080_),
    .C(_4115_),
    .D(_4148_),
    .X(_4149_));
 sg13g2_a21oi_1 _8909_ (.A1(_3895_),
    .A2(_4002_),
    .Y(_4150_),
    .B1(_4149_));
 sg13g2_buf_2 _8910_ (.A(_4150_),
    .X(_4151_));
 sg13g2_o21ai_1 _8911_ (.B1(net371),
    .Y(_4152_),
    .A1(_2016_),
    .A2(_2020_));
 sg13g2_a21oi_1 _8912_ (.A1(net387),
    .A2(_4152_),
    .Y(_4153_),
    .B1(net374));
 sg13g2_a21oi_1 _8913_ (.A1(_3702_),
    .A2(_4151_),
    .Y(_4154_),
    .B1(_4153_));
 sg13g2_nand2_1 _8914_ (.Y(_4155_),
    .A(net380),
    .B(_3679_));
 sg13g2_or3_1 _8915_ (.A(\num_neighbors[0] ),
    .B(_4155_),
    .C(_4151_),
    .X(_4156_));
 sg13g2_o21ai_1 _8916_ (.B1(_4156_),
    .Y(_1679_),
    .A1(_3294_),
    .A2(_4154_));
 sg13g2_nand3_1 _8917_ (.B(_3506_),
    .C(_3702_),
    .A(\num_neighbors[0] ),
    .Y(_4157_));
 sg13g2_nand2_1 _8918_ (.Y(_4158_),
    .A(\num_neighbors[1] ),
    .B(_4153_));
 sg13g2_o21ai_1 _8919_ (.B1(_4158_),
    .Y(_4159_),
    .A1(_4151_),
    .A2(_4157_));
 sg13g2_nor2_1 _8920_ (.A(_3506_),
    .B(_4155_),
    .Y(_4160_));
 sg13g2_o21ai_1 _8921_ (.B1(_4160_),
    .Y(_4161_),
    .A1(_3294_),
    .A2(_4151_));
 sg13g2_nand2b_1 _8922_ (.Y(_1680_),
    .B(_4161_),
    .A_N(_4159_));
 sg13g2_nand2_1 _8923_ (.Y(_4162_),
    .A(\num_neighbors[0] ),
    .B(\num_neighbors[1] ));
 sg13g2_or4_1 _8924_ (.A(_3507_),
    .B(_4155_),
    .C(_4151_),
    .D(_4162_),
    .X(_4163_));
 sg13g2_and2_1 _8925_ (.A(_3507_),
    .B(_3702_),
    .X(_4164_));
 sg13g2_o21ai_1 _8926_ (.B1(_4164_),
    .Y(_4165_),
    .A1(_4151_),
    .A2(_4162_));
 sg13g2_nand2_1 _8927_ (.Y(_4166_),
    .A(_3507_),
    .B(_4153_));
 sg13g2_nand3_1 _8928_ (.B(_4165_),
    .C(_4166_),
    .A(_4163_),
    .Y(_1681_));
 sg13g2_and3_1 _8929_ (.X(_4167_),
    .A(net372),
    .B(\num_neighbors[3] ),
    .C(_2022_));
 sg13g2_nand2_1 _8930_ (.Y(_4168_),
    .A(net372),
    .B(_2022_));
 sg13g2_nor2_1 _8931_ (.A(\num_neighbors[3] ),
    .B(_4168_),
    .Y(_4169_));
 sg13g2_nand3_1 _8932_ (.B(_3507_),
    .C(_4152_),
    .A(net387),
    .Y(_4170_));
 sg13g2_nor3_1 _8933_ (.A(_4151_),
    .B(_4162_),
    .C(_4170_),
    .Y(_4171_));
 sg13g2_mux2_1 _8934_ (.A0(_4167_),
    .A1(_4169_),
    .S(_4171_),
    .X(_1682_));
 sg13g2_inv_1 _8935_ (.Y(_4172_),
    .A(_1935_));
 sg13g2_nand2_1 _8936_ (.Y(_4173_),
    .A(_1980_),
    .B(_1979_));
 sg13g2_nor4_1 _8937_ (.A(_4172_),
    .B(_1936_),
    .C(_2060_),
    .D(_4173_),
    .Y(_4174_));
 sg13g2_o21ai_1 _8938_ (.B1(_4172_),
    .Y(_4175_),
    .A1(_1936_),
    .A2(net2));
 sg13g2_nand2b_1 _8939_ (.Y(_4176_),
    .B(_4175_),
    .A_N(_4174_));
 sg13g2_and2_1 _8940_ (.A(_2060_),
    .B(_2058_),
    .X(_4177_));
 sg13g2_o21ai_1 _8941_ (.B1(_1935_),
    .Y(_4178_),
    .A1(_4173_),
    .A2(_4177_));
 sg13g2_nand2_1 _8942_ (.Y(_4179_),
    .A(_1933_),
    .B(_4178_));
 sg13g2_a22oi_1 _8943_ (.Y(_4180_),
    .B1(_4179_),
    .B2(_1936_),
    .A2(_4176_),
    .A1(_1933_));
 sg13g2_nor2_1 _8944_ (.A(_3632_),
    .B(_4180_),
    .Y(_1683_));
 sg13g2_buf_1 _8945_ (.A(net330),
    .X(_4181_));
 sg13g2_nor2b_1 _8946_ (.A(net2),
    .B_N(_2057_),
    .Y(_4182_));
 sg13g2_and3_1 _8947_ (.X(_4183_),
    .A(_1979_),
    .B(_1982_),
    .C(_2084_));
 sg13g2_a21oi_1 _8948_ (.A1(_4172_),
    .A2(_4182_),
    .Y(_4184_),
    .B1(_4183_));
 sg13g2_nor2b_1 _8949_ (.A(_4179_),
    .B_N(_4184_),
    .Y(_4185_));
 sg13g2_buf_1 _8950_ (.A(_4185_),
    .X(_4186_));
 sg13g2_nand2_1 _8951_ (.Y(_4187_),
    .A(_1974_),
    .B(_1981_));
 sg13g2_nor2_1 _8952_ (.A(_2057_),
    .B(_4187_),
    .Y(_4188_));
 sg13g2_nand2_1 _8953_ (.Y(_4189_),
    .A(net216),
    .B(_4188_));
 sg13g2_mux2_1 _8954_ (.A0(_4189_),
    .A1(_4186_),
    .S(_1964_),
    .X(_4190_));
 sg13g2_nor2_1 _8955_ (.A(_4181_),
    .B(_4190_),
    .Y(_1684_));
 sg13g2_o21ai_1 _8956_ (.B1(net216),
    .Y(_4191_),
    .A1(_2057_),
    .A2(_4187_));
 sg13g2_nand2_1 _8957_ (.Y(_4192_),
    .A(_1796_),
    .B(_4191_));
 sg13g2_buf_1 _8958_ (.A(_4192_),
    .X(_4193_));
 sg13g2_buf_1 _8959_ (.A(_4193_),
    .X(_4194_));
 sg13g2_and4_1 _8960_ (.A(_1957_),
    .B(_1962_),
    .C(_1963_),
    .D(_1964_),
    .X(_4195_));
 sg13g2_nand3_1 _8961_ (.B(_1960_),
    .C(_4195_),
    .A(\timer[5] ),
    .Y(_4196_));
 sg13g2_inv_1 _8962_ (.Y(_4197_),
    .A(_4196_));
 sg13g2_nand4_1 _8963_ (.B(_4178_),
    .C(_4184_),
    .A(_1933_),
    .Y(_4198_),
    .D(_4197_));
 sg13g2_buf_2 _8964_ (.A(_4198_),
    .X(_4199_));
 sg13g2_nand3_1 _8965_ (.B(_1959_),
    .C(\timer[6] ),
    .A(\timer[8] ),
    .Y(_4200_));
 sg13g2_buf_1 _8966_ (.A(_4200_),
    .X(_4201_));
 sg13g2_nor2_2 _8967_ (.A(_4199_),
    .B(_4201_),
    .Y(_4202_));
 sg13g2_nand2_1 _8968_ (.Y(_4203_),
    .A(_1953_),
    .B(_4202_));
 sg13g2_xor2_1 _8969_ (.B(_4203_),
    .A(_1943_),
    .X(_4204_));
 sg13g2_nor2_1 _8970_ (.A(net68),
    .B(_4204_),
    .Y(_1685_));
 sg13g2_nand3_1 _8971_ (.B(_1953_),
    .C(_4202_),
    .A(_1943_),
    .Y(_4205_));
 sg13g2_xor2_1 _8972_ (.B(_4205_),
    .A(\timer[11] ),
    .X(_4206_));
 sg13g2_nor2_1 _8973_ (.A(net68),
    .B(_4206_),
    .Y(_1686_));
 sg13g2_inv_1 _8974_ (.Y(_4207_),
    .A(\timer[12] ));
 sg13g2_nand4_1 _8975_ (.B(_1943_),
    .C(_1953_),
    .A(\timer[11] ),
    .Y(_4208_),
    .D(_4202_));
 sg13g2_xnor2_1 _8976_ (.Y(_4209_),
    .A(_4207_),
    .B(_4208_));
 sg13g2_nor2_1 _8977_ (.A(net68),
    .B(_4209_),
    .Y(_1687_));
 sg13g2_or2_1 _8978_ (.X(_4210_),
    .B(_4208_),
    .A(_4207_));
 sg13g2_xor2_1 _8979_ (.B(_4210_),
    .A(\timer[13] ),
    .X(_4211_));
 sg13g2_nor2_1 _8980_ (.A(net68),
    .B(_4211_),
    .Y(_1688_));
 sg13g2_nand2_1 _8981_ (.Y(_4212_),
    .A(_1955_),
    .B(_4202_));
 sg13g2_xor2_1 _8982_ (.B(_4212_),
    .A(_1942_),
    .X(_4213_));
 sg13g2_nor2_1 _8983_ (.A(_4194_),
    .B(_4213_),
    .Y(_1689_));
 sg13g2_nand3_1 _8984_ (.B(_1955_),
    .C(_4202_),
    .A(_1942_),
    .Y(_4214_));
 sg13g2_xor2_1 _8985_ (.B(_4214_),
    .A(_1941_),
    .X(_4215_));
 sg13g2_nor2_1 _8986_ (.A(_4194_),
    .B(_4215_),
    .Y(_1690_));
 sg13g2_inv_1 _8987_ (.Y(_4216_),
    .A(_4201_));
 sg13g2_and4_1 _8988_ (.A(_1941_),
    .B(_1942_),
    .C(_1955_),
    .D(_4216_),
    .X(_4217_));
 sg13g2_nor2b_1 _8989_ (.A(_4199_),
    .B_N(_4217_),
    .Y(_4218_));
 sg13g2_xnor2_1 _8990_ (.Y(_4219_),
    .A(\timer[16] ),
    .B(_4218_));
 sg13g2_nor2_1 _8991_ (.A(net68),
    .B(_4219_),
    .Y(_1691_));
 sg13g2_nand2_1 _8992_ (.Y(_4220_),
    .A(\timer[16] ),
    .B(_4217_));
 sg13g2_nor2_1 _8993_ (.A(_4199_),
    .B(_4220_),
    .Y(_4221_));
 sg13g2_xnor2_1 _8994_ (.Y(_4222_),
    .A(_1947_),
    .B(_4221_));
 sg13g2_nor2_1 _8995_ (.A(net68),
    .B(_4222_),
    .Y(_1692_));
 sg13g2_inv_1 _8996_ (.Y(_4223_),
    .A(\timer[18] ));
 sg13g2_nand2_1 _8997_ (.Y(_4224_),
    .A(_1947_),
    .B(_4221_));
 sg13g2_xnor2_1 _8998_ (.Y(_4225_),
    .A(_4223_),
    .B(_4224_));
 sg13g2_nor2_1 _8999_ (.A(net68),
    .B(_4225_),
    .Y(_1693_));
 sg13g2_buf_1 _9000_ (.A(_4192_),
    .X(_4226_));
 sg13g2_inv_1 _9001_ (.Y(_4227_),
    .A(_1947_));
 sg13g2_nor4_2 _9002_ (.A(_4223_),
    .B(_4227_),
    .C(_4199_),
    .Y(_4228_),
    .D(_4220_));
 sg13g2_xnor2_1 _9003_ (.Y(_4229_),
    .A(_1939_),
    .B(_4228_));
 sg13g2_nor2_1 _9004_ (.A(net73),
    .B(_4229_),
    .Y(_1694_));
 sg13g2_nand2_1 _9005_ (.Y(_4230_),
    .A(_1964_),
    .B(_4186_));
 sg13g2_xor2_1 _9006_ (.B(_4230_),
    .A(_1963_),
    .X(_4231_));
 sg13g2_nor2_1 _9007_ (.A(net73),
    .B(_4231_),
    .Y(_1695_));
 sg13g2_nand2_1 _9008_ (.Y(_4232_),
    .A(_1939_),
    .B(_4228_));
 sg13g2_xor2_1 _9009_ (.B(_4232_),
    .A(_1950_),
    .X(_4233_));
 sg13g2_nor2_1 _9010_ (.A(net73),
    .B(_4233_),
    .Y(_1696_));
 sg13g2_nand3_1 _9011_ (.B(_1939_),
    .C(_4228_),
    .A(_1950_),
    .Y(_4234_));
 sg13g2_xor2_1 _9012_ (.B(_4234_),
    .A(\timer[21] ),
    .X(_4235_));
 sg13g2_nor2_1 _9013_ (.A(net73),
    .B(_4235_),
    .Y(_1697_));
 sg13g2_and4_1 _9014_ (.A(\timer[21] ),
    .B(_1950_),
    .C(_1939_),
    .D(_4228_),
    .X(_4236_));
 sg13g2_buf_8 _9015_ (.A(_4236_),
    .X(_4237_));
 sg13g2_nor2_1 _9016_ (.A(_1938_),
    .B(_4237_),
    .Y(_4238_));
 sg13g2_nor2_1 _9017_ (.A(net73),
    .B(_4238_),
    .Y(_1698_));
 sg13g2_a21oi_1 _9018_ (.A1(_1938_),
    .A2(_4237_),
    .Y(_4239_),
    .B1(_1966_));
 sg13g2_nor2_1 _9019_ (.A(net73),
    .B(_4239_),
    .Y(_1699_));
 sg13g2_inv_1 _9020_ (.Y(_4240_),
    .A(\timer[24] ));
 sg13g2_nand3_1 _9021_ (.B(_1938_),
    .C(_4237_),
    .A(_1966_),
    .Y(_4241_));
 sg13g2_a21oi_1 _9022_ (.A1(_4240_),
    .A2(_4241_),
    .Y(_1700_),
    .B1(_4193_));
 sg13g2_and4_1 _9023_ (.A(\timer[24] ),
    .B(_1966_),
    .C(_1938_),
    .D(_4237_),
    .X(_4242_));
 sg13g2_buf_8 _9024_ (.A(_4242_),
    .X(_4243_));
 sg13g2_nor2_1 _9025_ (.A(\timer[25] ),
    .B(_4243_),
    .Y(_4244_));
 sg13g2_nor2_1 _9026_ (.A(_4226_),
    .B(_4244_),
    .Y(_1701_));
 sg13g2_a21oi_1 _9027_ (.A1(\timer[25] ),
    .A2(_4243_),
    .Y(_4245_),
    .B1(\timer[26] ));
 sg13g2_nor2_1 _9028_ (.A(_4226_),
    .B(_4245_),
    .Y(_1702_));
 sg13g2_and3_1 _9029_ (.X(_4246_),
    .A(\timer[26] ),
    .B(\timer[25] ),
    .C(_4243_));
 sg13g2_nor2_1 _9030_ (.A(\timer[27] ),
    .B(_4246_),
    .Y(_4247_));
 sg13g2_nor2_1 _9031_ (.A(net73),
    .B(_4247_),
    .Y(_1703_));
 sg13g2_and2_1 _9032_ (.A(\timer[27] ),
    .B(_4246_),
    .X(_4248_));
 sg13g2_nor2_1 _9033_ (.A(\timer[28] ),
    .B(_4248_),
    .Y(_4249_));
 sg13g2_nor2_1 _9034_ (.A(net73),
    .B(_4249_),
    .Y(_1704_));
 sg13g2_and2_1 _9035_ (.A(\timer[28] ),
    .B(_4248_),
    .X(_4250_));
 sg13g2_buf_8 _9036_ (.A(_4250_),
    .X(_4251_));
 sg13g2_nor2_1 _9037_ (.A(\timer[29] ),
    .B(_4251_),
    .Y(_4252_));
 sg13g2_nor2_1 _9038_ (.A(net74),
    .B(_4252_),
    .Y(_1705_));
 sg13g2_nand3_1 _9039_ (.B(_1964_),
    .C(net216),
    .A(_1963_),
    .Y(_4253_));
 sg13g2_xor2_1 _9040_ (.B(_4253_),
    .A(_1962_),
    .X(_4254_));
 sg13g2_nor2_1 _9041_ (.A(net74),
    .B(_4254_),
    .Y(_1706_));
 sg13g2_a21o_1 _9042_ (.A2(_4251_),
    .A1(\timer[29] ),
    .B1(\timer[30] ),
    .X(_4255_));
 sg13g2_nor2b_1 _9043_ (.A(net68),
    .B_N(_4255_),
    .Y(_1707_));
 sg13g2_inv_1 _9044_ (.Y(_4256_),
    .A(\timer[31] ));
 sg13g2_nand3_1 _9045_ (.B(\timer[29] ),
    .C(_4251_),
    .A(\timer[30] ),
    .Y(_4257_));
 sg13g2_a21oi_1 _9046_ (.A1(_4256_),
    .A2(_4257_),
    .Y(_1708_),
    .B1(net74));
 sg13g2_nand4_1 _9047_ (.B(_1963_),
    .C(_1964_),
    .A(_1962_),
    .Y(_4258_),
    .D(net216));
 sg13g2_xor2_1 _9048_ (.B(_4258_),
    .A(_1957_),
    .X(_4259_));
 sg13g2_nor2_1 _9049_ (.A(net74),
    .B(_4259_),
    .Y(_1709_));
 sg13g2_nand4_1 _9050_ (.B(_1962_),
    .C(_1963_),
    .A(_1957_),
    .Y(_4260_),
    .D(_1964_));
 sg13g2_nand2_1 _9051_ (.Y(_4261_),
    .A(_4188_),
    .B(_4260_));
 sg13g2_inv_1 _9052_ (.Y(_4262_),
    .A(_1960_));
 sg13g2_a21oi_1 _9053_ (.A1(net216),
    .A2(_4261_),
    .Y(_4263_),
    .B1(_4262_));
 sg13g2_nor3_1 _9054_ (.A(_1960_),
    .B(_4189_),
    .C(_4260_),
    .Y(_4264_));
 sg13g2_o21ai_1 _9055_ (.B1(_2325_),
    .Y(_4265_),
    .A1(_4263_),
    .A2(_4264_));
 sg13g2_inv_1 _9056_ (.Y(_1710_),
    .A(_4265_));
 sg13g2_nand3_1 _9057_ (.B(net216),
    .C(_4195_),
    .A(_1960_),
    .Y(_4266_));
 sg13g2_xor2_1 _9058_ (.B(_4266_),
    .A(\timer[5] ),
    .X(_4267_));
 sg13g2_nor2_1 _9059_ (.A(net74),
    .B(_4267_),
    .Y(_1711_));
 sg13g2_inv_1 _9060_ (.Y(_4268_),
    .A(\timer[6] ));
 sg13g2_xnor2_1 _9061_ (.Y(_4269_),
    .A(_4268_),
    .B(_4199_));
 sg13g2_nor2_1 _9062_ (.A(net74),
    .B(_4269_),
    .Y(_1712_));
 sg13g2_nor2_1 _9063_ (.A(_4268_),
    .B(_4199_),
    .Y(_4270_));
 sg13g2_xnor2_1 _9064_ (.Y(_4271_),
    .A(_1959_),
    .B(_4270_));
 sg13g2_nor2_1 _9065_ (.A(net74),
    .B(_4271_),
    .Y(_1713_));
 sg13g2_nand2_1 _9066_ (.Y(_4272_),
    .A(_1959_),
    .B(_4270_));
 sg13g2_xor2_1 _9067_ (.B(_4272_),
    .A(\timer[8] ),
    .X(_4273_));
 sg13g2_nor2_1 _9068_ (.A(net74),
    .B(_4273_),
    .Y(_1714_));
 sg13g2_nand2b_1 _9069_ (.Y(_4274_),
    .B(_1953_),
    .A_N(net216));
 sg13g2_nor2_1 _9070_ (.A(_4196_),
    .B(_4201_),
    .Y(_4275_));
 sg13g2_xnor2_1 _9071_ (.Y(_4276_),
    .A(_0060_),
    .B(_4275_));
 sg13g2_nand3_1 _9072_ (.B(_4188_),
    .C(_4276_),
    .A(net216),
    .Y(_4277_));
 sg13g2_a21oi_1 _9073_ (.A1(_4274_),
    .A2(_4277_),
    .Y(_1715_),
    .B1(_2038_));
 sg13g2_a22oi_1 _9074_ (.Y(_4278_),
    .B1(_2172_),
    .B2(_2181_),
    .A2(_2167_),
    .A1(_1835_));
 sg13g2_nor2_1 _9075_ (.A(net264),
    .B(_4278_),
    .Y(_1716_));
 sg13g2_o21ai_1 _9076_ (.B1(_2183_),
    .Y(_4279_),
    .A1(_1835_),
    .A2(_2170_));
 sg13g2_a22oi_1 _9077_ (.Y(_4280_),
    .B1(_4279_),
    .B2(_1834_),
    .A2(_2172_),
    .A1(_1836_));
 sg13g2_nor2_1 _9078_ (.A(net264),
    .B(_4280_),
    .Y(_1717_));
 sg13g2_xnor2_1 _9079_ (.Y(_4281_),
    .A(_2193_),
    .B(_2174_));
 sg13g2_nor2_1 _9080_ (.A(_2167_),
    .B(_4281_),
    .Y(_4282_));
 sg13g2_a22oi_1 _9081_ (.Y(_4283_),
    .B1(_2177_),
    .B2(_4282_),
    .A2(_2167_),
    .A1(_1837_));
 sg13g2_nor2_1 _9082_ (.A(_4181_),
    .B(_4283_),
    .Y(_1718_));
 sg13g2_nand2b_1 _9083_ (.Y(_4284_),
    .B(_0067_),
    .A_N(net388));
 sg13g2_a21oi_1 _9084_ (.A1(_1870_),
    .A2(_1877_),
    .Y(_4285_),
    .B1(_1880_));
 sg13g2_nor2b_1 _9085_ (.A(_3600_),
    .B_N(_4285_),
    .Y(_4286_));
 sg13g2_buf_2 _9086_ (.A(_4286_),
    .X(_4287_));
 sg13g2_o21ai_1 _9087_ (.B1(_4287_),
    .Y(_4288_),
    .A1(_1870_),
    .A2(_4284_));
 sg13g2_buf_1 _9088_ (.A(_4288_),
    .X(_4289_));
 sg13g2_nor2_1 _9089_ (.A(_2067_),
    .B(_1882_),
    .Y(_4290_));
 sg13g2_a22oi_1 _9090_ (.Y(_4291_),
    .B1(_4290_),
    .B2(_4287_),
    .A2(_4289_),
    .A1(_1882_));
 sg13g2_nor2_1 _9091_ (.A(net264),
    .B(_4291_),
    .Y(_1722_));
 sg13g2_nand2b_1 _9092_ (.Y(_4292_),
    .B(_1882_),
    .A_N(_1881_));
 sg13g2_buf_1 _9093_ (.A(_4292_),
    .X(_4293_));
 sg13g2_nand2b_1 _9094_ (.Y(_4294_),
    .B(_1881_),
    .A_N(_1882_));
 sg13g2_o21ai_1 _9095_ (.B1(_4294_),
    .Y(_4295_),
    .A1(_4289_),
    .A2(_4293_));
 sg13g2_a22oi_1 _9096_ (.Y(_4296_),
    .B1(_4295_),
    .B2(net373),
    .A2(_4289_),
    .A1(_1881_));
 sg13g2_nor2_1 _9097_ (.A(net264),
    .B(_4296_),
    .Y(_1723_));
 sg13g2_buf_1 _9098_ (.A(\uart_rx_inst.bitIndex[2] ),
    .X(_4297_));
 sg13g2_nand2_1 _9099_ (.Y(_4298_),
    .A(net383),
    .B(_4289_));
 sg13g2_xor2_1 _9100_ (.B(_1883_),
    .A(_0059_),
    .X(_4299_));
 sg13g2_nand3_1 _9101_ (.B(_4287_),
    .C(_4299_),
    .A(_1871_),
    .Y(_4300_));
 sg13g2_a21oi_1 _9102_ (.A1(_4298_),
    .A2(_4300_),
    .Y(_1724_),
    .B1(net272));
 sg13g2_nand2_1 _9103_ (.Y(_4301_),
    .A(_2065_),
    .B(_4287_));
 sg13g2_buf_2 _9104_ (.A(_4301_),
    .X(_4302_));
 sg13g2_nor3_1 _9105_ (.A(_1881_),
    .B(_1882_),
    .C(net383),
    .Y(_4303_));
 sg13g2_nand2_1 _9106_ (.Y(_4304_),
    .A(_0595_),
    .B(_4303_));
 sg13g2_nand2_1 _9107_ (.Y(_4305_),
    .A(_1920_),
    .B(_1921_));
 sg13g2_o21ai_1 _9108_ (.B1(_1919_),
    .Y(_4306_),
    .A1(_1920_),
    .A2(_1921_));
 sg13g2_a21oi_2 _9109_ (.B1(_4302_),
    .Y(_4307_),
    .A2(_4306_),
    .A1(_4305_));
 sg13g2_a22oi_1 _9110_ (.Y(_4308_),
    .B1(_4307_),
    .B2(_4303_),
    .A2(_4304_),
    .A1(\uart_rx_inst.data[0] ));
 sg13g2_inv_1 _9111_ (.Y(_4309_),
    .A(_4308_));
 sg13g2_a22oi_1 _9112_ (.Y(_4310_),
    .B1(_4309_),
    .B2(_1871_),
    .A2(_4302_),
    .A1(\uart_rx_inst.data[0] ));
 sg13g2_nor2_1 _9113_ (.A(net264),
    .B(_4310_),
    .Y(_1725_));
 sg13g2_o21ai_1 _9114_ (.B1(_1870_),
    .Y(_4311_),
    .A1(net383),
    .A2(_4293_));
 sg13g2_nand3_1 _9115_ (.B(_4287_),
    .C(_4311_),
    .A(_2065_),
    .Y(_4312_));
 sg13g2_nor2_1 _9116_ (.A(_2067_),
    .B(_0595_),
    .Y(_4313_));
 sg13g2_and2_1 _9117_ (.A(_4307_),
    .B(_4313_),
    .X(_4314_));
 sg13g2_inv_1 _9118_ (.Y(_4315_),
    .A(_4314_));
 sg13g2_a21oi_1 _9119_ (.A1(_4294_),
    .A2(_4293_),
    .Y(_4316_),
    .B1(_4315_));
 sg13g2_inv_1 _9120_ (.Y(_4317_),
    .A(net383));
 sg13g2_a22oi_1 _9121_ (.Y(_4318_),
    .B1(_4316_),
    .B2(_4317_),
    .A2(_4312_),
    .A1(\uart_rx_inst.data[1] ));
 sg13g2_nor2_1 _9122_ (.A(net264),
    .B(_4318_),
    .Y(_1726_));
 sg13g2_inv_1 _9123_ (.Y(_4319_),
    .A(\uart_rx_inst.data[2] ));
 sg13g2_nor2_1 _9124_ (.A(net383),
    .B(_4294_),
    .Y(_4320_));
 sg13g2_nand2_1 _9125_ (.Y(_4321_),
    .A(_4307_),
    .B(_4320_));
 sg13g2_o21ai_1 _9126_ (.B1(_4321_),
    .Y(_4322_),
    .A1(_4319_),
    .A2(_4320_));
 sg13g2_a22oi_1 _9127_ (.Y(_4323_),
    .B1(_4322_),
    .B2(net373),
    .A2(_4302_),
    .A1(\uart_rx_inst.data[2] ));
 sg13g2_nor2_1 _9128_ (.A(net264),
    .B(_4323_),
    .Y(_1727_));
 sg13g2_o21ai_1 _9129_ (.B1(_1870_),
    .Y(_4324_),
    .A1(net383),
    .A2(_1883_));
 sg13g2_nand3_1 _9130_ (.B(_4287_),
    .C(_4324_),
    .A(_2065_),
    .Y(_4325_));
 sg13g2_or3_1 _9131_ (.A(_1881_),
    .B(_1882_),
    .C(_4317_),
    .X(_4326_));
 sg13g2_o21ai_1 _9132_ (.B1(_4326_),
    .Y(_4327_),
    .A1(net383),
    .A2(_1883_));
 sg13g2_a22oi_1 _9133_ (.Y(_4328_),
    .B1(_4327_),
    .B2(_4314_),
    .A2(_4325_),
    .A1(\uart_rx_inst.data[3] ));
 sg13g2_nor2_1 _9134_ (.A(net264),
    .B(_4328_),
    .Y(_1728_));
 sg13g2_buf_1 _9135_ (.A(net330),
    .X(_4329_));
 sg13g2_mux2_1 _9136_ (.A0(_4307_),
    .A1(\uart_rx_inst.data[4] ),
    .S(_4326_),
    .X(_4330_));
 sg13g2_a22oi_1 _9137_ (.Y(_4331_),
    .B1(_4330_),
    .B2(net373),
    .A2(_4302_),
    .A1(\uart_rx_inst.data[4] ));
 sg13g2_nor2_1 _9138_ (.A(net263),
    .B(_4331_),
    .Y(_1729_));
 sg13g2_o21ai_1 _9139_ (.B1(net373),
    .Y(_4332_),
    .A1(_4317_),
    .A2(_4293_));
 sg13g2_nand3_1 _9140_ (.B(_4287_),
    .C(_4332_),
    .A(net297),
    .Y(_4333_));
 sg13g2_a22oi_1 _9141_ (.Y(_4334_),
    .B1(_4333_),
    .B2(\uart_rx_inst.data[5] ),
    .A2(_4316_),
    .A1(net383));
 sg13g2_nor2_1 _9142_ (.A(net263),
    .B(_4334_),
    .Y(_1730_));
 sg13g2_nor2_1 _9143_ (.A(_4317_),
    .B(_4294_),
    .Y(_4335_));
 sg13g2_mux2_1 _9144_ (.A0(\uart_rx_inst.data[6] ),
    .A1(_4307_),
    .S(_4335_),
    .X(_4336_));
 sg13g2_a22oi_1 _9145_ (.Y(_4337_),
    .B1(_4336_),
    .B2(net373),
    .A2(_4302_),
    .A1(\uart_rx_inst.data[6] ));
 sg13g2_nor2_1 _9146_ (.A(net263),
    .B(_4337_),
    .Y(_1731_));
 sg13g2_nand3_1 _9147_ (.B(_1882_),
    .C(_4297_),
    .A(_1881_),
    .Y(_4338_));
 sg13g2_and2_1 _9148_ (.A(net373),
    .B(_4338_),
    .X(_4339_));
 sg13g2_o21ai_1 _9149_ (.B1(\uart_rx_inst.data[7] ),
    .Y(_4340_),
    .A1(_4302_),
    .A2(_4339_));
 sg13g2_or2_1 _9150_ (.X(_4341_),
    .B(_4338_),
    .A(_4315_));
 sg13g2_a21oi_1 _9151_ (.A1(_4340_),
    .A2(_4341_),
    .Y(_1732_),
    .B1(_2038_));
 sg13g2_nor2_1 _9152_ (.A(_1920_),
    .B(_1916_),
    .Y(_4342_));
 sg13g2_nor3_1 _9153_ (.A(net388),
    .B(net4),
    .C(net274),
    .Y(_4343_));
 sg13g2_o21ai_1 _9154_ (.B1(net329),
    .Y(_1733_),
    .A1(_4342_),
    .A2(_4343_));
 sg13g2_nor2_1 _9155_ (.A(_1919_),
    .B(_1916_),
    .Y(_4344_));
 sg13g2_nor3_1 _9156_ (.A(net388),
    .B(_1920_),
    .C(_1889_),
    .Y(_4345_));
 sg13g2_o21ai_1 _9157_ (.B1(_1913_),
    .Y(_1734_),
    .A1(_4344_),
    .A2(_4345_));
 sg13g2_nor2_1 _9158_ (.A(_1921_),
    .B(_1916_),
    .Y(_4346_));
 sg13g2_nor3_1 _9159_ (.A(_1914_),
    .B(_1919_),
    .C(net274),
    .Y(_4347_));
 sg13g2_o21ai_1 _9160_ (.B1(_1913_),
    .Y(_1735_),
    .A1(_4346_),
    .A2(_4347_));
 sg13g2_mux2_1 _9161_ (.A0(net388),
    .A1(_3604_),
    .S(_1917_),
    .X(_4348_));
 sg13g2_nand2_1 _9162_ (.Y(_4349_),
    .A(_1916_),
    .B(_4348_));
 sg13g2_buf_1 _9163_ (.A(_4349_),
    .X(_4350_));
 sg13g2_buf_1 _9164_ (.A(_4350_),
    .X(_4351_));
 sg13g2_inv_1 _9165_ (.Y(_4352_),
    .A(\uart_rx_inst.data[0] ));
 sg13g2_nor3_1 _9166_ (.A(net297),
    .B(_4352_),
    .C(net215),
    .Y(_4353_));
 sg13g2_a21oi_1 _9167_ (.A1(_1985_),
    .A2(net215),
    .Y(_4354_),
    .B1(_4353_));
 sg13g2_nor2_1 _9168_ (.A(net263),
    .B(_4354_),
    .Y(_1736_));
 sg13g2_inv_1 _9169_ (.Y(_4355_),
    .A(\uart_rx_inst.data[1] ));
 sg13g2_nor3_1 _9170_ (.A(net297),
    .B(_4355_),
    .C(net215),
    .Y(_4356_));
 sg13g2_a21oi_1 _9171_ (.A1(\uart_rx_data[1] ),
    .A2(net215),
    .Y(_4357_),
    .B1(_4356_));
 sg13g2_nor2_1 _9172_ (.A(net263),
    .B(_4357_),
    .Y(_1737_));
 sg13g2_nor3_1 _9173_ (.A(net297),
    .B(_4319_),
    .C(_4350_),
    .Y(_4358_));
 sg13g2_a21oi_1 _9174_ (.A1(\uart_rx_data[2] ),
    .A2(net215),
    .Y(_4359_),
    .B1(_4358_));
 sg13g2_nor2_1 _9175_ (.A(net263),
    .B(_4359_),
    .Y(_1738_));
 sg13g2_inv_1 _9176_ (.Y(_4360_),
    .A(\uart_rx_inst.data[3] ));
 sg13g2_nor3_1 _9177_ (.A(net297),
    .B(_4360_),
    .C(_4350_),
    .Y(_4361_));
 sg13g2_a21oi_1 _9178_ (.A1(\uart_rx_data[3] ),
    .A2(net215),
    .Y(_4362_),
    .B1(_4361_));
 sg13g2_nor2_1 _9179_ (.A(net263),
    .B(_4362_),
    .Y(_1739_));
 sg13g2_inv_1 _9180_ (.Y(_4363_),
    .A(\uart_rx_inst.data[4] ));
 sg13g2_nor3_1 _9181_ (.A(_3599_),
    .B(_4363_),
    .C(_4350_),
    .Y(_4364_));
 sg13g2_a21oi_1 _9182_ (.A1(_1986_),
    .A2(_4351_),
    .Y(_4365_),
    .B1(_4364_));
 sg13g2_nor2_1 _9183_ (.A(_4329_),
    .B(_4365_),
    .Y(_1740_));
 sg13g2_inv_1 _9184_ (.Y(_4366_),
    .A(\uart_rx_inst.data[5] ));
 sg13g2_nor3_1 _9185_ (.A(net297),
    .B(_4366_),
    .C(_4350_),
    .Y(_4367_));
 sg13g2_a21oi_1 _9186_ (.A1(\uart_rx_data[5] ),
    .A2(net215),
    .Y(_4368_),
    .B1(_4367_));
 sg13g2_nor2_1 _9187_ (.A(_4329_),
    .B(_4368_),
    .Y(_1741_));
 sg13g2_inv_1 _9188_ (.Y(_4369_),
    .A(\uart_rx_inst.data[6] ));
 sg13g2_nor3_1 _9189_ (.A(net297),
    .B(_4369_),
    .C(_4350_),
    .Y(_4370_));
 sg13g2_a21oi_1 _9190_ (.A1(\uart_rx_data[6] ),
    .A2(_4351_),
    .Y(_4371_),
    .B1(_4370_));
 sg13g2_nor2_1 _9191_ (.A(net263),
    .B(_4371_),
    .Y(_1742_));
 sg13g2_inv_1 _9192_ (.Y(_4372_),
    .A(\uart_rx_inst.data[7] ));
 sg13g2_nor3_1 _9193_ (.A(_3599_),
    .B(_4372_),
    .C(_4350_),
    .Y(_4373_));
 sg13g2_a21oi_1 _9194_ (.A1(\uart_rx_data[7] ),
    .A2(net215),
    .Y(_4374_),
    .B1(_4373_));
 sg13g2_nor2_1 _9195_ (.A(net273),
    .B(_4374_),
    .Y(_1743_));
 sg13g2_and3_1 _9196_ (.X(_1745_),
    .A(net322),
    .B(_0599_),
    .C(_1889_));
 sg13g2_xnor2_1 _9197_ (.Y(_4375_),
    .A(\uart_rx_inst.rxCounter[1] ),
    .B(\uart_rx_inst.rxCounter[0] ));
 sg13g2_nor3_1 _9198_ (.A(_2072_),
    .B(_1916_),
    .C(_4375_),
    .Y(_1746_));
 sg13g2_nand2b_1 _9199_ (.Y(_4376_),
    .B(_1878_),
    .A_N(\uart_rx_inst.rxCounter[3] ));
 sg13g2_nand2_1 _9200_ (.Y(_4377_),
    .A(\uart_rx_inst.rxCounter[1] ),
    .B(\uart_rx_inst.rxCounter[0] ));
 sg13g2_mux2_1 _9201_ (.A0(_1878_),
    .A1(_4376_),
    .S(_4377_),
    .X(_4378_));
 sg13g2_nor2_1 _9202_ (.A(net273),
    .B(_4378_),
    .Y(_1747_));
 sg13g2_nand2b_1 _9203_ (.Y(_4379_),
    .B(\uart_rx_inst.rxCounter[3] ),
    .A_N(_1878_));
 sg13g2_o21ai_1 _9204_ (.B1(_4379_),
    .Y(_4380_),
    .A1(_4377_),
    .A2(_4376_));
 sg13g2_and2_1 _9205_ (.A(net322),
    .B(_4380_),
    .X(_1748_));
 sg13g2_nor4_1 _9206_ (.A(_1872_),
    .B(_0067_),
    .C(_1927_),
    .D(_1925_),
    .Y(_4381_));
 sg13g2_nor4_1 _9207_ (.A(_1870_),
    .B(_1887_),
    .C(net388),
    .D(_1917_),
    .Y(_4382_));
 sg13g2_or3_1 _9208_ (.A(_1880_),
    .B(_4381_),
    .C(_4382_),
    .X(_4383_));
 sg13g2_buf_2 _9209_ (.A(_4383_),
    .X(_4384_));
 sg13g2_nor3_1 _9210_ (.A(_1870_),
    .B(_1917_),
    .C(_3600_),
    .Y(_4385_));
 sg13g2_nor3_1 _9211_ (.A(net389),
    .B(_4384_),
    .C(_4385_),
    .Y(_4386_));
 sg13g2_a21oi_1 _9212_ (.A1(net389),
    .A2(_4384_),
    .Y(_4387_),
    .B1(_4386_));
 sg13g2_nor2_1 _9213_ (.A(net273),
    .B(_4387_),
    .Y(_1749_));
 sg13g2_a21oi_1 _9214_ (.A1(_1917_),
    .A2(_2064_),
    .Y(_4388_),
    .B1(_1887_));
 sg13g2_a21oi_1 _9215_ (.A1(_0068_),
    .A2(_1886_),
    .Y(_4389_),
    .B1(_4388_));
 sg13g2_nor2_1 _9216_ (.A(net373),
    .B(_4389_),
    .Y(_4390_));
 sg13g2_inv_1 _9217_ (.Y(_4391_),
    .A(_4390_));
 sg13g2_nand2b_1 _9218_ (.Y(_4392_),
    .B(net389),
    .A_N(_1874_));
 sg13g2_nand2b_1 _9219_ (.Y(_4393_),
    .B(_1874_),
    .A_N(net389));
 sg13g2_o21ai_1 _9220_ (.B1(_4393_),
    .Y(_4394_),
    .A1(_4384_),
    .A2(_4392_));
 sg13g2_a22oi_1 _9221_ (.Y(_4395_),
    .B1(_4391_),
    .B2(_4394_),
    .A2(_4384_),
    .A1(_1874_));
 sg13g2_nor2_1 _9222_ (.A(net273),
    .B(_4395_),
    .Y(_1750_));
 sg13g2_nand2_1 _9223_ (.Y(_4396_),
    .A(_1874_),
    .B(_1875_));
 sg13g2_nor3_1 _9224_ (.A(_1873_),
    .B(_4396_),
    .C(_4384_),
    .Y(_4397_));
 sg13g2_a21o_1 _9225_ (.A2(_4396_),
    .A1(_1873_),
    .B1(_4397_),
    .X(_4398_));
 sg13g2_a22oi_1 _9226_ (.Y(_4399_),
    .B1(_4391_),
    .B2(_4398_),
    .A2(_4384_),
    .A1(_1873_));
 sg13g2_nor2_1 _9227_ (.A(net273),
    .B(_4399_),
    .Y(_1751_));
 sg13g2_o21ai_1 _9228_ (.B1(_2064_),
    .Y(_4400_),
    .A1(_1887_),
    .A2(_1917_));
 sg13g2_nand3_1 _9229_ (.B(_1874_),
    .C(net389),
    .A(_1873_),
    .Y(_4401_));
 sg13g2_nor3_1 _9230_ (.A(_1872_),
    .B(_4401_),
    .C(_4384_),
    .Y(_4402_));
 sg13g2_a21oi_1 _9231_ (.A1(_1872_),
    .A2(_4401_),
    .Y(_4403_),
    .B1(_4402_));
 sg13g2_a21oi_1 _9232_ (.A1(_2067_),
    .A2(_4400_),
    .Y(_4404_),
    .B1(_4403_));
 sg13g2_a21oi_1 _9233_ (.A1(_1872_),
    .A2(_4384_),
    .Y(_4405_),
    .B1(_4404_));
 sg13g2_nor2_1 _9234_ (.A(net273),
    .B(_4405_),
    .Y(_1752_));
 sg13g2_nor2_1 _9235_ (.A(_1980_),
    .B(_4172_),
    .Y(_4406_));
 sg13g2_o21ai_1 _9236_ (.B1(net274),
    .Y(_4407_),
    .A1(\uart_rx_inst.out_latched ),
    .A2(_4406_));
 sg13g2_nand3b_1 _9237_ (.B(_1935_),
    .C(_1916_),
    .Y(_4408_),
    .A_N(net388));
 sg13g2_a21oi_1 _9238_ (.A1(_4407_),
    .A2(_4408_),
    .Y(_1753_),
    .B1(net272));
 sg13g2_nor2b_1 _9239_ (.A(_2057_),
    .B_N(_1933_),
    .Y(_4409_));
 sg13g2_o21ai_1 _9240_ (.B1(_4409_),
    .Y(_4410_),
    .A1(_1937_),
    .A2(_4187_));
 sg13g2_a21oi_1 _9241_ (.A1(_4172_),
    .A2(_4410_),
    .Y(_4411_),
    .B1(_2332_));
 sg13g2_mux2_1 _9242_ (.A0(\action[0] ),
    .A1(_1935_),
    .S(_1933_),
    .X(_4412_));
 sg13g2_o21ai_1 _9243_ (.B1(_2325_),
    .Y(_4413_),
    .A1(_1980_),
    .A2(_4412_));
 sg13g2_a21oi_1 _9244_ (.A1(_1980_),
    .A2(_4411_),
    .Y(_1754_),
    .B1(_4413_));
 sg13g2_nor3_1 _9245_ (.A(_2040_),
    .B(_1906_),
    .C(_3505_),
    .Y(_4414_));
 sg13g2_nand2_1 _9246_ (.Y(_4415_),
    .A(net392),
    .B(net391));
 sg13g2_nand2_1 _9247_ (.Y(_4416_),
    .A(_2043_),
    .B(_4415_));
 sg13g2_nand2b_1 _9248_ (.Y(_4417_),
    .B(_2041_),
    .A_N(net392));
 sg13g2_nor2_1 _9249_ (.A(_2040_),
    .B(_1906_),
    .Y(_4418_));
 sg13g2_or4_1 _9250_ (.A(net391),
    .B(_0066_),
    .C(_4417_),
    .D(_4418_),
    .X(_4419_));
 sg13g2_nand2_1 _9251_ (.Y(_4420_),
    .A(_4416_),
    .B(_4419_));
 sg13g2_nor2_1 _9252_ (.A(_4414_),
    .B(_4420_),
    .Y(_4421_));
 sg13g2_nand2_1 _9253_ (.Y(_4422_),
    .A(net382),
    .B(_0046_));
 sg13g2_o21ai_1 _9254_ (.B1(_4422_),
    .Y(_4423_),
    .A1(_1790_),
    .A2(_4421_));
 sg13g2_o21ai_1 _9255_ (.B1(_3607_),
    .Y(_4424_),
    .A1(_1998_),
    .A2(_4418_));
 sg13g2_o21ai_1 _9256_ (.B1(_4424_),
    .Y(_4425_),
    .A1(_1909_),
    .A2(_2048_));
 sg13g2_nand2_2 _9257_ (.Y(_4426_),
    .A(net381),
    .B(_4425_));
 sg13g2_nand2_1 _9258_ (.Y(_4427_),
    .A(_1833_),
    .B(_1844_));
 sg13g2_a21oi_2 _9259_ (.B1(_1791_),
    .Y(_4428_),
    .A2(_4427_),
    .A1(net382));
 sg13g2_nand2_1 _9260_ (.Y(_4429_),
    .A(_4426_),
    .B(_4428_));
 sg13g2_buf_1 _9261_ (.A(_4429_),
    .X(_4430_));
 sg13g2_mux2_1 _9262_ (.A0(_4423_),
    .A1(\uart_tx_data[0] ),
    .S(net214),
    .X(_4431_));
 sg13g2_and2_1 _9263_ (.A(net322),
    .B(_4431_),
    .X(_1755_));
 sg13g2_inv_1 _9264_ (.Y(_4432_),
    .A(_0047_));
 sg13g2_a21oi_1 _9265_ (.A1(net328),
    .A2(_4432_),
    .Y(_4433_),
    .B1(net214));
 sg13g2_a21oi_1 _9266_ (.A1(\uart_tx_data[1] ),
    .A2(net214),
    .Y(_4434_),
    .B1(_4433_));
 sg13g2_nor3_2 _9267_ (.A(net382),
    .B(_4429_),
    .C(_4414_),
    .Y(_4435_));
 sg13g2_o21ai_1 _9268_ (.B1(_1906_),
    .Y(_4436_),
    .A1(net391),
    .A2(_4417_));
 sg13g2_and3_1 _9269_ (.X(_4437_),
    .A(_4416_),
    .B(_4435_),
    .C(_4436_));
 sg13g2_nor3_1 _9270_ (.A(net271),
    .B(_4434_),
    .C(_4437_),
    .Y(_1756_));
 sg13g2_nand2_1 _9271_ (.Y(_4438_),
    .A(\uart_tx_data[2] ),
    .B(net214));
 sg13g2_nand2b_1 _9272_ (.Y(_4439_),
    .B(net328),
    .A_N(_0048_));
 sg13g2_nand3_1 _9273_ (.B(_4428_),
    .C(_4439_),
    .A(_4426_),
    .Y(_4440_));
 sg13g2_a221oi_1 _9274_ (.B2(_4440_),
    .C1(net272),
    .B1(_4438_),
    .A1(_4419_),
    .Y(_1757_),
    .A2(_4435_));
 sg13g2_nand2_1 _9275_ (.Y(_4441_),
    .A(\uart_tx_data[3] ),
    .B(net214));
 sg13g2_nand2b_1 _9276_ (.Y(_4442_),
    .B(net328),
    .A_N(_0049_));
 sg13g2_nand3_1 _9277_ (.B(_4428_),
    .C(_4442_),
    .A(_4426_),
    .Y(_4443_));
 sg13g2_nor2_1 _9278_ (.A(_1906_),
    .B(_2043_),
    .Y(_4444_));
 sg13g2_a221oi_1 _9279_ (.B2(_4435_),
    .C1(net272),
    .B1(_4444_),
    .A1(_4441_),
    .Y(_1758_),
    .A2(_4443_));
 sg13g2_a21oi_1 _9280_ (.A1(_4426_),
    .A2(_4428_),
    .Y(_4445_),
    .B1(\uart_tx_data[4] ));
 sg13g2_nand2_1 _9281_ (.Y(_4446_),
    .A(net328),
    .B(_0050_));
 sg13g2_o21ai_1 _9282_ (.B1(_4446_),
    .Y(_4447_),
    .A1(net328),
    .A2(_4416_));
 sg13g2_nor2_1 _9283_ (.A(net214),
    .B(_4447_),
    .Y(_4448_));
 sg13g2_nor3_1 _9284_ (.A(net271),
    .B(_4445_),
    .C(_4448_),
    .Y(_1759_));
 sg13g2_inv_1 _9285_ (.Y(_4449_),
    .A(_0051_));
 sg13g2_a21oi_1 _9286_ (.A1(net328),
    .A2(_4449_),
    .Y(_4450_),
    .B1(_4430_));
 sg13g2_a21oi_1 _9287_ (.A1(\uart_tx_data[5] ),
    .A2(_4430_),
    .Y(_4451_),
    .B1(_4450_));
 sg13g2_nand2_1 _9288_ (.Y(_4452_),
    .A(net392),
    .B(_3642_));
 sg13g2_nor4_1 _9289_ (.A(net391),
    .B(_1908_),
    .C(_4418_),
    .D(_4452_),
    .Y(_4453_));
 sg13g2_and2_1 _9290_ (.A(_4418_),
    .B(_3505_),
    .X(_4454_));
 sg13g2_nor4_1 _9291_ (.A(_1994_),
    .B(net214),
    .C(_4453_),
    .D(_4454_),
    .Y(_4455_));
 sg13g2_nor3_1 _9292_ (.A(net271),
    .B(_4451_),
    .C(_4455_),
    .Y(_1760_));
 sg13g2_nand2_1 _9293_ (.Y(_4456_),
    .A(\uart_tx_data[6] ),
    .B(net214));
 sg13g2_nand2b_1 _9294_ (.Y(_4457_),
    .B(_1994_),
    .A_N(_0052_));
 sg13g2_nand3_1 _9295_ (.B(_4428_),
    .C(_4457_),
    .A(_4426_),
    .Y(_4458_));
 sg13g2_nand2_1 _9296_ (.Y(_4459_),
    .A(net391),
    .B(_2043_));
 sg13g2_a221oi_1 _9297_ (.B2(_4435_),
    .C1(net271),
    .B1(_4459_),
    .A1(_4456_),
    .Y(_1761_),
    .A2(_4458_));
 sg13g2_and2_1 _9298_ (.A(_1857_),
    .B(net262),
    .X(_4460_));
 sg13g2_o21ai_1 _9299_ (.B1(_4460_),
    .Y(_4461_),
    .A1(_1867_),
    .A2(_2070_));
 sg13g2_inv_1 _9300_ (.Y(_4462_),
    .A(_1867_));
 sg13g2_nand2_2 _9301_ (.Y(_4463_),
    .A(_1857_),
    .B(_1855_));
 sg13g2_nor3_1 _9302_ (.A(_4462_),
    .B(net390),
    .C(_4463_),
    .Y(_4464_));
 sg13g2_a21oi_1 _9303_ (.A1(net390),
    .A2(_4461_),
    .Y(_4465_),
    .B1(_4464_));
 sg13g2_nor2_1 _9304_ (.A(_2025_),
    .B(_4465_),
    .Y(_1762_));
 sg13g2_nand2b_1 _9305_ (.Y(_4466_),
    .B(net390),
    .A_N(_1862_));
 sg13g2_nand2b_1 _9306_ (.Y(_4467_),
    .B(_1862_),
    .A_N(_1863_));
 sg13g2_o21ai_1 _9307_ (.B1(_4467_),
    .Y(_4468_),
    .A1(_4463_),
    .A2(_4466_));
 sg13g2_a22oi_1 _9308_ (.Y(_4469_),
    .B1(_4468_),
    .B2(_1867_),
    .A2(_4461_),
    .A1(_1862_));
 sg13g2_nor2_1 _9309_ (.A(net273),
    .B(_4469_),
    .Y(_1763_));
 sg13g2_nor2_1 _9310_ (.A(_4462_),
    .B(_4463_),
    .Y(_4470_));
 sg13g2_xor2_1 _9311_ (.B(_1864_),
    .A(_0057_),
    .X(_4471_));
 sg13g2_a22oi_1 _9312_ (.Y(_4472_),
    .B1(_4470_),
    .B2(_4471_),
    .A2(_4461_),
    .A1(\uart_tx_inst.bitIndex[2] ));
 sg13g2_nor2_1 _9313_ (.A(_2025_),
    .B(_4472_),
    .Y(_1764_));
 sg13g2_a21oi_1 _9314_ (.A1(_2070_),
    .A2(net262),
    .Y(_4473_),
    .B1(_1858_));
 sg13g2_buf_2 _9315_ (.A(_4473_),
    .X(_4474_));
 sg13g2_a22oi_1 _9316_ (.Y(_4475_),
    .B1(_4474_),
    .B2(\uart_tx_inst.data[0] ),
    .A2(net261),
    .A1(\uart_tx_data[0] ));
 sg13g2_inv_1 _9317_ (.Y(_1765_),
    .A(_4475_));
 sg13g2_a22oi_1 _9318_ (.Y(_4476_),
    .B1(_4474_),
    .B2(\uart_tx_inst.data[1] ),
    .A2(net261),
    .A1(\uart_tx_data[1] ));
 sg13g2_inv_1 _9319_ (.Y(_1766_),
    .A(_4476_));
 sg13g2_a22oi_1 _9320_ (.Y(_4477_),
    .B1(_4474_),
    .B2(\uart_tx_inst.data[2] ),
    .A2(net261),
    .A1(\uart_tx_data[2] ));
 sg13g2_inv_1 _9321_ (.Y(_1767_),
    .A(_4477_));
 sg13g2_a22oi_1 _9322_ (.Y(_4478_),
    .B1(_4474_),
    .B2(\uart_tx_inst.data[3] ),
    .A2(net261),
    .A1(\uart_tx_data[3] ));
 sg13g2_inv_1 _9323_ (.Y(_1768_),
    .A(_4478_));
 sg13g2_a22oi_1 _9324_ (.Y(_4479_),
    .B1(_4474_),
    .B2(\uart_tx_inst.data[4] ),
    .A2(net261),
    .A1(\uart_tx_data[4] ));
 sg13g2_inv_1 _9325_ (.Y(_1769_),
    .A(_4479_));
 sg13g2_a22oi_1 _9326_ (.Y(_4480_),
    .B1(_4474_),
    .B2(\uart_tx_inst.data[5] ),
    .A2(net261),
    .A1(\uart_tx_data[5] ));
 sg13g2_inv_1 _9327_ (.Y(_1770_),
    .A(_4480_));
 sg13g2_a22oi_1 _9328_ (.Y(_4481_),
    .B1(_4474_),
    .B2(\uart_tx_inst.data[6] ),
    .A2(net261),
    .A1(\uart_tx_data[6] ));
 sg13g2_inv_1 _9329_ (.Y(_1771_),
    .A(_4481_));
 sg13g2_nor2_1 _9330_ (.A(uart_tx),
    .B(_4460_),
    .Y(_4482_));
 sg13g2_nor2b_1 _9331_ (.A(net390),
    .B_N(\uart_tx_inst.data[4] ),
    .Y(_4483_));
 sg13g2_a21oi_1 _9332_ (.A1(net390),
    .A2(\uart_tx_inst.data[5] ),
    .Y(_4484_),
    .B1(_4483_));
 sg13g2_nand3b_1 _9333_ (.B(\uart_tx_inst.data[6] ),
    .C(_1862_),
    .Y(_4485_),
    .A_N(net390));
 sg13g2_o21ai_1 _9334_ (.B1(_4485_),
    .Y(_4486_),
    .A1(_1862_),
    .A2(_4484_));
 sg13g2_mux4_1 _9335_ (.S0(net390),
    .A0(\uart_tx_inst.data[0] ),
    .A1(\uart_tx_inst.data[1] ),
    .A2(\uart_tx_inst.data[2] ),
    .A3(\uart_tx_inst.data[3] ),
    .S1(_1862_),
    .X(_4487_));
 sg13g2_nor2b_1 _9336_ (.A(\uart_tx_inst.bitIndex[2] ),
    .B_N(_4487_),
    .Y(_4488_));
 sg13g2_a21oi_1 _9337_ (.A1(\uart_tx_inst.bitIndex[2] ),
    .A2(_4486_),
    .Y(_4489_),
    .B1(_4488_));
 sg13g2_nor2_1 _9338_ (.A(_0596_),
    .B(_4489_),
    .Y(_4490_));
 sg13g2_nor4_1 _9339_ (.A(_2070_),
    .B(\uart_tx_inst.state[3] ),
    .C(_4463_),
    .D(_4490_),
    .Y(_4491_));
 sg13g2_o21ai_1 _9340_ (.B1(net329),
    .Y(_1772_),
    .A1(_4482_),
    .A2(_4491_));
 sg13g2_or2_1 _9341_ (.X(_4492_),
    .B(_1858_),
    .A(_1854_));
 sg13g2_buf_1 _9342_ (.A(_4492_),
    .X(_4493_));
 sg13g2_nand2_1 _9343_ (.Y(_4494_),
    .A(_1849_),
    .B(_1861_));
 sg13g2_o21ai_1 _9344_ (.B1(_4494_),
    .Y(_1774_),
    .A1(_1849_),
    .A2(_4493_));
 sg13g2_nand2_2 _9345_ (.Y(_4495_),
    .A(net372),
    .B(_4463_));
 sg13g2_nand2_1 _9346_ (.Y(_4496_),
    .A(_1849_),
    .B(_1857_));
 sg13g2_xor2_1 _9347_ (.B(_4496_),
    .A(_1848_),
    .X(_4497_));
 sg13g2_nor2_1 _9348_ (.A(_4495_),
    .B(_4497_),
    .Y(_1775_));
 sg13g2_nand3_1 _9349_ (.B(_1849_),
    .C(_1859_),
    .A(_1848_),
    .Y(_4498_));
 sg13g2_a21oi_1 _9350_ (.A1(_1848_),
    .A2(_1849_),
    .Y(_4499_),
    .B1(_4493_));
 sg13g2_o21ai_1 _9351_ (.B1(\uart_tx_inst.txCounter[2] ),
    .Y(_4500_),
    .A1(net261),
    .A2(_4499_));
 sg13g2_o21ai_1 _9352_ (.B1(_4500_),
    .Y(_1776_),
    .A1(\uart_tx_inst.txCounter[2] ),
    .A2(_4498_));
 sg13g2_and4_1 _9353_ (.A(\uart_tx_inst.txCounter[2] ),
    .B(_1848_),
    .C(_1849_),
    .D(_1857_),
    .X(_4501_));
 sg13g2_xnor2_1 _9354_ (.Y(_4502_),
    .A(\uart_tx_inst.txCounter[3] ),
    .B(_4501_));
 sg13g2_nor2_1 _9355_ (.A(_4495_),
    .B(_4502_),
    .Y(_1777_));
 sg13g2_a21o_1 _9356_ (.A2(_1859_),
    .A1(_1851_),
    .B1(_1860_),
    .X(_4503_));
 sg13g2_nor3_1 _9357_ (.A(\uart_tx_inst.txCounter[4] ),
    .B(_1851_),
    .C(_4493_),
    .Y(_4504_));
 sg13g2_a21o_1 _9358_ (.A2(_4503_),
    .A1(\uart_tx_inst.txCounter[4] ),
    .B1(_4504_),
    .X(_1778_));
 sg13g2_inv_1 _9359_ (.Y(_4505_),
    .A(\uart_tx_inst.txCounter[5] ));
 sg13g2_nand3_1 _9360_ (.B(\uart_tx_inst.txCounter[3] ),
    .C(_4501_),
    .A(\uart_tx_inst.txCounter[4] ),
    .Y(_4506_));
 sg13g2_xnor2_1 _9361_ (.Y(_4507_),
    .A(_4505_),
    .B(_4506_));
 sg13g2_nor2_1 _9362_ (.A(_4495_),
    .B(_4507_),
    .Y(_1779_));
 sg13g2_nor2_1 _9363_ (.A(_4505_),
    .B(_4506_),
    .Y(_4508_));
 sg13g2_xnor2_1 _9364_ (.Y(_4509_),
    .A(\uart_tx_inst.txCounter[6] ),
    .B(_4508_));
 sg13g2_nor2_1 _9365_ (.A(_4495_),
    .B(_4509_),
    .Y(_1780_));
 sg13g2_a21oi_1 _9366_ (.A1(\uart_tx_inst.txCounter[6] ),
    .A2(_4508_),
    .Y(_4510_),
    .B1(\uart_tx_inst.txCounter[7] ));
 sg13g2_nor2_1 _9367_ (.A(_4495_),
    .B(_4510_),
    .Y(_1781_));
 sg13g2_nor4_1 _9368_ (.A(_1892_),
    .B(\txstate[3] ),
    .C(\txstate[4] ),
    .D(\txstate[5] ),
    .Y(_4511_));
 sg13g2_nor2b_1 _9369_ (.A(_1783_),
    .B_N(net382),
    .Y(_4512_));
 sg13g2_nor3_1 _9370_ (.A(_1791_),
    .B(_4511_),
    .C(_4512_),
    .Y(_4513_));
 sg13g2_mux2_1 _9371_ (.A0(net398),
    .A1(net397),
    .S(_4513_),
    .X(_4514_));
 sg13g2_and2_1 _9372_ (.A(net322),
    .B(_4514_),
    .X(_1782_));
 sg13g2_nand2_1 _9373_ (.Y(_4515_),
    .A(_2114_),
    .B(_0071_));
 sg13g2_nor3_1 _9374_ (.A(net366),
    .B(net323),
    .C(\cell_index[4] ),
    .Y(_4516_));
 sg13g2_mux2_1 _9375_ (.A0(_2114_),
    .A1(_4515_),
    .S(_4516_),
    .X(_4517_));
 sg13g2_nand3_1 _9376_ (.B(_2095_),
    .C(_2093_),
    .A(_2092_),
    .Y(_4518_));
 sg13g2_nand2b_1 _9377_ (.Y(_4519_),
    .B(_4518_),
    .A_N(_2099_));
 sg13g2_xnor2_1 _9378_ (.Y(_4520_),
    .A(_2090_),
    .B(_4519_));
 sg13g2_nor3_2 _9379_ (.A(\hvsync_inst.vpos[9] ),
    .B(_4517_),
    .C(_4520_),
    .Y(net9));
 sg13g2_buf_2 _9380_ (.A(_2102_),
    .X(_4521_));
 sg13g2_buf_1 _9381_ (.A(net368),
    .X(_4522_));
 sg13g2_mux4_1 _9382_ (.S0(_4521_),
    .A0(\board_state[16] ),
    .A1(\board_state[17] ),
    .A2(\board_state[18] ),
    .A3(\board_state[19] ),
    .S1(net293),
    .X(_4523_));
 sg13g2_mux4_1 _9383_ (.S0(net325),
    .A0(\board_state[24] ),
    .A1(\board_state[25] ),
    .A2(\board_state[26] ),
    .A3(\board_state[27] ),
    .S1(net293),
    .X(_4524_));
 sg13g2_buf_2 _9384_ (.A(_2102_),
    .X(_4525_));
 sg13g2_buf_2 _9385_ (.A(net368),
    .X(_4526_));
 sg13g2_mux4_1 _9386_ (.S0(net292),
    .A0(\board_state[20] ),
    .A1(\board_state[21] ),
    .A2(\board_state[22] ),
    .A3(\board_state[23] ),
    .S1(net291),
    .X(_4527_));
 sg13g2_buf_2 _9387_ (.A(_2102_),
    .X(_4528_));
 sg13g2_mux4_1 _9388_ (.S0(net290),
    .A0(\board_state[28] ),
    .A1(\board_state[29] ),
    .A2(\board_state[30] ),
    .A3(\board_state[31] ),
    .S1(net291),
    .X(_4529_));
 sg13g2_mux4_1 _9389_ (.S0(net366),
    .A0(_4523_),
    .A1(_4524_),
    .A2(_4527_),
    .A3(_4529_),
    .S1(net323),
    .X(_4530_));
 sg13g2_mux4_1 _9390_ (.S0(net325),
    .A0(\board_state[0] ),
    .A1(\board_state[1] ),
    .A2(\board_state[2] ),
    .A3(\board_state[3] ),
    .S1(_4522_),
    .X(_4531_));
 sg13g2_mux4_1 _9391_ (.S0(net325),
    .A0(\board_state[8] ),
    .A1(\board_state[9] ),
    .A2(\board_state[10] ),
    .A3(\board_state[11] ),
    .S1(net324),
    .X(_4532_));
 sg13g2_buf_1 _9392_ (.A(net368),
    .X(_4533_));
 sg13g2_mux4_1 _9393_ (.S0(net290),
    .A0(\board_state[4] ),
    .A1(\board_state[5] ),
    .A2(\board_state[6] ),
    .A3(\board_state[7] ),
    .S1(net289),
    .X(_4534_));
 sg13g2_buf_2 _9394_ (.A(_2102_),
    .X(_4535_));
 sg13g2_mux4_1 _9395_ (.S0(_4535_),
    .A0(\board_state[12] ),
    .A1(\board_state[13] ),
    .A2(\board_state[14] ),
    .A3(\board_state[15] ),
    .S1(_4533_),
    .X(_4536_));
 sg13g2_mux4_1 _9396_ (.S0(net366),
    .A0(_4531_),
    .A1(_4532_),
    .A2(_4534_),
    .A3(_4536_),
    .S1(net323),
    .X(_4537_));
 sg13g2_mux4_1 _9397_ (.S0(_4525_),
    .A0(\board_state[48] ),
    .A1(\board_state[49] ),
    .A2(\board_state[50] ),
    .A3(\board_state[51] ),
    .S1(net291),
    .X(_4538_));
 sg13g2_mux4_1 _9398_ (.S0(_4528_),
    .A0(\board_state[56] ),
    .A1(\board_state[57] ),
    .A2(\board_state[58] ),
    .A3(\board_state[59] ),
    .S1(net289),
    .X(_4539_));
 sg13g2_buf_2 _9399_ (.A(_2101_),
    .X(_4540_));
 sg13g2_buf_1 _9400_ (.A(_2104_),
    .X(_4541_));
 sg13g2_buf_1 _9401_ (.A(_4541_),
    .X(_4542_));
 sg13g2_mux4_1 _9402_ (.S0(net342),
    .A0(\board_state[52] ),
    .A1(\board_state[53] ),
    .A2(\board_state[54] ),
    .A3(\board_state[55] ),
    .S1(net287),
    .X(_4543_));
 sg13g2_buf_1 _9403_ (.A(_4541_),
    .X(_4544_));
 sg13g2_mux4_1 _9404_ (.S0(net342),
    .A0(\board_state[60] ),
    .A1(\board_state[61] ),
    .A2(\board_state[62] ),
    .A3(\board_state[63] ),
    .S1(net286),
    .X(_4545_));
 sg13g2_buf_2 _9405_ (.A(net385),
    .X(_4546_));
 sg13g2_buf_2 _9406_ (.A(_2107_),
    .X(_4547_));
 sg13g2_mux4_1 _9407_ (.S0(_4546_),
    .A0(_4538_),
    .A1(_4539_),
    .A2(_4543_),
    .A3(_4545_),
    .S1(_4547_),
    .X(_4548_));
 sg13g2_mux4_1 _9408_ (.S0(_4528_),
    .A0(\board_state[32] ),
    .A1(\board_state[33] ),
    .A2(\board_state[34] ),
    .A3(\board_state[35] ),
    .S1(net291),
    .X(_4549_));
 sg13g2_mux4_1 _9409_ (.S0(net288),
    .A0(\board_state[40] ),
    .A1(\board_state[41] ),
    .A2(\board_state[42] ),
    .A3(\board_state[43] ),
    .S1(net289),
    .X(_4550_));
 sg13g2_mux4_1 _9410_ (.S0(net342),
    .A0(\board_state[36] ),
    .A1(\board_state[37] ),
    .A2(\board_state[38] ),
    .A3(\board_state[39] ),
    .S1(net287),
    .X(_4551_));
 sg13g2_buf_2 _9411_ (.A(_2101_),
    .X(_4552_));
 sg13g2_mux4_1 _9412_ (.S0(_4552_),
    .A0(\board_state[44] ),
    .A1(\board_state[45] ),
    .A2(\board_state[46] ),
    .A3(\board_state[47] ),
    .S1(_4544_),
    .X(_4553_));
 sg13g2_buf_1 _9413_ (.A(net367),
    .X(_4554_));
 sg13g2_mux4_1 _9414_ (.S0(net341),
    .A0(_4549_),
    .A1(_4550_),
    .A2(_4551_),
    .A3(_4553_),
    .S1(net285),
    .X(_4555_));
 sg13g2_mux4_1 _9415_ (.S0(net346),
    .A0(_4530_),
    .A1(_4537_),
    .A2(_4548_),
    .A3(_4555_),
    .S1(net347),
    .X(_4556_));
 sg13g2_mux4_1 _9416_ (.S0(net325),
    .A0(\board_state[80] ),
    .A1(\board_state[81] ),
    .A2(\board_state[82] ),
    .A3(\board_state[83] ),
    .S1(_4522_),
    .X(_4557_));
 sg13g2_mux4_1 _9417_ (.S0(_2103_),
    .A0(\board_state[88] ),
    .A1(\board_state[89] ),
    .A2(\board_state[90] ),
    .A3(\board_state[91] ),
    .S1(net324),
    .X(_4558_));
 sg13g2_mux4_1 _9418_ (.S0(net290),
    .A0(\board_state[84] ),
    .A1(\board_state[85] ),
    .A2(\board_state[86] ),
    .A3(\board_state[87] ),
    .S1(net289),
    .X(_4559_));
 sg13g2_mux4_1 _9419_ (.S0(net288),
    .A0(\board_state[92] ),
    .A1(\board_state[93] ),
    .A2(\board_state[94] ),
    .A3(\board_state[95] ),
    .S1(_4533_),
    .X(_4560_));
 sg13g2_mux4_1 _9420_ (.S0(_2113_),
    .A0(_4557_),
    .A1(_4558_),
    .A2(_4559_),
    .A3(_4560_),
    .S1(_2109_),
    .X(_4561_));
 sg13g2_mux4_1 _9421_ (.S0(_2103_),
    .A0(\board_state[64] ),
    .A1(\board_state[65] ),
    .A2(\board_state[66] ),
    .A3(\board_state[67] ),
    .S1(_2106_),
    .X(_4562_));
 sg13g2_mux4_1 _9422_ (.S0(net325),
    .A0(\board_state[72] ),
    .A1(\board_state[73] ),
    .A2(\board_state[74] ),
    .A3(\board_state[75] ),
    .S1(_2106_),
    .X(_4563_));
 sg13g2_buf_1 _9423_ (.A(net368),
    .X(_4564_));
 sg13g2_mux4_1 _9424_ (.S0(net288),
    .A0(\board_state[68] ),
    .A1(\board_state[69] ),
    .A2(\board_state[70] ),
    .A3(\board_state[71] ),
    .S1(net284),
    .X(_4565_));
 sg13g2_mux4_1 _9425_ (.S0(net288),
    .A0(\board_state[76] ),
    .A1(\board_state[77] ),
    .A2(\board_state[78] ),
    .A3(\board_state[79] ),
    .S1(_4564_),
    .X(_4566_));
 sg13g2_mux4_1 _9426_ (.S0(_2113_),
    .A0(_4562_),
    .A1(_4563_),
    .A2(_4565_),
    .A3(_4566_),
    .S1(_2109_),
    .X(_4567_));
 sg13g2_mux4_1 _9427_ (.S0(net290),
    .A0(\board_state[112] ),
    .A1(\board_state[113] ),
    .A2(\board_state[114] ),
    .A3(\board_state[115] ),
    .S1(net289),
    .X(_4568_));
 sg13g2_mux4_1 _9428_ (.S0(_4535_),
    .A0(\board_state[120] ),
    .A1(\board_state[121] ),
    .A2(\board_state[122] ),
    .A3(\board_state[123] ),
    .S1(net284),
    .X(_4569_));
 sg13g2_mux4_1 _9429_ (.S0(_4540_),
    .A0(\board_state[116] ),
    .A1(\board_state[117] ),
    .A2(\board_state[118] ),
    .A3(\board_state[119] ),
    .S1(_4544_),
    .X(_4570_));
 sg13g2_buf_1 _9430_ (.A(_4541_),
    .X(_4571_));
 sg13g2_mux4_1 _9431_ (.S0(_4552_),
    .A0(\board_state[124] ),
    .A1(\board_state[125] ),
    .A2(\board_state[126] ),
    .A3(\board_state[127] ),
    .S1(_4571_),
    .X(_4572_));
 sg13g2_mux4_1 _9432_ (.S0(net341),
    .A0(_4568_),
    .A1(_4569_),
    .A2(_4570_),
    .A3(_4572_),
    .S1(net285),
    .X(_4573_));
 sg13g2_mux4_1 _9433_ (.S0(net288),
    .A0(\board_state[96] ),
    .A1(\board_state[97] ),
    .A2(\board_state[98] ),
    .A3(\board_state[99] ),
    .S1(net289),
    .X(_4574_));
 sg13g2_mux4_1 _9434_ (.S0(_4521_),
    .A0(\board_state[104] ),
    .A1(\board_state[105] ),
    .A2(\board_state[106] ),
    .A3(\board_state[107] ),
    .S1(_4564_),
    .X(_4575_));
 sg13g2_mux4_1 _9435_ (.S0(net339),
    .A0(\board_state[100] ),
    .A1(\board_state[101] ),
    .A2(\board_state[102] ),
    .A3(\board_state[103] ),
    .S1(_4571_),
    .X(_4576_));
 sg13g2_buf_2 _9436_ (.A(_2102_),
    .X(_4577_));
 sg13g2_mux4_1 _9437_ (.S0(_4577_),
    .A0(\board_state[108] ),
    .A1(\board_state[109] ),
    .A2(\board_state[110] ),
    .A3(\board_state[111] ),
    .S1(net283),
    .X(_4578_));
 sg13g2_mux4_1 _9438_ (.S0(_4546_),
    .A0(_4574_),
    .A1(_4575_),
    .A2(_4576_),
    .A3(_4578_),
    .S1(net285),
    .X(_4579_));
 sg13g2_mux4_1 _9439_ (.S0(net346),
    .A0(_4561_),
    .A1(_4567_),
    .A2(_4573_),
    .A3(_4579_),
    .S1(_3575_),
    .X(_4580_));
 sg13g2_mux4_1 _9440_ (.S0(net290),
    .A0(\board_state[144] ),
    .A1(\board_state[145] ),
    .A2(\board_state[146] ),
    .A3(\board_state[147] ),
    .S1(_4526_),
    .X(_4581_));
 sg13g2_mux4_1 _9441_ (.S0(net290),
    .A0(\board_state[152] ),
    .A1(\board_state[153] ),
    .A2(\board_state[154] ),
    .A3(\board_state[155] ),
    .S1(net289),
    .X(_4582_));
 sg13g2_mux4_1 _9442_ (.S0(net342),
    .A0(\board_state[148] ),
    .A1(\board_state[149] ),
    .A2(\board_state[150] ),
    .A3(\board_state[151] ),
    .S1(_4542_),
    .X(_4583_));
 sg13g2_mux4_1 _9443_ (.S0(net342),
    .A0(\board_state[156] ),
    .A1(\board_state[157] ),
    .A2(\board_state[158] ),
    .A3(\board_state[159] ),
    .S1(net286),
    .X(_4584_));
 sg13g2_mux4_1 _9444_ (.S0(net341),
    .A0(_4581_),
    .A1(_4582_),
    .A2(_4583_),
    .A3(_4584_),
    .S1(_4547_),
    .X(_4585_));
 sg13g2_mux4_1 _9445_ (.S0(net290),
    .A0(\board_state[128] ),
    .A1(\board_state[129] ),
    .A2(\board_state[130] ),
    .A3(\board_state[131] ),
    .S1(net289),
    .X(_4586_));
 sg13g2_mux4_1 _9446_ (.S0(net288),
    .A0(\board_state[136] ),
    .A1(\board_state[137] ),
    .A2(\board_state[138] ),
    .A3(\board_state[139] ),
    .S1(net284),
    .X(_4587_));
 sg13g2_mux4_1 _9447_ (.S0(net339),
    .A0(\board_state[132] ),
    .A1(\board_state[133] ),
    .A2(\board_state[134] ),
    .A3(\board_state[135] ),
    .S1(net286),
    .X(_4588_));
 sg13g2_mux4_1 _9448_ (.S0(net282),
    .A0(\board_state[140] ),
    .A1(\board_state[141] ),
    .A2(\board_state[142] ),
    .A3(\board_state[143] ),
    .S1(net283),
    .X(_4589_));
 sg13g2_mux4_1 _9449_ (.S0(net341),
    .A0(_4586_),
    .A1(_4587_),
    .A2(_4588_),
    .A3(_4589_),
    .S1(net285),
    .X(_4590_));
 sg13g2_mux4_1 _9450_ (.S0(_4540_),
    .A0(\board_state[176] ),
    .A1(\board_state[177] ),
    .A2(\board_state[178] ),
    .A3(\board_state[179] ),
    .S1(_4542_),
    .X(_4591_));
 sg13g2_mux4_1 _9451_ (.S0(net339),
    .A0(\board_state[184] ),
    .A1(\board_state[185] ),
    .A2(\board_state[186] ),
    .A3(\board_state[187] ),
    .S1(net286),
    .X(_4592_));
 sg13g2_buf_2 _9452_ (.A(_2101_),
    .X(_4593_));
 sg13g2_buf_1 _9453_ (.A(_2104_),
    .X(_4594_));
 sg13g2_mux4_1 _9454_ (.S0(net338),
    .A0(\board_state[180] ),
    .A1(\board_state[181] ),
    .A2(\board_state[182] ),
    .A3(\board_state[183] ),
    .S1(net337),
    .X(_4595_));
 sg13g2_buf_2 _9455_ (.A(_2101_),
    .X(_4596_));
 sg13g2_mux4_1 _9456_ (.S0(net336),
    .A0(\board_state[188] ),
    .A1(\board_state[189] ),
    .A2(\board_state[190] ),
    .A3(\board_state[191] ),
    .S1(net337),
    .X(_4597_));
 sg13g2_mux4_1 _9457_ (.S0(net385),
    .A0(_4591_),
    .A1(_4592_),
    .A2(_4595_),
    .A3(_4597_),
    .S1(net367),
    .X(_4598_));
 sg13g2_mux4_1 _9458_ (.S0(net342),
    .A0(\board_state[160] ),
    .A1(\board_state[161] ),
    .A2(\board_state[162] ),
    .A3(\board_state[163] ),
    .S1(net286),
    .X(_4599_));
 sg13g2_mux4_1 _9459_ (.S0(net339),
    .A0(\board_state[168] ),
    .A1(\board_state[169] ),
    .A2(\board_state[170] ),
    .A3(\board_state[171] ),
    .S1(net283),
    .X(_4600_));
 sg13g2_mux4_1 _9460_ (.S0(net336),
    .A0(\board_state[164] ),
    .A1(\board_state[165] ),
    .A2(\board_state[166] ),
    .A3(\board_state[167] ),
    .S1(net337),
    .X(_4601_));
 sg13g2_buf_1 _9461_ (.A(_4541_),
    .X(_4602_));
 sg13g2_mux4_1 _9462_ (.S0(net336),
    .A0(\board_state[172] ),
    .A1(\board_state[173] ),
    .A2(\board_state[174] ),
    .A3(\board_state[175] ),
    .S1(_4602_),
    .X(_4603_));
 sg13g2_buf_2 _9463_ (.A(net385),
    .X(_4604_));
 sg13g2_mux4_1 _9464_ (.S0(_4604_),
    .A0(_4599_),
    .A1(_4600_),
    .A2(_4601_),
    .A3(_4603_),
    .S1(net367),
    .X(_4605_));
 sg13g2_mux4_1 _9465_ (.S0(_3669_),
    .A0(_4585_),
    .A1(_4590_),
    .A2(_4598_),
    .A3(_4605_),
    .S1(net347),
    .X(_4606_));
 sg13g2_mux4_1 _9466_ (.S0(net290),
    .A0(\board_state[208] ),
    .A1(\board_state[209] ),
    .A2(\board_state[210] ),
    .A3(\board_state[211] ),
    .S1(_4526_),
    .X(_4607_));
 sg13g2_mux4_1 _9467_ (.S0(net288),
    .A0(\board_state[216] ),
    .A1(\board_state[217] ),
    .A2(\board_state[218] ),
    .A3(\board_state[219] ),
    .S1(net284),
    .X(_4608_));
 sg13g2_mux4_1 _9468_ (.S0(net342),
    .A0(\board_state[212] ),
    .A1(\board_state[213] ),
    .A2(\board_state[214] ),
    .A3(\board_state[215] ),
    .S1(net286),
    .X(_4609_));
 sg13g2_mux4_1 _9469_ (.S0(net339),
    .A0(\board_state[220] ),
    .A1(\board_state[221] ),
    .A2(\board_state[222] ),
    .A3(\board_state[223] ),
    .S1(net283),
    .X(_4610_));
 sg13g2_mux4_1 _9470_ (.S0(net341),
    .A0(_4607_),
    .A1(_4608_),
    .A2(_4609_),
    .A3(_4610_),
    .S1(_4554_),
    .X(_4611_));
 sg13g2_mux4_1 _9471_ (.S0(net288),
    .A0(\board_state[192] ),
    .A1(\board_state[193] ),
    .A2(\board_state[194] ),
    .A3(\board_state[195] ),
    .S1(net284),
    .X(_4612_));
 sg13g2_mux4_1 _9472_ (.S0(net294),
    .A0(\board_state[200] ),
    .A1(\board_state[201] ),
    .A2(\board_state[202] ),
    .A3(\board_state[203] ),
    .S1(net284),
    .X(_4613_));
 sg13g2_mux4_1 _9473_ (.S0(net339),
    .A0(\board_state[196] ),
    .A1(\board_state[197] ),
    .A2(\board_state[198] ),
    .A3(\board_state[199] ),
    .S1(net283),
    .X(_4614_));
 sg13g2_mux4_1 _9474_ (.S0(net282),
    .A0(\board_state[204] ),
    .A1(\board_state[205] ),
    .A2(\board_state[206] ),
    .A3(\board_state[207] ),
    .S1(net283),
    .X(_4615_));
 sg13g2_mux4_1 _9475_ (.S0(net341),
    .A0(_4612_),
    .A1(_4613_),
    .A2(_4614_),
    .A3(_4615_),
    .S1(_4554_),
    .X(_4616_));
 sg13g2_mux4_1 _9476_ (.S0(net342),
    .A0(\board_state[240] ),
    .A1(\board_state[241] ),
    .A2(\board_state[242] ),
    .A3(\board_state[243] ),
    .S1(net286),
    .X(_4617_));
 sg13g2_mux4_1 _9477_ (.S0(net339),
    .A0(\board_state[248] ),
    .A1(\board_state[249] ),
    .A2(\board_state[250] ),
    .A3(\board_state[251] ),
    .S1(net283),
    .X(_4618_));
 sg13g2_mux4_1 _9478_ (.S0(net338),
    .A0(\board_state[244] ),
    .A1(\board_state[245] ),
    .A2(\board_state[246] ),
    .A3(\board_state[247] ),
    .S1(net337),
    .X(_4619_));
 sg13g2_mux4_1 _9479_ (.S0(net336),
    .A0(\board_state[252] ),
    .A1(\board_state[253] ),
    .A2(\board_state[254] ),
    .A3(\board_state[255] ),
    .S1(net337),
    .X(_4620_));
 sg13g2_mux4_1 _9480_ (.S0(net385),
    .A0(_4617_),
    .A1(_4618_),
    .A2(_4619_),
    .A3(_4620_),
    .S1(net367),
    .X(_4621_));
 sg13g2_mux4_1 _9481_ (.S0(net339),
    .A0(\board_state[224] ),
    .A1(\board_state[225] ),
    .A2(\board_state[226] ),
    .A3(\board_state[227] ),
    .S1(net286),
    .X(_4622_));
 sg13g2_mux4_1 _9482_ (.S0(_4577_),
    .A0(\board_state[232] ),
    .A1(\board_state[233] ),
    .A2(\board_state[234] ),
    .A3(\board_state[235] ),
    .S1(net283),
    .X(_4623_));
 sg13g2_mux4_1 _9483_ (.S0(_4596_),
    .A0(\board_state[228] ),
    .A1(\board_state[229] ),
    .A2(\board_state[230] ),
    .A3(\board_state[231] ),
    .S1(net337),
    .X(_4624_));
 sg13g2_mux4_1 _9484_ (.S0(_4596_),
    .A0(\board_state[236] ),
    .A1(\board_state[237] ),
    .A2(\board_state[238] ),
    .A3(\board_state[239] ),
    .S1(_4602_),
    .X(_4625_));
 sg13g2_mux4_1 _9485_ (.S0(_4604_),
    .A0(_4622_),
    .A1(_4623_),
    .A2(_4624_),
    .A3(_4625_),
    .S1(net367),
    .X(_4626_));
 sg13g2_mux4_1 _9486_ (.S0(_3669_),
    .A0(_4611_),
    .A1(_4616_),
    .A2(_4621_),
    .A3(_4626_),
    .S1(_3575_),
    .X(_4627_));
 sg13g2_mux4_1 _9487_ (.S0(_2092_),
    .A0(_4556_),
    .A1(_4580_),
    .A2(_4606_),
    .A3(_4627_),
    .S1(_2093_),
    .X(_4628_));
 sg13g2_mux4_1 _9488_ (.S0(net294),
    .A0(\board_state[272] ),
    .A1(\board_state[273] ),
    .A2(\board_state[274] ),
    .A3(\board_state[275] ),
    .S1(net284),
    .X(_4629_));
 sg13g2_mux4_1 _9489_ (.S0(net294),
    .A0(\board_state[280] ),
    .A1(\board_state[281] ),
    .A2(\board_state[282] ),
    .A3(\board_state[283] ),
    .S1(net284),
    .X(_4630_));
 sg13g2_buf_1 _9490_ (.A(_4541_),
    .X(_4631_));
 sg13g2_mux4_1 _9491_ (.S0(net282),
    .A0(\board_state[276] ),
    .A1(\board_state[277] ),
    .A2(\board_state[278] ),
    .A3(\board_state[279] ),
    .S1(net280),
    .X(_4632_));
 sg13g2_mux4_1 _9492_ (.S0(net282),
    .A0(\board_state[284] ),
    .A1(\board_state[285] ),
    .A2(\board_state[286] ),
    .A3(\board_state[287] ),
    .S1(net280),
    .X(_4633_));
 sg13g2_mux4_1 _9493_ (.S0(net341),
    .A0(_4629_),
    .A1(_4630_),
    .A2(_4632_),
    .A3(_4633_),
    .S1(net285),
    .X(_4634_));
 sg13g2_mux4_1 _9494_ (.S0(net294),
    .A0(\board_state[256] ),
    .A1(\board_state[257] ),
    .A2(\board_state[258] ),
    .A3(\board_state[259] ),
    .S1(net293),
    .X(_4635_));
 sg13g2_mux4_1 _9495_ (.S0(net294),
    .A0(\board_state[264] ),
    .A1(\board_state[265] ),
    .A2(\board_state[266] ),
    .A3(\board_state[267] ),
    .S1(net293),
    .X(_4636_));
 sg13g2_buf_2 _9496_ (.A(_2102_),
    .X(_4637_));
 sg13g2_mux4_1 _9497_ (.S0(net279),
    .A0(\board_state[260] ),
    .A1(\board_state[261] ),
    .A2(\board_state[262] ),
    .A3(\board_state[263] ),
    .S1(net280),
    .X(_4638_));
 sg13g2_buf_1 _9498_ (.A(_4541_),
    .X(_4639_));
 sg13g2_mux4_1 _9499_ (.S0(net279),
    .A0(\board_state[268] ),
    .A1(\board_state[269] ),
    .A2(\board_state[270] ),
    .A3(\board_state[271] ),
    .S1(net278),
    .X(_4640_));
 sg13g2_mux4_1 _9500_ (.S0(net341),
    .A0(_4635_),
    .A1(_4636_),
    .A2(_4638_),
    .A3(_4640_),
    .S1(net285),
    .X(_4641_));
 sg13g2_mux4_1 _9501_ (.S0(net282),
    .A0(\board_state[304] ),
    .A1(\board_state[305] ),
    .A2(\board_state[306] ),
    .A3(\board_state[307] ),
    .S1(net280),
    .X(_4642_));
 sg13g2_mux4_1 _9502_ (.S0(net279),
    .A0(\board_state[312] ),
    .A1(\board_state[313] ),
    .A2(\board_state[314] ),
    .A3(\board_state[315] ),
    .S1(net280),
    .X(_4643_));
 sg13g2_mux4_1 _9503_ (.S0(net336),
    .A0(\board_state[308] ),
    .A1(\board_state[309] ),
    .A2(\board_state[310] ),
    .A3(\board_state[311] ),
    .S1(net281),
    .X(_4644_));
 sg13g2_buf_2 _9504_ (.A(_2101_),
    .X(_4645_));
 sg13g2_mux4_1 _9505_ (.S0(net334),
    .A0(\board_state[316] ),
    .A1(\board_state[317] ),
    .A2(\board_state[318] ),
    .A3(\board_state[319] ),
    .S1(net281),
    .X(_4646_));
 sg13g2_mux4_1 _9506_ (.S0(net335),
    .A0(_4642_),
    .A1(_4643_),
    .A2(_4644_),
    .A3(_4646_),
    .S1(net340),
    .X(_4647_));
 sg13g2_mux4_1 _9507_ (.S0(net282),
    .A0(\board_state[288] ),
    .A1(\board_state[289] ),
    .A2(\board_state[290] ),
    .A3(\board_state[291] ),
    .S1(net280),
    .X(_4648_));
 sg13g2_mux4_1 _9508_ (.S0(net279),
    .A0(\board_state[296] ),
    .A1(\board_state[297] ),
    .A2(\board_state[298] ),
    .A3(\board_state[299] ),
    .S1(net278),
    .X(_4649_));
 sg13g2_mux4_1 _9509_ (.S0(net336),
    .A0(\board_state[292] ),
    .A1(\board_state[293] ),
    .A2(\board_state[294] ),
    .A3(\board_state[295] ),
    .S1(net281),
    .X(_4650_));
 sg13g2_buf_1 _9510_ (.A(_4541_),
    .X(_4651_));
 sg13g2_mux4_1 _9511_ (.S0(net334),
    .A0(\board_state[300] ),
    .A1(\board_state[301] ),
    .A2(\board_state[302] ),
    .A3(\board_state[303] ),
    .S1(net277),
    .X(_4652_));
 sg13g2_mux4_1 _9512_ (.S0(net335),
    .A0(_4648_),
    .A1(_4649_),
    .A2(_4650_),
    .A3(_4652_),
    .S1(net340),
    .X(_4653_));
 sg13g2_mux4_1 _9513_ (.S0(net346),
    .A0(_4634_),
    .A1(_4641_),
    .A2(_4647_),
    .A3(_4653_),
    .S1(net347),
    .X(_4654_));
 sg13g2_mux4_1 _9514_ (.S0(net294),
    .A0(\board_state[336] ),
    .A1(\board_state[337] ),
    .A2(\board_state[338] ),
    .A3(\board_state[339] ),
    .S1(net293),
    .X(_4655_));
 sg13g2_mux4_1 _9515_ (.S0(net294),
    .A0(\board_state[344] ),
    .A1(\board_state[345] ),
    .A2(\board_state[346] ),
    .A3(\board_state[347] ),
    .S1(net293),
    .X(_4656_));
 sg13g2_mux4_1 _9516_ (.S0(net279),
    .A0(\board_state[340] ),
    .A1(\board_state[341] ),
    .A2(\board_state[342] ),
    .A3(\board_state[343] ),
    .S1(net280),
    .X(_4657_));
 sg13g2_mux4_1 _9517_ (.S0(net279),
    .A0(\board_state[348] ),
    .A1(\board_state[349] ),
    .A2(\board_state[350] ),
    .A3(\board_state[351] ),
    .S1(net278),
    .X(_4658_));
 sg13g2_mux4_1 _9518_ (.S0(net366),
    .A0(_4655_),
    .A1(_4656_),
    .A2(_4657_),
    .A3(_4658_),
    .S1(net285),
    .X(_4659_));
 sg13g2_mux4_1 _9519_ (.S0(net294),
    .A0(\board_state[320] ),
    .A1(\board_state[321] ),
    .A2(\board_state[322] ),
    .A3(\board_state[323] ),
    .S1(net293),
    .X(_4660_));
 sg13g2_mux4_1 _9520_ (.S0(net325),
    .A0(\board_state[328] ),
    .A1(\board_state[329] ),
    .A2(\board_state[330] ),
    .A3(\board_state[331] ),
    .S1(net293),
    .X(_4661_));
 sg13g2_mux4_1 _9521_ (.S0(net292),
    .A0(\board_state[324] ),
    .A1(\board_state[325] ),
    .A2(\board_state[326] ),
    .A3(\board_state[327] ),
    .S1(net278),
    .X(_4662_));
 sg13g2_mux4_1 _9522_ (.S0(net292),
    .A0(\board_state[332] ),
    .A1(\board_state[333] ),
    .A2(\board_state[334] ),
    .A3(\board_state[335] ),
    .S1(net291),
    .X(_4663_));
 sg13g2_mux4_1 _9523_ (.S0(net366),
    .A0(_4660_),
    .A1(_4661_),
    .A2(_4662_),
    .A3(_4663_),
    .S1(net285),
    .X(_4664_));
 sg13g2_mux4_1 _9524_ (.S0(_4637_),
    .A0(\board_state[368] ),
    .A1(\board_state[369] ),
    .A2(\board_state[370] ),
    .A3(\board_state[371] ),
    .S1(net280),
    .X(_4665_));
 sg13g2_mux4_1 _9525_ (.S0(net292),
    .A0(\board_state[376] ),
    .A1(\board_state[377] ),
    .A2(\board_state[378] ),
    .A3(\board_state[379] ),
    .S1(net278),
    .X(_4666_));
 sg13g2_mux4_1 _9526_ (.S0(net334),
    .A0(\board_state[372] ),
    .A1(\board_state[373] ),
    .A2(\board_state[374] ),
    .A3(\board_state[375] ),
    .S1(net277),
    .X(_4667_));
 sg13g2_buf_2 _9527_ (.A(_2101_),
    .X(_4668_));
 sg13g2_mux4_1 _9528_ (.S0(net333),
    .A0(\board_state[380] ),
    .A1(\board_state[381] ),
    .A2(\board_state[382] ),
    .A3(\board_state[383] ),
    .S1(net277),
    .X(_4669_));
 sg13g2_mux4_1 _9529_ (.S0(net335),
    .A0(_4665_),
    .A1(_4666_),
    .A2(_4667_),
    .A3(_4669_),
    .S1(net340),
    .X(_4670_));
 sg13g2_mux4_1 _9530_ (.S0(net279),
    .A0(\board_state[352] ),
    .A1(\board_state[353] ),
    .A2(\board_state[354] ),
    .A3(\board_state[355] ),
    .S1(net278),
    .X(_4671_));
 sg13g2_mux4_1 _9531_ (.S0(net292),
    .A0(\board_state[360] ),
    .A1(\board_state[361] ),
    .A2(\board_state[362] ),
    .A3(\board_state[363] ),
    .S1(net291),
    .X(_4672_));
 sg13g2_mux4_1 _9532_ (.S0(net333),
    .A0(\board_state[356] ),
    .A1(\board_state[357] ),
    .A2(\board_state[358] ),
    .A3(\board_state[359] ),
    .S1(net277),
    .X(_4673_));
 sg13g2_mux4_1 _9533_ (.S0(net333),
    .A0(\board_state[364] ),
    .A1(\board_state[365] ),
    .A2(\board_state[366] ),
    .A3(\board_state[367] ),
    .S1(net287),
    .X(_4674_));
 sg13g2_mux4_1 _9534_ (.S0(net335),
    .A0(_4671_),
    .A1(_4672_),
    .A2(_4673_),
    .A3(_4674_),
    .S1(net340),
    .X(_4675_));
 sg13g2_mux4_1 _9535_ (.S0(net346),
    .A0(_4659_),
    .A1(_4664_),
    .A2(_4670_),
    .A3(_4675_),
    .S1(net347),
    .X(_4676_));
 sg13g2_mux4_1 _9536_ (.S0(net282),
    .A0(\board_state[400] ),
    .A1(\board_state[401] ),
    .A2(\board_state[402] ),
    .A3(\board_state[403] ),
    .S1(_4631_),
    .X(_4677_));
 sg13g2_mux4_1 _9537_ (.S0(_4637_),
    .A0(\board_state[408] ),
    .A1(\board_state[409] ),
    .A2(\board_state[410] ),
    .A3(\board_state[411] ),
    .S1(net278),
    .X(_4678_));
 sg13g2_mux4_1 _9538_ (.S0(net336),
    .A0(\board_state[404] ),
    .A1(\board_state[405] ),
    .A2(\board_state[406] ),
    .A3(\board_state[407] ),
    .S1(net281),
    .X(_4679_));
 sg13g2_mux4_1 _9539_ (.S0(net334),
    .A0(\board_state[412] ),
    .A1(\board_state[413] ),
    .A2(\board_state[414] ),
    .A3(\board_state[415] ),
    .S1(net277),
    .X(_4680_));
 sg13g2_mux4_1 _9540_ (.S0(net335),
    .A0(_4677_),
    .A1(_4678_),
    .A2(_4679_),
    .A3(_4680_),
    .S1(net340),
    .X(_4681_));
 sg13g2_mux4_1 _9541_ (.S0(net279),
    .A0(\board_state[384] ),
    .A1(\board_state[385] ),
    .A2(\board_state[386] ),
    .A3(\board_state[387] ),
    .S1(net278),
    .X(_4682_));
 sg13g2_mux4_1 _9542_ (.S0(net292),
    .A0(\board_state[392] ),
    .A1(\board_state[393] ),
    .A2(\board_state[394] ),
    .A3(\board_state[395] ),
    .S1(net291),
    .X(_4683_));
 sg13g2_mux4_1 _9543_ (.S0(net334),
    .A0(\board_state[388] ),
    .A1(\board_state[389] ),
    .A2(\board_state[390] ),
    .A3(\board_state[391] ),
    .S1(net277),
    .X(_4684_));
 sg13g2_mux4_1 _9544_ (.S0(net333),
    .A0(\board_state[396] ),
    .A1(\board_state[397] ),
    .A2(\board_state[398] ),
    .A3(\board_state[399] ),
    .S1(net287),
    .X(_4685_));
 sg13g2_mux4_1 _9545_ (.S0(net335),
    .A0(_4682_),
    .A1(_4683_),
    .A2(_4684_),
    .A3(_4685_),
    .S1(net340),
    .X(_4686_));
 sg13g2_mux4_1 _9546_ (.S0(net336),
    .A0(\board_state[432] ),
    .A1(\board_state[433] ),
    .A2(\board_state[434] ),
    .A3(\board_state[435] ),
    .S1(net281),
    .X(_4687_));
 sg13g2_mux4_1 _9547_ (.S0(net334),
    .A0(\board_state[440] ),
    .A1(\board_state[441] ),
    .A2(\board_state[442] ),
    .A3(\board_state[443] ),
    .S1(net277),
    .X(_4688_));
 sg13g2_mux4_1 _9548_ (.S0(net338),
    .A0(\board_state[436] ),
    .A1(\board_state[437] ),
    .A2(\board_state[438] ),
    .A3(\board_state[439] ),
    .S1(net368),
    .X(_4689_));
 sg13g2_mux4_1 _9549_ (.S0(net338),
    .A0(\board_state[444] ),
    .A1(\board_state[445] ),
    .A2(\board_state[446] ),
    .A3(\board_state[447] ),
    .S1(net368),
    .X(_4690_));
 sg13g2_mux4_1 _9550_ (.S0(net385),
    .A0(_4687_),
    .A1(_4688_),
    .A2(_4689_),
    .A3(_4690_),
    .S1(net367),
    .X(_4691_));
 sg13g2_mux4_1 _9551_ (.S0(net334),
    .A0(\board_state[416] ),
    .A1(\board_state[417] ),
    .A2(\board_state[418] ),
    .A3(\board_state[419] ),
    .S1(net281),
    .X(_4692_));
 sg13g2_mux4_1 _9552_ (.S0(_4668_),
    .A0(\board_state[424] ),
    .A1(\board_state[425] ),
    .A2(\board_state[426] ),
    .A3(\board_state[427] ),
    .S1(net287),
    .X(_4693_));
 sg13g2_mux4_1 _9553_ (.S0(net338),
    .A0(\board_state[420] ),
    .A1(\board_state[421] ),
    .A2(\board_state[422] ),
    .A3(\board_state[423] ),
    .S1(net368),
    .X(_4694_));
 sg13g2_mux4_1 _9554_ (.S0(net338),
    .A0(\board_state[428] ),
    .A1(\board_state[429] ),
    .A2(\board_state[430] ),
    .A3(\board_state[431] ),
    .S1(net337),
    .X(_4695_));
 sg13g2_mux4_1 _9555_ (.S0(net385),
    .A0(_4692_),
    .A1(_4693_),
    .A2(_4694_),
    .A3(_4695_),
    .S1(net367),
    .X(_4696_));
 sg13g2_mux4_1 _9556_ (.S0(net346),
    .A0(_4681_),
    .A1(_4686_),
    .A2(_4691_),
    .A3(_4696_),
    .S1(_2095_),
    .X(_4697_));
 sg13g2_mux4_1 _9557_ (.S0(net282),
    .A0(\board_state[464] ),
    .A1(\board_state[465] ),
    .A2(\board_state[466] ),
    .A3(\board_state[467] ),
    .S1(_4631_),
    .X(_4698_));
 sg13g2_mux4_1 _9558_ (.S0(net292),
    .A0(\board_state[472] ),
    .A1(\board_state[473] ),
    .A2(\board_state[474] ),
    .A3(\board_state[475] ),
    .S1(_4639_),
    .X(_4699_));
 sg13g2_mux4_1 _9559_ (.S0(net334),
    .A0(\board_state[468] ),
    .A1(\board_state[469] ),
    .A2(\board_state[470] ),
    .A3(\board_state[471] ),
    .S1(net281),
    .X(_4700_));
 sg13g2_mux4_1 _9560_ (.S0(net333),
    .A0(\board_state[476] ),
    .A1(\board_state[477] ),
    .A2(\board_state[478] ),
    .A3(\board_state[479] ),
    .S1(net277),
    .X(_4701_));
 sg13g2_mux4_1 _9561_ (.S0(net335),
    .A0(_4698_),
    .A1(_4699_),
    .A2(_4700_),
    .A3(_4701_),
    .S1(net340),
    .X(_4702_));
 sg13g2_mux4_1 _9562_ (.S0(net292),
    .A0(\board_state[448] ),
    .A1(\board_state[449] ),
    .A2(\board_state[450] ),
    .A3(\board_state[451] ),
    .S1(_4639_),
    .X(_4703_));
 sg13g2_mux4_1 _9563_ (.S0(_4525_),
    .A0(\board_state[456] ),
    .A1(\board_state[457] ),
    .A2(\board_state[458] ),
    .A3(\board_state[459] ),
    .S1(net291),
    .X(_4704_));
 sg13g2_mux4_1 _9564_ (.S0(net333),
    .A0(\board_state[452] ),
    .A1(\board_state[453] ),
    .A2(\board_state[454] ),
    .A3(\board_state[455] ),
    .S1(net287),
    .X(_4705_));
 sg13g2_mux4_1 _9565_ (.S0(net333),
    .A0(\board_state[460] ),
    .A1(\board_state[461] ),
    .A2(\board_state[462] ),
    .A3(\board_state[463] ),
    .S1(net287),
    .X(_4706_));
 sg13g2_mux4_1 _9566_ (.S0(net335),
    .A0(_4703_),
    .A1(_4704_),
    .A2(_4705_),
    .A3(_4706_),
    .S1(net340),
    .X(_4707_));
 sg13g2_mux4_1 _9567_ (.S0(_4645_),
    .A0(\board_state[496] ),
    .A1(\board_state[497] ),
    .A2(\board_state[498] ),
    .A3(\board_state[499] ),
    .S1(net281),
    .X(_4708_));
 sg13g2_mux4_1 _9568_ (.S0(net333),
    .A0(\board_state[504] ),
    .A1(\board_state[505] ),
    .A2(\board_state[506] ),
    .A3(\board_state[507] ),
    .S1(_4651_),
    .X(_4709_));
 sg13g2_mux4_1 _9569_ (.S0(net338),
    .A0(\board_state[500] ),
    .A1(\board_state[501] ),
    .A2(\board_state[502] ),
    .A3(\board_state[503] ),
    .S1(net368),
    .X(_4710_));
 sg13g2_mux4_1 _9570_ (.S0(net338),
    .A0(\board_state[508] ),
    .A1(\board_state[509] ),
    .A2(\board_state[510] ),
    .A3(\board_state[511] ),
    .S1(net337),
    .X(_4711_));
 sg13g2_mux4_1 _9571_ (.S0(net385),
    .A0(_4708_),
    .A1(_4709_),
    .A2(_4710_),
    .A3(_4711_),
    .S1(_2108_),
    .X(_4712_));
 sg13g2_mux4_1 _9572_ (.S0(_4645_),
    .A0(\board_state[480] ),
    .A1(\board_state[481] ),
    .A2(\board_state[482] ),
    .A3(\board_state[483] ),
    .S1(_4651_),
    .X(_4713_));
 sg13g2_mux4_1 _9573_ (.S0(_4668_),
    .A0(\board_state[488] ),
    .A1(\board_state[489] ),
    .A2(\board_state[490] ),
    .A3(\board_state[491] ),
    .S1(net287),
    .X(_4714_));
 sg13g2_mux4_1 _9574_ (.S0(_4593_),
    .A0(\board_state[484] ),
    .A1(\board_state[485] ),
    .A2(\board_state[486] ),
    .A3(\board_state[487] ),
    .S1(_4594_),
    .X(_4715_));
 sg13g2_mux4_1 _9575_ (.S0(_4593_),
    .A0(\board_state[492] ),
    .A1(\board_state[493] ),
    .A2(\board_state[494] ),
    .A3(\board_state[495] ),
    .S1(_4594_),
    .X(_4716_));
 sg13g2_mux4_1 _9576_ (.S0(_2112_),
    .A0(_4713_),
    .A1(_4714_),
    .A2(_4715_),
    .A3(_4716_),
    .S1(_2108_),
    .X(_4717_));
 sg13g2_mux4_1 _9577_ (.S0(net346),
    .A0(_4702_),
    .A1(_4707_),
    .A2(_4712_),
    .A3(_4717_),
    .S1(net347),
    .X(_4718_));
 sg13g2_mux4_1 _9578_ (.S0(_2092_),
    .A0(_4654_),
    .A1(_4676_),
    .A2(_4697_),
    .A3(_4718_),
    .S1(_2093_),
    .X(_4719_));
 sg13g2_mux2_1 _9579_ (.A0(_4628_),
    .A1(_4719_),
    .S(_2099_),
    .X(_4720_));
 sg13g2_inv_1 _9580_ (.Y(_4721_),
    .A(_2119_));
 sg13g2_nor2b_1 _9581_ (.A(_2120_),
    .B_N(_4734_),
    .Y(_4722_));
 sg13g2_a21oi_1 _9582_ (.A1(_2120_),
    .A2(_4735_),
    .Y(_4723_),
    .B1(_4722_));
 sg13g2_nor2_1 _9583_ (.A(_2117_),
    .B(_4736_),
    .Y(_4724_));
 sg13g2_a21oi_1 _9584_ (.A1(_2117_),
    .A2(_4723_),
    .Y(_4725_),
    .B1(_4724_));
 sg13g2_nor2_1 _9585_ (.A(_4721_),
    .B(_2117_),
    .Y(_4726_));
 sg13g2_a22oi_1 _9586_ (.Y(_4727_),
    .B1(_4726_),
    .B2(_4733_),
    .A2(_4725_),
    .A1(_4721_));
 sg13g2_mux2_1 _9587_ (.A0(_4735_),
    .A1(_4734_),
    .S(_2120_),
    .X(_4728_));
 sg13g2_nor2_1 _9588_ (.A(_2117_),
    .B(_0072_),
    .Y(_4729_));
 sg13g2_mux2_1 _9589_ (.A0(_4733_),
    .A1(_4736_),
    .S(_2119_),
    .X(_4730_));
 sg13g2_a221oi_1 _9590_ (.B2(_2117_),
    .C1(_2118_),
    .B1(_4730_),
    .A1(_4728_),
    .Y(_4731_),
    .A2(_4729_));
 sg13g2_a21oi_1 _9591_ (.A1(_2118_),
    .A2(_4727_),
    .Y(_4732_),
    .B1(_4731_));
 sg13g2_and3_1 _9592_ (.X(net6),
    .A(net9),
    .B(_4720_),
    .C(_4732_));
 sg13g2_dfrbp_1 _9593_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net417),
    .D(_0600_),
    .Q_N(_5388_),
    .Q(_0000_));
 sg13g2_dfrbp_1 _9594_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net418),
    .D(_0601_),
    .Q_N(_5387_),
    .Q(_0001_));
 sg13g2_dfrbp_1 _9595_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net419),
    .D(_0602_),
    .Q_N(_5386_),
    .Q(_0002_));
 sg13g2_dfrbp_1 _9596_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net420),
    .D(_0603_),
    .Q_N(_5385_),
    .Q(_0003_));
 sg13g2_dfrbp_1 _9597_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net421),
    .D(_0604_),
    .Q_N(_5384_),
    .Q(_0004_));
 sg13g2_dfrbp_1 _9598_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net422),
    .D(_0605_),
    .Q_N(_5383_),
    .Q(_0005_));
 sg13g2_dfrbp_1 _9599_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net423),
    .D(_0606_),
    .Q_N(_5382_),
    .Q(_0006_));
 sg13g2_dfrbp_1 _9600_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net424),
    .D(_0607_),
    .Q_N(_5381_),
    .Q(_0007_));
 sg13g2_dfrbp_1 _9601_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net425),
    .D(_0608_),
    .Q_N(_5389_),
    .Q(_0008_));
 sg13g2_dfrbp_1 _9602_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net426),
    .D(_0009_),
    .Q_N(_5390_),
    .Q(_4735_));
 sg13g2_dfrbp_1 _9603_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net427),
    .D(_0012_),
    .Q_N(_5391_),
    .Q(_4736_));
 sg13g2_dfrbp_1 _9604_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net428),
    .D(_0011_),
    .Q_N(_5392_),
    .Q(_4733_));
 sg13g2_dfrbp_1 _9605_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net429),
    .D(_0010_),
    .Q_N(_5393_),
    .Q(_4734_));
 sg13g2_dfrbp_1 _9606_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net430),
    .D(_0013_),
    .Q_N(_5394_),
    .Q(_0046_));
 sg13g2_dfrbp_1 _9607_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net431),
    .D(_0014_),
    .Q_N(_5395_),
    .Q(_0047_));
 sg13g2_dfrbp_1 _9608_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net432),
    .D(_0015_),
    .Q_N(_5396_),
    .Q(_0048_));
 sg13g2_dfrbp_1 _9609_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net433),
    .D(_0016_),
    .Q_N(_5397_),
    .Q(_0049_));
 sg13g2_dfrbp_1 _9610_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net434),
    .D(_0017_),
    .Q_N(_5398_),
    .Q(_0050_));
 sg13g2_dfrbp_1 _9611_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net435),
    .D(_0018_),
    .Q_N(_5399_),
    .Q(_0051_));
 sg13g2_dfrbp_1 _9612_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net436),
    .D(_0019_),
    .Q_N(_5400_),
    .Q(_0052_));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_tiehi _9593__417 (.L_HI(net417));
 sg13g2_buf_1 _9615_ (.A(net437),
    .X(uio_oe[0]));
 sg13g2_buf_1 _9616_ (.A(net402),
    .X(uio_oe[1]));
 sg13g2_buf_1 _9617_ (.A(net403),
    .X(uio_oe[2]));
 sg13g2_buf_1 _9618_ (.A(net404),
    .X(uio_oe[3]));
 sg13g2_buf_1 _9619_ (.A(net405),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9620_ (.A(net406),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9621_ (.A(net407),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9622_ (.A(net408),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9623_ (.A(net6),
    .X(net5));
 sg13g2_buf_1 _9624_ (.A(net409),
    .X(uio_out[2]));
 sg13g2_buf_1 _9625_ (.A(\hvsync_inst.vsync ),
    .X(net7));
 sg13g2_buf_1 _9626_ (.A(net9),
    .X(net8));
 sg13g2_buf_1 _9627_ (.A(net438),
    .X(uio_out[6]));
 sg13g2_buf_1 _9628_ (.A(hsync),
    .X(net10));
 sg13g2_buf_1 _9629_ (.A(net410),
    .X(uo_out[0]));
 sg13g2_buf_1 _9630_ (.A(net411),
    .X(uo_out[1]));
 sg13g2_buf_1 _9631_ (.A(net412),
    .X(uo_out[2]));
 sg13g2_buf_1 _9632_ (.A(net413),
    .X(uo_out[3]));
 sg13g2_buf_1 _9633_ (.A(uart_tx),
    .X(net11));
 sg13g2_buf_1 _9634_ (.A(net414),
    .X(uo_out[5]));
 sg13g2_buf_1 _9635_ (.A(net415),
    .X(uo_out[6]));
 sg13g2_buf_1 _9636_ (.A(net416),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \action[0]$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net439),
    .D(_0020_),
    .Q_N(_5401_),
    .Q(\action[0] ));
 sg13g2_dfrbp_1 \action[1]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net440),
    .D(_0021_),
    .Q_N(_5402_),
    .Q(\action[1] ));
 sg13g2_dfrbp_1 \action[2]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net441),
    .D(_0022_),
    .Q_N(_5403_),
    .Q(\action[2] ));
 sg13g2_dfrbp_1 \action[3]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net442),
    .D(_0023_),
    .Q_N(_0055_),
    .Q(\action[3] ));
 sg13g2_dfrbp_1 \action[4]$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net443),
    .D(_0024_),
    .Q_N(_5404_),
    .Q(\action[4] ));
 sg13g2_dfrbp_1 \action[5]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net444),
    .D(_0025_),
    .Q_N(_5405_),
    .Q(\action[5] ));
 sg13g2_dfrbp_1 \action[6]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net445),
    .D(_0026_),
    .Q_N(_0058_),
    .Q(\action[6] ));
 sg13g2_dfrbp_1 \action[7]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net446),
    .D(_0027_),
    .Q_N(_0053_),
    .Q(\action[7] ));
 sg13g2_dfrbp_1 \board_state[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net447),
    .D(_0609_),
    .Q_N(_0082_),
    .Q(\board_state[0] ));
 sg13g2_dfrbp_1 \board_state[100]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net448),
    .D(_0610_),
    .Q_N(_0183_),
    .Q(\board_state[100] ));
 sg13g2_dfrbp_1 \board_state[101]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net449),
    .D(_0611_),
    .Q_N(_0184_),
    .Q(\board_state[101] ));
 sg13g2_dfrbp_1 \board_state[102]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net450),
    .D(_0612_),
    .Q_N(_0185_),
    .Q(\board_state[102] ));
 sg13g2_dfrbp_1 \board_state[103]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net451),
    .D(_0613_),
    .Q_N(_0186_),
    .Q(\board_state[103] ));
 sg13g2_dfrbp_1 \board_state[104]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net452),
    .D(_0614_),
    .Q_N(_0187_),
    .Q(\board_state[104] ));
 sg13g2_dfrbp_1 \board_state[105]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net453),
    .D(_0615_),
    .Q_N(_0188_),
    .Q(\board_state[105] ));
 sg13g2_dfrbp_1 \board_state[106]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net454),
    .D(_0616_),
    .Q_N(_0189_),
    .Q(\board_state[106] ));
 sg13g2_dfrbp_1 \board_state[107]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net455),
    .D(_0617_),
    .Q_N(_0190_),
    .Q(\board_state[107] ));
 sg13g2_dfrbp_1 \board_state[108]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net456),
    .D(_0618_),
    .Q_N(_0191_),
    .Q(\board_state[108] ));
 sg13g2_dfrbp_1 \board_state[109]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net457),
    .D(_0619_),
    .Q_N(_0192_),
    .Q(\board_state[109] ));
 sg13g2_dfrbp_1 \board_state[10]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net458),
    .D(_0620_),
    .Q_N(_0093_),
    .Q(\board_state[10] ));
 sg13g2_dfrbp_1 \board_state[110]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net459),
    .D(_0621_),
    .Q_N(_0193_),
    .Q(\board_state[110] ));
 sg13g2_dfrbp_1 \board_state[111]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net460),
    .D(_0622_),
    .Q_N(_0194_),
    .Q(\board_state[111] ));
 sg13g2_dfrbp_1 \board_state[112]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net461),
    .D(_0623_),
    .Q_N(_0195_),
    .Q(\board_state[112] ));
 sg13g2_dfrbp_1 \board_state[113]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net462),
    .D(_0624_),
    .Q_N(_0196_),
    .Q(\board_state[113] ));
 sg13g2_dfrbp_1 \board_state[114]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net463),
    .D(_0625_),
    .Q_N(_0197_),
    .Q(\board_state[114] ));
 sg13g2_dfrbp_1 \board_state[115]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net464),
    .D(_0626_),
    .Q_N(_0198_),
    .Q(\board_state[115] ));
 sg13g2_dfrbp_1 \board_state[116]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net465),
    .D(_0627_),
    .Q_N(_0199_),
    .Q(\board_state[116] ));
 sg13g2_dfrbp_1 \board_state[117]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net466),
    .D(_0628_),
    .Q_N(_0200_),
    .Q(\board_state[117] ));
 sg13g2_dfrbp_1 \board_state[118]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net467),
    .D(_0629_),
    .Q_N(_0201_),
    .Q(\board_state[118] ));
 sg13g2_dfrbp_1 \board_state[119]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net468),
    .D(_0630_),
    .Q_N(_0202_),
    .Q(\board_state[119] ));
 sg13g2_dfrbp_1 \board_state[11]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net469),
    .D(_0631_),
    .Q_N(_0094_),
    .Q(\board_state[11] ));
 sg13g2_dfrbp_1 \board_state[120]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net470),
    .D(_0632_),
    .Q_N(_0203_),
    .Q(\board_state[120] ));
 sg13g2_dfrbp_1 \board_state[121]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net471),
    .D(_0633_),
    .Q_N(_0204_),
    .Q(\board_state[121] ));
 sg13g2_dfrbp_1 \board_state[122]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net472),
    .D(_0634_),
    .Q_N(_0205_),
    .Q(\board_state[122] ));
 sg13g2_dfrbp_1 \board_state[123]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net473),
    .D(_0635_),
    .Q_N(_0206_),
    .Q(\board_state[123] ));
 sg13g2_dfrbp_1 \board_state[124]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net474),
    .D(_0636_),
    .Q_N(_0207_),
    .Q(\board_state[124] ));
 sg13g2_dfrbp_1 \board_state[125]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net475),
    .D(_0637_),
    .Q_N(_0208_),
    .Q(\board_state[125] ));
 sg13g2_dfrbp_1 \board_state[126]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net476),
    .D(_0638_),
    .Q_N(_0209_),
    .Q(\board_state[126] ));
 sg13g2_dfrbp_1 \board_state[127]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net477),
    .D(_0639_),
    .Q_N(_0210_),
    .Q(\board_state[127] ));
 sg13g2_dfrbp_1 \board_state[128]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net478),
    .D(_0640_),
    .Q_N(_0211_),
    .Q(\board_state[128] ));
 sg13g2_dfrbp_1 \board_state[129]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net479),
    .D(_0641_),
    .Q_N(_0212_),
    .Q(\board_state[129] ));
 sg13g2_dfrbp_1 \board_state[12]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net480),
    .D(_0642_),
    .Q_N(_0095_),
    .Q(\board_state[12] ));
 sg13g2_dfrbp_1 \board_state[130]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net481),
    .D(_0643_),
    .Q_N(_0213_),
    .Q(\board_state[130] ));
 sg13g2_dfrbp_1 \board_state[131]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net482),
    .D(_0644_),
    .Q_N(_0214_),
    .Q(\board_state[131] ));
 sg13g2_dfrbp_1 \board_state[132]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net483),
    .D(_0645_),
    .Q_N(_0215_),
    .Q(\board_state[132] ));
 sg13g2_dfrbp_1 \board_state[133]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net484),
    .D(_0646_),
    .Q_N(_0216_),
    .Q(\board_state[133] ));
 sg13g2_dfrbp_1 \board_state[134]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net485),
    .D(_0647_),
    .Q_N(_0217_),
    .Q(\board_state[134] ));
 sg13g2_dfrbp_1 \board_state[135]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net486),
    .D(_0648_),
    .Q_N(_0218_),
    .Q(\board_state[135] ));
 sg13g2_dfrbp_1 \board_state[136]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net487),
    .D(_0649_),
    .Q_N(_0219_),
    .Q(\board_state[136] ));
 sg13g2_dfrbp_1 \board_state[137]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net488),
    .D(_0650_),
    .Q_N(_0220_),
    .Q(\board_state[137] ));
 sg13g2_dfrbp_1 \board_state[138]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net489),
    .D(_0651_),
    .Q_N(_0221_),
    .Q(\board_state[138] ));
 sg13g2_dfrbp_1 \board_state[139]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net490),
    .D(_0652_),
    .Q_N(_0222_),
    .Q(\board_state[139] ));
 sg13g2_dfrbp_1 \board_state[13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net491),
    .D(_0653_),
    .Q_N(_0096_),
    .Q(\board_state[13] ));
 sg13g2_dfrbp_1 \board_state[140]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net492),
    .D(_0654_),
    .Q_N(_0223_),
    .Q(\board_state[140] ));
 sg13g2_dfrbp_1 \board_state[141]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net493),
    .D(_0655_),
    .Q_N(_0224_),
    .Q(\board_state[141] ));
 sg13g2_dfrbp_1 \board_state[142]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net494),
    .D(_0656_),
    .Q_N(_0225_),
    .Q(\board_state[142] ));
 sg13g2_dfrbp_1 \board_state[143]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net495),
    .D(_0657_),
    .Q_N(_0226_),
    .Q(\board_state[143] ));
 sg13g2_dfrbp_1 \board_state[144]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net496),
    .D(_0658_),
    .Q_N(_0227_),
    .Q(\board_state[144] ));
 sg13g2_dfrbp_1 \board_state[145]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net497),
    .D(_0659_),
    .Q_N(_0228_),
    .Q(\board_state[145] ));
 sg13g2_dfrbp_1 \board_state[146]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net498),
    .D(_0660_),
    .Q_N(_0229_),
    .Q(\board_state[146] ));
 sg13g2_dfrbp_1 \board_state[147]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net499),
    .D(_0661_),
    .Q_N(_0230_),
    .Q(\board_state[147] ));
 sg13g2_dfrbp_1 \board_state[148]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net500),
    .D(_0662_),
    .Q_N(_0231_),
    .Q(\board_state[148] ));
 sg13g2_dfrbp_1 \board_state[149]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net501),
    .D(_0663_),
    .Q_N(_0232_),
    .Q(\board_state[149] ));
 sg13g2_dfrbp_1 \board_state[14]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net502),
    .D(_0664_),
    .Q_N(_0097_),
    .Q(\board_state[14] ));
 sg13g2_dfrbp_1 \board_state[150]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net503),
    .D(_0665_),
    .Q_N(_0233_),
    .Q(\board_state[150] ));
 sg13g2_dfrbp_1 \board_state[151]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net504),
    .D(_0666_),
    .Q_N(_0234_),
    .Q(\board_state[151] ));
 sg13g2_dfrbp_1 \board_state[152]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net505),
    .D(_0667_),
    .Q_N(_0235_),
    .Q(\board_state[152] ));
 sg13g2_dfrbp_1 \board_state[153]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net506),
    .D(_0668_),
    .Q_N(_0236_),
    .Q(\board_state[153] ));
 sg13g2_dfrbp_1 \board_state[154]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net507),
    .D(_0669_),
    .Q_N(_0237_),
    .Q(\board_state[154] ));
 sg13g2_dfrbp_1 \board_state[155]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net508),
    .D(_0670_),
    .Q_N(_0238_),
    .Q(\board_state[155] ));
 sg13g2_dfrbp_1 \board_state[156]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net509),
    .D(_0671_),
    .Q_N(_0239_),
    .Q(\board_state[156] ));
 sg13g2_dfrbp_1 \board_state[157]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net510),
    .D(_0672_),
    .Q_N(_0240_),
    .Q(\board_state[157] ));
 sg13g2_dfrbp_1 \board_state[158]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net511),
    .D(_0673_),
    .Q_N(_0241_),
    .Q(\board_state[158] ));
 sg13g2_dfrbp_1 \board_state[159]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net512),
    .D(_0674_),
    .Q_N(_0242_),
    .Q(\board_state[159] ));
 sg13g2_dfrbp_1 \board_state[15]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net513),
    .D(_0675_),
    .Q_N(_0098_),
    .Q(\board_state[15] ));
 sg13g2_dfrbp_1 \board_state[160]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net514),
    .D(_0676_),
    .Q_N(_0243_),
    .Q(\board_state[160] ));
 sg13g2_dfrbp_1 \board_state[161]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net515),
    .D(_0677_),
    .Q_N(_0244_),
    .Q(\board_state[161] ));
 sg13g2_dfrbp_1 \board_state[162]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net516),
    .D(_0678_),
    .Q_N(_0245_),
    .Q(\board_state[162] ));
 sg13g2_dfrbp_1 \board_state[163]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net517),
    .D(_0679_),
    .Q_N(_0246_),
    .Q(\board_state[163] ));
 sg13g2_dfrbp_1 \board_state[164]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net518),
    .D(_0680_),
    .Q_N(_0247_),
    .Q(\board_state[164] ));
 sg13g2_dfrbp_1 \board_state[165]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net519),
    .D(_0681_),
    .Q_N(_0248_),
    .Q(\board_state[165] ));
 sg13g2_dfrbp_1 \board_state[166]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net520),
    .D(_0682_),
    .Q_N(_0249_),
    .Q(\board_state[166] ));
 sg13g2_dfrbp_1 \board_state[167]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net521),
    .D(_0683_),
    .Q_N(_0250_),
    .Q(\board_state[167] ));
 sg13g2_dfrbp_1 \board_state[168]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net522),
    .D(_0684_),
    .Q_N(_0251_),
    .Q(\board_state[168] ));
 sg13g2_dfrbp_1 \board_state[169]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net523),
    .D(_0685_),
    .Q_N(_0252_),
    .Q(\board_state[169] ));
 sg13g2_dfrbp_1 \board_state[16]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net524),
    .D(_0686_),
    .Q_N(_0099_),
    .Q(\board_state[16] ));
 sg13g2_dfrbp_1 \board_state[170]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net525),
    .D(_0687_),
    .Q_N(_0253_),
    .Q(\board_state[170] ));
 sg13g2_dfrbp_1 \board_state[171]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net526),
    .D(_0688_),
    .Q_N(_0254_),
    .Q(\board_state[171] ));
 sg13g2_dfrbp_1 \board_state[172]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net527),
    .D(_0689_),
    .Q_N(_0255_),
    .Q(\board_state[172] ));
 sg13g2_dfrbp_1 \board_state[173]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net528),
    .D(_0690_),
    .Q_N(_0256_),
    .Q(\board_state[173] ));
 sg13g2_dfrbp_1 \board_state[174]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net529),
    .D(_0691_),
    .Q_N(_0257_),
    .Q(\board_state[174] ));
 sg13g2_dfrbp_1 \board_state[175]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net530),
    .D(_0692_),
    .Q_N(_0258_),
    .Q(\board_state[175] ));
 sg13g2_dfrbp_1 \board_state[176]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net531),
    .D(_0693_),
    .Q_N(_0259_),
    .Q(\board_state[176] ));
 sg13g2_dfrbp_1 \board_state[177]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net532),
    .D(_0694_),
    .Q_N(_0260_),
    .Q(\board_state[177] ));
 sg13g2_dfrbp_1 \board_state[178]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net533),
    .D(_0695_),
    .Q_N(_0261_),
    .Q(\board_state[178] ));
 sg13g2_dfrbp_1 \board_state[179]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net534),
    .D(_0696_),
    .Q_N(_0262_),
    .Q(\board_state[179] ));
 sg13g2_dfrbp_1 \board_state[17]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net535),
    .D(_0697_),
    .Q_N(_0100_),
    .Q(\board_state[17] ));
 sg13g2_dfrbp_1 \board_state[180]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net536),
    .D(_0698_),
    .Q_N(_0263_),
    .Q(\board_state[180] ));
 sg13g2_dfrbp_1 \board_state[181]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net537),
    .D(_0699_),
    .Q_N(_0264_),
    .Q(\board_state[181] ));
 sg13g2_dfrbp_1 \board_state[182]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net538),
    .D(_0700_),
    .Q_N(_0265_),
    .Q(\board_state[182] ));
 sg13g2_dfrbp_1 \board_state[183]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net539),
    .D(_0701_),
    .Q_N(_0266_),
    .Q(\board_state[183] ));
 sg13g2_dfrbp_1 \board_state[184]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net540),
    .D(_0702_),
    .Q_N(_0267_),
    .Q(\board_state[184] ));
 sg13g2_dfrbp_1 \board_state[185]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net541),
    .D(_0703_),
    .Q_N(_0268_),
    .Q(\board_state[185] ));
 sg13g2_dfrbp_1 \board_state[186]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net542),
    .D(_0704_),
    .Q_N(_0269_),
    .Q(\board_state[186] ));
 sg13g2_dfrbp_1 \board_state[187]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net543),
    .D(_0705_),
    .Q_N(_0270_),
    .Q(\board_state[187] ));
 sg13g2_dfrbp_1 \board_state[188]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net544),
    .D(_0706_),
    .Q_N(_0271_),
    .Q(\board_state[188] ));
 sg13g2_dfrbp_1 \board_state[189]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net545),
    .D(_0707_),
    .Q_N(_0272_),
    .Q(\board_state[189] ));
 sg13g2_dfrbp_1 \board_state[18]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net546),
    .D(_0708_),
    .Q_N(_0101_),
    .Q(\board_state[18] ));
 sg13g2_dfrbp_1 \board_state[190]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net547),
    .D(_0709_),
    .Q_N(_0273_),
    .Q(\board_state[190] ));
 sg13g2_dfrbp_1 \board_state[191]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net548),
    .D(_0710_),
    .Q_N(_0274_),
    .Q(\board_state[191] ));
 sg13g2_dfrbp_1 \board_state[192]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net549),
    .D(_0711_),
    .Q_N(_0275_),
    .Q(\board_state[192] ));
 sg13g2_dfrbp_1 \board_state[193]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net550),
    .D(_0712_),
    .Q_N(_0276_),
    .Q(\board_state[193] ));
 sg13g2_dfrbp_1 \board_state[194]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net551),
    .D(_0713_),
    .Q_N(_0277_),
    .Q(\board_state[194] ));
 sg13g2_dfrbp_1 \board_state[195]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net552),
    .D(_0714_),
    .Q_N(_0278_),
    .Q(\board_state[195] ));
 sg13g2_dfrbp_1 \board_state[196]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net553),
    .D(_0715_),
    .Q_N(_0279_),
    .Q(\board_state[196] ));
 sg13g2_dfrbp_1 \board_state[197]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net554),
    .D(_0716_),
    .Q_N(_0280_),
    .Q(\board_state[197] ));
 sg13g2_dfrbp_1 \board_state[198]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net555),
    .D(_0717_),
    .Q_N(_0281_),
    .Q(\board_state[198] ));
 sg13g2_dfrbp_1 \board_state[199]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net556),
    .D(_0718_),
    .Q_N(_0282_),
    .Q(\board_state[199] ));
 sg13g2_dfrbp_1 \board_state[19]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net557),
    .D(_0719_),
    .Q_N(_0102_),
    .Q(\board_state[19] ));
 sg13g2_dfrbp_1 \board_state[1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net558),
    .D(_0720_),
    .Q_N(_0083_),
    .Q(\board_state[1] ));
 sg13g2_dfrbp_1 \board_state[200]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net559),
    .D(_0721_),
    .Q_N(_0283_),
    .Q(\board_state[200] ));
 sg13g2_dfrbp_1 \board_state[201]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net560),
    .D(_0722_),
    .Q_N(_0284_),
    .Q(\board_state[201] ));
 sg13g2_dfrbp_1 \board_state[202]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net561),
    .D(_0723_),
    .Q_N(_0285_),
    .Q(\board_state[202] ));
 sg13g2_dfrbp_1 \board_state[203]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net562),
    .D(_0724_),
    .Q_N(_0286_),
    .Q(\board_state[203] ));
 sg13g2_dfrbp_1 \board_state[204]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net563),
    .D(_0725_),
    .Q_N(_0287_),
    .Q(\board_state[204] ));
 sg13g2_dfrbp_1 \board_state[205]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net564),
    .D(_0726_),
    .Q_N(_0288_),
    .Q(\board_state[205] ));
 sg13g2_dfrbp_1 \board_state[206]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net565),
    .D(_0727_),
    .Q_N(_0289_),
    .Q(\board_state[206] ));
 sg13g2_dfrbp_1 \board_state[207]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net566),
    .D(_0728_),
    .Q_N(_0290_),
    .Q(\board_state[207] ));
 sg13g2_dfrbp_1 \board_state[208]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net567),
    .D(_0729_),
    .Q_N(_0291_),
    .Q(\board_state[208] ));
 sg13g2_dfrbp_1 \board_state[209]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net568),
    .D(_0730_),
    .Q_N(_0292_),
    .Q(\board_state[209] ));
 sg13g2_dfrbp_1 \board_state[20]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net569),
    .D(_0731_),
    .Q_N(_0103_),
    .Q(\board_state[20] ));
 sg13g2_dfrbp_1 \board_state[210]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net570),
    .D(_0732_),
    .Q_N(_0293_),
    .Q(\board_state[210] ));
 sg13g2_dfrbp_1 \board_state[211]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net571),
    .D(_0733_),
    .Q_N(_0294_),
    .Q(\board_state[211] ));
 sg13g2_dfrbp_1 \board_state[212]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net572),
    .D(_0734_),
    .Q_N(_0295_),
    .Q(\board_state[212] ));
 sg13g2_dfrbp_1 \board_state[213]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net573),
    .D(_0735_),
    .Q_N(_0296_),
    .Q(\board_state[213] ));
 sg13g2_dfrbp_1 \board_state[214]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net574),
    .D(_0736_),
    .Q_N(_0297_),
    .Q(\board_state[214] ));
 sg13g2_dfrbp_1 \board_state[215]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net575),
    .D(_0737_),
    .Q_N(_0298_),
    .Q(\board_state[215] ));
 sg13g2_dfrbp_1 \board_state[216]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net576),
    .D(_0738_),
    .Q_N(_0299_),
    .Q(\board_state[216] ));
 sg13g2_dfrbp_1 \board_state[217]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net577),
    .D(_0739_),
    .Q_N(_0300_),
    .Q(\board_state[217] ));
 sg13g2_dfrbp_1 \board_state[218]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net578),
    .D(_0740_),
    .Q_N(_0301_),
    .Q(\board_state[218] ));
 sg13g2_dfrbp_1 \board_state[219]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net579),
    .D(_0741_),
    .Q_N(_0302_),
    .Q(\board_state[219] ));
 sg13g2_dfrbp_1 \board_state[21]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net580),
    .D(_0742_),
    .Q_N(_0104_),
    .Q(\board_state[21] ));
 sg13g2_dfrbp_1 \board_state[220]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net581),
    .D(_0743_),
    .Q_N(_0303_),
    .Q(\board_state[220] ));
 sg13g2_dfrbp_1 \board_state[221]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net582),
    .D(_0744_),
    .Q_N(_0304_),
    .Q(\board_state[221] ));
 sg13g2_dfrbp_1 \board_state[222]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net583),
    .D(_0745_),
    .Q_N(_0305_),
    .Q(\board_state[222] ));
 sg13g2_dfrbp_1 \board_state[223]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net584),
    .D(_0746_),
    .Q_N(_0306_),
    .Q(\board_state[223] ));
 sg13g2_dfrbp_1 \board_state[224]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net585),
    .D(_0747_),
    .Q_N(_0307_),
    .Q(\board_state[224] ));
 sg13g2_dfrbp_1 \board_state[225]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net586),
    .D(_0748_),
    .Q_N(_0308_),
    .Q(\board_state[225] ));
 sg13g2_dfrbp_1 \board_state[226]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net587),
    .D(_0749_),
    .Q_N(_0309_),
    .Q(\board_state[226] ));
 sg13g2_dfrbp_1 \board_state[227]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net588),
    .D(_0750_),
    .Q_N(_0310_),
    .Q(\board_state[227] ));
 sg13g2_dfrbp_1 \board_state[228]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net589),
    .D(_0751_),
    .Q_N(_0311_),
    .Q(\board_state[228] ));
 sg13g2_dfrbp_1 \board_state[229]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net590),
    .D(_0752_),
    .Q_N(_0312_),
    .Q(\board_state[229] ));
 sg13g2_dfrbp_1 \board_state[22]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net591),
    .D(_0753_),
    .Q_N(_0105_),
    .Q(\board_state[22] ));
 sg13g2_dfrbp_1 \board_state[230]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net592),
    .D(_0754_),
    .Q_N(_0313_),
    .Q(\board_state[230] ));
 sg13g2_dfrbp_1 \board_state[231]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net593),
    .D(_0755_),
    .Q_N(_0314_),
    .Q(\board_state[231] ));
 sg13g2_dfrbp_1 \board_state[232]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net594),
    .D(_0756_),
    .Q_N(_0315_),
    .Q(\board_state[232] ));
 sg13g2_dfrbp_1 \board_state[233]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net595),
    .D(_0757_),
    .Q_N(_0316_),
    .Q(\board_state[233] ));
 sg13g2_dfrbp_1 \board_state[234]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net596),
    .D(_0758_),
    .Q_N(_0317_),
    .Q(\board_state[234] ));
 sg13g2_dfrbp_1 \board_state[235]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net597),
    .D(_0759_),
    .Q_N(_0318_),
    .Q(\board_state[235] ));
 sg13g2_dfrbp_1 \board_state[236]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net598),
    .D(_0760_),
    .Q_N(_0319_),
    .Q(\board_state[236] ));
 sg13g2_dfrbp_1 \board_state[237]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net599),
    .D(_0761_),
    .Q_N(_0320_),
    .Q(\board_state[237] ));
 sg13g2_dfrbp_1 \board_state[238]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net600),
    .D(_0762_),
    .Q_N(_0321_),
    .Q(\board_state[238] ));
 sg13g2_dfrbp_1 \board_state[239]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net601),
    .D(_0763_),
    .Q_N(_0322_),
    .Q(\board_state[239] ));
 sg13g2_dfrbp_1 \board_state[23]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net602),
    .D(_0764_),
    .Q_N(_0106_),
    .Q(\board_state[23] ));
 sg13g2_dfrbp_1 \board_state[240]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net603),
    .D(_0765_),
    .Q_N(_0323_),
    .Q(\board_state[240] ));
 sg13g2_dfrbp_1 \board_state[241]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net604),
    .D(_0766_),
    .Q_N(_0324_),
    .Q(\board_state[241] ));
 sg13g2_dfrbp_1 \board_state[242]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net605),
    .D(_0767_),
    .Q_N(_0325_),
    .Q(\board_state[242] ));
 sg13g2_dfrbp_1 \board_state[243]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net606),
    .D(_0768_),
    .Q_N(_0326_),
    .Q(\board_state[243] ));
 sg13g2_dfrbp_1 \board_state[244]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net607),
    .D(_0769_),
    .Q_N(_0327_),
    .Q(\board_state[244] ));
 sg13g2_dfrbp_1 \board_state[245]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net608),
    .D(_0770_),
    .Q_N(_0328_),
    .Q(\board_state[245] ));
 sg13g2_dfrbp_1 \board_state[246]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net609),
    .D(_0771_),
    .Q_N(_0329_),
    .Q(\board_state[246] ));
 sg13g2_dfrbp_1 \board_state[247]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net610),
    .D(_0772_),
    .Q_N(_0330_),
    .Q(\board_state[247] ));
 sg13g2_dfrbp_1 \board_state[248]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net611),
    .D(_0773_),
    .Q_N(_0331_),
    .Q(\board_state[248] ));
 sg13g2_dfrbp_1 \board_state[249]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net612),
    .D(_0774_),
    .Q_N(_0332_),
    .Q(\board_state[249] ));
 sg13g2_dfrbp_1 \board_state[24]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net613),
    .D(_0775_),
    .Q_N(_0107_),
    .Q(\board_state[24] ));
 sg13g2_dfrbp_1 \board_state[250]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net614),
    .D(_0776_),
    .Q_N(_0333_),
    .Q(\board_state[250] ));
 sg13g2_dfrbp_1 \board_state[251]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net615),
    .D(_0777_),
    .Q_N(_0334_),
    .Q(\board_state[251] ));
 sg13g2_dfrbp_1 \board_state[252]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net616),
    .D(_0778_),
    .Q_N(_0335_),
    .Q(\board_state[252] ));
 sg13g2_dfrbp_1 \board_state[253]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net617),
    .D(_0779_),
    .Q_N(_0336_),
    .Q(\board_state[253] ));
 sg13g2_dfrbp_1 \board_state[254]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net618),
    .D(_0780_),
    .Q_N(_0337_),
    .Q(\board_state[254] ));
 sg13g2_dfrbp_1 \board_state[255]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net619),
    .D(_0781_),
    .Q_N(_0338_),
    .Q(\board_state[255] ));
 sg13g2_dfrbp_1 \board_state[256]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net620),
    .D(_0782_),
    .Q_N(_0339_),
    .Q(\board_state[256] ));
 sg13g2_dfrbp_1 \board_state[257]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net621),
    .D(_0783_),
    .Q_N(_0340_),
    .Q(\board_state[257] ));
 sg13g2_dfrbp_1 \board_state[258]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net622),
    .D(_0784_),
    .Q_N(_0341_),
    .Q(\board_state[258] ));
 sg13g2_dfrbp_1 \board_state[259]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net623),
    .D(_0785_),
    .Q_N(_0342_),
    .Q(\board_state[259] ));
 sg13g2_dfrbp_1 \board_state[25]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net624),
    .D(_0786_),
    .Q_N(_0108_),
    .Q(\board_state[25] ));
 sg13g2_dfrbp_1 \board_state[260]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net625),
    .D(_0787_),
    .Q_N(_0343_),
    .Q(\board_state[260] ));
 sg13g2_dfrbp_1 \board_state[261]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net626),
    .D(_0788_),
    .Q_N(_0344_),
    .Q(\board_state[261] ));
 sg13g2_dfrbp_1 \board_state[262]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net627),
    .D(_0789_),
    .Q_N(_0345_),
    .Q(\board_state[262] ));
 sg13g2_dfrbp_1 \board_state[263]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net628),
    .D(_0790_),
    .Q_N(_0346_),
    .Q(\board_state[263] ));
 sg13g2_dfrbp_1 \board_state[264]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net629),
    .D(_0791_),
    .Q_N(_0347_),
    .Q(\board_state[264] ));
 sg13g2_dfrbp_1 \board_state[265]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net630),
    .D(_0792_),
    .Q_N(_0348_),
    .Q(\board_state[265] ));
 sg13g2_dfrbp_1 \board_state[266]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net631),
    .D(_0793_),
    .Q_N(_0349_),
    .Q(\board_state[266] ));
 sg13g2_dfrbp_1 \board_state[267]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net632),
    .D(_0794_),
    .Q_N(_0350_),
    .Q(\board_state[267] ));
 sg13g2_dfrbp_1 \board_state[268]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net633),
    .D(_0795_),
    .Q_N(_0351_),
    .Q(\board_state[268] ));
 sg13g2_dfrbp_1 \board_state[269]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net634),
    .D(_0796_),
    .Q_N(_0352_),
    .Q(\board_state[269] ));
 sg13g2_dfrbp_1 \board_state[26]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net635),
    .D(_0797_),
    .Q_N(_0109_),
    .Q(\board_state[26] ));
 sg13g2_dfrbp_1 \board_state[270]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net636),
    .D(_0798_),
    .Q_N(_0353_),
    .Q(\board_state[270] ));
 sg13g2_dfrbp_1 \board_state[271]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net637),
    .D(_0799_),
    .Q_N(_0354_),
    .Q(\board_state[271] ));
 sg13g2_dfrbp_1 \board_state[272]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net638),
    .D(_0800_),
    .Q_N(_0355_),
    .Q(\board_state[272] ));
 sg13g2_dfrbp_1 \board_state[273]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net639),
    .D(_0801_),
    .Q_N(_0356_),
    .Q(\board_state[273] ));
 sg13g2_dfrbp_1 \board_state[274]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net640),
    .D(_0802_),
    .Q_N(_0357_),
    .Q(\board_state[274] ));
 sg13g2_dfrbp_1 \board_state[275]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net641),
    .D(_0803_),
    .Q_N(_0358_),
    .Q(\board_state[275] ));
 sg13g2_dfrbp_1 \board_state[276]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net642),
    .D(_0804_),
    .Q_N(_0359_),
    .Q(\board_state[276] ));
 sg13g2_dfrbp_1 \board_state[277]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net643),
    .D(_0805_),
    .Q_N(_0360_),
    .Q(\board_state[277] ));
 sg13g2_dfrbp_1 \board_state[278]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net644),
    .D(_0806_),
    .Q_N(_0361_),
    .Q(\board_state[278] ));
 sg13g2_dfrbp_1 \board_state[279]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net645),
    .D(_0807_),
    .Q_N(_0362_),
    .Q(\board_state[279] ));
 sg13g2_dfrbp_1 \board_state[27]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net646),
    .D(_0808_),
    .Q_N(_0110_),
    .Q(\board_state[27] ));
 sg13g2_dfrbp_1 \board_state[280]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net647),
    .D(_0809_),
    .Q_N(_0363_),
    .Q(\board_state[280] ));
 sg13g2_dfrbp_1 \board_state[281]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net648),
    .D(_0810_),
    .Q_N(_0364_),
    .Q(\board_state[281] ));
 sg13g2_dfrbp_1 \board_state[282]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net649),
    .D(_0811_),
    .Q_N(_0365_),
    .Q(\board_state[282] ));
 sg13g2_dfrbp_1 \board_state[283]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net650),
    .D(_0812_),
    .Q_N(_0366_),
    .Q(\board_state[283] ));
 sg13g2_dfrbp_1 \board_state[284]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net651),
    .D(_0813_),
    .Q_N(_0367_),
    .Q(\board_state[284] ));
 sg13g2_dfrbp_1 \board_state[285]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net652),
    .D(_0814_),
    .Q_N(_0368_),
    .Q(\board_state[285] ));
 sg13g2_dfrbp_1 \board_state[286]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net653),
    .D(_0815_),
    .Q_N(_0369_),
    .Q(\board_state[286] ));
 sg13g2_dfrbp_1 \board_state[287]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net654),
    .D(_0816_),
    .Q_N(_0370_),
    .Q(\board_state[287] ));
 sg13g2_dfrbp_1 \board_state[288]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net655),
    .D(_0817_),
    .Q_N(_0371_),
    .Q(\board_state[288] ));
 sg13g2_dfrbp_1 \board_state[289]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net656),
    .D(_0818_),
    .Q_N(_0372_),
    .Q(\board_state[289] ));
 sg13g2_dfrbp_1 \board_state[28]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net657),
    .D(_0819_),
    .Q_N(_0111_),
    .Q(\board_state[28] ));
 sg13g2_dfrbp_1 \board_state[290]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net658),
    .D(_0820_),
    .Q_N(_0373_),
    .Q(\board_state[290] ));
 sg13g2_dfrbp_1 \board_state[291]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net659),
    .D(_0821_),
    .Q_N(_0374_),
    .Q(\board_state[291] ));
 sg13g2_dfrbp_1 \board_state[292]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net660),
    .D(_0822_),
    .Q_N(_0375_),
    .Q(\board_state[292] ));
 sg13g2_dfrbp_1 \board_state[293]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net661),
    .D(_0823_),
    .Q_N(_0376_),
    .Q(\board_state[293] ));
 sg13g2_dfrbp_1 \board_state[294]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net662),
    .D(_0824_),
    .Q_N(_0377_),
    .Q(\board_state[294] ));
 sg13g2_dfrbp_1 \board_state[295]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net663),
    .D(_0825_),
    .Q_N(_0378_),
    .Q(\board_state[295] ));
 sg13g2_dfrbp_1 \board_state[296]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net664),
    .D(_0826_),
    .Q_N(_0379_),
    .Q(\board_state[296] ));
 sg13g2_dfrbp_1 \board_state[297]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net665),
    .D(_0827_),
    .Q_N(_0380_),
    .Q(\board_state[297] ));
 sg13g2_dfrbp_1 \board_state[298]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net666),
    .D(_0828_),
    .Q_N(_0381_),
    .Q(\board_state[298] ));
 sg13g2_dfrbp_1 \board_state[299]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net667),
    .D(_0829_),
    .Q_N(_0382_),
    .Q(\board_state[299] ));
 sg13g2_dfrbp_1 \board_state[29]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net668),
    .D(_0830_),
    .Q_N(_0112_),
    .Q(\board_state[29] ));
 sg13g2_dfrbp_1 \board_state[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net669),
    .D(_0831_),
    .Q_N(_0085_),
    .Q(\board_state[2] ));
 sg13g2_dfrbp_1 \board_state[300]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net670),
    .D(_0832_),
    .Q_N(_0383_),
    .Q(\board_state[300] ));
 sg13g2_dfrbp_1 \board_state[301]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net671),
    .D(_0833_),
    .Q_N(_0384_),
    .Q(\board_state[301] ));
 sg13g2_dfrbp_1 \board_state[302]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net672),
    .D(_0834_),
    .Q_N(_0385_),
    .Q(\board_state[302] ));
 sg13g2_dfrbp_1 \board_state[303]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net673),
    .D(_0835_),
    .Q_N(_0386_),
    .Q(\board_state[303] ));
 sg13g2_dfrbp_1 \board_state[304]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net674),
    .D(_0836_),
    .Q_N(_0387_),
    .Q(\board_state[304] ));
 sg13g2_dfrbp_1 \board_state[305]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net675),
    .D(_0837_),
    .Q_N(_0388_),
    .Q(\board_state[305] ));
 sg13g2_dfrbp_1 \board_state[306]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net676),
    .D(_0838_),
    .Q_N(_0389_),
    .Q(\board_state[306] ));
 sg13g2_dfrbp_1 \board_state[307]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net677),
    .D(_0839_),
    .Q_N(_0390_),
    .Q(\board_state[307] ));
 sg13g2_dfrbp_1 \board_state[308]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net678),
    .D(_0840_),
    .Q_N(_0391_),
    .Q(\board_state[308] ));
 sg13g2_dfrbp_1 \board_state[309]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net679),
    .D(_0841_),
    .Q_N(_0392_),
    .Q(\board_state[309] ));
 sg13g2_dfrbp_1 \board_state[30]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net680),
    .D(_0842_),
    .Q_N(_0113_),
    .Q(\board_state[30] ));
 sg13g2_dfrbp_1 \board_state[310]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net681),
    .D(_0843_),
    .Q_N(_0393_),
    .Q(\board_state[310] ));
 sg13g2_dfrbp_1 \board_state[311]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net682),
    .D(_0844_),
    .Q_N(_0394_),
    .Q(\board_state[311] ));
 sg13g2_dfrbp_1 \board_state[312]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net683),
    .D(_0845_),
    .Q_N(_0395_),
    .Q(\board_state[312] ));
 sg13g2_dfrbp_1 \board_state[313]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net684),
    .D(_0846_),
    .Q_N(_0396_),
    .Q(\board_state[313] ));
 sg13g2_dfrbp_1 \board_state[314]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net685),
    .D(_0847_),
    .Q_N(_0397_),
    .Q(\board_state[314] ));
 sg13g2_dfrbp_1 \board_state[315]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net686),
    .D(_0848_),
    .Q_N(_0398_),
    .Q(\board_state[315] ));
 sg13g2_dfrbp_1 \board_state[316]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net687),
    .D(_0849_),
    .Q_N(_0399_),
    .Q(\board_state[316] ));
 sg13g2_dfrbp_1 \board_state[317]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net688),
    .D(_0850_),
    .Q_N(_0400_),
    .Q(\board_state[317] ));
 sg13g2_dfrbp_1 \board_state[318]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net689),
    .D(_0851_),
    .Q_N(_0401_),
    .Q(\board_state[318] ));
 sg13g2_dfrbp_1 \board_state[319]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net690),
    .D(_0852_),
    .Q_N(_0402_),
    .Q(\board_state[319] ));
 sg13g2_dfrbp_1 \board_state[31]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net691),
    .D(_0853_),
    .Q_N(_0114_),
    .Q(\board_state[31] ));
 sg13g2_dfrbp_1 \board_state[320]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net692),
    .D(_0854_),
    .Q_N(_0403_),
    .Q(\board_state[320] ));
 sg13g2_dfrbp_1 \board_state[321]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net693),
    .D(_0855_),
    .Q_N(_0404_),
    .Q(\board_state[321] ));
 sg13g2_dfrbp_1 \board_state[322]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net694),
    .D(_0856_),
    .Q_N(_0405_),
    .Q(\board_state[322] ));
 sg13g2_dfrbp_1 \board_state[323]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net695),
    .D(_0857_),
    .Q_N(_0406_),
    .Q(\board_state[323] ));
 sg13g2_dfrbp_1 \board_state[324]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net696),
    .D(_0858_),
    .Q_N(_0407_),
    .Q(\board_state[324] ));
 sg13g2_dfrbp_1 \board_state[325]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net697),
    .D(_0859_),
    .Q_N(_0408_),
    .Q(\board_state[325] ));
 sg13g2_dfrbp_1 \board_state[326]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net698),
    .D(_0860_),
    .Q_N(_0409_),
    .Q(\board_state[326] ));
 sg13g2_dfrbp_1 \board_state[327]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net699),
    .D(_0861_),
    .Q_N(_0410_),
    .Q(\board_state[327] ));
 sg13g2_dfrbp_1 \board_state[328]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net700),
    .D(_0862_),
    .Q_N(_0411_),
    .Q(\board_state[328] ));
 sg13g2_dfrbp_1 \board_state[329]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net701),
    .D(_0863_),
    .Q_N(_0412_),
    .Q(\board_state[329] ));
 sg13g2_dfrbp_1 \board_state[32]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net702),
    .D(_0864_),
    .Q_N(_0115_),
    .Q(\board_state[32] ));
 sg13g2_dfrbp_1 \board_state[330]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net703),
    .D(_0865_),
    .Q_N(_0413_),
    .Q(\board_state[330] ));
 sg13g2_dfrbp_1 \board_state[331]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net704),
    .D(_0866_),
    .Q_N(_0414_),
    .Q(\board_state[331] ));
 sg13g2_dfrbp_1 \board_state[332]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net705),
    .D(_0867_),
    .Q_N(_0415_),
    .Q(\board_state[332] ));
 sg13g2_dfrbp_1 \board_state[333]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net706),
    .D(_0868_),
    .Q_N(_0416_),
    .Q(\board_state[333] ));
 sg13g2_dfrbp_1 \board_state[334]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net707),
    .D(_0869_),
    .Q_N(_0417_),
    .Q(\board_state[334] ));
 sg13g2_dfrbp_1 \board_state[335]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net708),
    .D(_0870_),
    .Q_N(_0418_),
    .Q(\board_state[335] ));
 sg13g2_dfrbp_1 \board_state[336]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net709),
    .D(_0871_),
    .Q_N(_0419_),
    .Q(\board_state[336] ));
 sg13g2_dfrbp_1 \board_state[337]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net710),
    .D(_0872_),
    .Q_N(_0420_),
    .Q(\board_state[337] ));
 sg13g2_dfrbp_1 \board_state[338]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net711),
    .D(_0873_),
    .Q_N(_0421_),
    .Q(\board_state[338] ));
 sg13g2_dfrbp_1 \board_state[339]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net712),
    .D(_0874_),
    .Q_N(_0422_),
    .Q(\board_state[339] ));
 sg13g2_dfrbp_1 \board_state[33]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net713),
    .D(_0875_),
    .Q_N(_0116_),
    .Q(\board_state[33] ));
 sg13g2_dfrbp_1 \board_state[340]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net714),
    .D(_0876_),
    .Q_N(_0423_),
    .Q(\board_state[340] ));
 sg13g2_dfrbp_1 \board_state[341]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net715),
    .D(_0877_),
    .Q_N(_0424_),
    .Q(\board_state[341] ));
 sg13g2_dfrbp_1 \board_state[342]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net716),
    .D(_0878_),
    .Q_N(_0425_),
    .Q(\board_state[342] ));
 sg13g2_dfrbp_1 \board_state[343]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net717),
    .D(_0879_),
    .Q_N(_0426_),
    .Q(\board_state[343] ));
 sg13g2_dfrbp_1 \board_state[344]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net718),
    .D(_0880_),
    .Q_N(_0427_),
    .Q(\board_state[344] ));
 sg13g2_dfrbp_1 \board_state[345]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net719),
    .D(_0881_),
    .Q_N(_0428_),
    .Q(\board_state[345] ));
 sg13g2_dfrbp_1 \board_state[346]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net720),
    .D(_0882_),
    .Q_N(_0429_),
    .Q(\board_state[346] ));
 sg13g2_dfrbp_1 \board_state[347]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net721),
    .D(_0883_),
    .Q_N(_0430_),
    .Q(\board_state[347] ));
 sg13g2_dfrbp_1 \board_state[348]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net722),
    .D(_0884_),
    .Q_N(_0431_),
    .Q(\board_state[348] ));
 sg13g2_dfrbp_1 \board_state[349]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net723),
    .D(_0885_),
    .Q_N(_0432_),
    .Q(\board_state[349] ));
 sg13g2_dfrbp_1 \board_state[34]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net724),
    .D(_0886_),
    .Q_N(_0117_),
    .Q(\board_state[34] ));
 sg13g2_dfrbp_1 \board_state[350]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net725),
    .D(_0887_),
    .Q_N(_0433_),
    .Q(\board_state[350] ));
 sg13g2_dfrbp_1 \board_state[351]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net726),
    .D(_0888_),
    .Q_N(_0434_),
    .Q(\board_state[351] ));
 sg13g2_dfrbp_1 \board_state[352]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net727),
    .D(_0889_),
    .Q_N(_0435_),
    .Q(\board_state[352] ));
 sg13g2_dfrbp_1 \board_state[353]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net728),
    .D(_0890_),
    .Q_N(_0436_),
    .Q(\board_state[353] ));
 sg13g2_dfrbp_1 \board_state[354]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net729),
    .D(_0891_),
    .Q_N(_0437_),
    .Q(\board_state[354] ));
 sg13g2_dfrbp_1 \board_state[355]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net730),
    .D(_0892_),
    .Q_N(_0438_),
    .Q(\board_state[355] ));
 sg13g2_dfrbp_1 \board_state[356]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net731),
    .D(_0893_),
    .Q_N(_0439_),
    .Q(\board_state[356] ));
 sg13g2_dfrbp_1 \board_state[357]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net732),
    .D(_0894_),
    .Q_N(_0440_),
    .Q(\board_state[357] ));
 sg13g2_dfrbp_1 \board_state[358]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net733),
    .D(_0895_),
    .Q_N(_0441_),
    .Q(\board_state[358] ));
 sg13g2_dfrbp_1 \board_state[359]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net734),
    .D(_0896_),
    .Q_N(_0442_),
    .Q(\board_state[359] ));
 sg13g2_dfrbp_1 \board_state[35]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net735),
    .D(_0897_),
    .Q_N(_0118_),
    .Q(\board_state[35] ));
 sg13g2_dfrbp_1 \board_state[360]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net736),
    .D(_0898_),
    .Q_N(_0443_),
    .Q(\board_state[360] ));
 sg13g2_dfrbp_1 \board_state[361]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net737),
    .D(_0899_),
    .Q_N(_0444_),
    .Q(\board_state[361] ));
 sg13g2_dfrbp_1 \board_state[362]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net738),
    .D(_0900_),
    .Q_N(_0445_),
    .Q(\board_state[362] ));
 sg13g2_dfrbp_1 \board_state[363]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net739),
    .D(_0901_),
    .Q_N(_0446_),
    .Q(\board_state[363] ));
 sg13g2_dfrbp_1 \board_state[364]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net740),
    .D(_0902_),
    .Q_N(_0447_),
    .Q(\board_state[364] ));
 sg13g2_dfrbp_1 \board_state[365]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net741),
    .D(_0903_),
    .Q_N(_0448_),
    .Q(\board_state[365] ));
 sg13g2_dfrbp_1 \board_state[366]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net742),
    .D(_0904_),
    .Q_N(_0449_),
    .Q(\board_state[366] ));
 sg13g2_dfrbp_1 \board_state[367]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net743),
    .D(_0905_),
    .Q_N(_0450_),
    .Q(\board_state[367] ));
 sg13g2_dfrbp_1 \board_state[368]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net744),
    .D(_0906_),
    .Q_N(_0451_),
    .Q(\board_state[368] ));
 sg13g2_dfrbp_1 \board_state[369]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net745),
    .D(_0907_),
    .Q_N(_0452_),
    .Q(\board_state[369] ));
 sg13g2_dfrbp_1 \board_state[36]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net746),
    .D(_0908_),
    .Q_N(_0119_),
    .Q(\board_state[36] ));
 sg13g2_dfrbp_1 \board_state[370]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net747),
    .D(_0909_),
    .Q_N(_0453_),
    .Q(\board_state[370] ));
 sg13g2_dfrbp_1 \board_state[371]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net748),
    .D(_0910_),
    .Q_N(_0454_),
    .Q(\board_state[371] ));
 sg13g2_dfrbp_1 \board_state[372]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net749),
    .D(_0911_),
    .Q_N(_0455_),
    .Q(\board_state[372] ));
 sg13g2_dfrbp_1 \board_state[373]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net750),
    .D(_0912_),
    .Q_N(_0456_),
    .Q(\board_state[373] ));
 sg13g2_dfrbp_1 \board_state[374]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net751),
    .D(_0913_),
    .Q_N(_0457_),
    .Q(\board_state[374] ));
 sg13g2_dfrbp_1 \board_state[375]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net752),
    .D(_0914_),
    .Q_N(_0458_),
    .Q(\board_state[375] ));
 sg13g2_dfrbp_1 \board_state[376]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net753),
    .D(_0915_),
    .Q_N(_0459_),
    .Q(\board_state[376] ));
 sg13g2_dfrbp_1 \board_state[377]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net754),
    .D(_0916_),
    .Q_N(_0460_),
    .Q(\board_state[377] ));
 sg13g2_dfrbp_1 \board_state[378]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net755),
    .D(_0917_),
    .Q_N(_0461_),
    .Q(\board_state[378] ));
 sg13g2_dfrbp_1 \board_state[379]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net756),
    .D(_0918_),
    .Q_N(_0462_),
    .Q(\board_state[379] ));
 sg13g2_dfrbp_1 \board_state[37]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net757),
    .D(_0919_),
    .Q_N(_0120_),
    .Q(\board_state[37] ));
 sg13g2_dfrbp_1 \board_state[380]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net758),
    .D(_0920_),
    .Q_N(_0463_),
    .Q(\board_state[380] ));
 sg13g2_dfrbp_1 \board_state[381]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net759),
    .D(_0921_),
    .Q_N(_0464_),
    .Q(\board_state[381] ));
 sg13g2_dfrbp_1 \board_state[382]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net760),
    .D(_0922_),
    .Q_N(_0465_),
    .Q(\board_state[382] ));
 sg13g2_dfrbp_1 \board_state[383]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net761),
    .D(_0923_),
    .Q_N(_0466_),
    .Q(\board_state[383] ));
 sg13g2_dfrbp_1 \board_state[384]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net762),
    .D(_0924_),
    .Q_N(_0467_),
    .Q(\board_state[384] ));
 sg13g2_dfrbp_1 \board_state[385]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net763),
    .D(_0925_),
    .Q_N(_0468_),
    .Q(\board_state[385] ));
 sg13g2_dfrbp_1 \board_state[386]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net764),
    .D(_0926_),
    .Q_N(_0469_),
    .Q(\board_state[386] ));
 sg13g2_dfrbp_1 \board_state[387]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net765),
    .D(_0927_),
    .Q_N(_0470_),
    .Q(\board_state[387] ));
 sg13g2_dfrbp_1 \board_state[388]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net766),
    .D(_0928_),
    .Q_N(_0471_),
    .Q(\board_state[388] ));
 sg13g2_dfrbp_1 \board_state[389]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net767),
    .D(_0929_),
    .Q_N(_0472_),
    .Q(\board_state[389] ));
 sg13g2_dfrbp_1 \board_state[38]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net768),
    .D(_0930_),
    .Q_N(_0121_),
    .Q(\board_state[38] ));
 sg13g2_dfrbp_1 \board_state[390]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net769),
    .D(_0931_),
    .Q_N(_0473_),
    .Q(\board_state[390] ));
 sg13g2_dfrbp_1 \board_state[391]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net770),
    .D(_0932_),
    .Q_N(_0474_),
    .Q(\board_state[391] ));
 sg13g2_dfrbp_1 \board_state[392]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net771),
    .D(_0933_),
    .Q_N(_0475_),
    .Q(\board_state[392] ));
 sg13g2_dfrbp_1 \board_state[393]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net772),
    .D(_0934_),
    .Q_N(_0476_),
    .Q(\board_state[393] ));
 sg13g2_dfrbp_1 \board_state[394]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net773),
    .D(_0935_),
    .Q_N(_0477_),
    .Q(\board_state[394] ));
 sg13g2_dfrbp_1 \board_state[395]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net774),
    .D(_0936_),
    .Q_N(_0478_),
    .Q(\board_state[395] ));
 sg13g2_dfrbp_1 \board_state[396]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net775),
    .D(_0937_),
    .Q_N(_0479_),
    .Q(\board_state[396] ));
 sg13g2_dfrbp_1 \board_state[397]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net776),
    .D(_0938_),
    .Q_N(_0480_),
    .Q(\board_state[397] ));
 sg13g2_dfrbp_1 \board_state[398]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net777),
    .D(_0939_),
    .Q_N(_0481_),
    .Q(\board_state[398] ));
 sg13g2_dfrbp_1 \board_state[399]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net778),
    .D(_0940_),
    .Q_N(_0482_),
    .Q(\board_state[399] ));
 sg13g2_dfrbp_1 \board_state[39]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net779),
    .D(_0941_),
    .Q_N(_0122_),
    .Q(\board_state[39] ));
 sg13g2_dfrbp_1 \board_state[3]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net780),
    .D(_0942_),
    .Q_N(_0086_),
    .Q(\board_state[3] ));
 sg13g2_dfrbp_1 \board_state[400]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net781),
    .D(_0943_),
    .Q_N(_0483_),
    .Q(\board_state[400] ));
 sg13g2_dfrbp_1 \board_state[401]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net782),
    .D(_0944_),
    .Q_N(_0484_),
    .Q(\board_state[401] ));
 sg13g2_dfrbp_1 \board_state[402]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net783),
    .D(_0945_),
    .Q_N(_0485_),
    .Q(\board_state[402] ));
 sg13g2_dfrbp_1 \board_state[403]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net784),
    .D(_0946_),
    .Q_N(_0486_),
    .Q(\board_state[403] ));
 sg13g2_dfrbp_1 \board_state[404]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net785),
    .D(_0947_),
    .Q_N(_0487_),
    .Q(\board_state[404] ));
 sg13g2_dfrbp_1 \board_state[405]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net786),
    .D(_0948_),
    .Q_N(_0488_),
    .Q(\board_state[405] ));
 sg13g2_dfrbp_1 \board_state[406]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net787),
    .D(_0949_),
    .Q_N(_0489_),
    .Q(\board_state[406] ));
 sg13g2_dfrbp_1 \board_state[407]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net788),
    .D(_0950_),
    .Q_N(_0490_),
    .Q(\board_state[407] ));
 sg13g2_dfrbp_1 \board_state[408]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net789),
    .D(_0951_),
    .Q_N(_0491_),
    .Q(\board_state[408] ));
 sg13g2_dfrbp_1 \board_state[409]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net790),
    .D(_0952_),
    .Q_N(_0492_),
    .Q(\board_state[409] ));
 sg13g2_dfrbp_1 \board_state[40]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net791),
    .D(_0953_),
    .Q_N(_0123_),
    .Q(\board_state[40] ));
 sg13g2_dfrbp_1 \board_state[410]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net792),
    .D(_0954_),
    .Q_N(_0493_),
    .Q(\board_state[410] ));
 sg13g2_dfrbp_1 \board_state[411]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net793),
    .D(_0955_),
    .Q_N(_0494_),
    .Q(\board_state[411] ));
 sg13g2_dfrbp_1 \board_state[412]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net794),
    .D(_0956_),
    .Q_N(_0495_),
    .Q(\board_state[412] ));
 sg13g2_dfrbp_1 \board_state[413]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net795),
    .D(_0957_),
    .Q_N(_0496_),
    .Q(\board_state[413] ));
 sg13g2_dfrbp_1 \board_state[414]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net796),
    .D(_0958_),
    .Q_N(_0497_),
    .Q(\board_state[414] ));
 sg13g2_dfrbp_1 \board_state[415]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net797),
    .D(_0959_),
    .Q_N(_0498_),
    .Q(\board_state[415] ));
 sg13g2_dfrbp_1 \board_state[416]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net798),
    .D(_0960_),
    .Q_N(_0499_),
    .Q(\board_state[416] ));
 sg13g2_dfrbp_1 \board_state[417]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net799),
    .D(_0961_),
    .Q_N(_0500_),
    .Q(\board_state[417] ));
 sg13g2_dfrbp_1 \board_state[418]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net800),
    .D(_0962_),
    .Q_N(_0501_),
    .Q(\board_state[418] ));
 sg13g2_dfrbp_1 \board_state[419]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net801),
    .D(_0963_),
    .Q_N(_0502_),
    .Q(\board_state[419] ));
 sg13g2_dfrbp_1 \board_state[41]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net802),
    .D(_0964_),
    .Q_N(_0124_),
    .Q(\board_state[41] ));
 sg13g2_dfrbp_1 \board_state[420]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net803),
    .D(_0965_),
    .Q_N(_0503_),
    .Q(\board_state[420] ));
 sg13g2_dfrbp_1 \board_state[421]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net804),
    .D(_0966_),
    .Q_N(_0504_),
    .Q(\board_state[421] ));
 sg13g2_dfrbp_1 \board_state[422]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net805),
    .D(_0967_),
    .Q_N(_0505_),
    .Q(\board_state[422] ));
 sg13g2_dfrbp_1 \board_state[423]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net806),
    .D(_0968_),
    .Q_N(_0506_),
    .Q(\board_state[423] ));
 sg13g2_dfrbp_1 \board_state[424]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net807),
    .D(_0969_),
    .Q_N(_0507_),
    .Q(\board_state[424] ));
 sg13g2_dfrbp_1 \board_state[425]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net808),
    .D(_0970_),
    .Q_N(_0508_),
    .Q(\board_state[425] ));
 sg13g2_dfrbp_1 \board_state[426]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net809),
    .D(_0971_),
    .Q_N(_0509_),
    .Q(\board_state[426] ));
 sg13g2_dfrbp_1 \board_state[427]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net810),
    .D(_0972_),
    .Q_N(_0510_),
    .Q(\board_state[427] ));
 sg13g2_dfrbp_1 \board_state[428]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net811),
    .D(_0973_),
    .Q_N(_0511_),
    .Q(\board_state[428] ));
 sg13g2_dfrbp_1 \board_state[429]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net812),
    .D(_0974_),
    .Q_N(_0512_),
    .Q(\board_state[429] ));
 sg13g2_dfrbp_1 \board_state[42]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net813),
    .D(_0975_),
    .Q_N(_0125_),
    .Q(\board_state[42] ));
 sg13g2_dfrbp_1 \board_state[430]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net814),
    .D(_0976_),
    .Q_N(_0513_),
    .Q(\board_state[430] ));
 sg13g2_dfrbp_1 \board_state[431]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net815),
    .D(_0977_),
    .Q_N(_0514_),
    .Q(\board_state[431] ));
 sg13g2_dfrbp_1 \board_state[432]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net816),
    .D(_0978_),
    .Q_N(_0515_),
    .Q(\board_state[432] ));
 sg13g2_dfrbp_1 \board_state[433]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net817),
    .D(_0979_),
    .Q_N(_0516_),
    .Q(\board_state[433] ));
 sg13g2_dfrbp_1 \board_state[434]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net818),
    .D(_0980_),
    .Q_N(_0517_),
    .Q(\board_state[434] ));
 sg13g2_dfrbp_1 \board_state[435]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net819),
    .D(_0981_),
    .Q_N(_0518_),
    .Q(\board_state[435] ));
 sg13g2_dfrbp_1 \board_state[436]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net820),
    .D(_0982_),
    .Q_N(_0519_),
    .Q(\board_state[436] ));
 sg13g2_dfrbp_1 \board_state[437]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net821),
    .D(_0983_),
    .Q_N(_0520_),
    .Q(\board_state[437] ));
 sg13g2_dfrbp_1 \board_state[438]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net822),
    .D(_0984_),
    .Q_N(_0521_),
    .Q(\board_state[438] ));
 sg13g2_dfrbp_1 \board_state[439]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net823),
    .D(_0985_),
    .Q_N(_0522_),
    .Q(\board_state[439] ));
 sg13g2_dfrbp_1 \board_state[43]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net824),
    .D(_0986_),
    .Q_N(_0126_),
    .Q(\board_state[43] ));
 sg13g2_dfrbp_1 \board_state[440]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net825),
    .D(_0987_),
    .Q_N(_0523_),
    .Q(\board_state[440] ));
 sg13g2_dfrbp_1 \board_state[441]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net826),
    .D(_0988_),
    .Q_N(_0524_),
    .Q(\board_state[441] ));
 sg13g2_dfrbp_1 \board_state[442]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net827),
    .D(_0989_),
    .Q_N(_0525_),
    .Q(\board_state[442] ));
 sg13g2_dfrbp_1 \board_state[443]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net828),
    .D(_0990_),
    .Q_N(_0526_),
    .Q(\board_state[443] ));
 sg13g2_dfrbp_1 \board_state[444]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net829),
    .D(_0991_),
    .Q_N(_0527_),
    .Q(\board_state[444] ));
 sg13g2_dfrbp_1 \board_state[445]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net830),
    .D(_0992_),
    .Q_N(_0528_),
    .Q(\board_state[445] ));
 sg13g2_dfrbp_1 \board_state[446]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net831),
    .D(_0993_),
    .Q_N(_0529_),
    .Q(\board_state[446] ));
 sg13g2_dfrbp_1 \board_state[447]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net832),
    .D(_0994_),
    .Q_N(_0530_),
    .Q(\board_state[447] ));
 sg13g2_dfrbp_1 \board_state[448]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net833),
    .D(_0995_),
    .Q_N(_0531_),
    .Q(\board_state[448] ));
 sg13g2_dfrbp_1 \board_state[449]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net834),
    .D(_0996_),
    .Q_N(_0532_),
    .Q(\board_state[449] ));
 sg13g2_dfrbp_1 \board_state[44]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net835),
    .D(_0997_),
    .Q_N(_0127_),
    .Q(\board_state[44] ));
 sg13g2_dfrbp_1 \board_state[450]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net836),
    .D(_0998_),
    .Q_N(_0533_),
    .Q(\board_state[450] ));
 sg13g2_dfrbp_1 \board_state[451]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net837),
    .D(_0999_),
    .Q_N(_0534_),
    .Q(\board_state[451] ));
 sg13g2_dfrbp_1 \board_state[452]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net838),
    .D(_1000_),
    .Q_N(_0535_),
    .Q(\board_state[452] ));
 sg13g2_dfrbp_1 \board_state[453]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net839),
    .D(_1001_),
    .Q_N(_0536_),
    .Q(\board_state[453] ));
 sg13g2_dfrbp_1 \board_state[454]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net840),
    .D(_1002_),
    .Q_N(_0537_),
    .Q(\board_state[454] ));
 sg13g2_dfrbp_1 \board_state[455]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net841),
    .D(_1003_),
    .Q_N(_0538_),
    .Q(\board_state[455] ));
 sg13g2_dfrbp_1 \board_state[456]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net842),
    .D(_1004_),
    .Q_N(_0539_),
    .Q(\board_state[456] ));
 sg13g2_dfrbp_1 \board_state[457]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net843),
    .D(_1005_),
    .Q_N(_0540_),
    .Q(\board_state[457] ));
 sg13g2_dfrbp_1 \board_state[458]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net844),
    .D(_1006_),
    .Q_N(_0541_),
    .Q(\board_state[458] ));
 sg13g2_dfrbp_1 \board_state[459]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net845),
    .D(_1007_),
    .Q_N(_0542_),
    .Q(\board_state[459] ));
 sg13g2_dfrbp_1 \board_state[45]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net846),
    .D(_1008_),
    .Q_N(_0128_),
    .Q(\board_state[45] ));
 sg13g2_dfrbp_1 \board_state[460]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net847),
    .D(_1009_),
    .Q_N(_0543_),
    .Q(\board_state[460] ));
 sg13g2_dfrbp_1 \board_state[461]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net848),
    .D(_1010_),
    .Q_N(_0544_),
    .Q(\board_state[461] ));
 sg13g2_dfrbp_1 \board_state[462]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net849),
    .D(_1011_),
    .Q_N(_0545_),
    .Q(\board_state[462] ));
 sg13g2_dfrbp_1 \board_state[463]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net850),
    .D(_1012_),
    .Q_N(_0546_),
    .Q(\board_state[463] ));
 sg13g2_dfrbp_1 \board_state[464]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net851),
    .D(_1013_),
    .Q_N(_0547_),
    .Q(\board_state[464] ));
 sg13g2_dfrbp_1 \board_state[465]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net852),
    .D(_1014_),
    .Q_N(_0548_),
    .Q(\board_state[465] ));
 sg13g2_dfrbp_1 \board_state[466]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net853),
    .D(_1015_),
    .Q_N(_0549_),
    .Q(\board_state[466] ));
 sg13g2_dfrbp_1 \board_state[467]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net854),
    .D(_1016_),
    .Q_N(_0550_),
    .Q(\board_state[467] ));
 sg13g2_dfrbp_1 \board_state[468]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net855),
    .D(_1017_),
    .Q_N(_0551_),
    .Q(\board_state[468] ));
 sg13g2_dfrbp_1 \board_state[469]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net856),
    .D(_1018_),
    .Q_N(_0552_),
    .Q(\board_state[469] ));
 sg13g2_dfrbp_1 \board_state[46]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net857),
    .D(_1019_),
    .Q_N(_0129_),
    .Q(\board_state[46] ));
 sg13g2_dfrbp_1 \board_state[470]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net858),
    .D(_1020_),
    .Q_N(_0553_),
    .Q(\board_state[470] ));
 sg13g2_dfrbp_1 \board_state[471]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net859),
    .D(_1021_),
    .Q_N(_0554_),
    .Q(\board_state[471] ));
 sg13g2_dfrbp_1 \board_state[472]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net860),
    .D(_1022_),
    .Q_N(_0555_),
    .Q(\board_state[472] ));
 sg13g2_dfrbp_1 \board_state[473]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net861),
    .D(_1023_),
    .Q_N(_0556_),
    .Q(\board_state[473] ));
 sg13g2_dfrbp_1 \board_state[474]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net862),
    .D(_1024_),
    .Q_N(_0557_),
    .Q(\board_state[474] ));
 sg13g2_dfrbp_1 \board_state[475]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net863),
    .D(_1025_),
    .Q_N(_0558_),
    .Q(\board_state[475] ));
 sg13g2_dfrbp_1 \board_state[476]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net864),
    .D(_1026_),
    .Q_N(_0559_),
    .Q(\board_state[476] ));
 sg13g2_dfrbp_1 \board_state[477]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net865),
    .D(_1027_),
    .Q_N(_0560_),
    .Q(\board_state[477] ));
 sg13g2_dfrbp_1 \board_state[478]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net866),
    .D(_1028_),
    .Q_N(_0561_),
    .Q(\board_state[478] ));
 sg13g2_dfrbp_1 \board_state[479]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net867),
    .D(_1029_),
    .Q_N(_0562_),
    .Q(\board_state[479] ));
 sg13g2_dfrbp_1 \board_state[47]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net868),
    .D(_1030_),
    .Q_N(_0130_),
    .Q(\board_state[47] ));
 sg13g2_dfrbp_1 \board_state[480]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net869),
    .D(_1031_),
    .Q_N(_0563_),
    .Q(\board_state[480] ));
 sg13g2_dfrbp_1 \board_state[481]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net870),
    .D(_1032_),
    .Q_N(_0564_),
    .Q(\board_state[481] ));
 sg13g2_dfrbp_1 \board_state[482]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net871),
    .D(_1033_),
    .Q_N(_0565_),
    .Q(\board_state[482] ));
 sg13g2_dfrbp_1 \board_state[483]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net872),
    .D(_1034_),
    .Q_N(_0566_),
    .Q(\board_state[483] ));
 sg13g2_dfrbp_1 \board_state[484]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net873),
    .D(_1035_),
    .Q_N(_0567_),
    .Q(\board_state[484] ));
 sg13g2_dfrbp_1 \board_state[485]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net874),
    .D(_1036_),
    .Q_N(_0568_),
    .Q(\board_state[485] ));
 sg13g2_dfrbp_1 \board_state[486]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net875),
    .D(_1037_),
    .Q_N(_0569_),
    .Q(\board_state[486] ));
 sg13g2_dfrbp_1 \board_state[487]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net876),
    .D(_1038_),
    .Q_N(_0570_),
    .Q(\board_state[487] ));
 sg13g2_dfrbp_1 \board_state[488]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net877),
    .D(_1039_),
    .Q_N(_0571_),
    .Q(\board_state[488] ));
 sg13g2_dfrbp_1 \board_state[489]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net878),
    .D(_1040_),
    .Q_N(_0572_),
    .Q(\board_state[489] ));
 sg13g2_dfrbp_1 \board_state[48]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net879),
    .D(_1041_),
    .Q_N(_0131_),
    .Q(\board_state[48] ));
 sg13g2_dfrbp_1 \board_state[490]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net880),
    .D(_1042_),
    .Q_N(_0573_),
    .Q(\board_state[490] ));
 sg13g2_dfrbp_1 \board_state[491]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net881),
    .D(_1043_),
    .Q_N(_0574_),
    .Q(\board_state[491] ));
 sg13g2_dfrbp_1 \board_state[492]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net882),
    .D(_1044_),
    .Q_N(_0575_),
    .Q(\board_state[492] ));
 sg13g2_dfrbp_1 \board_state[493]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net883),
    .D(_1045_),
    .Q_N(_0576_),
    .Q(\board_state[493] ));
 sg13g2_dfrbp_1 \board_state[494]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net884),
    .D(_1046_),
    .Q_N(_0577_),
    .Q(\board_state[494] ));
 sg13g2_dfrbp_1 \board_state[495]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net885),
    .D(_1047_),
    .Q_N(_0578_),
    .Q(\board_state[495] ));
 sg13g2_dfrbp_1 \board_state[496]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net886),
    .D(_1048_),
    .Q_N(_0579_),
    .Q(\board_state[496] ));
 sg13g2_dfrbp_1 \board_state[497]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net887),
    .D(_1049_),
    .Q_N(_0580_),
    .Q(\board_state[497] ));
 sg13g2_dfrbp_1 \board_state[498]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net888),
    .D(_1050_),
    .Q_N(_0581_),
    .Q(\board_state[498] ));
 sg13g2_dfrbp_1 \board_state[499]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net889),
    .D(_1051_),
    .Q_N(_0582_),
    .Q(\board_state[499] ));
 sg13g2_dfrbp_1 \board_state[49]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net890),
    .D(_1052_),
    .Q_N(_0132_),
    .Q(\board_state[49] ));
 sg13g2_dfrbp_1 \board_state[4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net891),
    .D(_1053_),
    .Q_N(_0087_),
    .Q(\board_state[4] ));
 sg13g2_dfrbp_1 \board_state[500]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net892),
    .D(_1054_),
    .Q_N(_0583_),
    .Q(\board_state[500] ));
 sg13g2_dfrbp_1 \board_state[501]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net893),
    .D(_1055_),
    .Q_N(_0584_),
    .Q(\board_state[501] ));
 sg13g2_dfrbp_1 \board_state[502]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net894),
    .D(_1056_),
    .Q_N(_0585_),
    .Q(\board_state[502] ));
 sg13g2_dfrbp_1 \board_state[503]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net895),
    .D(_1057_),
    .Q_N(_0586_),
    .Q(\board_state[503] ));
 sg13g2_dfrbp_1 \board_state[504]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net896),
    .D(_1058_),
    .Q_N(_0587_),
    .Q(\board_state[504] ));
 sg13g2_dfrbp_1 \board_state[505]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net897),
    .D(_1059_),
    .Q_N(_0588_),
    .Q(\board_state[505] ));
 sg13g2_dfrbp_1 \board_state[506]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net898),
    .D(_1060_),
    .Q_N(_0589_),
    .Q(\board_state[506] ));
 sg13g2_dfrbp_1 \board_state[507]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net899),
    .D(_1061_),
    .Q_N(_0590_),
    .Q(\board_state[507] ));
 sg13g2_dfrbp_1 \board_state[508]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net900),
    .D(_1062_),
    .Q_N(_0591_),
    .Q(\board_state[508] ));
 sg13g2_dfrbp_1 \board_state[509]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net901),
    .D(_1063_),
    .Q_N(_0592_),
    .Q(\board_state[509] ));
 sg13g2_dfrbp_1 \board_state[50]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net902),
    .D(_1064_),
    .Q_N(_0133_),
    .Q(\board_state[50] ));
 sg13g2_dfrbp_1 \board_state[510]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net903),
    .D(_1065_),
    .Q_N(_0593_),
    .Q(\board_state[510] ));
 sg13g2_dfrbp_1 \board_state[511]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net904),
    .D(_1066_),
    .Q_N(_0594_),
    .Q(\board_state[511] ));
 sg13g2_dfrbp_1 \board_state[51]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net905),
    .D(_1067_),
    .Q_N(_0134_),
    .Q(\board_state[51] ));
 sg13g2_dfrbp_1 \board_state[52]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net906),
    .D(_1068_),
    .Q_N(_0135_),
    .Q(\board_state[52] ));
 sg13g2_dfrbp_1 \board_state[53]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net907),
    .D(_1069_),
    .Q_N(_0136_),
    .Q(\board_state[53] ));
 sg13g2_dfrbp_1 \board_state[54]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net908),
    .D(_1070_),
    .Q_N(_0137_),
    .Q(\board_state[54] ));
 sg13g2_dfrbp_1 \board_state[55]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net909),
    .D(_1071_),
    .Q_N(_0138_),
    .Q(\board_state[55] ));
 sg13g2_dfrbp_1 \board_state[56]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net910),
    .D(_1072_),
    .Q_N(_0139_),
    .Q(\board_state[56] ));
 sg13g2_dfrbp_1 \board_state[57]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net911),
    .D(_1073_),
    .Q_N(_0140_),
    .Q(\board_state[57] ));
 sg13g2_dfrbp_1 \board_state[58]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net912),
    .D(_1074_),
    .Q_N(_0141_),
    .Q(\board_state[58] ));
 sg13g2_dfrbp_1 \board_state[59]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net913),
    .D(_1075_),
    .Q_N(_0142_),
    .Q(\board_state[59] ));
 sg13g2_dfrbp_1 \board_state[5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net914),
    .D(_1076_),
    .Q_N(_0088_),
    .Q(\board_state[5] ));
 sg13g2_dfrbp_1 \board_state[60]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net915),
    .D(_1077_),
    .Q_N(_0143_),
    .Q(\board_state[60] ));
 sg13g2_dfrbp_1 \board_state[61]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net916),
    .D(_1078_),
    .Q_N(_0144_),
    .Q(\board_state[61] ));
 sg13g2_dfrbp_1 \board_state[62]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net917),
    .D(_1079_),
    .Q_N(_0145_),
    .Q(\board_state[62] ));
 sg13g2_dfrbp_1 \board_state[63]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net918),
    .D(_1080_),
    .Q_N(_0146_),
    .Q(\board_state[63] ));
 sg13g2_dfrbp_1 \board_state[64]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net919),
    .D(_1081_),
    .Q_N(_0147_),
    .Q(\board_state[64] ));
 sg13g2_dfrbp_1 \board_state[65]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net920),
    .D(_1082_),
    .Q_N(_0148_),
    .Q(\board_state[65] ));
 sg13g2_dfrbp_1 \board_state[66]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net921),
    .D(_1083_),
    .Q_N(_0149_),
    .Q(\board_state[66] ));
 sg13g2_dfrbp_1 \board_state[67]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net922),
    .D(_1084_),
    .Q_N(_0150_),
    .Q(\board_state[67] ));
 sg13g2_dfrbp_1 \board_state[68]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net923),
    .D(_1085_),
    .Q_N(_0151_),
    .Q(\board_state[68] ));
 sg13g2_dfrbp_1 \board_state[69]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net924),
    .D(_1086_),
    .Q_N(_0152_),
    .Q(\board_state[69] ));
 sg13g2_dfrbp_1 \board_state[6]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net925),
    .D(_1087_),
    .Q_N(_0089_),
    .Q(\board_state[6] ));
 sg13g2_dfrbp_1 \board_state[70]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net926),
    .D(_1088_),
    .Q_N(_0153_),
    .Q(\board_state[70] ));
 sg13g2_dfrbp_1 \board_state[71]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net927),
    .D(_1089_),
    .Q_N(_0154_),
    .Q(\board_state[71] ));
 sg13g2_dfrbp_1 \board_state[72]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net928),
    .D(_1090_),
    .Q_N(_0155_),
    .Q(\board_state[72] ));
 sg13g2_dfrbp_1 \board_state[73]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net929),
    .D(_1091_),
    .Q_N(_0156_),
    .Q(\board_state[73] ));
 sg13g2_dfrbp_1 \board_state[74]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net930),
    .D(_1092_),
    .Q_N(_0157_),
    .Q(\board_state[74] ));
 sg13g2_dfrbp_1 \board_state[75]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net931),
    .D(_1093_),
    .Q_N(_0158_),
    .Q(\board_state[75] ));
 sg13g2_dfrbp_1 \board_state[76]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net932),
    .D(_1094_),
    .Q_N(_0159_),
    .Q(\board_state[76] ));
 sg13g2_dfrbp_1 \board_state[77]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net933),
    .D(_1095_),
    .Q_N(_0160_),
    .Q(\board_state[77] ));
 sg13g2_dfrbp_1 \board_state[78]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net934),
    .D(_1096_),
    .Q_N(_0161_),
    .Q(\board_state[78] ));
 sg13g2_dfrbp_1 \board_state[79]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net935),
    .D(_1097_),
    .Q_N(_0162_),
    .Q(\board_state[79] ));
 sg13g2_dfrbp_1 \board_state[7]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net936),
    .D(_1098_),
    .Q_N(_0090_),
    .Q(\board_state[7] ));
 sg13g2_dfrbp_1 \board_state[80]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net937),
    .D(_1099_),
    .Q_N(_0163_),
    .Q(\board_state[80] ));
 sg13g2_dfrbp_1 \board_state[81]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net938),
    .D(_1100_),
    .Q_N(_0164_),
    .Q(\board_state[81] ));
 sg13g2_dfrbp_1 \board_state[82]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net939),
    .D(_1101_),
    .Q_N(_0165_),
    .Q(\board_state[82] ));
 sg13g2_dfrbp_1 \board_state[83]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net940),
    .D(_1102_),
    .Q_N(_0166_),
    .Q(\board_state[83] ));
 sg13g2_dfrbp_1 \board_state[84]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net941),
    .D(_1103_),
    .Q_N(_0167_),
    .Q(\board_state[84] ));
 sg13g2_dfrbp_1 \board_state[85]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net942),
    .D(_1104_),
    .Q_N(_0168_),
    .Q(\board_state[85] ));
 sg13g2_dfrbp_1 \board_state[86]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net943),
    .D(_1105_),
    .Q_N(_0169_),
    .Q(\board_state[86] ));
 sg13g2_dfrbp_1 \board_state[87]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net944),
    .D(_1106_),
    .Q_N(_0170_),
    .Q(\board_state[87] ));
 sg13g2_dfrbp_1 \board_state[88]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net945),
    .D(_1107_),
    .Q_N(_0171_),
    .Q(\board_state[88] ));
 sg13g2_dfrbp_1 \board_state[89]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net946),
    .D(_1108_),
    .Q_N(_0172_),
    .Q(\board_state[89] ));
 sg13g2_dfrbp_1 \board_state[8]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net947),
    .D(_1109_),
    .Q_N(_0091_),
    .Q(\board_state[8] ));
 sg13g2_dfrbp_1 \board_state[90]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net948),
    .D(_1110_),
    .Q_N(_0173_),
    .Q(\board_state[90] ));
 sg13g2_dfrbp_1 \board_state[91]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net949),
    .D(_1111_),
    .Q_N(_0174_),
    .Q(\board_state[91] ));
 sg13g2_dfrbp_1 \board_state[92]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net950),
    .D(_1112_),
    .Q_N(_0175_),
    .Q(\board_state[92] ));
 sg13g2_dfrbp_1 \board_state[93]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net951),
    .D(_1113_),
    .Q_N(_0176_),
    .Q(\board_state[93] ));
 sg13g2_dfrbp_1 \board_state[94]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net952),
    .D(_1114_),
    .Q_N(_0177_),
    .Q(\board_state[94] ));
 sg13g2_dfrbp_1 \board_state[95]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net953),
    .D(_1115_),
    .Q_N(_0178_),
    .Q(\board_state[95] ));
 sg13g2_dfrbp_1 \board_state[96]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net954),
    .D(_1116_),
    .Q_N(_0179_),
    .Q(\board_state[96] ));
 sg13g2_dfrbp_1 \board_state[97]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net955),
    .D(_1117_),
    .Q_N(_0180_),
    .Q(\board_state[97] ));
 sg13g2_dfrbp_1 \board_state[98]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net956),
    .D(_1118_),
    .Q_N(_0181_),
    .Q(\board_state[98] ));
 sg13g2_dfrbp_1 \board_state[99]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net957),
    .D(_1119_),
    .Q_N(_0182_),
    .Q(\board_state[99] ));
 sg13g2_dfrbp_1 \board_state[9]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net958),
    .D(_1120_),
    .Q_N(_0092_),
    .Q(\board_state[9] ));
 sg13g2_dfrbp_1 \board_state_next[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net959),
    .D(_1121_),
    .Q_N(_5380_),
    .Q(\board_state_next[0] ));
 sg13g2_dfrbp_1 \board_state_next[100]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net960),
    .D(_1122_),
    .Q_N(_5379_),
    .Q(\board_state_next[100] ));
 sg13g2_dfrbp_1 \board_state_next[101]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net961),
    .D(_1123_),
    .Q_N(_5378_),
    .Q(\board_state_next[101] ));
 sg13g2_dfrbp_1 \board_state_next[102]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net962),
    .D(_1124_),
    .Q_N(_5377_),
    .Q(\board_state_next[102] ));
 sg13g2_dfrbp_1 \board_state_next[103]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net963),
    .D(_1125_),
    .Q_N(_5376_),
    .Q(\board_state_next[103] ));
 sg13g2_dfrbp_1 \board_state_next[104]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net964),
    .D(_1126_),
    .Q_N(_5375_),
    .Q(\board_state_next[104] ));
 sg13g2_dfrbp_1 \board_state_next[105]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net965),
    .D(_1127_),
    .Q_N(_5374_),
    .Q(\board_state_next[105] ));
 sg13g2_dfrbp_1 \board_state_next[106]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net966),
    .D(_1128_),
    .Q_N(_5373_),
    .Q(\board_state_next[106] ));
 sg13g2_dfrbp_1 \board_state_next[107]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net967),
    .D(_1129_),
    .Q_N(_5372_),
    .Q(\board_state_next[107] ));
 sg13g2_dfrbp_1 \board_state_next[108]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net968),
    .D(_1130_),
    .Q_N(_5371_),
    .Q(\board_state_next[108] ));
 sg13g2_dfrbp_1 \board_state_next[109]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net969),
    .D(_1131_),
    .Q_N(_5370_),
    .Q(\board_state_next[109] ));
 sg13g2_dfrbp_1 \board_state_next[10]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net970),
    .D(_1132_),
    .Q_N(_5369_),
    .Q(\board_state_next[10] ));
 sg13g2_dfrbp_1 \board_state_next[110]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net971),
    .D(_1133_),
    .Q_N(_5368_),
    .Q(\board_state_next[110] ));
 sg13g2_dfrbp_1 \board_state_next[111]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net972),
    .D(_1134_),
    .Q_N(_5367_),
    .Q(\board_state_next[111] ));
 sg13g2_dfrbp_1 \board_state_next[112]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net973),
    .D(_1135_),
    .Q_N(_5366_),
    .Q(\board_state_next[112] ));
 sg13g2_dfrbp_1 \board_state_next[113]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net974),
    .D(_1136_),
    .Q_N(_5365_),
    .Q(\board_state_next[113] ));
 sg13g2_dfrbp_1 \board_state_next[114]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net975),
    .D(_1137_),
    .Q_N(_5364_),
    .Q(\board_state_next[114] ));
 sg13g2_dfrbp_1 \board_state_next[115]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net976),
    .D(_1138_),
    .Q_N(_5363_),
    .Q(\board_state_next[115] ));
 sg13g2_dfrbp_1 \board_state_next[116]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net977),
    .D(_1139_),
    .Q_N(_5362_),
    .Q(\board_state_next[116] ));
 sg13g2_dfrbp_1 \board_state_next[117]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net978),
    .D(_1140_),
    .Q_N(_5361_),
    .Q(\board_state_next[117] ));
 sg13g2_dfrbp_1 \board_state_next[118]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net979),
    .D(_1141_),
    .Q_N(_5360_),
    .Q(\board_state_next[118] ));
 sg13g2_dfrbp_1 \board_state_next[119]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net980),
    .D(_1142_),
    .Q_N(_5359_),
    .Q(\board_state_next[119] ));
 sg13g2_dfrbp_1 \board_state_next[11]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net981),
    .D(_1143_),
    .Q_N(_5358_),
    .Q(\board_state_next[11] ));
 sg13g2_dfrbp_1 \board_state_next[120]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net982),
    .D(_1144_),
    .Q_N(_5357_),
    .Q(\board_state_next[120] ));
 sg13g2_dfrbp_1 \board_state_next[121]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net983),
    .D(_1145_),
    .Q_N(_5356_),
    .Q(\board_state_next[121] ));
 sg13g2_dfrbp_1 \board_state_next[122]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net984),
    .D(_1146_),
    .Q_N(_5355_),
    .Q(\board_state_next[122] ));
 sg13g2_dfrbp_1 \board_state_next[123]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net985),
    .D(_1147_),
    .Q_N(_5354_),
    .Q(\board_state_next[123] ));
 sg13g2_dfrbp_1 \board_state_next[124]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net986),
    .D(_1148_),
    .Q_N(_5353_),
    .Q(\board_state_next[124] ));
 sg13g2_dfrbp_1 \board_state_next[125]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net987),
    .D(_1149_),
    .Q_N(_5352_),
    .Q(\board_state_next[125] ));
 sg13g2_dfrbp_1 \board_state_next[126]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net988),
    .D(_1150_),
    .Q_N(_5351_),
    .Q(\board_state_next[126] ));
 sg13g2_dfrbp_1 \board_state_next[127]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net989),
    .D(_1151_),
    .Q_N(_5350_),
    .Q(\board_state_next[127] ));
 sg13g2_dfrbp_1 \board_state_next[128]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net990),
    .D(_1152_),
    .Q_N(_5349_),
    .Q(\board_state_next[128] ));
 sg13g2_dfrbp_1 \board_state_next[129]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net991),
    .D(_1153_),
    .Q_N(_5348_),
    .Q(\board_state_next[129] ));
 sg13g2_dfrbp_1 \board_state_next[12]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net992),
    .D(_1154_),
    .Q_N(_5347_),
    .Q(\board_state_next[12] ));
 sg13g2_dfrbp_1 \board_state_next[130]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net993),
    .D(_1155_),
    .Q_N(_5346_),
    .Q(\board_state_next[130] ));
 sg13g2_dfrbp_1 \board_state_next[131]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net994),
    .D(_1156_),
    .Q_N(_5345_),
    .Q(\board_state_next[131] ));
 sg13g2_dfrbp_1 \board_state_next[132]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net995),
    .D(_1157_),
    .Q_N(_5344_),
    .Q(\board_state_next[132] ));
 sg13g2_dfrbp_1 \board_state_next[133]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net996),
    .D(_1158_),
    .Q_N(_5343_),
    .Q(\board_state_next[133] ));
 sg13g2_dfrbp_1 \board_state_next[134]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net997),
    .D(_1159_),
    .Q_N(_5342_),
    .Q(\board_state_next[134] ));
 sg13g2_dfrbp_1 \board_state_next[135]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net998),
    .D(_1160_),
    .Q_N(_5341_),
    .Q(\board_state_next[135] ));
 sg13g2_dfrbp_1 \board_state_next[136]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net999),
    .D(_1161_),
    .Q_N(_5340_),
    .Q(\board_state_next[136] ));
 sg13g2_dfrbp_1 \board_state_next[137]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1000),
    .D(_1162_),
    .Q_N(_5339_),
    .Q(\board_state_next[137] ));
 sg13g2_dfrbp_1 \board_state_next[138]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1001),
    .D(_1163_),
    .Q_N(_5338_),
    .Q(\board_state_next[138] ));
 sg13g2_dfrbp_1 \board_state_next[139]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1002),
    .D(_1164_),
    .Q_N(_5337_),
    .Q(\board_state_next[139] ));
 sg13g2_dfrbp_1 \board_state_next[13]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1003),
    .D(_1165_),
    .Q_N(_5336_),
    .Q(\board_state_next[13] ));
 sg13g2_dfrbp_1 \board_state_next[140]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1004),
    .D(_1166_),
    .Q_N(_5335_),
    .Q(\board_state_next[140] ));
 sg13g2_dfrbp_1 \board_state_next[141]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1005),
    .D(_1167_),
    .Q_N(_5334_),
    .Q(\board_state_next[141] ));
 sg13g2_dfrbp_1 \board_state_next[142]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1006),
    .D(_1168_),
    .Q_N(_5333_),
    .Q(\board_state_next[142] ));
 sg13g2_dfrbp_1 \board_state_next[143]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1007),
    .D(_1169_),
    .Q_N(_5332_),
    .Q(\board_state_next[143] ));
 sg13g2_dfrbp_1 \board_state_next[144]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1008),
    .D(_1170_),
    .Q_N(_5331_),
    .Q(\board_state_next[144] ));
 sg13g2_dfrbp_1 \board_state_next[145]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1009),
    .D(_1171_),
    .Q_N(_5330_),
    .Q(\board_state_next[145] ));
 sg13g2_dfrbp_1 \board_state_next[146]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1010),
    .D(_1172_),
    .Q_N(_5329_),
    .Q(\board_state_next[146] ));
 sg13g2_dfrbp_1 \board_state_next[147]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1011),
    .D(_1173_),
    .Q_N(_5328_),
    .Q(\board_state_next[147] ));
 sg13g2_dfrbp_1 \board_state_next[148]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1012),
    .D(_1174_),
    .Q_N(_5327_),
    .Q(\board_state_next[148] ));
 sg13g2_dfrbp_1 \board_state_next[149]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1013),
    .D(_1175_),
    .Q_N(_5326_),
    .Q(\board_state_next[149] ));
 sg13g2_dfrbp_1 \board_state_next[14]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1014),
    .D(_1176_),
    .Q_N(_5325_),
    .Q(\board_state_next[14] ));
 sg13g2_dfrbp_1 \board_state_next[150]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1015),
    .D(_1177_),
    .Q_N(_5324_),
    .Q(\board_state_next[150] ));
 sg13g2_dfrbp_1 \board_state_next[151]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1016),
    .D(_1178_),
    .Q_N(_5323_),
    .Q(\board_state_next[151] ));
 sg13g2_dfrbp_1 \board_state_next[152]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1017),
    .D(_1179_),
    .Q_N(_5322_),
    .Q(\board_state_next[152] ));
 sg13g2_dfrbp_1 \board_state_next[153]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1018),
    .D(_1180_),
    .Q_N(_5321_),
    .Q(\board_state_next[153] ));
 sg13g2_dfrbp_1 \board_state_next[154]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1019),
    .D(_1181_),
    .Q_N(_5320_),
    .Q(\board_state_next[154] ));
 sg13g2_dfrbp_1 \board_state_next[155]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1020),
    .D(_1182_),
    .Q_N(_5319_),
    .Q(\board_state_next[155] ));
 sg13g2_dfrbp_1 \board_state_next[156]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1021),
    .D(_1183_),
    .Q_N(_5318_),
    .Q(\board_state_next[156] ));
 sg13g2_dfrbp_1 \board_state_next[157]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1022),
    .D(_1184_),
    .Q_N(_5317_),
    .Q(\board_state_next[157] ));
 sg13g2_dfrbp_1 \board_state_next[158]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1023),
    .D(_1185_),
    .Q_N(_5316_),
    .Q(\board_state_next[158] ));
 sg13g2_dfrbp_1 \board_state_next[159]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1024),
    .D(_1186_),
    .Q_N(_5315_),
    .Q(\board_state_next[159] ));
 sg13g2_dfrbp_1 \board_state_next[15]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1025),
    .D(_1187_),
    .Q_N(_5314_),
    .Q(\board_state_next[15] ));
 sg13g2_dfrbp_1 \board_state_next[160]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1026),
    .D(_1188_),
    .Q_N(_5313_),
    .Q(\board_state_next[160] ));
 sg13g2_dfrbp_1 \board_state_next[161]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1027),
    .D(_1189_),
    .Q_N(_5312_),
    .Q(\board_state_next[161] ));
 sg13g2_dfrbp_1 \board_state_next[162]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1028),
    .D(_1190_),
    .Q_N(_5311_),
    .Q(\board_state_next[162] ));
 sg13g2_dfrbp_1 \board_state_next[163]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1029),
    .D(_1191_),
    .Q_N(_5310_),
    .Q(\board_state_next[163] ));
 sg13g2_dfrbp_1 \board_state_next[164]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1030),
    .D(_1192_),
    .Q_N(_5309_),
    .Q(\board_state_next[164] ));
 sg13g2_dfrbp_1 \board_state_next[165]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1031),
    .D(_1193_),
    .Q_N(_5308_),
    .Q(\board_state_next[165] ));
 sg13g2_dfrbp_1 \board_state_next[166]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1032),
    .D(_1194_),
    .Q_N(_5307_),
    .Q(\board_state_next[166] ));
 sg13g2_dfrbp_1 \board_state_next[167]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1033),
    .D(_1195_),
    .Q_N(_5306_),
    .Q(\board_state_next[167] ));
 sg13g2_dfrbp_1 \board_state_next[168]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1034),
    .D(_1196_),
    .Q_N(_5305_),
    .Q(\board_state_next[168] ));
 sg13g2_dfrbp_1 \board_state_next[169]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1035),
    .D(_1197_),
    .Q_N(_5304_),
    .Q(\board_state_next[169] ));
 sg13g2_dfrbp_1 \board_state_next[16]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1036),
    .D(_1198_),
    .Q_N(_5303_),
    .Q(\board_state_next[16] ));
 sg13g2_dfrbp_1 \board_state_next[170]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1037),
    .D(_1199_),
    .Q_N(_5302_),
    .Q(\board_state_next[170] ));
 sg13g2_dfrbp_1 \board_state_next[171]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1038),
    .D(_1200_),
    .Q_N(_5301_),
    .Q(\board_state_next[171] ));
 sg13g2_dfrbp_1 \board_state_next[172]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1039),
    .D(_1201_),
    .Q_N(_5300_),
    .Q(\board_state_next[172] ));
 sg13g2_dfrbp_1 \board_state_next[173]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1040),
    .D(_1202_),
    .Q_N(_5299_),
    .Q(\board_state_next[173] ));
 sg13g2_dfrbp_1 \board_state_next[174]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1041),
    .D(_1203_),
    .Q_N(_5298_),
    .Q(\board_state_next[174] ));
 sg13g2_dfrbp_1 \board_state_next[175]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1042),
    .D(_1204_),
    .Q_N(_5297_),
    .Q(\board_state_next[175] ));
 sg13g2_dfrbp_1 \board_state_next[176]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1043),
    .D(_1205_),
    .Q_N(_5296_),
    .Q(\board_state_next[176] ));
 sg13g2_dfrbp_1 \board_state_next[177]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1044),
    .D(_1206_),
    .Q_N(_5295_),
    .Q(\board_state_next[177] ));
 sg13g2_dfrbp_1 \board_state_next[178]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1045),
    .D(_1207_),
    .Q_N(_5294_),
    .Q(\board_state_next[178] ));
 sg13g2_dfrbp_1 \board_state_next[179]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1046),
    .D(_1208_),
    .Q_N(_5293_),
    .Q(\board_state_next[179] ));
 sg13g2_dfrbp_1 \board_state_next[17]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1047),
    .D(_1209_),
    .Q_N(_5292_),
    .Q(\board_state_next[17] ));
 sg13g2_dfrbp_1 \board_state_next[180]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1048),
    .D(_1210_),
    .Q_N(_5291_),
    .Q(\board_state_next[180] ));
 sg13g2_dfrbp_1 \board_state_next[181]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1049),
    .D(_1211_),
    .Q_N(_5290_),
    .Q(\board_state_next[181] ));
 sg13g2_dfrbp_1 \board_state_next[182]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1050),
    .D(_1212_),
    .Q_N(_5289_),
    .Q(\board_state_next[182] ));
 sg13g2_dfrbp_1 \board_state_next[183]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1051),
    .D(_1213_),
    .Q_N(_5288_),
    .Q(\board_state_next[183] ));
 sg13g2_dfrbp_1 \board_state_next[184]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1052),
    .D(_1214_),
    .Q_N(_5287_),
    .Q(\board_state_next[184] ));
 sg13g2_dfrbp_1 \board_state_next[185]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1053),
    .D(_1215_),
    .Q_N(_5286_),
    .Q(\board_state_next[185] ));
 sg13g2_dfrbp_1 \board_state_next[186]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1054),
    .D(_1216_),
    .Q_N(_5285_),
    .Q(\board_state_next[186] ));
 sg13g2_dfrbp_1 \board_state_next[187]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1055),
    .D(_1217_),
    .Q_N(_5284_),
    .Q(\board_state_next[187] ));
 sg13g2_dfrbp_1 \board_state_next[188]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1056),
    .D(_1218_),
    .Q_N(_5283_),
    .Q(\board_state_next[188] ));
 sg13g2_dfrbp_1 \board_state_next[189]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1057),
    .D(_1219_),
    .Q_N(_5282_),
    .Q(\board_state_next[189] ));
 sg13g2_dfrbp_1 \board_state_next[18]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1058),
    .D(_1220_),
    .Q_N(_5281_),
    .Q(\board_state_next[18] ));
 sg13g2_dfrbp_1 \board_state_next[190]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1059),
    .D(_1221_),
    .Q_N(_5280_),
    .Q(\board_state_next[190] ));
 sg13g2_dfrbp_1 \board_state_next[191]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1060),
    .D(_1222_),
    .Q_N(_5279_),
    .Q(\board_state_next[191] ));
 sg13g2_dfrbp_1 \board_state_next[192]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1061),
    .D(_1223_),
    .Q_N(_5278_),
    .Q(\board_state_next[192] ));
 sg13g2_dfrbp_1 \board_state_next[193]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1062),
    .D(_1224_),
    .Q_N(_5277_),
    .Q(\board_state_next[193] ));
 sg13g2_dfrbp_1 \board_state_next[194]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1063),
    .D(_1225_),
    .Q_N(_5276_),
    .Q(\board_state_next[194] ));
 sg13g2_dfrbp_1 \board_state_next[195]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1064),
    .D(_1226_),
    .Q_N(_5275_),
    .Q(\board_state_next[195] ));
 sg13g2_dfrbp_1 \board_state_next[196]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1065),
    .D(_1227_),
    .Q_N(_5274_),
    .Q(\board_state_next[196] ));
 sg13g2_dfrbp_1 \board_state_next[197]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1066),
    .D(_1228_),
    .Q_N(_5273_),
    .Q(\board_state_next[197] ));
 sg13g2_dfrbp_1 \board_state_next[198]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1067),
    .D(_1229_),
    .Q_N(_5272_),
    .Q(\board_state_next[198] ));
 sg13g2_dfrbp_1 \board_state_next[199]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1068),
    .D(_1230_),
    .Q_N(_5271_),
    .Q(\board_state_next[199] ));
 sg13g2_dfrbp_1 \board_state_next[19]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1069),
    .D(_1231_),
    .Q_N(_5270_),
    .Q(\board_state_next[19] ));
 sg13g2_dfrbp_1 \board_state_next[1]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1070),
    .D(_1232_),
    .Q_N(_5269_),
    .Q(\board_state_next[1] ));
 sg13g2_dfrbp_1 \board_state_next[200]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1071),
    .D(_1233_),
    .Q_N(_5268_),
    .Q(\board_state_next[200] ));
 sg13g2_dfrbp_1 \board_state_next[201]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1072),
    .D(_1234_),
    .Q_N(_5267_),
    .Q(\board_state_next[201] ));
 sg13g2_dfrbp_1 \board_state_next[202]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1073),
    .D(_1235_),
    .Q_N(_5266_),
    .Q(\board_state_next[202] ));
 sg13g2_dfrbp_1 \board_state_next[203]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1074),
    .D(_1236_),
    .Q_N(_5265_),
    .Q(\board_state_next[203] ));
 sg13g2_dfrbp_1 \board_state_next[204]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1075),
    .D(_1237_),
    .Q_N(_5264_),
    .Q(\board_state_next[204] ));
 sg13g2_dfrbp_1 \board_state_next[205]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1076),
    .D(_1238_),
    .Q_N(_5263_),
    .Q(\board_state_next[205] ));
 sg13g2_dfrbp_1 \board_state_next[206]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1077),
    .D(_1239_),
    .Q_N(_5262_),
    .Q(\board_state_next[206] ));
 sg13g2_dfrbp_1 \board_state_next[207]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1078),
    .D(_1240_),
    .Q_N(_5261_),
    .Q(\board_state_next[207] ));
 sg13g2_dfrbp_1 \board_state_next[208]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1079),
    .D(_1241_),
    .Q_N(_5260_),
    .Q(\board_state_next[208] ));
 sg13g2_dfrbp_1 \board_state_next[209]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1080),
    .D(_1242_),
    .Q_N(_5259_),
    .Q(\board_state_next[209] ));
 sg13g2_dfrbp_1 \board_state_next[20]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1081),
    .D(_1243_),
    .Q_N(_5258_),
    .Q(\board_state_next[20] ));
 sg13g2_dfrbp_1 \board_state_next[210]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1082),
    .D(_1244_),
    .Q_N(_5257_),
    .Q(\board_state_next[210] ));
 sg13g2_dfrbp_1 \board_state_next[211]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1083),
    .D(_1245_),
    .Q_N(_5256_),
    .Q(\board_state_next[211] ));
 sg13g2_dfrbp_1 \board_state_next[212]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1084),
    .D(_1246_),
    .Q_N(_5255_),
    .Q(\board_state_next[212] ));
 sg13g2_dfrbp_1 \board_state_next[213]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1085),
    .D(_1247_),
    .Q_N(_5254_),
    .Q(\board_state_next[213] ));
 sg13g2_dfrbp_1 \board_state_next[214]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1086),
    .D(_1248_),
    .Q_N(_5253_),
    .Q(\board_state_next[214] ));
 sg13g2_dfrbp_1 \board_state_next[215]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1087),
    .D(_1249_),
    .Q_N(_5252_),
    .Q(\board_state_next[215] ));
 sg13g2_dfrbp_1 \board_state_next[216]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1088),
    .D(_1250_),
    .Q_N(_5251_),
    .Q(\board_state_next[216] ));
 sg13g2_dfrbp_1 \board_state_next[217]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1089),
    .D(_1251_),
    .Q_N(_5250_),
    .Q(\board_state_next[217] ));
 sg13g2_dfrbp_1 \board_state_next[218]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1090),
    .D(_1252_),
    .Q_N(_5249_),
    .Q(\board_state_next[218] ));
 sg13g2_dfrbp_1 \board_state_next[219]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1091),
    .D(_1253_),
    .Q_N(_5248_),
    .Q(\board_state_next[219] ));
 sg13g2_dfrbp_1 \board_state_next[21]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1092),
    .D(_1254_),
    .Q_N(_5247_),
    .Q(\board_state_next[21] ));
 sg13g2_dfrbp_1 \board_state_next[220]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1093),
    .D(_1255_),
    .Q_N(_5246_),
    .Q(\board_state_next[220] ));
 sg13g2_dfrbp_1 \board_state_next[221]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1094),
    .D(_1256_),
    .Q_N(_5245_),
    .Q(\board_state_next[221] ));
 sg13g2_dfrbp_1 \board_state_next[222]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1095),
    .D(_1257_),
    .Q_N(_5244_),
    .Q(\board_state_next[222] ));
 sg13g2_dfrbp_1 \board_state_next[223]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1096),
    .D(_1258_),
    .Q_N(_5243_),
    .Q(\board_state_next[223] ));
 sg13g2_dfrbp_1 \board_state_next[224]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1097),
    .D(_1259_),
    .Q_N(_5242_),
    .Q(\board_state_next[224] ));
 sg13g2_dfrbp_1 \board_state_next[225]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1098),
    .D(_1260_),
    .Q_N(_5241_),
    .Q(\board_state_next[225] ));
 sg13g2_dfrbp_1 \board_state_next[226]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1099),
    .D(_1261_),
    .Q_N(_5240_),
    .Q(\board_state_next[226] ));
 sg13g2_dfrbp_1 \board_state_next[227]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1100),
    .D(_1262_),
    .Q_N(_5239_),
    .Q(\board_state_next[227] ));
 sg13g2_dfrbp_1 \board_state_next[228]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1101),
    .D(_1263_),
    .Q_N(_5238_),
    .Q(\board_state_next[228] ));
 sg13g2_dfrbp_1 \board_state_next[229]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1102),
    .D(_1264_),
    .Q_N(_5237_),
    .Q(\board_state_next[229] ));
 sg13g2_dfrbp_1 \board_state_next[22]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1103),
    .D(_1265_),
    .Q_N(_5236_),
    .Q(\board_state_next[22] ));
 sg13g2_dfrbp_1 \board_state_next[230]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1104),
    .D(_1266_),
    .Q_N(_5235_),
    .Q(\board_state_next[230] ));
 sg13g2_dfrbp_1 \board_state_next[231]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1105),
    .D(_1267_),
    .Q_N(_5234_),
    .Q(\board_state_next[231] ));
 sg13g2_dfrbp_1 \board_state_next[232]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1106),
    .D(_1268_),
    .Q_N(_5233_),
    .Q(\board_state_next[232] ));
 sg13g2_dfrbp_1 \board_state_next[233]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1107),
    .D(_1269_),
    .Q_N(_5232_),
    .Q(\board_state_next[233] ));
 sg13g2_dfrbp_1 \board_state_next[234]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1108),
    .D(_1270_),
    .Q_N(_5231_),
    .Q(\board_state_next[234] ));
 sg13g2_dfrbp_1 \board_state_next[235]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1109),
    .D(_1271_),
    .Q_N(_5230_),
    .Q(\board_state_next[235] ));
 sg13g2_dfrbp_1 \board_state_next[236]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1110),
    .D(_1272_),
    .Q_N(_5229_),
    .Q(\board_state_next[236] ));
 sg13g2_dfrbp_1 \board_state_next[237]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1111),
    .D(_1273_),
    .Q_N(_5228_),
    .Q(\board_state_next[237] ));
 sg13g2_dfrbp_1 \board_state_next[238]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1112),
    .D(_1274_),
    .Q_N(_5227_),
    .Q(\board_state_next[238] ));
 sg13g2_dfrbp_1 \board_state_next[239]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1113),
    .D(_1275_),
    .Q_N(_5226_),
    .Q(\board_state_next[239] ));
 sg13g2_dfrbp_1 \board_state_next[23]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1114),
    .D(_1276_),
    .Q_N(_5225_),
    .Q(\board_state_next[23] ));
 sg13g2_dfrbp_1 \board_state_next[240]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1115),
    .D(_1277_),
    .Q_N(_5224_),
    .Q(\board_state_next[240] ));
 sg13g2_dfrbp_1 \board_state_next[241]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1116),
    .D(_1278_),
    .Q_N(_5223_),
    .Q(\board_state_next[241] ));
 sg13g2_dfrbp_1 \board_state_next[242]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1117),
    .D(_1279_),
    .Q_N(_5222_),
    .Q(\board_state_next[242] ));
 sg13g2_dfrbp_1 \board_state_next[243]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1118),
    .D(_1280_),
    .Q_N(_5221_),
    .Q(\board_state_next[243] ));
 sg13g2_dfrbp_1 \board_state_next[244]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1119),
    .D(_1281_),
    .Q_N(_5220_),
    .Q(\board_state_next[244] ));
 sg13g2_dfrbp_1 \board_state_next[245]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1120),
    .D(_1282_),
    .Q_N(_5219_),
    .Q(\board_state_next[245] ));
 sg13g2_dfrbp_1 \board_state_next[246]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1121),
    .D(_1283_),
    .Q_N(_5218_),
    .Q(\board_state_next[246] ));
 sg13g2_dfrbp_1 \board_state_next[247]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1122),
    .D(_1284_),
    .Q_N(_5217_),
    .Q(\board_state_next[247] ));
 sg13g2_dfrbp_1 \board_state_next[248]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1123),
    .D(_1285_),
    .Q_N(_5216_),
    .Q(\board_state_next[248] ));
 sg13g2_dfrbp_1 \board_state_next[249]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1124),
    .D(_1286_),
    .Q_N(_5215_),
    .Q(\board_state_next[249] ));
 sg13g2_dfrbp_1 \board_state_next[24]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1125),
    .D(_1287_),
    .Q_N(_5214_),
    .Q(\board_state_next[24] ));
 sg13g2_dfrbp_1 \board_state_next[250]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1126),
    .D(_1288_),
    .Q_N(_5213_),
    .Q(\board_state_next[250] ));
 sg13g2_dfrbp_1 \board_state_next[251]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1127),
    .D(_1289_),
    .Q_N(_5212_),
    .Q(\board_state_next[251] ));
 sg13g2_dfrbp_1 \board_state_next[252]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1128),
    .D(_1290_),
    .Q_N(_5211_),
    .Q(\board_state_next[252] ));
 sg13g2_dfrbp_1 \board_state_next[253]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1129),
    .D(_1291_),
    .Q_N(_5210_),
    .Q(\board_state_next[253] ));
 sg13g2_dfrbp_1 \board_state_next[254]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1130),
    .D(_1292_),
    .Q_N(_5209_),
    .Q(\board_state_next[254] ));
 sg13g2_dfrbp_1 \board_state_next[255]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1131),
    .D(_1293_),
    .Q_N(_5208_),
    .Q(\board_state_next[255] ));
 sg13g2_dfrbp_1 \board_state_next[256]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1132),
    .D(_1294_),
    .Q_N(_5207_),
    .Q(\board_state_next[256] ));
 sg13g2_dfrbp_1 \board_state_next[257]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1133),
    .D(_1295_),
    .Q_N(_5206_),
    .Q(\board_state_next[257] ));
 sg13g2_dfrbp_1 \board_state_next[258]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1134),
    .D(_1296_),
    .Q_N(_5205_),
    .Q(\board_state_next[258] ));
 sg13g2_dfrbp_1 \board_state_next[259]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1135),
    .D(_1297_),
    .Q_N(_5204_),
    .Q(\board_state_next[259] ));
 sg13g2_dfrbp_1 \board_state_next[25]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1136),
    .D(_1298_),
    .Q_N(_5203_),
    .Q(\board_state_next[25] ));
 sg13g2_dfrbp_1 \board_state_next[260]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1137),
    .D(_1299_),
    .Q_N(_5202_),
    .Q(\board_state_next[260] ));
 sg13g2_dfrbp_1 \board_state_next[261]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1138),
    .D(_1300_),
    .Q_N(_5201_),
    .Q(\board_state_next[261] ));
 sg13g2_dfrbp_1 \board_state_next[262]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1139),
    .D(_1301_),
    .Q_N(_5200_),
    .Q(\board_state_next[262] ));
 sg13g2_dfrbp_1 \board_state_next[263]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1140),
    .D(_1302_),
    .Q_N(_5199_),
    .Q(\board_state_next[263] ));
 sg13g2_dfrbp_1 \board_state_next[264]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1141),
    .D(_1303_),
    .Q_N(_5198_),
    .Q(\board_state_next[264] ));
 sg13g2_dfrbp_1 \board_state_next[265]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1142),
    .D(_1304_),
    .Q_N(_5197_),
    .Q(\board_state_next[265] ));
 sg13g2_dfrbp_1 \board_state_next[266]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1143),
    .D(_1305_),
    .Q_N(_5196_),
    .Q(\board_state_next[266] ));
 sg13g2_dfrbp_1 \board_state_next[267]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1144),
    .D(_1306_),
    .Q_N(_5195_),
    .Q(\board_state_next[267] ));
 sg13g2_dfrbp_1 \board_state_next[268]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1145),
    .D(_1307_),
    .Q_N(_5194_),
    .Q(\board_state_next[268] ));
 sg13g2_dfrbp_1 \board_state_next[269]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1146),
    .D(_1308_),
    .Q_N(_5193_),
    .Q(\board_state_next[269] ));
 sg13g2_dfrbp_1 \board_state_next[26]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1147),
    .D(_1309_),
    .Q_N(_5192_),
    .Q(\board_state_next[26] ));
 sg13g2_dfrbp_1 \board_state_next[270]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1148),
    .D(_1310_),
    .Q_N(_5191_),
    .Q(\board_state_next[270] ));
 sg13g2_dfrbp_1 \board_state_next[271]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1149),
    .D(_1311_),
    .Q_N(_5190_),
    .Q(\board_state_next[271] ));
 sg13g2_dfrbp_1 \board_state_next[272]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1150),
    .D(_1312_),
    .Q_N(_5189_),
    .Q(\board_state_next[272] ));
 sg13g2_dfrbp_1 \board_state_next[273]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1151),
    .D(_1313_),
    .Q_N(_5188_),
    .Q(\board_state_next[273] ));
 sg13g2_dfrbp_1 \board_state_next[274]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1152),
    .D(_1314_),
    .Q_N(_5187_),
    .Q(\board_state_next[274] ));
 sg13g2_dfrbp_1 \board_state_next[275]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1153),
    .D(_1315_),
    .Q_N(_5186_),
    .Q(\board_state_next[275] ));
 sg13g2_dfrbp_1 \board_state_next[276]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1154),
    .D(_1316_),
    .Q_N(_5185_),
    .Q(\board_state_next[276] ));
 sg13g2_dfrbp_1 \board_state_next[277]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1155),
    .D(_1317_),
    .Q_N(_5184_),
    .Q(\board_state_next[277] ));
 sg13g2_dfrbp_1 \board_state_next[278]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1156),
    .D(_1318_),
    .Q_N(_5183_),
    .Q(\board_state_next[278] ));
 sg13g2_dfrbp_1 \board_state_next[279]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1157),
    .D(_1319_),
    .Q_N(_5182_),
    .Q(\board_state_next[279] ));
 sg13g2_dfrbp_1 \board_state_next[27]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1158),
    .D(_1320_),
    .Q_N(_5181_),
    .Q(\board_state_next[27] ));
 sg13g2_dfrbp_1 \board_state_next[280]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1159),
    .D(_1321_),
    .Q_N(_5180_),
    .Q(\board_state_next[280] ));
 sg13g2_dfrbp_1 \board_state_next[281]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1160),
    .D(_1322_),
    .Q_N(_5179_),
    .Q(\board_state_next[281] ));
 sg13g2_dfrbp_1 \board_state_next[282]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1161),
    .D(_1323_),
    .Q_N(_5178_),
    .Q(\board_state_next[282] ));
 sg13g2_dfrbp_1 \board_state_next[283]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1162),
    .D(_1324_),
    .Q_N(_5177_),
    .Q(\board_state_next[283] ));
 sg13g2_dfrbp_1 \board_state_next[284]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1163),
    .D(_1325_),
    .Q_N(_5176_),
    .Q(\board_state_next[284] ));
 sg13g2_dfrbp_1 \board_state_next[285]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1164),
    .D(_1326_),
    .Q_N(_5175_),
    .Q(\board_state_next[285] ));
 sg13g2_dfrbp_1 \board_state_next[286]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1165),
    .D(_1327_),
    .Q_N(_5174_),
    .Q(\board_state_next[286] ));
 sg13g2_dfrbp_1 \board_state_next[287]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1166),
    .D(_1328_),
    .Q_N(_5173_),
    .Q(\board_state_next[287] ));
 sg13g2_dfrbp_1 \board_state_next[288]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1167),
    .D(_1329_),
    .Q_N(_5172_),
    .Q(\board_state_next[288] ));
 sg13g2_dfrbp_1 \board_state_next[289]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1168),
    .D(_1330_),
    .Q_N(_5171_),
    .Q(\board_state_next[289] ));
 sg13g2_dfrbp_1 \board_state_next[28]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1169),
    .D(_1331_),
    .Q_N(_5170_),
    .Q(\board_state_next[28] ));
 sg13g2_dfrbp_1 \board_state_next[290]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1170),
    .D(_1332_),
    .Q_N(_5169_),
    .Q(\board_state_next[290] ));
 sg13g2_dfrbp_1 \board_state_next[291]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1171),
    .D(_1333_),
    .Q_N(_5168_),
    .Q(\board_state_next[291] ));
 sg13g2_dfrbp_1 \board_state_next[292]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1172),
    .D(_1334_),
    .Q_N(_5167_),
    .Q(\board_state_next[292] ));
 sg13g2_dfrbp_1 \board_state_next[293]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1173),
    .D(_1335_),
    .Q_N(_5166_),
    .Q(\board_state_next[293] ));
 sg13g2_dfrbp_1 \board_state_next[294]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1174),
    .D(_1336_),
    .Q_N(_5165_),
    .Q(\board_state_next[294] ));
 sg13g2_dfrbp_1 \board_state_next[295]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1175),
    .D(_1337_),
    .Q_N(_5164_),
    .Q(\board_state_next[295] ));
 sg13g2_dfrbp_1 \board_state_next[296]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1176),
    .D(_1338_),
    .Q_N(_5163_),
    .Q(\board_state_next[296] ));
 sg13g2_dfrbp_1 \board_state_next[297]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1177),
    .D(_1339_),
    .Q_N(_5162_),
    .Q(\board_state_next[297] ));
 sg13g2_dfrbp_1 \board_state_next[298]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1178),
    .D(_1340_),
    .Q_N(_5161_),
    .Q(\board_state_next[298] ));
 sg13g2_dfrbp_1 \board_state_next[299]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1179),
    .D(_1341_),
    .Q_N(_5160_),
    .Q(\board_state_next[299] ));
 sg13g2_dfrbp_1 \board_state_next[29]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1180),
    .D(_1342_),
    .Q_N(_5159_),
    .Q(\board_state_next[29] ));
 sg13g2_dfrbp_1 \board_state_next[2]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1181),
    .D(_1343_),
    .Q_N(_5158_),
    .Q(\board_state_next[2] ));
 sg13g2_dfrbp_1 \board_state_next[300]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1182),
    .D(_1344_),
    .Q_N(_5157_),
    .Q(\board_state_next[300] ));
 sg13g2_dfrbp_1 \board_state_next[301]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1183),
    .D(_1345_),
    .Q_N(_5156_),
    .Q(\board_state_next[301] ));
 sg13g2_dfrbp_1 \board_state_next[302]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1184),
    .D(_1346_),
    .Q_N(_5155_),
    .Q(\board_state_next[302] ));
 sg13g2_dfrbp_1 \board_state_next[303]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1185),
    .D(_1347_),
    .Q_N(_5154_),
    .Q(\board_state_next[303] ));
 sg13g2_dfrbp_1 \board_state_next[304]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1186),
    .D(_1348_),
    .Q_N(_5153_),
    .Q(\board_state_next[304] ));
 sg13g2_dfrbp_1 \board_state_next[305]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1187),
    .D(_1349_),
    .Q_N(_5152_),
    .Q(\board_state_next[305] ));
 sg13g2_dfrbp_1 \board_state_next[306]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1188),
    .D(_1350_),
    .Q_N(_5151_),
    .Q(\board_state_next[306] ));
 sg13g2_dfrbp_1 \board_state_next[307]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1189),
    .D(_1351_),
    .Q_N(_5150_),
    .Q(\board_state_next[307] ));
 sg13g2_dfrbp_1 \board_state_next[308]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1190),
    .D(_1352_),
    .Q_N(_5149_),
    .Q(\board_state_next[308] ));
 sg13g2_dfrbp_1 \board_state_next[309]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1191),
    .D(_1353_),
    .Q_N(_5148_),
    .Q(\board_state_next[309] ));
 sg13g2_dfrbp_1 \board_state_next[30]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1192),
    .D(_1354_),
    .Q_N(_5147_),
    .Q(\board_state_next[30] ));
 sg13g2_dfrbp_1 \board_state_next[310]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1193),
    .D(_1355_),
    .Q_N(_5146_),
    .Q(\board_state_next[310] ));
 sg13g2_dfrbp_1 \board_state_next[311]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1194),
    .D(_1356_),
    .Q_N(_5145_),
    .Q(\board_state_next[311] ));
 sg13g2_dfrbp_1 \board_state_next[312]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1195),
    .D(_1357_),
    .Q_N(_5144_),
    .Q(\board_state_next[312] ));
 sg13g2_dfrbp_1 \board_state_next[313]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1196),
    .D(_1358_),
    .Q_N(_5143_),
    .Q(\board_state_next[313] ));
 sg13g2_dfrbp_1 \board_state_next[314]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1197),
    .D(_1359_),
    .Q_N(_5142_),
    .Q(\board_state_next[314] ));
 sg13g2_dfrbp_1 \board_state_next[315]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1198),
    .D(_1360_),
    .Q_N(_5141_),
    .Q(\board_state_next[315] ));
 sg13g2_dfrbp_1 \board_state_next[316]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1199),
    .D(_1361_),
    .Q_N(_5140_),
    .Q(\board_state_next[316] ));
 sg13g2_dfrbp_1 \board_state_next[317]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1200),
    .D(_1362_),
    .Q_N(_5139_),
    .Q(\board_state_next[317] ));
 sg13g2_dfrbp_1 \board_state_next[318]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1201),
    .D(_1363_),
    .Q_N(_5138_),
    .Q(\board_state_next[318] ));
 sg13g2_dfrbp_1 \board_state_next[319]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1202),
    .D(_1364_),
    .Q_N(_5137_),
    .Q(\board_state_next[319] ));
 sg13g2_dfrbp_1 \board_state_next[31]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1203),
    .D(_1365_),
    .Q_N(_5136_),
    .Q(\board_state_next[31] ));
 sg13g2_dfrbp_1 \board_state_next[320]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1204),
    .D(_1366_),
    .Q_N(_5135_),
    .Q(\board_state_next[320] ));
 sg13g2_dfrbp_1 \board_state_next[321]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1205),
    .D(_1367_),
    .Q_N(_5134_),
    .Q(\board_state_next[321] ));
 sg13g2_dfrbp_1 \board_state_next[322]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1206),
    .D(_1368_),
    .Q_N(_5133_),
    .Q(\board_state_next[322] ));
 sg13g2_dfrbp_1 \board_state_next[323]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1207),
    .D(_1369_),
    .Q_N(_5132_),
    .Q(\board_state_next[323] ));
 sg13g2_dfrbp_1 \board_state_next[324]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1208),
    .D(_1370_),
    .Q_N(_5131_),
    .Q(\board_state_next[324] ));
 sg13g2_dfrbp_1 \board_state_next[325]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1209),
    .D(_1371_),
    .Q_N(_5130_),
    .Q(\board_state_next[325] ));
 sg13g2_dfrbp_1 \board_state_next[326]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1210),
    .D(_1372_),
    .Q_N(_5129_),
    .Q(\board_state_next[326] ));
 sg13g2_dfrbp_1 \board_state_next[327]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1211),
    .D(_1373_),
    .Q_N(_5128_),
    .Q(\board_state_next[327] ));
 sg13g2_dfrbp_1 \board_state_next[328]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1212),
    .D(_1374_),
    .Q_N(_5127_),
    .Q(\board_state_next[328] ));
 sg13g2_dfrbp_1 \board_state_next[329]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1213),
    .D(_1375_),
    .Q_N(_5126_),
    .Q(\board_state_next[329] ));
 sg13g2_dfrbp_1 \board_state_next[32]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1214),
    .D(_1376_),
    .Q_N(_5125_),
    .Q(\board_state_next[32] ));
 sg13g2_dfrbp_1 \board_state_next[330]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1215),
    .D(_1377_),
    .Q_N(_5124_),
    .Q(\board_state_next[330] ));
 sg13g2_dfrbp_1 \board_state_next[331]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1216),
    .D(_1378_),
    .Q_N(_5123_),
    .Q(\board_state_next[331] ));
 sg13g2_dfrbp_1 \board_state_next[332]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1217),
    .D(_1379_),
    .Q_N(_5122_),
    .Q(\board_state_next[332] ));
 sg13g2_dfrbp_1 \board_state_next[333]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1218),
    .D(_1380_),
    .Q_N(_5121_),
    .Q(\board_state_next[333] ));
 sg13g2_dfrbp_1 \board_state_next[334]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1219),
    .D(_1381_),
    .Q_N(_5120_),
    .Q(\board_state_next[334] ));
 sg13g2_dfrbp_1 \board_state_next[335]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1220),
    .D(_1382_),
    .Q_N(_5119_),
    .Q(\board_state_next[335] ));
 sg13g2_dfrbp_1 \board_state_next[336]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1221),
    .D(_1383_),
    .Q_N(_5118_),
    .Q(\board_state_next[336] ));
 sg13g2_dfrbp_1 \board_state_next[337]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1222),
    .D(_1384_),
    .Q_N(_5117_),
    .Q(\board_state_next[337] ));
 sg13g2_dfrbp_1 \board_state_next[338]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1223),
    .D(_1385_),
    .Q_N(_5116_),
    .Q(\board_state_next[338] ));
 sg13g2_dfrbp_1 \board_state_next[339]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1224),
    .D(_1386_),
    .Q_N(_5115_),
    .Q(\board_state_next[339] ));
 sg13g2_dfrbp_1 \board_state_next[33]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1225),
    .D(_1387_),
    .Q_N(_5114_),
    .Q(\board_state_next[33] ));
 sg13g2_dfrbp_1 \board_state_next[340]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1226),
    .D(_1388_),
    .Q_N(_5113_),
    .Q(\board_state_next[340] ));
 sg13g2_dfrbp_1 \board_state_next[341]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1227),
    .D(_1389_),
    .Q_N(_5112_),
    .Q(\board_state_next[341] ));
 sg13g2_dfrbp_1 \board_state_next[342]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1228),
    .D(_1390_),
    .Q_N(_5111_),
    .Q(\board_state_next[342] ));
 sg13g2_dfrbp_1 \board_state_next[343]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1229),
    .D(_1391_),
    .Q_N(_5110_),
    .Q(\board_state_next[343] ));
 sg13g2_dfrbp_1 \board_state_next[344]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1230),
    .D(_1392_),
    .Q_N(_5109_),
    .Q(\board_state_next[344] ));
 sg13g2_dfrbp_1 \board_state_next[345]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1231),
    .D(_1393_),
    .Q_N(_5108_),
    .Q(\board_state_next[345] ));
 sg13g2_dfrbp_1 \board_state_next[346]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1232),
    .D(_1394_),
    .Q_N(_5107_),
    .Q(\board_state_next[346] ));
 sg13g2_dfrbp_1 \board_state_next[347]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1233),
    .D(_1395_),
    .Q_N(_5106_),
    .Q(\board_state_next[347] ));
 sg13g2_dfrbp_1 \board_state_next[348]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1234),
    .D(_1396_),
    .Q_N(_5105_),
    .Q(\board_state_next[348] ));
 sg13g2_dfrbp_1 \board_state_next[349]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1235),
    .D(_1397_),
    .Q_N(_5104_),
    .Q(\board_state_next[349] ));
 sg13g2_dfrbp_1 \board_state_next[34]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1236),
    .D(_1398_),
    .Q_N(_5103_),
    .Q(\board_state_next[34] ));
 sg13g2_dfrbp_1 \board_state_next[350]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1237),
    .D(_1399_),
    .Q_N(_5102_),
    .Q(\board_state_next[350] ));
 sg13g2_dfrbp_1 \board_state_next[351]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1238),
    .D(_1400_),
    .Q_N(_5101_),
    .Q(\board_state_next[351] ));
 sg13g2_dfrbp_1 \board_state_next[352]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1239),
    .D(_1401_),
    .Q_N(_5100_),
    .Q(\board_state_next[352] ));
 sg13g2_dfrbp_1 \board_state_next[353]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1240),
    .D(_1402_),
    .Q_N(_5099_),
    .Q(\board_state_next[353] ));
 sg13g2_dfrbp_1 \board_state_next[354]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1241),
    .D(_1403_),
    .Q_N(_5098_),
    .Q(\board_state_next[354] ));
 sg13g2_dfrbp_1 \board_state_next[355]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1242),
    .D(_1404_),
    .Q_N(_5097_),
    .Q(\board_state_next[355] ));
 sg13g2_dfrbp_1 \board_state_next[356]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1243),
    .D(_1405_),
    .Q_N(_5096_),
    .Q(\board_state_next[356] ));
 sg13g2_dfrbp_1 \board_state_next[357]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1244),
    .D(_1406_),
    .Q_N(_5095_),
    .Q(\board_state_next[357] ));
 sg13g2_dfrbp_1 \board_state_next[358]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1245),
    .D(_1407_),
    .Q_N(_5094_),
    .Q(\board_state_next[358] ));
 sg13g2_dfrbp_1 \board_state_next[359]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1246),
    .D(_1408_),
    .Q_N(_5093_),
    .Q(\board_state_next[359] ));
 sg13g2_dfrbp_1 \board_state_next[35]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1247),
    .D(_1409_),
    .Q_N(_5092_),
    .Q(\board_state_next[35] ));
 sg13g2_dfrbp_1 \board_state_next[360]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1248),
    .D(_1410_),
    .Q_N(_5091_),
    .Q(\board_state_next[360] ));
 sg13g2_dfrbp_1 \board_state_next[361]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1249),
    .D(_1411_),
    .Q_N(_5090_),
    .Q(\board_state_next[361] ));
 sg13g2_dfrbp_1 \board_state_next[362]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1250),
    .D(_1412_),
    .Q_N(_5089_),
    .Q(\board_state_next[362] ));
 sg13g2_dfrbp_1 \board_state_next[363]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1251),
    .D(_1413_),
    .Q_N(_5088_),
    .Q(\board_state_next[363] ));
 sg13g2_dfrbp_1 \board_state_next[364]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1252),
    .D(_1414_),
    .Q_N(_5087_),
    .Q(\board_state_next[364] ));
 sg13g2_dfrbp_1 \board_state_next[365]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1253),
    .D(_1415_),
    .Q_N(_5086_),
    .Q(\board_state_next[365] ));
 sg13g2_dfrbp_1 \board_state_next[366]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1254),
    .D(_1416_),
    .Q_N(_5085_),
    .Q(\board_state_next[366] ));
 sg13g2_dfrbp_1 \board_state_next[367]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1255),
    .D(_1417_),
    .Q_N(_5084_),
    .Q(\board_state_next[367] ));
 sg13g2_dfrbp_1 \board_state_next[368]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1256),
    .D(_1418_),
    .Q_N(_5083_),
    .Q(\board_state_next[368] ));
 sg13g2_dfrbp_1 \board_state_next[369]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1257),
    .D(_1419_),
    .Q_N(_5082_),
    .Q(\board_state_next[369] ));
 sg13g2_dfrbp_1 \board_state_next[36]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1258),
    .D(_1420_),
    .Q_N(_5081_),
    .Q(\board_state_next[36] ));
 sg13g2_dfrbp_1 \board_state_next[370]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1259),
    .D(_1421_),
    .Q_N(_5080_),
    .Q(\board_state_next[370] ));
 sg13g2_dfrbp_1 \board_state_next[371]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1260),
    .D(_1422_),
    .Q_N(_5079_),
    .Q(\board_state_next[371] ));
 sg13g2_dfrbp_1 \board_state_next[372]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1261),
    .D(_1423_),
    .Q_N(_5078_),
    .Q(\board_state_next[372] ));
 sg13g2_dfrbp_1 \board_state_next[373]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1262),
    .D(_1424_),
    .Q_N(_5077_),
    .Q(\board_state_next[373] ));
 sg13g2_dfrbp_1 \board_state_next[374]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1263),
    .D(_1425_),
    .Q_N(_5076_),
    .Q(\board_state_next[374] ));
 sg13g2_dfrbp_1 \board_state_next[375]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1264),
    .D(_1426_),
    .Q_N(_5075_),
    .Q(\board_state_next[375] ));
 sg13g2_dfrbp_1 \board_state_next[376]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1265),
    .D(_1427_),
    .Q_N(_5074_),
    .Q(\board_state_next[376] ));
 sg13g2_dfrbp_1 \board_state_next[377]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1266),
    .D(_1428_),
    .Q_N(_5073_),
    .Q(\board_state_next[377] ));
 sg13g2_dfrbp_1 \board_state_next[378]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1267),
    .D(_1429_),
    .Q_N(_5072_),
    .Q(\board_state_next[378] ));
 sg13g2_dfrbp_1 \board_state_next[379]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1268),
    .D(_1430_),
    .Q_N(_5071_),
    .Q(\board_state_next[379] ));
 sg13g2_dfrbp_1 \board_state_next[37]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1269),
    .D(_1431_),
    .Q_N(_5070_),
    .Q(\board_state_next[37] ));
 sg13g2_dfrbp_1 \board_state_next[380]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1270),
    .D(_1432_),
    .Q_N(_5069_),
    .Q(\board_state_next[380] ));
 sg13g2_dfrbp_1 \board_state_next[381]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1271),
    .D(_1433_),
    .Q_N(_5068_),
    .Q(\board_state_next[381] ));
 sg13g2_dfrbp_1 \board_state_next[382]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1272),
    .D(_1434_),
    .Q_N(_5067_),
    .Q(\board_state_next[382] ));
 sg13g2_dfrbp_1 \board_state_next[383]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1273),
    .D(_1435_),
    .Q_N(_5066_),
    .Q(\board_state_next[383] ));
 sg13g2_dfrbp_1 \board_state_next[384]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1274),
    .D(_1436_),
    .Q_N(_5065_),
    .Q(\board_state_next[384] ));
 sg13g2_dfrbp_1 \board_state_next[385]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1275),
    .D(_1437_),
    .Q_N(_5064_),
    .Q(\board_state_next[385] ));
 sg13g2_dfrbp_1 \board_state_next[386]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1276),
    .D(_1438_),
    .Q_N(_5063_),
    .Q(\board_state_next[386] ));
 sg13g2_dfrbp_1 \board_state_next[387]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1277),
    .D(_1439_),
    .Q_N(_5062_),
    .Q(\board_state_next[387] ));
 sg13g2_dfrbp_1 \board_state_next[388]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1278),
    .D(_1440_),
    .Q_N(_5061_),
    .Q(\board_state_next[388] ));
 sg13g2_dfrbp_1 \board_state_next[389]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1279),
    .D(_1441_),
    .Q_N(_5060_),
    .Q(\board_state_next[389] ));
 sg13g2_dfrbp_1 \board_state_next[38]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1280),
    .D(_1442_),
    .Q_N(_5059_),
    .Q(\board_state_next[38] ));
 sg13g2_dfrbp_1 \board_state_next[390]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1281),
    .D(_1443_),
    .Q_N(_5058_),
    .Q(\board_state_next[390] ));
 sg13g2_dfrbp_1 \board_state_next[391]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1282),
    .D(_1444_),
    .Q_N(_5057_),
    .Q(\board_state_next[391] ));
 sg13g2_dfrbp_1 \board_state_next[392]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1283),
    .D(_1445_),
    .Q_N(_5056_),
    .Q(\board_state_next[392] ));
 sg13g2_dfrbp_1 \board_state_next[393]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1284),
    .D(_1446_),
    .Q_N(_5055_),
    .Q(\board_state_next[393] ));
 sg13g2_dfrbp_1 \board_state_next[394]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1285),
    .D(_1447_),
    .Q_N(_5054_),
    .Q(\board_state_next[394] ));
 sg13g2_dfrbp_1 \board_state_next[395]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1286),
    .D(_1448_),
    .Q_N(_5053_),
    .Q(\board_state_next[395] ));
 sg13g2_dfrbp_1 \board_state_next[396]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1287),
    .D(_1449_),
    .Q_N(_5052_),
    .Q(\board_state_next[396] ));
 sg13g2_dfrbp_1 \board_state_next[397]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1288),
    .D(_1450_),
    .Q_N(_5051_),
    .Q(\board_state_next[397] ));
 sg13g2_dfrbp_1 \board_state_next[398]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1289),
    .D(_1451_),
    .Q_N(_5050_),
    .Q(\board_state_next[398] ));
 sg13g2_dfrbp_1 \board_state_next[399]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1290),
    .D(_1452_),
    .Q_N(_5049_),
    .Q(\board_state_next[399] ));
 sg13g2_dfrbp_1 \board_state_next[39]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1291),
    .D(_1453_),
    .Q_N(_5048_),
    .Q(\board_state_next[39] ));
 sg13g2_dfrbp_1 \board_state_next[3]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1292),
    .D(_1454_),
    .Q_N(_5047_),
    .Q(\board_state_next[3] ));
 sg13g2_dfrbp_1 \board_state_next[400]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1293),
    .D(_1455_),
    .Q_N(_5046_),
    .Q(\board_state_next[400] ));
 sg13g2_dfrbp_1 \board_state_next[401]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1294),
    .D(_1456_),
    .Q_N(_5045_),
    .Q(\board_state_next[401] ));
 sg13g2_dfrbp_1 \board_state_next[402]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1295),
    .D(_1457_),
    .Q_N(_5044_),
    .Q(\board_state_next[402] ));
 sg13g2_dfrbp_1 \board_state_next[403]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1296),
    .D(_1458_),
    .Q_N(_5043_),
    .Q(\board_state_next[403] ));
 sg13g2_dfrbp_1 \board_state_next[404]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1297),
    .D(_1459_),
    .Q_N(_5042_),
    .Q(\board_state_next[404] ));
 sg13g2_dfrbp_1 \board_state_next[405]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1298),
    .D(_1460_),
    .Q_N(_5041_),
    .Q(\board_state_next[405] ));
 sg13g2_dfrbp_1 \board_state_next[406]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1299),
    .D(_1461_),
    .Q_N(_5040_),
    .Q(\board_state_next[406] ));
 sg13g2_dfrbp_1 \board_state_next[407]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1300),
    .D(_1462_),
    .Q_N(_5039_),
    .Q(\board_state_next[407] ));
 sg13g2_dfrbp_1 \board_state_next[408]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1301),
    .D(_1463_),
    .Q_N(_5038_),
    .Q(\board_state_next[408] ));
 sg13g2_dfrbp_1 \board_state_next[409]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1302),
    .D(_1464_),
    .Q_N(_5037_),
    .Q(\board_state_next[409] ));
 sg13g2_dfrbp_1 \board_state_next[40]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1303),
    .D(_1465_),
    .Q_N(_5036_),
    .Q(\board_state_next[40] ));
 sg13g2_dfrbp_1 \board_state_next[410]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1304),
    .D(_1466_),
    .Q_N(_5035_),
    .Q(\board_state_next[410] ));
 sg13g2_dfrbp_1 \board_state_next[411]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1305),
    .D(_1467_),
    .Q_N(_5034_),
    .Q(\board_state_next[411] ));
 sg13g2_dfrbp_1 \board_state_next[412]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1306),
    .D(_1468_),
    .Q_N(_5033_),
    .Q(\board_state_next[412] ));
 sg13g2_dfrbp_1 \board_state_next[413]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1307),
    .D(_1469_),
    .Q_N(_5032_),
    .Q(\board_state_next[413] ));
 sg13g2_dfrbp_1 \board_state_next[414]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1308),
    .D(_1470_),
    .Q_N(_5031_),
    .Q(\board_state_next[414] ));
 sg13g2_dfrbp_1 \board_state_next[415]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1309),
    .D(_1471_),
    .Q_N(_5030_),
    .Q(\board_state_next[415] ));
 sg13g2_dfrbp_1 \board_state_next[416]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1310),
    .D(_1472_),
    .Q_N(_5029_),
    .Q(\board_state_next[416] ));
 sg13g2_dfrbp_1 \board_state_next[417]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1311),
    .D(_1473_),
    .Q_N(_5028_),
    .Q(\board_state_next[417] ));
 sg13g2_dfrbp_1 \board_state_next[418]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1312),
    .D(_1474_),
    .Q_N(_5027_),
    .Q(\board_state_next[418] ));
 sg13g2_dfrbp_1 \board_state_next[419]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1313),
    .D(_1475_),
    .Q_N(_5026_),
    .Q(\board_state_next[419] ));
 sg13g2_dfrbp_1 \board_state_next[41]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1314),
    .D(_1476_),
    .Q_N(_5025_),
    .Q(\board_state_next[41] ));
 sg13g2_dfrbp_1 \board_state_next[420]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1315),
    .D(_1477_),
    .Q_N(_5024_),
    .Q(\board_state_next[420] ));
 sg13g2_dfrbp_1 \board_state_next[421]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1316),
    .D(_1478_),
    .Q_N(_5023_),
    .Q(\board_state_next[421] ));
 sg13g2_dfrbp_1 \board_state_next[422]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1317),
    .D(_1479_),
    .Q_N(_5022_),
    .Q(\board_state_next[422] ));
 sg13g2_dfrbp_1 \board_state_next[423]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1318),
    .D(_1480_),
    .Q_N(_5021_),
    .Q(\board_state_next[423] ));
 sg13g2_dfrbp_1 \board_state_next[424]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1319),
    .D(_1481_),
    .Q_N(_5020_),
    .Q(\board_state_next[424] ));
 sg13g2_dfrbp_1 \board_state_next[425]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1320),
    .D(_1482_),
    .Q_N(_5019_),
    .Q(\board_state_next[425] ));
 sg13g2_dfrbp_1 \board_state_next[426]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1321),
    .D(_1483_),
    .Q_N(_5018_),
    .Q(\board_state_next[426] ));
 sg13g2_dfrbp_1 \board_state_next[427]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1322),
    .D(_1484_),
    .Q_N(_5017_),
    .Q(\board_state_next[427] ));
 sg13g2_dfrbp_1 \board_state_next[428]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1323),
    .D(_1485_),
    .Q_N(_5016_),
    .Q(\board_state_next[428] ));
 sg13g2_dfrbp_1 \board_state_next[429]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1324),
    .D(_1486_),
    .Q_N(_5015_),
    .Q(\board_state_next[429] ));
 sg13g2_dfrbp_1 \board_state_next[42]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1325),
    .D(_1487_),
    .Q_N(_5014_),
    .Q(\board_state_next[42] ));
 sg13g2_dfrbp_1 \board_state_next[430]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1326),
    .D(_1488_),
    .Q_N(_5013_),
    .Q(\board_state_next[430] ));
 sg13g2_dfrbp_1 \board_state_next[431]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1327),
    .D(_1489_),
    .Q_N(_5012_),
    .Q(\board_state_next[431] ));
 sg13g2_dfrbp_1 \board_state_next[432]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1328),
    .D(_1490_),
    .Q_N(_5011_),
    .Q(\board_state_next[432] ));
 sg13g2_dfrbp_1 \board_state_next[433]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1329),
    .D(_1491_),
    .Q_N(_5010_),
    .Q(\board_state_next[433] ));
 sg13g2_dfrbp_1 \board_state_next[434]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1330),
    .D(_1492_),
    .Q_N(_5009_),
    .Q(\board_state_next[434] ));
 sg13g2_dfrbp_1 \board_state_next[435]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1331),
    .D(_1493_),
    .Q_N(_5008_),
    .Q(\board_state_next[435] ));
 sg13g2_dfrbp_1 \board_state_next[436]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1332),
    .D(_1494_),
    .Q_N(_5007_),
    .Q(\board_state_next[436] ));
 sg13g2_dfrbp_1 \board_state_next[437]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1333),
    .D(_1495_),
    .Q_N(_5006_),
    .Q(\board_state_next[437] ));
 sg13g2_dfrbp_1 \board_state_next[438]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1334),
    .D(_1496_),
    .Q_N(_5005_),
    .Q(\board_state_next[438] ));
 sg13g2_dfrbp_1 \board_state_next[439]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1335),
    .D(_1497_),
    .Q_N(_5004_),
    .Q(\board_state_next[439] ));
 sg13g2_dfrbp_1 \board_state_next[43]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1336),
    .D(_1498_),
    .Q_N(_5003_),
    .Q(\board_state_next[43] ));
 sg13g2_dfrbp_1 \board_state_next[440]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1337),
    .D(_1499_),
    .Q_N(_5002_),
    .Q(\board_state_next[440] ));
 sg13g2_dfrbp_1 \board_state_next[441]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1338),
    .D(_1500_),
    .Q_N(_5001_),
    .Q(\board_state_next[441] ));
 sg13g2_dfrbp_1 \board_state_next[442]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1339),
    .D(_1501_),
    .Q_N(_5000_),
    .Q(\board_state_next[442] ));
 sg13g2_dfrbp_1 \board_state_next[443]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1340),
    .D(_1502_),
    .Q_N(_4999_),
    .Q(\board_state_next[443] ));
 sg13g2_dfrbp_1 \board_state_next[444]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1341),
    .D(_1503_),
    .Q_N(_4998_),
    .Q(\board_state_next[444] ));
 sg13g2_dfrbp_1 \board_state_next[445]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1342),
    .D(_1504_),
    .Q_N(_4997_),
    .Q(\board_state_next[445] ));
 sg13g2_dfrbp_1 \board_state_next[446]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1343),
    .D(_1505_),
    .Q_N(_4996_),
    .Q(\board_state_next[446] ));
 sg13g2_dfrbp_1 \board_state_next[447]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1344),
    .D(_1506_),
    .Q_N(_4995_),
    .Q(\board_state_next[447] ));
 sg13g2_dfrbp_1 \board_state_next[448]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1345),
    .D(_1507_),
    .Q_N(_4994_),
    .Q(\board_state_next[448] ));
 sg13g2_dfrbp_1 \board_state_next[449]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1346),
    .D(_1508_),
    .Q_N(_4993_),
    .Q(\board_state_next[449] ));
 sg13g2_dfrbp_1 \board_state_next[44]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1347),
    .D(_1509_),
    .Q_N(_4992_),
    .Q(\board_state_next[44] ));
 sg13g2_dfrbp_1 \board_state_next[450]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1348),
    .D(_1510_),
    .Q_N(_4991_),
    .Q(\board_state_next[450] ));
 sg13g2_dfrbp_1 \board_state_next[451]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1349),
    .D(_1511_),
    .Q_N(_4990_),
    .Q(\board_state_next[451] ));
 sg13g2_dfrbp_1 \board_state_next[452]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1350),
    .D(_1512_),
    .Q_N(_4989_),
    .Q(\board_state_next[452] ));
 sg13g2_dfrbp_1 \board_state_next[453]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1351),
    .D(_1513_),
    .Q_N(_4988_),
    .Q(\board_state_next[453] ));
 sg13g2_dfrbp_1 \board_state_next[454]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1352),
    .D(_1514_),
    .Q_N(_4987_),
    .Q(\board_state_next[454] ));
 sg13g2_dfrbp_1 \board_state_next[455]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1353),
    .D(_1515_),
    .Q_N(_4986_),
    .Q(\board_state_next[455] ));
 sg13g2_dfrbp_1 \board_state_next[456]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1354),
    .D(_1516_),
    .Q_N(_4985_),
    .Q(\board_state_next[456] ));
 sg13g2_dfrbp_1 \board_state_next[457]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1355),
    .D(_1517_),
    .Q_N(_4984_),
    .Q(\board_state_next[457] ));
 sg13g2_dfrbp_1 \board_state_next[458]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1356),
    .D(_1518_),
    .Q_N(_4983_),
    .Q(\board_state_next[458] ));
 sg13g2_dfrbp_1 \board_state_next[459]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1357),
    .D(_1519_),
    .Q_N(_4982_),
    .Q(\board_state_next[459] ));
 sg13g2_dfrbp_1 \board_state_next[45]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1358),
    .D(_1520_),
    .Q_N(_4981_),
    .Q(\board_state_next[45] ));
 sg13g2_dfrbp_1 \board_state_next[460]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1359),
    .D(_1521_),
    .Q_N(_4980_),
    .Q(\board_state_next[460] ));
 sg13g2_dfrbp_1 \board_state_next[461]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1360),
    .D(_1522_),
    .Q_N(_4979_),
    .Q(\board_state_next[461] ));
 sg13g2_dfrbp_1 \board_state_next[462]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1361),
    .D(_1523_),
    .Q_N(_4978_),
    .Q(\board_state_next[462] ));
 sg13g2_dfrbp_1 \board_state_next[463]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1362),
    .D(_1524_),
    .Q_N(_4977_),
    .Q(\board_state_next[463] ));
 sg13g2_dfrbp_1 \board_state_next[464]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1363),
    .D(_1525_),
    .Q_N(_4976_),
    .Q(\board_state_next[464] ));
 sg13g2_dfrbp_1 \board_state_next[465]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1364),
    .D(_1526_),
    .Q_N(_4975_),
    .Q(\board_state_next[465] ));
 sg13g2_dfrbp_1 \board_state_next[466]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1365),
    .D(_1527_),
    .Q_N(_4974_),
    .Q(\board_state_next[466] ));
 sg13g2_dfrbp_1 \board_state_next[467]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1366),
    .D(_1528_),
    .Q_N(_4973_),
    .Q(\board_state_next[467] ));
 sg13g2_dfrbp_1 \board_state_next[468]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1367),
    .D(_1529_),
    .Q_N(_4972_),
    .Q(\board_state_next[468] ));
 sg13g2_dfrbp_1 \board_state_next[469]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1368),
    .D(_1530_),
    .Q_N(_4971_),
    .Q(\board_state_next[469] ));
 sg13g2_dfrbp_1 \board_state_next[46]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1369),
    .D(_1531_),
    .Q_N(_4970_),
    .Q(\board_state_next[46] ));
 sg13g2_dfrbp_1 \board_state_next[470]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1370),
    .D(_1532_),
    .Q_N(_4969_),
    .Q(\board_state_next[470] ));
 sg13g2_dfrbp_1 \board_state_next[471]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1371),
    .D(_1533_),
    .Q_N(_4968_),
    .Q(\board_state_next[471] ));
 sg13g2_dfrbp_1 \board_state_next[472]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1372),
    .D(_1534_),
    .Q_N(_4967_),
    .Q(\board_state_next[472] ));
 sg13g2_dfrbp_1 \board_state_next[473]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1373),
    .D(_1535_),
    .Q_N(_4966_),
    .Q(\board_state_next[473] ));
 sg13g2_dfrbp_1 \board_state_next[474]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1374),
    .D(_1536_),
    .Q_N(_4965_),
    .Q(\board_state_next[474] ));
 sg13g2_dfrbp_1 \board_state_next[475]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1375),
    .D(_1537_),
    .Q_N(_4964_),
    .Q(\board_state_next[475] ));
 sg13g2_dfrbp_1 \board_state_next[476]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1376),
    .D(_1538_),
    .Q_N(_4963_),
    .Q(\board_state_next[476] ));
 sg13g2_dfrbp_1 \board_state_next[477]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1377),
    .D(_1539_),
    .Q_N(_4962_),
    .Q(\board_state_next[477] ));
 sg13g2_dfrbp_1 \board_state_next[478]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1378),
    .D(_1540_),
    .Q_N(_4961_),
    .Q(\board_state_next[478] ));
 sg13g2_dfrbp_1 \board_state_next[479]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1379),
    .D(_1541_),
    .Q_N(_4960_),
    .Q(\board_state_next[479] ));
 sg13g2_dfrbp_1 \board_state_next[47]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1380),
    .D(_1542_),
    .Q_N(_4959_),
    .Q(\board_state_next[47] ));
 sg13g2_dfrbp_1 \board_state_next[480]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1381),
    .D(_1543_),
    .Q_N(_4958_),
    .Q(\board_state_next[480] ));
 sg13g2_dfrbp_1 \board_state_next[481]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1382),
    .D(_1544_),
    .Q_N(_4957_),
    .Q(\board_state_next[481] ));
 sg13g2_dfrbp_1 \board_state_next[482]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1383),
    .D(_1545_),
    .Q_N(_4956_),
    .Q(\board_state_next[482] ));
 sg13g2_dfrbp_1 \board_state_next[483]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1384),
    .D(_1546_),
    .Q_N(_4955_),
    .Q(\board_state_next[483] ));
 sg13g2_dfrbp_1 \board_state_next[484]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1385),
    .D(_1547_),
    .Q_N(_4954_),
    .Q(\board_state_next[484] ));
 sg13g2_dfrbp_1 \board_state_next[485]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1386),
    .D(_1548_),
    .Q_N(_4953_),
    .Q(\board_state_next[485] ));
 sg13g2_dfrbp_1 \board_state_next[486]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1387),
    .D(_1549_),
    .Q_N(_4952_),
    .Q(\board_state_next[486] ));
 sg13g2_dfrbp_1 \board_state_next[487]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1388),
    .D(_1550_),
    .Q_N(_4951_),
    .Q(\board_state_next[487] ));
 sg13g2_dfrbp_1 \board_state_next[488]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1389),
    .D(_1551_),
    .Q_N(_4950_),
    .Q(\board_state_next[488] ));
 sg13g2_dfrbp_1 \board_state_next[489]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1390),
    .D(_1552_),
    .Q_N(_4949_),
    .Q(\board_state_next[489] ));
 sg13g2_dfrbp_1 \board_state_next[48]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1391),
    .D(_1553_),
    .Q_N(_4948_),
    .Q(\board_state_next[48] ));
 sg13g2_dfrbp_1 \board_state_next[490]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1392),
    .D(_1554_),
    .Q_N(_4947_),
    .Q(\board_state_next[490] ));
 sg13g2_dfrbp_1 \board_state_next[491]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1393),
    .D(_1555_),
    .Q_N(_4946_),
    .Q(\board_state_next[491] ));
 sg13g2_dfrbp_1 \board_state_next[492]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1394),
    .D(_1556_),
    .Q_N(_4945_),
    .Q(\board_state_next[492] ));
 sg13g2_dfrbp_1 \board_state_next[493]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1395),
    .D(_1557_),
    .Q_N(_4944_),
    .Q(\board_state_next[493] ));
 sg13g2_dfrbp_1 \board_state_next[494]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1396),
    .D(_1558_),
    .Q_N(_4943_),
    .Q(\board_state_next[494] ));
 sg13g2_dfrbp_1 \board_state_next[495]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1397),
    .D(_1559_),
    .Q_N(_4942_),
    .Q(\board_state_next[495] ));
 sg13g2_dfrbp_1 \board_state_next[496]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1398),
    .D(_1560_),
    .Q_N(_4941_),
    .Q(\board_state_next[496] ));
 sg13g2_dfrbp_1 \board_state_next[497]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1399),
    .D(_1561_),
    .Q_N(_4940_),
    .Q(\board_state_next[497] ));
 sg13g2_dfrbp_1 \board_state_next[498]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1400),
    .D(_1562_),
    .Q_N(_4939_),
    .Q(\board_state_next[498] ));
 sg13g2_dfrbp_1 \board_state_next[499]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1401),
    .D(_1563_),
    .Q_N(_4938_),
    .Q(\board_state_next[499] ));
 sg13g2_dfrbp_1 \board_state_next[49]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1402),
    .D(_1564_),
    .Q_N(_4937_),
    .Q(\board_state_next[49] ));
 sg13g2_dfrbp_1 \board_state_next[4]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1403),
    .D(_1565_),
    .Q_N(_4936_),
    .Q(\board_state_next[4] ));
 sg13g2_dfrbp_1 \board_state_next[500]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1404),
    .D(_1566_),
    .Q_N(_4935_),
    .Q(\board_state_next[500] ));
 sg13g2_dfrbp_1 \board_state_next[501]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1405),
    .D(_1567_),
    .Q_N(_4934_),
    .Q(\board_state_next[501] ));
 sg13g2_dfrbp_1 \board_state_next[502]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1406),
    .D(_1568_),
    .Q_N(_4933_),
    .Q(\board_state_next[502] ));
 sg13g2_dfrbp_1 \board_state_next[503]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1407),
    .D(_1569_),
    .Q_N(_4932_),
    .Q(\board_state_next[503] ));
 sg13g2_dfrbp_1 \board_state_next[504]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1408),
    .D(_1570_),
    .Q_N(_4931_),
    .Q(\board_state_next[504] ));
 sg13g2_dfrbp_1 \board_state_next[505]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1409),
    .D(_1571_),
    .Q_N(_4930_),
    .Q(\board_state_next[505] ));
 sg13g2_dfrbp_1 \board_state_next[506]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1410),
    .D(_1572_),
    .Q_N(_4929_),
    .Q(\board_state_next[506] ));
 sg13g2_dfrbp_1 \board_state_next[507]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1411),
    .D(_1573_),
    .Q_N(_4928_),
    .Q(\board_state_next[507] ));
 sg13g2_dfrbp_1 \board_state_next[508]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1412),
    .D(_1574_),
    .Q_N(_4927_),
    .Q(\board_state_next[508] ));
 sg13g2_dfrbp_1 \board_state_next[509]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1413),
    .D(_1575_),
    .Q_N(_4926_),
    .Q(\board_state_next[509] ));
 sg13g2_dfrbp_1 \board_state_next[50]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1414),
    .D(_1576_),
    .Q_N(_4925_),
    .Q(\board_state_next[50] ));
 sg13g2_dfrbp_1 \board_state_next[510]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1415),
    .D(_1577_),
    .Q_N(_4924_),
    .Q(\board_state_next[510] ));
 sg13g2_dfrbp_1 \board_state_next[511]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1416),
    .D(_1578_),
    .Q_N(_4923_),
    .Q(\board_state_next[511] ));
 sg13g2_dfrbp_1 \board_state_next[51]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1417),
    .D(_1579_),
    .Q_N(_4922_),
    .Q(\board_state_next[51] ));
 sg13g2_dfrbp_1 \board_state_next[52]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1418),
    .D(_1580_),
    .Q_N(_4921_),
    .Q(\board_state_next[52] ));
 sg13g2_dfrbp_1 \board_state_next[53]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1419),
    .D(_1581_),
    .Q_N(_4920_),
    .Q(\board_state_next[53] ));
 sg13g2_dfrbp_1 \board_state_next[54]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1420),
    .D(_1582_),
    .Q_N(_4919_),
    .Q(\board_state_next[54] ));
 sg13g2_dfrbp_1 \board_state_next[55]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1421),
    .D(_1583_),
    .Q_N(_4918_),
    .Q(\board_state_next[55] ));
 sg13g2_dfrbp_1 \board_state_next[56]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1422),
    .D(_1584_),
    .Q_N(_4917_),
    .Q(\board_state_next[56] ));
 sg13g2_dfrbp_1 \board_state_next[57]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1423),
    .D(_1585_),
    .Q_N(_4916_),
    .Q(\board_state_next[57] ));
 sg13g2_dfrbp_1 \board_state_next[58]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1424),
    .D(_1586_),
    .Q_N(_4915_),
    .Q(\board_state_next[58] ));
 sg13g2_dfrbp_1 \board_state_next[59]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1425),
    .D(_1587_),
    .Q_N(_4914_),
    .Q(\board_state_next[59] ));
 sg13g2_dfrbp_1 \board_state_next[5]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1426),
    .D(_1588_),
    .Q_N(_4913_),
    .Q(\board_state_next[5] ));
 sg13g2_dfrbp_1 \board_state_next[60]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1427),
    .D(_1589_),
    .Q_N(_4912_),
    .Q(\board_state_next[60] ));
 sg13g2_dfrbp_1 \board_state_next[61]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1428),
    .D(_1590_),
    .Q_N(_4911_),
    .Q(\board_state_next[61] ));
 sg13g2_dfrbp_1 \board_state_next[62]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1429),
    .D(_1591_),
    .Q_N(_4910_),
    .Q(\board_state_next[62] ));
 sg13g2_dfrbp_1 \board_state_next[63]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1430),
    .D(_1592_),
    .Q_N(_4909_),
    .Q(\board_state_next[63] ));
 sg13g2_dfrbp_1 \board_state_next[64]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1431),
    .D(_1593_),
    .Q_N(_4908_),
    .Q(\board_state_next[64] ));
 sg13g2_dfrbp_1 \board_state_next[65]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1432),
    .D(_1594_),
    .Q_N(_4907_),
    .Q(\board_state_next[65] ));
 sg13g2_dfrbp_1 \board_state_next[66]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1433),
    .D(_1595_),
    .Q_N(_4906_),
    .Q(\board_state_next[66] ));
 sg13g2_dfrbp_1 \board_state_next[67]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1434),
    .D(_1596_),
    .Q_N(_4905_),
    .Q(\board_state_next[67] ));
 sg13g2_dfrbp_1 \board_state_next[68]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1435),
    .D(_1597_),
    .Q_N(_4904_),
    .Q(\board_state_next[68] ));
 sg13g2_dfrbp_1 \board_state_next[69]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1436),
    .D(_1598_),
    .Q_N(_4903_),
    .Q(\board_state_next[69] ));
 sg13g2_dfrbp_1 \board_state_next[6]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1437),
    .D(_1599_),
    .Q_N(_4902_),
    .Q(\board_state_next[6] ));
 sg13g2_dfrbp_1 \board_state_next[70]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1438),
    .D(_1600_),
    .Q_N(_4901_),
    .Q(\board_state_next[70] ));
 sg13g2_dfrbp_1 \board_state_next[71]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1439),
    .D(_1601_),
    .Q_N(_4900_),
    .Q(\board_state_next[71] ));
 sg13g2_dfrbp_1 \board_state_next[72]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1440),
    .D(_1602_),
    .Q_N(_4899_),
    .Q(\board_state_next[72] ));
 sg13g2_dfrbp_1 \board_state_next[73]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1441),
    .D(_1603_),
    .Q_N(_4898_),
    .Q(\board_state_next[73] ));
 sg13g2_dfrbp_1 \board_state_next[74]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1442),
    .D(_1604_),
    .Q_N(_4897_),
    .Q(\board_state_next[74] ));
 sg13g2_dfrbp_1 \board_state_next[75]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1443),
    .D(_1605_),
    .Q_N(_4896_),
    .Q(\board_state_next[75] ));
 sg13g2_dfrbp_1 \board_state_next[76]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1444),
    .D(_1606_),
    .Q_N(_4895_),
    .Q(\board_state_next[76] ));
 sg13g2_dfrbp_1 \board_state_next[77]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1445),
    .D(_1607_),
    .Q_N(_4894_),
    .Q(\board_state_next[77] ));
 sg13g2_dfrbp_1 \board_state_next[78]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1446),
    .D(_1608_),
    .Q_N(_4893_),
    .Q(\board_state_next[78] ));
 sg13g2_dfrbp_1 \board_state_next[79]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1447),
    .D(_1609_),
    .Q_N(_4892_),
    .Q(\board_state_next[79] ));
 sg13g2_dfrbp_1 \board_state_next[7]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1448),
    .D(_1610_),
    .Q_N(_4891_),
    .Q(\board_state_next[7] ));
 sg13g2_dfrbp_1 \board_state_next[80]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1449),
    .D(_1611_),
    .Q_N(_4890_),
    .Q(\board_state_next[80] ));
 sg13g2_dfrbp_1 \board_state_next[81]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1450),
    .D(_1612_),
    .Q_N(_4889_),
    .Q(\board_state_next[81] ));
 sg13g2_dfrbp_1 \board_state_next[82]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1451),
    .D(_1613_),
    .Q_N(_4888_),
    .Q(\board_state_next[82] ));
 sg13g2_dfrbp_1 \board_state_next[83]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1452),
    .D(_1614_),
    .Q_N(_4887_),
    .Q(\board_state_next[83] ));
 sg13g2_dfrbp_1 \board_state_next[84]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1453),
    .D(_1615_),
    .Q_N(_4886_),
    .Q(\board_state_next[84] ));
 sg13g2_dfrbp_1 \board_state_next[85]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1454),
    .D(_1616_),
    .Q_N(_4885_),
    .Q(\board_state_next[85] ));
 sg13g2_dfrbp_1 \board_state_next[86]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1455),
    .D(_1617_),
    .Q_N(_4884_),
    .Q(\board_state_next[86] ));
 sg13g2_dfrbp_1 \board_state_next[87]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1456),
    .D(_1618_),
    .Q_N(_4883_),
    .Q(\board_state_next[87] ));
 sg13g2_dfrbp_1 \board_state_next[88]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1457),
    .D(_1619_),
    .Q_N(_4882_),
    .Q(\board_state_next[88] ));
 sg13g2_dfrbp_1 \board_state_next[89]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1458),
    .D(_1620_),
    .Q_N(_4881_),
    .Q(\board_state_next[89] ));
 sg13g2_dfrbp_1 \board_state_next[8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1459),
    .D(_1621_),
    .Q_N(_4880_),
    .Q(\board_state_next[8] ));
 sg13g2_dfrbp_1 \board_state_next[90]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1460),
    .D(_1622_),
    .Q_N(_4879_),
    .Q(\board_state_next[90] ));
 sg13g2_dfrbp_1 \board_state_next[91]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1461),
    .D(_1623_),
    .Q_N(_4878_),
    .Q(\board_state_next[91] ));
 sg13g2_dfrbp_1 \board_state_next[92]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1462),
    .D(_1624_),
    .Q_N(_4877_),
    .Q(\board_state_next[92] ));
 sg13g2_dfrbp_1 \board_state_next[93]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1463),
    .D(_1625_),
    .Q_N(_4876_),
    .Q(\board_state_next[93] ));
 sg13g2_dfrbp_1 \board_state_next[94]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1464),
    .D(_1626_),
    .Q_N(_4875_),
    .Q(\board_state_next[94] ));
 sg13g2_dfrbp_1 \board_state_next[95]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1465),
    .D(_1627_),
    .Q_N(_4874_),
    .Q(\board_state_next[95] ));
 sg13g2_dfrbp_1 \board_state_next[96]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1466),
    .D(_1628_),
    .Q_N(_4873_),
    .Q(\board_state_next[96] ));
 sg13g2_dfrbp_1 \board_state_next[97]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1467),
    .D(_1629_),
    .Q_N(_4872_),
    .Q(\board_state_next[97] ));
 sg13g2_dfrbp_1 \board_state_next[98]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1468),
    .D(_1630_),
    .Q_N(_4871_),
    .Q(\board_state_next[98] ));
 sg13g2_dfrbp_1 \board_state_next[99]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1469),
    .D(_1631_),
    .Q_N(_4870_),
    .Q(\board_state_next[99] ));
 sg13g2_dfrbp_1 \board_state_next[9]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1470),
    .D(_1632_),
    .Q_N(_4869_),
    .Q(\board_state_next[9] ));
 sg13g2_dfrbp_1 \colindex[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1471),
    .D(_1633_),
    .Q_N(_4868_),
    .Q(\colindex[0] ));
 sg13g2_dfrbp_1 \colindex[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1472),
    .D(_1634_),
    .Q_N(_4867_),
    .Q(\colindex[1] ));
 sg13g2_dfrbp_1 \colindex[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1473),
    .D(_1635_),
    .Q_N(_4866_),
    .Q(\colindex[2] ));
 sg13g2_dfrbp_1 \colindex[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1474),
    .D(_1636_),
    .Q_N(_4865_),
    .Q(\colindex[3] ));
 sg13g2_dfrbp_1 \colindex[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1475),
    .D(_1637_),
    .Q_N(_4864_),
    .Q(\colindex[4] ));
 sg13g2_dfrbp_1 \colindex[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1476),
    .D(_1638_),
    .Q_N(_4863_),
    .Q(\colindex[5] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[0]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1477),
    .D(_1639_),
    .Q_N(_0598_),
    .Q(\hvsync_inst.hpos[0] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[1]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1478),
    .D(_1640_),
    .Q_N(_0072_),
    .Q(\hvsync_inst.hpos[1] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[2]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1479),
    .D(_1641_),
    .Q_N(_4862_),
    .Q(\hvsync_inst.hpos[2] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[3]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1480),
    .D(_1642_),
    .Q_N(_4861_),
    .Q(\hvsync_inst.hpos[3] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[4]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1481),
    .D(_1643_),
    .Q_N(_4860_),
    .Q(\cell_index[0] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[5]$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1482),
    .D(_1644_),
    .Q_N(_4859_),
    .Q(\cell_index[1] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[6]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1483),
    .D(_1645_),
    .Q_N(_4858_),
    .Q(\cell_index[2] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[7]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1484),
    .D(_1646_),
    .Q_N(_0071_),
    .Q(\cell_index[3] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[8]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1485),
    .D(_1647_),
    .Q_N(_4857_),
    .Q(\cell_index[4] ));
 sg13g2_dfrbp_1 \hvsync_inst.hpos[9]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1486),
    .D(_1648_),
    .Q_N(_5406_),
    .Q(\hvsync_inst.hpos[9] ));
 sg13g2_dfrbp_1 \hvsync_inst.hsync$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1487),
    .D(_0044_),
    .Q_N(_4856_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[0]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1488),
    .D(_1649_),
    .Q_N(_0597_),
    .Q(\hvsync_inst.vpos[0] ));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[1]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1489),
    .D(_1650_),
    .Q_N(_4855_),
    .Q(\hvsync_inst.vpos[1] ));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[2]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1490),
    .D(_1651_),
    .Q_N(_0069_),
    .Q(\hvsync_inst.vpos[2] ));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[3]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1491),
    .D(_1652_),
    .Q_N(_0070_),
    .Q(\hvsync_inst.vpos[3] ));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[4]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1492),
    .D(_1653_),
    .Q_N(_4854_),
    .Q(\cell_index[5] ));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[5]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1493),
    .D(_1654_),
    .Q_N(_4853_),
    .Q(\cell_index[6] ));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[6]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1494),
    .D(_1655_),
    .Q_N(_4852_),
    .Q(\cell_index[7] ));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[7]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1495),
    .D(_1656_),
    .Q_N(_4851_),
    .Q(\cell_index[8] ));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[8]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1496),
    .D(_1657_),
    .Q_N(_4850_),
    .Q(\hvsync_inst.vpos[8] ));
 sg13g2_dfrbp_1 \hvsync_inst.vpos[9]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1497),
    .D(_1658_),
    .Q_N(_5407_),
    .Q(\hvsync_inst.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_inst.vsync$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1498),
    .D(_0045_),
    .Q_N(_0064_),
    .Q(\hvsync_inst.vsync ));
 sg13g2_dfrbp_1 \index[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1499),
    .D(_0600_),
    .Q_N(_0054_),
    .Q(\cell_x[0] ));
 sg13g2_dfrbp_1 \index[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1500),
    .D(_0601_),
    .Q_N(_0084_),
    .Q(\cell_x[1] ));
 sg13g2_dfrbp_1 \index[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1501),
    .D(_0602_),
    .Q_N(_0073_),
    .Q(\cell_x[2] ));
 sg13g2_dfrbp_1 \index[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1502),
    .D(_0603_),
    .Q_N(_0074_),
    .Q(\cell_x[3] ));
 sg13g2_dfrbp_1 \index[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1503),
    .D(_0604_),
    .Q_N(_0075_),
    .Q(\cell_x[4] ));
 sg13g2_dfrbp_1 \index[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1504),
    .D(_0605_),
    .Q_N(_0076_),
    .Q(\cell_y[0] ));
 sg13g2_dfrbp_1 \index[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1505),
    .D(_0606_),
    .Q_N(_0077_),
    .Q(\cell_y[1] ));
 sg13g2_dfrbp_1 \index[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1506),
    .D(_0607_),
    .Q_N(_0078_),
    .Q(\cell_y[2] ));
 sg13g2_dfrbp_1 \index[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1507),
    .D(_0608_),
    .Q_N(_0065_),
    .Q(\cell_y[3] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[0]$_SDFF_PN1_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1508),
    .D(_1659_),
    .Q_N(_4849_),
    .Q(\lfsr.lfsr_reg[0] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[10]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1509),
    .D(_1660_),
    .Q_N(_4848_),
    .Q(\lfsr.lfsr_reg[10] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[11]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1510),
    .D(_1661_),
    .Q_N(_4847_),
    .Q(\lfsr.lfsr_reg[11] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[12]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1511),
    .D(_1662_),
    .Q_N(_4846_),
    .Q(\lfsr.lfsr_reg[12] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[13]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1512),
    .D(_1663_),
    .Q_N(_4845_),
    .Q(\lfsr.lfsr_reg[13] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[14]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1513),
    .D(_1664_),
    .Q_N(_4844_),
    .Q(\lfsr.lfsr_reg[14] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[15]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1514),
    .D(_1665_),
    .Q_N(_4843_),
    .Q(\lfsr.lfsr_reg[15] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[1]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1515),
    .D(_1666_),
    .Q_N(_4842_),
    .Q(\lfsr.lfsr_reg[1] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[2]$_SDFF_PN0_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1516),
    .D(_1667_),
    .Q_N(_4841_),
    .Q(\lfsr.lfsr_reg[2] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[3]$_SDFF_PN0_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1517),
    .D(_1668_),
    .Q_N(_4840_),
    .Q(\lfsr.lfsr_reg[3] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[4]$_SDFF_PN0_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1518),
    .D(_1669_),
    .Q_N(_4839_),
    .Q(\lfsr.lfsr_reg[4] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[5]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1519),
    .D(_1670_),
    .Q_N(_4838_),
    .Q(\lfsr.lfsr_reg[5] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[6]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1520),
    .D(_1671_),
    .Q_N(_4837_),
    .Q(\lfsr.lfsr_reg[6] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[7]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1521),
    .D(_1672_),
    .Q_N(_4836_),
    .Q(\lfsr.lfsr_reg[7] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[8]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1522),
    .D(_1673_),
    .Q_N(_4835_),
    .Q(\lfsr.lfsr_reg[8] ));
 sg13g2_dfrbp_1 \lfsr.lfsr_reg[9]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1523),
    .D(_1674_),
    .Q_N(_4834_),
    .Q(\lfsr.lfsr_reg[9] ));
 sg13g2_dfrbp_1 \neigh_index[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1524),
    .D(_1675_),
    .Q_N(_4833_),
    .Q(\neigh_index[0] ));
 sg13g2_dfrbp_1 \neigh_index[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1525),
    .D(_1676_),
    .Q_N(_4832_),
    .Q(\neigh_index[1] ));
 sg13g2_dfrbp_1 \neigh_index[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1526),
    .D(_1677_),
    .Q_N(_4831_),
    .Q(\neigh_index[2] ));
 sg13g2_dfrbp_1 \neigh_index[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1527),
    .D(_1678_),
    .Q_N(_4830_),
    .Q(\neigh_index[3] ));
 sg13g2_dfrbp_1 \num_neighbors[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1528),
    .D(_1679_),
    .Q_N(_4829_),
    .Q(\num_neighbors[0] ));
 sg13g2_dfrbp_1 \num_neighbors[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1529),
    .D(_1680_),
    .Q_N(_4828_),
    .Q(\num_neighbors[1] ));
 sg13g2_dfrbp_1 \num_neighbors[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1530),
    .D(_1681_),
    .Q_N(_4827_),
    .Q(\num_neighbors[2] ));
 sg13g2_dfrbp_1 \num_neighbors[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1531),
    .D(_1682_),
    .Q_N(_4826_),
    .Q(\num_neighbors[3] ));
 sg13g2_dfrbp_1 \running$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1532),
    .D(_1683_),
    .Q_N(_0062_),
    .Q(running));
 sg13g2_dfrbp_1 \timer[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1533),
    .D(_1684_),
    .Q_N(_4825_),
    .Q(\timer[0] ));
 sg13g2_dfrbp_1 \timer[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1534),
    .D(_1685_),
    .Q_N(_4824_),
    .Q(\timer[10] ));
 sg13g2_dfrbp_1 \timer[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1535),
    .D(_1686_),
    .Q_N(_4823_),
    .Q(\timer[11] ));
 sg13g2_dfrbp_1 \timer[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1536),
    .D(_1687_),
    .Q_N(_4822_),
    .Q(\timer[12] ));
 sg13g2_dfrbp_1 \timer[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1537),
    .D(_1688_),
    .Q_N(_4821_),
    .Q(\timer[13] ));
 sg13g2_dfrbp_1 \timer[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1538),
    .D(_1689_),
    .Q_N(_4820_),
    .Q(\timer[14] ));
 sg13g2_dfrbp_1 \timer[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1539),
    .D(_1690_),
    .Q_N(_4819_),
    .Q(\timer[15] ));
 sg13g2_dfrbp_1 \timer[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1540),
    .D(_1691_),
    .Q_N(_4818_),
    .Q(\timer[16] ));
 sg13g2_dfrbp_1 \timer[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1541),
    .D(_1692_),
    .Q_N(_4817_),
    .Q(\timer[17] ));
 sg13g2_dfrbp_1 \timer[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1542),
    .D(_1693_),
    .Q_N(_4816_),
    .Q(\timer[18] ));
 sg13g2_dfrbp_1 \timer[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1543),
    .D(_1694_),
    .Q_N(_4815_),
    .Q(\timer[19] ));
 sg13g2_dfrbp_1 \timer[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1544),
    .D(_1695_),
    .Q_N(_4814_),
    .Q(\timer[1] ));
 sg13g2_dfrbp_1 \timer[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1545),
    .D(_1696_),
    .Q_N(_4813_),
    .Q(\timer[20] ));
 sg13g2_dfrbp_1 \timer[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1546),
    .D(_1697_),
    .Q_N(_4812_),
    .Q(\timer[21] ));
 sg13g2_dfrbp_1 \timer[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1547),
    .D(_1698_),
    .Q_N(_4811_),
    .Q(\timer[22] ));
 sg13g2_dfrbp_1 \timer[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1548),
    .D(_1699_),
    .Q_N(_4810_),
    .Q(\timer[23] ));
 sg13g2_dfrbp_1 \timer[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1549),
    .D(_1700_),
    .Q_N(_4809_),
    .Q(\timer[24] ));
 sg13g2_dfrbp_1 \timer[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1550),
    .D(_1701_),
    .Q_N(_4808_),
    .Q(\timer[25] ));
 sg13g2_dfrbp_1 \timer[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1551),
    .D(_1702_),
    .Q_N(_4807_),
    .Q(\timer[26] ));
 sg13g2_dfrbp_1 \timer[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1552),
    .D(_1703_),
    .Q_N(_4806_),
    .Q(\timer[27] ));
 sg13g2_dfrbp_1 \timer[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1553),
    .D(_1704_),
    .Q_N(_4805_),
    .Q(\timer[28] ));
 sg13g2_dfrbp_1 \timer[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1554),
    .D(_1705_),
    .Q_N(_4804_),
    .Q(\timer[29] ));
 sg13g2_dfrbp_1 \timer[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1555),
    .D(_1706_),
    .Q_N(_4803_),
    .Q(\timer[2] ));
 sg13g2_dfrbp_1 \timer[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1556),
    .D(_1707_),
    .Q_N(_4802_),
    .Q(\timer[30] ));
 sg13g2_dfrbp_1 \timer[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1557),
    .D(_1708_),
    .Q_N(_4801_),
    .Q(\timer[31] ));
 sg13g2_dfrbp_1 \timer[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1558),
    .D(_1709_),
    .Q_N(_4800_),
    .Q(\timer[3] ));
 sg13g2_dfrbp_1 \timer[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1559),
    .D(_1710_),
    .Q_N(_4799_),
    .Q(\timer[4] ));
 sg13g2_dfrbp_1 \timer[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1560),
    .D(_1711_),
    .Q_N(_4798_),
    .Q(\timer[5] ));
 sg13g2_dfrbp_1 \timer[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1561),
    .D(_1712_),
    .Q_N(_4797_),
    .Q(\timer[6] ));
 sg13g2_dfrbp_1 \timer[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1562),
    .D(_1713_),
    .Q_N(_4796_),
    .Q(\timer[7] ));
 sg13g2_dfrbp_1 \timer[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1563),
    .D(_1714_),
    .Q_N(_4795_),
    .Q(\timer[8] ));
 sg13g2_dfrbp_1 \timer[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1564),
    .D(_1715_),
    .Q_N(_0060_),
    .Q(\timer[9] ));
 sg13g2_dfrbp_1 \txindex[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1565),
    .D(_1716_),
    .Q_N(_0080_),
    .Q(\txindex[0] ));
 sg13g2_dfrbp_1 \txindex[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1566),
    .D(_1717_),
    .Q_N(_0056_),
    .Q(\txindex[1] ));
 sg13g2_dfrbp_1 \txindex[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1567),
    .D(_1718_),
    .Q_N(_0081_),
    .Q(\txindex[2] ));
 sg13g2_dfrbp_1 \txindex[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1568),
    .D(net168),
    .Q_N(_4794_),
    .Q(\txindex[3] ));
 sg13g2_dfrbp_1 \txindex[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1569),
    .D(_1720_),
    .Q_N(_4793_),
    .Q(\txindex[4] ));
 sg13g2_dfrbp_1 \txindex[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1570),
    .D(_1721_),
    .Q_N(_5408_),
    .Q(\txindex[5] ));
 sg13g2_dfrbp_1 \txstate[0]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1571),
    .D(_0028_),
    .Q_N(_0061_),
    .Q(\txstate[0] ));
 sg13g2_dfrbp_1 \txstate[2]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1572),
    .D(_0029_),
    .Q_N(_5409_),
    .Q(\txstate[2] ));
 sg13g2_dfrbp_1 \txstate[3]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1573),
    .D(_0030_),
    .Q_N(_5410_),
    .Q(\txstate[3] ));
 sg13g2_dfrbp_1 \txstate[4]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1574),
    .D(_0031_),
    .Q_N(_0063_),
    .Q(\txstate[4] ));
 sg13g2_dfrbp_1 \txstate[5]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1575),
    .D(_0032_),
    .Q_N(_5411_),
    .Q(\txstate[5] ));
 sg13g2_dfrbp_1 \txstate[6]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1576),
    .D(_0033_),
    .Q_N(_5412_),
    .Q(\txstate[6] ));
 sg13g2_dfrbp_1 \txstate[7]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1577),
    .D(_0034_),
    .Q_N(_0079_),
    .Q(\txstate[7] ));
 sg13g2_dfrbp_1 \txstate[8]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1578),
    .D(_0035_),
    .Q_N(_0066_),
    .Q(\txstate[8] ));
 sg13g2_dfrbp_1 \uart_rx_inst.bitIndex[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1579),
    .D(_1722_),
    .Q_N(_0595_),
    .Q(\uart_rx_inst.bitIndex[0] ));
 sg13g2_dfrbp_1 \uart_rx_inst.bitIndex[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1580),
    .D(_1723_),
    .Q_N(_4792_),
    .Q(\uart_rx_inst.bitIndex[1] ));
 sg13g2_dfrbp_1 \uart_rx_inst.bitIndex[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1581),
    .D(_1724_),
    .Q_N(_0059_),
    .Q(\uart_rx_inst.bitIndex[2] ));
 sg13g2_dfrbp_1 \uart_rx_inst.data[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1582),
    .D(_1725_),
    .Q_N(_4791_),
    .Q(\uart_rx_inst.data[0] ));
 sg13g2_dfrbp_1 \uart_rx_inst.data[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1583),
    .D(_1726_),
    .Q_N(_4790_),
    .Q(\uart_rx_inst.data[1] ));
 sg13g2_dfrbp_1 \uart_rx_inst.data[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1584),
    .D(_1727_),
    .Q_N(_4789_),
    .Q(\uart_rx_inst.data[2] ));
 sg13g2_dfrbp_1 \uart_rx_inst.data[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1585),
    .D(_1728_),
    .Q_N(_4788_),
    .Q(\uart_rx_inst.data[3] ));
 sg13g2_dfrbp_1 \uart_rx_inst.data[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1586),
    .D(_1729_),
    .Q_N(_4787_),
    .Q(\uart_rx_inst.data[4] ));
 sg13g2_dfrbp_1 \uart_rx_inst.data[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1587),
    .D(_1730_),
    .Q_N(_4786_),
    .Q(\uart_rx_inst.data[5] ));
 sg13g2_dfrbp_1 \uart_rx_inst.data[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1588),
    .D(_1731_),
    .Q_N(_4785_),
    .Q(\uart_rx_inst.data[6] ));
 sg13g2_dfrbp_1 \uart_rx_inst.data[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1589),
    .D(_1732_),
    .Q_N(_4784_),
    .Q(\uart_rx_inst.data[7] ));
 sg13g2_dfrbp_1 \uart_rx_inst.inputReg[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1590),
    .D(_1733_),
    .Q_N(_4783_),
    .Q(\uart_rx_inst.inputReg[0] ));
 sg13g2_dfrbp_1 \uart_rx_inst.inputReg[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1591),
    .D(_1734_),
    .Q_N(_4782_),
    .Q(\uart_rx_inst.inputReg[1] ));
 sg13g2_dfrbp_1 \uart_rx_inst.inputReg[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1592),
    .D(_1735_),
    .Q_N(_4781_),
    .Q(\uart_rx_inst.inputReg[2] ));
 sg13g2_dfrbp_1 \uart_rx_inst.out[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1593),
    .D(_1736_),
    .Q_N(_4780_),
    .Q(\uart_rx_data[0] ));
 sg13g2_dfrbp_1 \uart_rx_inst.out[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1594),
    .D(_1737_),
    .Q_N(_4779_),
    .Q(\uart_rx_data[1] ));
 sg13g2_dfrbp_1 \uart_rx_inst.out[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1595),
    .D(_1738_),
    .Q_N(_4778_),
    .Q(\uart_rx_data[2] ));
 sg13g2_dfrbp_1 \uart_rx_inst.out[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1596),
    .D(_1739_),
    .Q_N(_4777_),
    .Q(\uart_rx_data[3] ));
 sg13g2_dfrbp_1 \uart_rx_inst.out[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1597),
    .D(_1740_),
    .Q_N(_4776_),
    .Q(\uart_rx_data[4] ));
 sg13g2_dfrbp_1 \uart_rx_inst.out[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1598),
    .D(_1741_),
    .Q_N(_4775_),
    .Q(\uart_rx_data[5] ));
 sg13g2_dfrbp_1 \uart_rx_inst.out[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1599),
    .D(_1742_),
    .Q_N(_4774_),
    .Q(\uart_rx_data[6] ));
 sg13g2_dfrbp_1 \uart_rx_inst.out[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1600),
    .D(_1743_),
    .Q_N(_4773_),
    .Q(\uart_rx_data[7] ));
 sg13g2_dfrbp_1 \uart_rx_inst.out_latched$_SDFFE_PP0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1601),
    .D(_1744_),
    .Q_N(_4772_),
    .Q(\uart_rx_inst.out_latched ));
 sg13g2_dfrbp_1 \uart_rx_inst.rxCounter[0]$_SDFF_PN0_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1602),
    .D(_1745_),
    .Q_N(_0599_),
    .Q(\uart_rx_inst.rxCounter[0] ));
 sg13g2_dfrbp_1 \uart_rx_inst.rxCounter[1]$_SDFF_PN0_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1603),
    .D(_1746_),
    .Q_N(_4771_),
    .Q(\uart_rx_inst.rxCounter[1] ));
 sg13g2_dfrbp_1 \uart_rx_inst.rxCounter[2]$_SDFF_PN0_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1604),
    .D(_1747_),
    .Q_N(_4770_),
    .Q(\uart_rx_inst.rxCounter[2] ));
 sg13g2_dfrbp_1 \uart_rx_inst.rxCounter[3]$_SDFF_PN0_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1605),
    .D(_1748_),
    .Q_N(_4769_),
    .Q(\uart_rx_inst.rxCounter[3] ));
 sg13g2_dfrbp_1 \uart_rx_inst.sampleCount[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1606),
    .D(_1749_),
    .Q_N(_4768_),
    .Q(\uart_rx_inst.sampleCount[0] ));
 sg13g2_dfrbp_1 \uart_rx_inst.sampleCount[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1607),
    .D(_1750_),
    .Q_N(_4767_),
    .Q(\uart_rx_inst.sampleCount[1] ));
 sg13g2_dfrbp_1 \uart_rx_inst.sampleCount[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1608),
    .D(_1751_),
    .Q_N(_4766_),
    .Q(\uart_rx_inst.sampleCount[2] ));
 sg13g2_dfrbp_1 \uart_rx_inst.sampleCount[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1609),
    .D(_1752_),
    .Q_N(_5413_),
    .Q(\uart_rx_inst.sampleCount[3] ));
 sg13g2_dfrbp_1 \uart_rx_inst.state[0]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1610),
    .D(_0036_),
    .Q_N(_5414_),
    .Q(\uart_rx_inst.state[0] ));
 sg13g2_dfrbp_1 \uart_rx_inst.state[1]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1611),
    .D(_0037_),
    .Q_N(_5415_),
    .Q(\uart_rx_inst.state[1] ));
 sg13g2_dfrbp_1 \uart_rx_inst.state[2]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1612),
    .D(_0038_),
    .Q_N(_0067_),
    .Q(\uart_rx_inst.state[2] ));
 sg13g2_dfrbp_1 \uart_rx_inst.state[3]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1613),
    .D(_0039_),
    .Q_N(_0068_),
    .Q(\uart_rx_inst.state[3] ));
 sg13g2_dfrbp_1 \uart_rx_inst.valid$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1614),
    .D(_1753_),
    .Q_N(_4765_),
    .Q(\uart_rx_inst.valid ));
 sg13g2_dfrbp_1 \uart_rx_ready$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1615),
    .D(_1754_),
    .Q_N(_4764_),
    .Q(\uart_rx_inst.ready ));
 sg13g2_dfrbp_1 \uart_tx_data[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1616),
    .D(_1755_),
    .Q_N(_4763_),
    .Q(\uart_tx_data[0] ));
 sg13g2_dfrbp_1 \uart_tx_data[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1617),
    .D(_1756_),
    .Q_N(_4762_),
    .Q(\uart_tx_data[1] ));
 sg13g2_dfrbp_1 \uart_tx_data[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1618),
    .D(_1757_),
    .Q_N(_4761_),
    .Q(\uart_tx_data[2] ));
 sg13g2_dfrbp_1 \uart_tx_data[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1619),
    .D(_1758_),
    .Q_N(_4760_),
    .Q(\uart_tx_data[3] ));
 sg13g2_dfrbp_1 \uart_tx_data[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1620),
    .D(_1759_),
    .Q_N(_4759_),
    .Q(\uart_tx_data[4] ));
 sg13g2_dfrbp_1 \uart_tx_data[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1621),
    .D(_1760_),
    .Q_N(_4758_),
    .Q(\uart_tx_data[5] ));
 sg13g2_dfrbp_1 \uart_tx_data[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1622),
    .D(_1761_),
    .Q_N(_4757_),
    .Q(\uart_tx_data[6] ));
 sg13g2_dfrbp_1 \uart_tx_inst.bitIndex[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1623),
    .D(_1762_),
    .Q_N(_4756_),
    .Q(\uart_tx_inst.bitIndex[0] ));
 sg13g2_dfrbp_1 \uart_tx_inst.bitIndex[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1624),
    .D(_1763_),
    .Q_N(_4755_),
    .Q(\uart_tx_inst.bitIndex[1] ));
 sg13g2_dfrbp_1 \uart_tx_inst.bitIndex[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1625),
    .D(_1764_),
    .Q_N(_0057_),
    .Q(\uart_tx_inst.bitIndex[2] ));
 sg13g2_dfrbp_1 \uart_tx_inst.data[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1626),
    .D(_1765_),
    .Q_N(_4754_),
    .Q(\uart_tx_inst.data[0] ));
 sg13g2_dfrbp_1 \uart_tx_inst.data[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1627),
    .D(_1766_),
    .Q_N(_4753_),
    .Q(\uart_tx_inst.data[1] ));
 sg13g2_dfrbp_1 \uart_tx_inst.data[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1628),
    .D(_1767_),
    .Q_N(_4752_),
    .Q(\uart_tx_inst.data[2] ));
 sg13g2_dfrbp_1 \uart_tx_inst.data[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1629),
    .D(_1768_),
    .Q_N(_4751_),
    .Q(\uart_tx_inst.data[3] ));
 sg13g2_dfrbp_1 \uart_tx_inst.data[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1630),
    .D(_1769_),
    .Q_N(_4750_),
    .Q(\uart_tx_inst.data[4] ));
 sg13g2_dfrbp_1 \uart_tx_inst.data[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1631),
    .D(_1770_),
    .Q_N(_4749_),
    .Q(\uart_tx_inst.data[5] ));
 sg13g2_dfrbp_1 \uart_tx_inst.data[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1632),
    .D(_1771_),
    .Q_N(_4748_),
    .Q(\uart_tx_inst.data[6] ));
 sg13g2_dfrbp_1 \uart_tx_inst.out$_SDFFE_PN1P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1633),
    .D(_1772_),
    .Q_N(_4747_),
    .Q(uart_tx));
 sg13g2_dfrbp_1 \uart_tx_inst.ready$_SDFFE_PP0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1634),
    .D(_1773_),
    .Q_N(_5416_),
    .Q(\uart_tx_inst.ready ));
 sg13g2_dfrbp_1 \uart_tx_inst.state[0]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1635),
    .D(_0040_),
    .Q_N(_5417_),
    .Q(\uart_tx_inst.state[0] ));
 sg13g2_dfrbp_1 \uart_tx_inst.state[1]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1636),
    .D(_0041_),
    .Q_N(_0596_),
    .Q(\uart_tx_inst.state[1] ));
 sg13g2_dfrbp_1 \uart_tx_inst.state[2]$_DFF_P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1637),
    .D(_0042_),
    .Q_N(_5418_),
    .Q(\uart_tx_inst.state[2] ));
 sg13g2_dfrbp_1 \uart_tx_inst.state[3]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1638),
    .D(_0043_),
    .Q_N(_4746_),
    .Q(\uart_tx_inst.state[3] ));
 sg13g2_dfrbp_1 \uart_tx_inst.txCounter[0]$_SDFFE_PN0N_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1639),
    .D(_1774_),
    .Q_N(_4745_),
    .Q(\uart_tx_inst.txCounter[0] ));
 sg13g2_dfrbp_1 \uart_tx_inst.txCounter[1]$_SDFFE_PN0N_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1640),
    .D(_1775_),
    .Q_N(_4744_),
    .Q(\uart_tx_inst.txCounter[1] ));
 sg13g2_dfrbp_1 \uart_tx_inst.txCounter[2]$_SDFFE_PN0N_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1641),
    .D(_1776_),
    .Q_N(_4743_),
    .Q(\uart_tx_inst.txCounter[2] ));
 sg13g2_dfrbp_1 \uart_tx_inst.txCounter[3]$_SDFFE_PN0N_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1642),
    .D(_1777_),
    .Q_N(_4742_),
    .Q(\uart_tx_inst.txCounter[3] ));
 sg13g2_dfrbp_1 \uart_tx_inst.txCounter[4]$_SDFFE_PN0N_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1643),
    .D(_1778_),
    .Q_N(_4741_),
    .Q(\uart_tx_inst.txCounter[4] ));
 sg13g2_dfrbp_1 \uart_tx_inst.txCounter[5]$_SDFFE_PN0N_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1644),
    .D(_1779_),
    .Q_N(_4740_),
    .Q(\uart_tx_inst.txCounter[5] ));
 sg13g2_dfrbp_1 \uart_tx_inst.txCounter[6]$_SDFFE_PN0N_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1645),
    .D(_1780_),
    .Q_N(_4739_),
    .Q(\uart_tx_inst.txCounter[6] ));
 sg13g2_dfrbp_1 \uart_tx_inst.txCounter[7]$_SDFFE_PN0N_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1646),
    .D(_1781_),
    .Q_N(_4738_),
    .Q(\uart_tx_inst.txCounter[7] ));
 sg13g2_dfrbp_1 \uart_tx_valid$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1647),
    .D(_1782_),
    .Q_N(_4737_),
    .Q(\uart_tx_inst.valid ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[0]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[1]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[3]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[4]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[5]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[4]));
 sg13g2_buf_2 fanout12 (.A(_3242_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_3231_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_3220_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_3209_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_3192_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_3178_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_3167_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_3153_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_3142_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_3127_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_3115_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_3101_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_3086_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_3068_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_3053_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_3040_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_3024_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_3011_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_2996_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_2982_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_2970_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_2956_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_2942_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_2927_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_2916_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_2902_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_2891_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_2877_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_2862_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_2846_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_2830_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_2814_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_2799_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_2786_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_2771_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_2757_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2746_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_2731_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_2720_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_2706_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_2691_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2677_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2666_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2652_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_2635_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2600_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2549_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_2535_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_3281_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_3267_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_3256_),
    .X(net62));
 sg13g2_buf_1 fanout63 (.A(_3126_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_2981_),
    .X(net64));
 sg13g2_buf_1 fanout65 (.A(_2845_),
    .X(net65));
 sg13g2_buf_1 fanout66 (.A(_2705_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_2534_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_4194_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_3844_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_3829_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_3795_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_3743_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_4226_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_4193_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_3791_),
    .X(net75));
 sg13g2_buf_4 fanout76 (.X(net76),
    .A(_3545_));
 sg13g2_buf_4 fanout77 (.X(net77),
    .A(_3544_));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(_3543_));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(_3542_));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_3541_));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(_3540_));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_3539_));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_3537_));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(_3536_));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_3535_));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(_3534_));
 sg13g2_buf_4 fanout87 (.X(net87),
    .A(_3533_));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(_3532_));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(_3531_));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(_3529_));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(_3528_));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(_3527_));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(_3526_));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(_3525_));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(_3524_));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(_3523_));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(_3521_));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(_3520_));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(_3519_));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(_3518_));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(_3517_));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(_3516_));
 sg13g2_buf_2 fanout103 (.A(_2210_),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(_3959_));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(_3942_));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_3896_));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(_3839_));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(_3837_));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(_3834_));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_3802_));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(_3790_));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(_3769_));
 sg13g2_buf_8 fanout113 (.A(_3758_),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(_3572_));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(_3571_));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_3570_));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(_3569_));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(_3568_));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(_3567_));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(_3566_));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(_3565_));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(_3564_));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(_3563_));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(_3561_));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(_3560_));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_3559_));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_3558_));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(_3557_));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(_3556_));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_3555_));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(_3553_));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(_3552_));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(_3551_));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(_3550_));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(_3549_));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(_3548_));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(_3547_));
 sg13g2_buf_2 fanout138 (.A(_3087_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_3082_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_3078_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_3076_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_3073_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_3071_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_3056_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_3044_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_3041_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_3038_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_2863_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_2857_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_2853_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_2851_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_2841_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_2825_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_2821_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_2819_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_2817_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_2815_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_2638_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_2629_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_2619_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_2615_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_2611_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_2607_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_2603_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_2598_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_2594_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_2571_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_1719_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_2247_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_2228_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_2221_),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(_4055_),
    .X(net172));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(_3989_));
 sg13g2_buf_8 fanout174 (.A(_3972_),
    .X(net174));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(_3950_));
 sg13g2_buf_8 fanout176 (.A(_3906_),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(_3870_),
    .X(net177));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(_3862_));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(_3859_));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(_3847_));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(_3836_));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(_3833_));
 sg13g2_buf_8 fanout183 (.A(_3831_),
    .X(net183));
 sg13g2_buf_8 fanout184 (.A(_3800_),
    .X(net184));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(_3798_));
 sg13g2_buf_8 fanout186 (.A(_3796_),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(_3768_));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(_3757_));
 sg13g2_buf_2 fanout189 (.A(_3084_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_3080_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_3030_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_3014_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_3012_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_3008_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_2860_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_2855_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_2806_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_2789_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_2787_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_2784_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_2633_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_2625_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_2590_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_2586_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_2582_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_2556_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_2547_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_2263_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_2231_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_2226_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_2220_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_2209_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_2140_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_4430_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_4351_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_4186_),
    .X(net216));
 sg13g2_buf_8 fanout217 (.A(_3939_),
    .X(net217));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(_3905_));
 sg13g2_buf_2 fanout219 (.A(_3832_),
    .X(net219));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(_3830_));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(_3797_));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(_3767_));
 sg13g2_buf_2 fanout223 (.A(_3613_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_3270_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_3207_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_3197_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_3160_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_3113_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_3061_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_3006_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_2961_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_2912_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_2867_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_2809_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_2760_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_2713_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_2701_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_2664_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_2578_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_2192_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_2950_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_2782_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_2737_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_2687_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_2642_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_2568_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_2540_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_3247_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_3183_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_3137_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_3091_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_3033_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_2985_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_2936_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_2888_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_2836_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_2421_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_2412_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_2374_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_2340_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_1861_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_1855_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_4329_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_4181_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_3632_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_2387_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_2364_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_2357_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_2346_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_2336_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_2072_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_2038_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_2025_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_1889_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_1869_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_1817_),
    .X(net276));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(_4651_));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(_4639_));
 sg13g2_buf_8 fanout279 (.A(_4637_),
    .X(net279));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(_4631_));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(_4602_));
 sg13g2_buf_8 fanout282 (.A(_4577_),
    .X(net282));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_4571_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_4564_));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_4554_));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(_4544_));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_4542_));
 sg13g2_buf_8 fanout288 (.A(_4535_),
    .X(net288));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(_4533_));
 sg13g2_buf_8 fanout290 (.A(_4528_),
    .X(net290));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(_4526_));
 sg13g2_buf_8 fanout292 (.A(_4525_),
    .X(net292));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(_4522_));
 sg13g2_buf_8 fanout294 (.A(_4521_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_3687_),
    .X(net295));
 sg13g2_buf_1 fanout296 (.A(_3677_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_3599_),
    .X(net297));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(_3423_));
 sg13g2_buf_8 fanout299 (.A(_3422_),
    .X(net299));
 sg13g2_buf_8 fanout300 (.A(_3420_),
    .X(net300));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(_3415_));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(_3361_));
 sg13g2_buf_8 fanout303 (.A(_3360_),
    .X(net303));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(_3349_));
 sg13g2_buf_8 fanout305 (.A(_3348_),
    .X(net305));
 sg13g2_buf_4 fanout306 (.X(net306),
    .A(_3334_));
 sg13g2_buf_8 fanout307 (.A(_3333_),
    .X(net307));
 sg13g2_buf_4 fanout308 (.X(net308),
    .A(_3324_));
 sg13g2_buf_8 fanout309 (.A(_3323_),
    .X(net309));
 sg13g2_buf_4 fanout310 (.X(net310),
    .A(_3318_));
 sg13g2_buf_8 fanout311 (.A(_3317_),
    .X(net311));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(_3306_));
 sg13g2_buf_8 fanout313 (.A(_3304_),
    .X(net313));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(_3300_));
 sg13g2_buf_8 fanout315 (.A(_3297_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_2462_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_2403_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_2371_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_2349_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_2341_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_2338_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_2325_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_2109_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_2106_),
    .X(net324));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_2103_));
 sg13g2_buf_2 fanout326 (.A(_2031_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_2016_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_1994_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_1913_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_1832_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_1816_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_1813_),
    .X(net332));
 sg13g2_buf_8 fanout333 (.A(_4668_),
    .X(net333));
 sg13g2_buf_8 fanout334 (.A(_4645_),
    .X(net334));
 sg13g2_buf_8 fanout335 (.A(_4604_),
    .X(net335));
 sg13g2_buf_8 fanout336 (.A(_4596_),
    .X(net336));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(_4594_));
 sg13g2_buf_8 fanout338 (.A(_4593_),
    .X(net338));
 sg13g2_buf_8 fanout339 (.A(_4552_),
    .X(net339));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(_4547_));
 sg13g2_buf_8 fanout341 (.A(_4546_),
    .X(net341));
 sg13g2_buf_8 fanout342 (.A(_4540_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_3686_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_3682_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_3678_),
    .X(net345));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(_3669_));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_3575_));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(_3437_));
 sg13g2_buf_8 fanout349 (.A(_3436_),
    .X(net349));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(_3430_));
 sg13g2_buf_8 fanout351 (.A(_3429_),
    .X(net351));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(_3382_));
 sg13g2_buf_8 fanout353 (.A(_3381_),
    .X(net353));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(_3378_));
 sg13g2_buf_8 fanout355 (.A(_3377_),
    .X(net355));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(_3328_));
 sg13g2_buf_8 fanout357 (.A(_3327_),
    .X(net357));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(_3312_));
 sg13g2_buf_8 fanout359 (.A(_3310_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_3299_),
    .X(net360));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(_3296_));
 sg13g2_buf_2 fanout362 (.A(_2481_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_2402_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_2367_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_2345_),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(_2113_));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(_2108_));
 sg13g2_buf_2 fanout368 (.A(_2105_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_2028_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_2015_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_2013_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_1912_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_1871_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_1831_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_1824_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_1822_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_1815_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_1812_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_1809_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_1798_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_1795_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_1790_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_4297_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_2378_),
    .X(net384));
 sg13g2_buf_4 fanout385 (.X(net385),
    .A(_2112_));
 sg13g2_buf_2 fanout386 (.A(_2018_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_2011_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_1914_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_1875_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_1863_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_1835_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_1834_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_1823_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_1819_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_1807_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_1806_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_1800_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_1799_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_1796_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_1786_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_1793_),
    .X(net401));
 sg13g2_tielo _9616__402 (.L_LO(net402));
 sg13g2_tielo _9617__403 (.L_LO(net403));
 sg13g2_tielo _9618__404 (.L_LO(net404));
 sg13g2_tielo _9619__405 (.L_LO(net405));
 sg13g2_tielo _9620__406 (.L_LO(net406));
 sg13g2_tielo _9621__407 (.L_LO(net407));
 sg13g2_tielo _9622__408 (.L_LO(net408));
 sg13g2_tielo _9624__409 (.L_LO(net409));
 sg13g2_tielo _9629__410 (.L_LO(net410));
 sg13g2_tielo _9630__411 (.L_LO(net411));
 sg13g2_tielo _9631__412 (.L_LO(net412));
 sg13g2_tielo _9632__413 (.L_LO(net413));
 sg13g2_tielo _9634__414 (.L_LO(net414));
 sg13g2_tielo _9635__415 (.L_LO(net415));
 sg13g2_tielo _9636__416 (.L_LO(net416));
 sg13g2_tiehi _9594__418 (.L_HI(net418));
 sg13g2_tiehi _9595__419 (.L_HI(net419));
 sg13g2_tiehi _9596__420 (.L_HI(net420));
 sg13g2_tiehi _9597__421 (.L_HI(net421));
 sg13g2_tiehi _9598__422 (.L_HI(net422));
 sg13g2_tiehi _9599__423 (.L_HI(net423));
 sg13g2_tiehi _9600__424 (.L_HI(net424));
 sg13g2_tiehi _9601__425 (.L_HI(net425));
 sg13g2_tiehi _9602__426 (.L_HI(net426));
 sg13g2_tiehi _9603__427 (.L_HI(net427));
 sg13g2_tiehi _9604__428 (.L_HI(net428));
 sg13g2_tiehi _9605__429 (.L_HI(net429));
 sg13g2_tiehi _9606__430 (.L_HI(net430));
 sg13g2_tiehi _9607__431 (.L_HI(net431));
 sg13g2_tiehi _9608__432 (.L_HI(net432));
 sg13g2_tiehi _9609__433 (.L_HI(net433));
 sg13g2_tiehi _9610__434 (.L_HI(net434));
 sg13g2_tiehi _9611__435 (.L_HI(net435));
 sg13g2_tiehi _9612__436 (.L_HI(net436));
 sg13g2_tiehi _9615__437 (.L_HI(net437));
 sg13g2_tiehi _9627__438 (.L_HI(net438));
 sg13g2_tiehi \action[0]$_DFF_P__439  (.L_HI(net439));
 sg13g2_tiehi \action[1]$_DFF_P__440  (.L_HI(net440));
 sg13g2_tiehi \action[2]$_DFF_P__441  (.L_HI(net441));
 sg13g2_tiehi \action[3]$_DFF_P__442  (.L_HI(net442));
 sg13g2_tiehi \action[4]$_DFF_P__443  (.L_HI(net443));
 sg13g2_tiehi \action[5]$_DFF_P__444  (.L_HI(net444));
 sg13g2_tiehi \action[6]$_DFF_P__445  (.L_HI(net445));
 sg13g2_tiehi \action[7]$_DFF_P__446  (.L_HI(net446));
 sg13g2_tiehi \board_state[0]$_DFFE_PP__447  (.L_HI(net447));
 sg13g2_tiehi \board_state[100]$_DFFE_PP__448  (.L_HI(net448));
 sg13g2_tiehi \board_state[101]$_DFFE_PP__449  (.L_HI(net449));
 sg13g2_tiehi \board_state[102]$_DFFE_PP__450  (.L_HI(net450));
 sg13g2_tiehi \board_state[103]$_DFFE_PP__451  (.L_HI(net451));
 sg13g2_tiehi \board_state[104]$_DFFE_PP__452  (.L_HI(net452));
 sg13g2_tiehi \board_state[105]$_DFFE_PP__453  (.L_HI(net453));
 sg13g2_tiehi \board_state[106]$_DFFE_PP__454  (.L_HI(net454));
 sg13g2_tiehi \board_state[107]$_DFFE_PP__455  (.L_HI(net455));
 sg13g2_tiehi \board_state[108]$_DFFE_PP__456  (.L_HI(net456));
 sg13g2_tiehi \board_state[109]$_DFFE_PP__457  (.L_HI(net457));
 sg13g2_tiehi \board_state[10]$_DFFE_PP__458  (.L_HI(net458));
 sg13g2_tiehi \board_state[110]$_DFFE_PP__459  (.L_HI(net459));
 sg13g2_tiehi \board_state[111]$_DFFE_PP__460  (.L_HI(net460));
 sg13g2_tiehi \board_state[112]$_DFFE_PP__461  (.L_HI(net461));
 sg13g2_tiehi \board_state[113]$_DFFE_PP__462  (.L_HI(net462));
 sg13g2_tiehi \board_state[114]$_DFFE_PP__463  (.L_HI(net463));
 sg13g2_tiehi \board_state[115]$_DFFE_PP__464  (.L_HI(net464));
 sg13g2_tiehi \board_state[116]$_DFFE_PP__465  (.L_HI(net465));
 sg13g2_tiehi \board_state[117]$_DFFE_PP__466  (.L_HI(net466));
 sg13g2_tiehi \board_state[118]$_DFFE_PP__467  (.L_HI(net467));
 sg13g2_tiehi \board_state[119]$_DFFE_PP__468  (.L_HI(net468));
 sg13g2_tiehi \board_state[11]$_DFFE_PP__469  (.L_HI(net469));
 sg13g2_tiehi \board_state[120]$_DFFE_PP__470  (.L_HI(net470));
 sg13g2_tiehi \board_state[121]$_DFFE_PP__471  (.L_HI(net471));
 sg13g2_tiehi \board_state[122]$_DFFE_PP__472  (.L_HI(net472));
 sg13g2_tiehi \board_state[123]$_DFFE_PP__473  (.L_HI(net473));
 sg13g2_tiehi \board_state[124]$_DFFE_PP__474  (.L_HI(net474));
 sg13g2_tiehi \board_state[125]$_DFFE_PP__475  (.L_HI(net475));
 sg13g2_tiehi \board_state[126]$_DFFE_PP__476  (.L_HI(net476));
 sg13g2_tiehi \board_state[127]$_DFFE_PP__477  (.L_HI(net477));
 sg13g2_tiehi \board_state[128]$_DFFE_PP__478  (.L_HI(net478));
 sg13g2_tiehi \board_state[129]$_DFFE_PP__479  (.L_HI(net479));
 sg13g2_tiehi \board_state[12]$_DFFE_PP__480  (.L_HI(net480));
 sg13g2_tiehi \board_state[130]$_DFFE_PP__481  (.L_HI(net481));
 sg13g2_tiehi \board_state[131]$_DFFE_PP__482  (.L_HI(net482));
 sg13g2_tiehi \board_state[132]$_DFFE_PP__483  (.L_HI(net483));
 sg13g2_tiehi \board_state[133]$_DFFE_PP__484  (.L_HI(net484));
 sg13g2_tiehi \board_state[134]$_DFFE_PP__485  (.L_HI(net485));
 sg13g2_tiehi \board_state[135]$_DFFE_PP__486  (.L_HI(net486));
 sg13g2_tiehi \board_state[136]$_DFFE_PP__487  (.L_HI(net487));
 sg13g2_tiehi \board_state[137]$_DFFE_PP__488  (.L_HI(net488));
 sg13g2_tiehi \board_state[138]$_DFFE_PP__489  (.L_HI(net489));
 sg13g2_tiehi \board_state[139]$_DFFE_PP__490  (.L_HI(net490));
 sg13g2_tiehi \board_state[13]$_DFFE_PP__491  (.L_HI(net491));
 sg13g2_tiehi \board_state[140]$_DFFE_PP__492  (.L_HI(net492));
 sg13g2_tiehi \board_state[141]$_DFFE_PP__493  (.L_HI(net493));
 sg13g2_tiehi \board_state[142]$_DFFE_PP__494  (.L_HI(net494));
 sg13g2_tiehi \board_state[143]$_DFFE_PP__495  (.L_HI(net495));
 sg13g2_tiehi \board_state[144]$_DFFE_PP__496  (.L_HI(net496));
 sg13g2_tiehi \board_state[145]$_DFFE_PP__497  (.L_HI(net497));
 sg13g2_tiehi \board_state[146]$_DFFE_PP__498  (.L_HI(net498));
 sg13g2_tiehi \board_state[147]$_DFFE_PP__499  (.L_HI(net499));
 sg13g2_tiehi \board_state[148]$_DFFE_PP__500  (.L_HI(net500));
 sg13g2_tiehi \board_state[149]$_DFFE_PP__501  (.L_HI(net501));
 sg13g2_tiehi \board_state[14]$_DFFE_PP__502  (.L_HI(net502));
 sg13g2_tiehi \board_state[150]$_DFFE_PP__503  (.L_HI(net503));
 sg13g2_tiehi \board_state[151]$_DFFE_PP__504  (.L_HI(net504));
 sg13g2_tiehi \board_state[152]$_DFFE_PP__505  (.L_HI(net505));
 sg13g2_tiehi \board_state[153]$_DFFE_PP__506  (.L_HI(net506));
 sg13g2_tiehi \board_state[154]$_DFFE_PP__507  (.L_HI(net507));
 sg13g2_tiehi \board_state[155]$_DFFE_PP__508  (.L_HI(net508));
 sg13g2_tiehi \board_state[156]$_DFFE_PP__509  (.L_HI(net509));
 sg13g2_tiehi \board_state[157]$_DFFE_PP__510  (.L_HI(net510));
 sg13g2_tiehi \board_state[158]$_DFFE_PP__511  (.L_HI(net511));
 sg13g2_tiehi \board_state[159]$_DFFE_PP__512  (.L_HI(net512));
 sg13g2_tiehi \board_state[15]$_DFFE_PP__513  (.L_HI(net513));
 sg13g2_tiehi \board_state[160]$_DFFE_PP__514  (.L_HI(net514));
 sg13g2_tiehi \board_state[161]$_DFFE_PP__515  (.L_HI(net515));
 sg13g2_tiehi \board_state[162]$_DFFE_PP__516  (.L_HI(net516));
 sg13g2_tiehi \board_state[163]$_DFFE_PP__517  (.L_HI(net517));
 sg13g2_tiehi \board_state[164]$_DFFE_PP__518  (.L_HI(net518));
 sg13g2_tiehi \board_state[165]$_DFFE_PP__519  (.L_HI(net519));
 sg13g2_tiehi \board_state[166]$_DFFE_PP__520  (.L_HI(net520));
 sg13g2_tiehi \board_state[167]$_DFFE_PP__521  (.L_HI(net521));
 sg13g2_tiehi \board_state[168]$_DFFE_PP__522  (.L_HI(net522));
 sg13g2_tiehi \board_state[169]$_DFFE_PP__523  (.L_HI(net523));
 sg13g2_tiehi \board_state[16]$_DFFE_PP__524  (.L_HI(net524));
 sg13g2_tiehi \board_state[170]$_DFFE_PP__525  (.L_HI(net525));
 sg13g2_tiehi \board_state[171]$_DFFE_PP__526  (.L_HI(net526));
 sg13g2_tiehi \board_state[172]$_DFFE_PP__527  (.L_HI(net527));
 sg13g2_tiehi \board_state[173]$_DFFE_PP__528  (.L_HI(net528));
 sg13g2_tiehi \board_state[174]$_DFFE_PP__529  (.L_HI(net529));
 sg13g2_tiehi \board_state[175]$_DFFE_PP__530  (.L_HI(net530));
 sg13g2_tiehi \board_state[176]$_DFFE_PP__531  (.L_HI(net531));
 sg13g2_tiehi \board_state[177]$_DFFE_PP__532  (.L_HI(net532));
 sg13g2_tiehi \board_state[178]$_DFFE_PP__533  (.L_HI(net533));
 sg13g2_tiehi \board_state[179]$_DFFE_PP__534  (.L_HI(net534));
 sg13g2_tiehi \board_state[17]$_DFFE_PP__535  (.L_HI(net535));
 sg13g2_tiehi \board_state[180]$_DFFE_PP__536  (.L_HI(net536));
 sg13g2_tiehi \board_state[181]$_DFFE_PP__537  (.L_HI(net537));
 sg13g2_tiehi \board_state[182]$_DFFE_PP__538  (.L_HI(net538));
 sg13g2_tiehi \board_state[183]$_DFFE_PP__539  (.L_HI(net539));
 sg13g2_tiehi \board_state[184]$_DFFE_PP__540  (.L_HI(net540));
 sg13g2_tiehi \board_state[185]$_DFFE_PP__541  (.L_HI(net541));
 sg13g2_tiehi \board_state[186]$_DFFE_PP__542  (.L_HI(net542));
 sg13g2_tiehi \board_state[187]$_DFFE_PP__543  (.L_HI(net543));
 sg13g2_tiehi \board_state[188]$_DFFE_PP__544  (.L_HI(net544));
 sg13g2_tiehi \board_state[189]$_DFFE_PP__545  (.L_HI(net545));
 sg13g2_tiehi \board_state[18]$_DFFE_PP__546  (.L_HI(net546));
 sg13g2_tiehi \board_state[190]$_DFFE_PP__547  (.L_HI(net547));
 sg13g2_tiehi \board_state[191]$_DFFE_PP__548  (.L_HI(net548));
 sg13g2_tiehi \board_state[192]$_DFFE_PP__549  (.L_HI(net549));
 sg13g2_tiehi \board_state[193]$_DFFE_PP__550  (.L_HI(net550));
 sg13g2_tiehi \board_state[194]$_DFFE_PP__551  (.L_HI(net551));
 sg13g2_tiehi \board_state[195]$_DFFE_PP__552  (.L_HI(net552));
 sg13g2_tiehi \board_state[196]$_DFFE_PP__553  (.L_HI(net553));
 sg13g2_tiehi \board_state[197]$_DFFE_PP__554  (.L_HI(net554));
 sg13g2_tiehi \board_state[198]$_DFFE_PP__555  (.L_HI(net555));
 sg13g2_tiehi \board_state[199]$_DFFE_PP__556  (.L_HI(net556));
 sg13g2_tiehi \board_state[19]$_DFFE_PP__557  (.L_HI(net557));
 sg13g2_tiehi \board_state[1]$_DFFE_PP__558  (.L_HI(net558));
 sg13g2_tiehi \board_state[200]$_DFFE_PP__559  (.L_HI(net559));
 sg13g2_tiehi \board_state[201]$_DFFE_PP__560  (.L_HI(net560));
 sg13g2_tiehi \board_state[202]$_DFFE_PP__561  (.L_HI(net561));
 sg13g2_tiehi \board_state[203]$_DFFE_PP__562  (.L_HI(net562));
 sg13g2_tiehi \board_state[204]$_DFFE_PP__563  (.L_HI(net563));
 sg13g2_tiehi \board_state[205]$_DFFE_PP__564  (.L_HI(net564));
 sg13g2_tiehi \board_state[206]$_DFFE_PP__565  (.L_HI(net565));
 sg13g2_tiehi \board_state[207]$_DFFE_PP__566  (.L_HI(net566));
 sg13g2_tiehi \board_state[208]$_DFFE_PP__567  (.L_HI(net567));
 sg13g2_tiehi \board_state[209]$_DFFE_PP__568  (.L_HI(net568));
 sg13g2_tiehi \board_state[20]$_DFFE_PP__569  (.L_HI(net569));
 sg13g2_tiehi \board_state[210]$_DFFE_PP__570  (.L_HI(net570));
 sg13g2_tiehi \board_state[211]$_DFFE_PP__571  (.L_HI(net571));
 sg13g2_tiehi \board_state[212]$_DFFE_PP__572  (.L_HI(net572));
 sg13g2_tiehi \board_state[213]$_DFFE_PP__573  (.L_HI(net573));
 sg13g2_tiehi \board_state[214]$_DFFE_PP__574  (.L_HI(net574));
 sg13g2_tiehi \board_state[215]$_DFFE_PP__575  (.L_HI(net575));
 sg13g2_tiehi \board_state[216]$_DFFE_PP__576  (.L_HI(net576));
 sg13g2_tiehi \board_state[217]$_DFFE_PP__577  (.L_HI(net577));
 sg13g2_tiehi \board_state[218]$_DFFE_PP__578  (.L_HI(net578));
 sg13g2_tiehi \board_state[219]$_DFFE_PP__579  (.L_HI(net579));
 sg13g2_tiehi \board_state[21]$_DFFE_PP__580  (.L_HI(net580));
 sg13g2_tiehi \board_state[220]$_DFFE_PP__581  (.L_HI(net581));
 sg13g2_tiehi \board_state[221]$_DFFE_PP__582  (.L_HI(net582));
 sg13g2_tiehi \board_state[222]$_DFFE_PP__583  (.L_HI(net583));
 sg13g2_tiehi \board_state[223]$_DFFE_PP__584  (.L_HI(net584));
 sg13g2_tiehi \board_state[224]$_DFFE_PP__585  (.L_HI(net585));
 sg13g2_tiehi \board_state[225]$_DFFE_PP__586  (.L_HI(net586));
 sg13g2_tiehi \board_state[226]$_DFFE_PP__587  (.L_HI(net587));
 sg13g2_tiehi \board_state[227]$_DFFE_PP__588  (.L_HI(net588));
 sg13g2_tiehi \board_state[228]$_DFFE_PP__589  (.L_HI(net589));
 sg13g2_tiehi \board_state[229]$_DFFE_PP__590  (.L_HI(net590));
 sg13g2_tiehi \board_state[22]$_DFFE_PP__591  (.L_HI(net591));
 sg13g2_tiehi \board_state[230]$_DFFE_PP__592  (.L_HI(net592));
 sg13g2_tiehi \board_state[231]$_DFFE_PP__593  (.L_HI(net593));
 sg13g2_tiehi \board_state[232]$_DFFE_PP__594  (.L_HI(net594));
 sg13g2_tiehi \board_state[233]$_DFFE_PP__595  (.L_HI(net595));
 sg13g2_tiehi \board_state[234]$_DFFE_PP__596  (.L_HI(net596));
 sg13g2_tiehi \board_state[235]$_DFFE_PP__597  (.L_HI(net597));
 sg13g2_tiehi \board_state[236]$_DFFE_PP__598  (.L_HI(net598));
 sg13g2_tiehi \board_state[237]$_DFFE_PP__599  (.L_HI(net599));
 sg13g2_tiehi \board_state[238]$_DFFE_PP__600  (.L_HI(net600));
 sg13g2_tiehi \board_state[239]$_DFFE_PP__601  (.L_HI(net601));
 sg13g2_tiehi \board_state[23]$_DFFE_PP__602  (.L_HI(net602));
 sg13g2_tiehi \board_state[240]$_DFFE_PP__603  (.L_HI(net603));
 sg13g2_tiehi \board_state[241]$_DFFE_PP__604  (.L_HI(net604));
 sg13g2_tiehi \board_state[242]$_DFFE_PP__605  (.L_HI(net605));
 sg13g2_tiehi \board_state[243]$_DFFE_PP__606  (.L_HI(net606));
 sg13g2_tiehi \board_state[244]$_DFFE_PP__607  (.L_HI(net607));
 sg13g2_tiehi \board_state[245]$_DFFE_PP__608  (.L_HI(net608));
 sg13g2_tiehi \board_state[246]$_DFFE_PP__609  (.L_HI(net609));
 sg13g2_tiehi \board_state[247]$_DFFE_PP__610  (.L_HI(net610));
 sg13g2_tiehi \board_state[248]$_DFFE_PP__611  (.L_HI(net611));
 sg13g2_tiehi \board_state[249]$_DFFE_PP__612  (.L_HI(net612));
 sg13g2_tiehi \board_state[24]$_DFFE_PP__613  (.L_HI(net613));
 sg13g2_tiehi \board_state[250]$_DFFE_PP__614  (.L_HI(net614));
 sg13g2_tiehi \board_state[251]$_DFFE_PP__615  (.L_HI(net615));
 sg13g2_tiehi \board_state[252]$_DFFE_PP__616  (.L_HI(net616));
 sg13g2_tiehi \board_state[253]$_DFFE_PP__617  (.L_HI(net617));
 sg13g2_tiehi \board_state[254]$_DFFE_PP__618  (.L_HI(net618));
 sg13g2_tiehi \board_state[255]$_DFFE_PP__619  (.L_HI(net619));
 sg13g2_tiehi \board_state[256]$_DFFE_PP__620  (.L_HI(net620));
 sg13g2_tiehi \board_state[257]$_DFFE_PP__621  (.L_HI(net621));
 sg13g2_tiehi \board_state[258]$_DFFE_PP__622  (.L_HI(net622));
 sg13g2_tiehi \board_state[259]$_DFFE_PP__623  (.L_HI(net623));
 sg13g2_tiehi \board_state[25]$_DFFE_PP__624  (.L_HI(net624));
 sg13g2_tiehi \board_state[260]$_DFFE_PP__625  (.L_HI(net625));
 sg13g2_tiehi \board_state[261]$_DFFE_PP__626  (.L_HI(net626));
 sg13g2_tiehi \board_state[262]$_DFFE_PP__627  (.L_HI(net627));
 sg13g2_tiehi \board_state[263]$_DFFE_PP__628  (.L_HI(net628));
 sg13g2_tiehi \board_state[264]$_DFFE_PP__629  (.L_HI(net629));
 sg13g2_tiehi \board_state[265]$_DFFE_PP__630  (.L_HI(net630));
 sg13g2_tiehi \board_state[266]$_DFFE_PP__631  (.L_HI(net631));
 sg13g2_tiehi \board_state[267]$_DFFE_PP__632  (.L_HI(net632));
 sg13g2_tiehi \board_state[268]$_DFFE_PP__633  (.L_HI(net633));
 sg13g2_tiehi \board_state[269]$_DFFE_PP__634  (.L_HI(net634));
 sg13g2_tiehi \board_state[26]$_DFFE_PP__635  (.L_HI(net635));
 sg13g2_tiehi \board_state[270]$_DFFE_PP__636  (.L_HI(net636));
 sg13g2_tiehi \board_state[271]$_DFFE_PP__637  (.L_HI(net637));
 sg13g2_tiehi \board_state[272]$_DFFE_PP__638  (.L_HI(net638));
 sg13g2_tiehi \board_state[273]$_DFFE_PP__639  (.L_HI(net639));
 sg13g2_tiehi \board_state[274]$_DFFE_PP__640  (.L_HI(net640));
 sg13g2_tiehi \board_state[275]$_DFFE_PP__641  (.L_HI(net641));
 sg13g2_tiehi \board_state[276]$_DFFE_PP__642  (.L_HI(net642));
 sg13g2_tiehi \board_state[277]$_DFFE_PP__643  (.L_HI(net643));
 sg13g2_tiehi \board_state[278]$_DFFE_PP__644  (.L_HI(net644));
 sg13g2_tiehi \board_state[279]$_DFFE_PP__645  (.L_HI(net645));
 sg13g2_tiehi \board_state[27]$_DFFE_PP__646  (.L_HI(net646));
 sg13g2_tiehi \board_state[280]$_DFFE_PP__647  (.L_HI(net647));
 sg13g2_tiehi \board_state[281]$_DFFE_PP__648  (.L_HI(net648));
 sg13g2_tiehi \board_state[282]$_DFFE_PP__649  (.L_HI(net649));
 sg13g2_tiehi \board_state[283]$_DFFE_PP__650  (.L_HI(net650));
 sg13g2_tiehi \board_state[284]$_DFFE_PP__651  (.L_HI(net651));
 sg13g2_tiehi \board_state[285]$_DFFE_PP__652  (.L_HI(net652));
 sg13g2_tiehi \board_state[286]$_DFFE_PP__653  (.L_HI(net653));
 sg13g2_tiehi \board_state[287]$_DFFE_PP__654  (.L_HI(net654));
 sg13g2_tiehi \board_state[288]$_DFFE_PP__655  (.L_HI(net655));
 sg13g2_tiehi \board_state[289]$_DFFE_PP__656  (.L_HI(net656));
 sg13g2_tiehi \board_state[28]$_DFFE_PP__657  (.L_HI(net657));
 sg13g2_tiehi \board_state[290]$_DFFE_PP__658  (.L_HI(net658));
 sg13g2_tiehi \board_state[291]$_DFFE_PP__659  (.L_HI(net659));
 sg13g2_tiehi \board_state[292]$_DFFE_PP__660  (.L_HI(net660));
 sg13g2_tiehi \board_state[293]$_DFFE_PP__661  (.L_HI(net661));
 sg13g2_tiehi \board_state[294]$_DFFE_PP__662  (.L_HI(net662));
 sg13g2_tiehi \board_state[295]$_DFFE_PP__663  (.L_HI(net663));
 sg13g2_tiehi \board_state[296]$_DFFE_PP__664  (.L_HI(net664));
 sg13g2_tiehi \board_state[297]$_DFFE_PP__665  (.L_HI(net665));
 sg13g2_tiehi \board_state[298]$_DFFE_PP__666  (.L_HI(net666));
 sg13g2_tiehi \board_state[299]$_DFFE_PP__667  (.L_HI(net667));
 sg13g2_tiehi \board_state[29]$_DFFE_PP__668  (.L_HI(net668));
 sg13g2_tiehi \board_state[2]$_DFFE_PP__669  (.L_HI(net669));
 sg13g2_tiehi \board_state[300]$_DFFE_PP__670  (.L_HI(net670));
 sg13g2_tiehi \board_state[301]$_DFFE_PP__671  (.L_HI(net671));
 sg13g2_tiehi \board_state[302]$_DFFE_PP__672  (.L_HI(net672));
 sg13g2_tiehi \board_state[303]$_DFFE_PP__673  (.L_HI(net673));
 sg13g2_tiehi \board_state[304]$_DFFE_PP__674  (.L_HI(net674));
 sg13g2_tiehi \board_state[305]$_DFFE_PP__675  (.L_HI(net675));
 sg13g2_tiehi \board_state[306]$_DFFE_PP__676  (.L_HI(net676));
 sg13g2_tiehi \board_state[307]$_DFFE_PP__677  (.L_HI(net677));
 sg13g2_tiehi \board_state[308]$_DFFE_PP__678  (.L_HI(net678));
 sg13g2_tiehi \board_state[309]$_DFFE_PP__679  (.L_HI(net679));
 sg13g2_tiehi \board_state[30]$_DFFE_PP__680  (.L_HI(net680));
 sg13g2_tiehi \board_state[310]$_DFFE_PP__681  (.L_HI(net681));
 sg13g2_tiehi \board_state[311]$_DFFE_PP__682  (.L_HI(net682));
 sg13g2_tiehi \board_state[312]$_DFFE_PP__683  (.L_HI(net683));
 sg13g2_tiehi \board_state[313]$_DFFE_PP__684  (.L_HI(net684));
 sg13g2_tiehi \board_state[314]$_DFFE_PP__685  (.L_HI(net685));
 sg13g2_tiehi \board_state[315]$_DFFE_PP__686  (.L_HI(net686));
 sg13g2_tiehi \board_state[316]$_DFFE_PP__687  (.L_HI(net687));
 sg13g2_tiehi \board_state[317]$_DFFE_PP__688  (.L_HI(net688));
 sg13g2_tiehi \board_state[318]$_DFFE_PP__689  (.L_HI(net689));
 sg13g2_tiehi \board_state[319]$_DFFE_PP__690  (.L_HI(net690));
 sg13g2_tiehi \board_state[31]$_DFFE_PP__691  (.L_HI(net691));
 sg13g2_tiehi \board_state[320]$_DFFE_PP__692  (.L_HI(net692));
 sg13g2_tiehi \board_state[321]$_DFFE_PP__693  (.L_HI(net693));
 sg13g2_tiehi \board_state[322]$_DFFE_PP__694  (.L_HI(net694));
 sg13g2_tiehi \board_state[323]$_DFFE_PP__695  (.L_HI(net695));
 sg13g2_tiehi \board_state[324]$_DFFE_PP__696  (.L_HI(net696));
 sg13g2_tiehi \board_state[325]$_DFFE_PP__697  (.L_HI(net697));
 sg13g2_tiehi \board_state[326]$_DFFE_PP__698  (.L_HI(net698));
 sg13g2_tiehi \board_state[327]$_DFFE_PP__699  (.L_HI(net699));
 sg13g2_tiehi \board_state[328]$_DFFE_PP__700  (.L_HI(net700));
 sg13g2_tiehi \board_state[329]$_DFFE_PP__701  (.L_HI(net701));
 sg13g2_tiehi \board_state[32]$_DFFE_PP__702  (.L_HI(net702));
 sg13g2_tiehi \board_state[330]$_DFFE_PP__703  (.L_HI(net703));
 sg13g2_tiehi \board_state[331]$_DFFE_PP__704  (.L_HI(net704));
 sg13g2_tiehi \board_state[332]$_DFFE_PP__705  (.L_HI(net705));
 sg13g2_tiehi \board_state[333]$_DFFE_PP__706  (.L_HI(net706));
 sg13g2_tiehi \board_state[334]$_DFFE_PP__707  (.L_HI(net707));
 sg13g2_tiehi \board_state[335]$_DFFE_PP__708  (.L_HI(net708));
 sg13g2_tiehi \board_state[336]$_DFFE_PP__709  (.L_HI(net709));
 sg13g2_tiehi \board_state[337]$_DFFE_PP__710  (.L_HI(net710));
 sg13g2_tiehi \board_state[338]$_DFFE_PP__711  (.L_HI(net711));
 sg13g2_tiehi \board_state[339]$_DFFE_PP__712  (.L_HI(net712));
 sg13g2_tiehi \board_state[33]$_DFFE_PP__713  (.L_HI(net713));
 sg13g2_tiehi \board_state[340]$_DFFE_PP__714  (.L_HI(net714));
 sg13g2_tiehi \board_state[341]$_DFFE_PP__715  (.L_HI(net715));
 sg13g2_tiehi \board_state[342]$_DFFE_PP__716  (.L_HI(net716));
 sg13g2_tiehi \board_state[343]$_DFFE_PP__717  (.L_HI(net717));
 sg13g2_tiehi \board_state[344]$_DFFE_PP__718  (.L_HI(net718));
 sg13g2_tiehi \board_state[345]$_DFFE_PP__719  (.L_HI(net719));
 sg13g2_tiehi \board_state[346]$_DFFE_PP__720  (.L_HI(net720));
 sg13g2_tiehi \board_state[347]$_DFFE_PP__721  (.L_HI(net721));
 sg13g2_tiehi \board_state[348]$_DFFE_PP__722  (.L_HI(net722));
 sg13g2_tiehi \board_state[349]$_DFFE_PP__723  (.L_HI(net723));
 sg13g2_tiehi \board_state[34]$_DFFE_PP__724  (.L_HI(net724));
 sg13g2_tiehi \board_state[350]$_DFFE_PP__725  (.L_HI(net725));
 sg13g2_tiehi \board_state[351]$_DFFE_PP__726  (.L_HI(net726));
 sg13g2_tiehi \board_state[352]$_DFFE_PP__727  (.L_HI(net727));
 sg13g2_tiehi \board_state[353]$_DFFE_PP__728  (.L_HI(net728));
 sg13g2_tiehi \board_state[354]$_DFFE_PP__729  (.L_HI(net729));
 sg13g2_tiehi \board_state[355]$_DFFE_PP__730  (.L_HI(net730));
 sg13g2_tiehi \board_state[356]$_DFFE_PP__731  (.L_HI(net731));
 sg13g2_tiehi \board_state[357]$_DFFE_PP__732  (.L_HI(net732));
 sg13g2_tiehi \board_state[358]$_DFFE_PP__733  (.L_HI(net733));
 sg13g2_tiehi \board_state[359]$_DFFE_PP__734  (.L_HI(net734));
 sg13g2_tiehi \board_state[35]$_DFFE_PP__735  (.L_HI(net735));
 sg13g2_tiehi \board_state[360]$_DFFE_PP__736  (.L_HI(net736));
 sg13g2_tiehi \board_state[361]$_DFFE_PP__737  (.L_HI(net737));
 sg13g2_tiehi \board_state[362]$_DFFE_PP__738  (.L_HI(net738));
 sg13g2_tiehi \board_state[363]$_DFFE_PP__739  (.L_HI(net739));
 sg13g2_tiehi \board_state[364]$_DFFE_PP__740  (.L_HI(net740));
 sg13g2_tiehi \board_state[365]$_DFFE_PP__741  (.L_HI(net741));
 sg13g2_tiehi \board_state[366]$_DFFE_PP__742  (.L_HI(net742));
 sg13g2_tiehi \board_state[367]$_DFFE_PP__743  (.L_HI(net743));
 sg13g2_tiehi \board_state[368]$_DFFE_PP__744  (.L_HI(net744));
 sg13g2_tiehi \board_state[369]$_DFFE_PP__745  (.L_HI(net745));
 sg13g2_tiehi \board_state[36]$_DFFE_PP__746  (.L_HI(net746));
 sg13g2_tiehi \board_state[370]$_DFFE_PP__747  (.L_HI(net747));
 sg13g2_tiehi \board_state[371]$_DFFE_PP__748  (.L_HI(net748));
 sg13g2_tiehi \board_state[372]$_DFFE_PP__749  (.L_HI(net749));
 sg13g2_tiehi \board_state[373]$_DFFE_PP__750  (.L_HI(net750));
 sg13g2_tiehi \board_state[374]$_DFFE_PP__751  (.L_HI(net751));
 sg13g2_tiehi \board_state[375]$_DFFE_PP__752  (.L_HI(net752));
 sg13g2_tiehi \board_state[376]$_DFFE_PP__753  (.L_HI(net753));
 sg13g2_tiehi \board_state[377]$_DFFE_PP__754  (.L_HI(net754));
 sg13g2_tiehi \board_state[378]$_DFFE_PP__755  (.L_HI(net755));
 sg13g2_tiehi \board_state[379]$_DFFE_PP__756  (.L_HI(net756));
 sg13g2_tiehi \board_state[37]$_DFFE_PP__757  (.L_HI(net757));
 sg13g2_tiehi \board_state[380]$_DFFE_PP__758  (.L_HI(net758));
 sg13g2_tiehi \board_state[381]$_DFFE_PP__759  (.L_HI(net759));
 sg13g2_tiehi \board_state[382]$_DFFE_PP__760  (.L_HI(net760));
 sg13g2_tiehi \board_state[383]$_DFFE_PP__761  (.L_HI(net761));
 sg13g2_tiehi \board_state[384]$_DFFE_PP__762  (.L_HI(net762));
 sg13g2_tiehi \board_state[385]$_DFFE_PP__763  (.L_HI(net763));
 sg13g2_tiehi \board_state[386]$_DFFE_PP__764  (.L_HI(net764));
 sg13g2_tiehi \board_state[387]$_DFFE_PP__765  (.L_HI(net765));
 sg13g2_tiehi \board_state[388]$_DFFE_PP__766  (.L_HI(net766));
 sg13g2_tiehi \board_state[389]$_DFFE_PP__767  (.L_HI(net767));
 sg13g2_tiehi \board_state[38]$_DFFE_PP__768  (.L_HI(net768));
 sg13g2_tiehi \board_state[390]$_DFFE_PP__769  (.L_HI(net769));
 sg13g2_tiehi \board_state[391]$_DFFE_PP__770  (.L_HI(net770));
 sg13g2_tiehi \board_state[392]$_DFFE_PP__771  (.L_HI(net771));
 sg13g2_tiehi \board_state[393]$_DFFE_PP__772  (.L_HI(net772));
 sg13g2_tiehi \board_state[394]$_DFFE_PP__773  (.L_HI(net773));
 sg13g2_tiehi \board_state[395]$_DFFE_PP__774  (.L_HI(net774));
 sg13g2_tiehi \board_state[396]$_DFFE_PP__775  (.L_HI(net775));
 sg13g2_tiehi \board_state[397]$_DFFE_PP__776  (.L_HI(net776));
 sg13g2_tiehi \board_state[398]$_DFFE_PP__777  (.L_HI(net777));
 sg13g2_tiehi \board_state[399]$_DFFE_PP__778  (.L_HI(net778));
 sg13g2_tiehi \board_state[39]$_DFFE_PP__779  (.L_HI(net779));
 sg13g2_tiehi \board_state[3]$_DFFE_PP__780  (.L_HI(net780));
 sg13g2_tiehi \board_state[400]$_DFFE_PP__781  (.L_HI(net781));
 sg13g2_tiehi \board_state[401]$_DFFE_PP__782  (.L_HI(net782));
 sg13g2_tiehi \board_state[402]$_DFFE_PP__783  (.L_HI(net783));
 sg13g2_tiehi \board_state[403]$_DFFE_PP__784  (.L_HI(net784));
 sg13g2_tiehi \board_state[404]$_DFFE_PP__785  (.L_HI(net785));
 sg13g2_tiehi \board_state[405]$_DFFE_PP__786  (.L_HI(net786));
 sg13g2_tiehi \board_state[406]$_DFFE_PP__787  (.L_HI(net787));
 sg13g2_tiehi \board_state[407]$_DFFE_PP__788  (.L_HI(net788));
 sg13g2_tiehi \board_state[408]$_DFFE_PP__789  (.L_HI(net789));
 sg13g2_tiehi \board_state[409]$_DFFE_PP__790  (.L_HI(net790));
 sg13g2_tiehi \board_state[40]$_DFFE_PP__791  (.L_HI(net791));
 sg13g2_tiehi \board_state[410]$_DFFE_PP__792  (.L_HI(net792));
 sg13g2_tiehi \board_state[411]$_DFFE_PP__793  (.L_HI(net793));
 sg13g2_tiehi \board_state[412]$_DFFE_PP__794  (.L_HI(net794));
 sg13g2_tiehi \board_state[413]$_DFFE_PP__795  (.L_HI(net795));
 sg13g2_tiehi \board_state[414]$_DFFE_PP__796  (.L_HI(net796));
 sg13g2_tiehi \board_state[415]$_DFFE_PP__797  (.L_HI(net797));
 sg13g2_tiehi \board_state[416]$_DFFE_PP__798  (.L_HI(net798));
 sg13g2_tiehi \board_state[417]$_DFFE_PP__799  (.L_HI(net799));
 sg13g2_tiehi \board_state[418]$_DFFE_PP__800  (.L_HI(net800));
 sg13g2_tiehi \board_state[419]$_DFFE_PP__801  (.L_HI(net801));
 sg13g2_tiehi \board_state[41]$_DFFE_PP__802  (.L_HI(net802));
 sg13g2_tiehi \board_state[420]$_DFFE_PP__803  (.L_HI(net803));
 sg13g2_tiehi \board_state[421]$_DFFE_PP__804  (.L_HI(net804));
 sg13g2_tiehi \board_state[422]$_DFFE_PP__805  (.L_HI(net805));
 sg13g2_tiehi \board_state[423]$_DFFE_PP__806  (.L_HI(net806));
 sg13g2_tiehi \board_state[424]$_DFFE_PP__807  (.L_HI(net807));
 sg13g2_tiehi \board_state[425]$_DFFE_PP__808  (.L_HI(net808));
 sg13g2_tiehi \board_state[426]$_DFFE_PP__809  (.L_HI(net809));
 sg13g2_tiehi \board_state[427]$_DFFE_PP__810  (.L_HI(net810));
 sg13g2_tiehi \board_state[428]$_DFFE_PP__811  (.L_HI(net811));
 sg13g2_tiehi \board_state[429]$_DFFE_PP__812  (.L_HI(net812));
 sg13g2_tiehi \board_state[42]$_DFFE_PP__813  (.L_HI(net813));
 sg13g2_tiehi \board_state[430]$_DFFE_PP__814  (.L_HI(net814));
 sg13g2_tiehi \board_state[431]$_DFFE_PP__815  (.L_HI(net815));
 sg13g2_tiehi \board_state[432]$_DFFE_PP__816  (.L_HI(net816));
 sg13g2_tiehi \board_state[433]$_DFFE_PP__817  (.L_HI(net817));
 sg13g2_tiehi \board_state[434]$_DFFE_PP__818  (.L_HI(net818));
 sg13g2_tiehi \board_state[435]$_DFFE_PP__819  (.L_HI(net819));
 sg13g2_tiehi \board_state[436]$_DFFE_PP__820  (.L_HI(net820));
 sg13g2_tiehi \board_state[437]$_DFFE_PP__821  (.L_HI(net821));
 sg13g2_tiehi \board_state[438]$_DFFE_PP__822  (.L_HI(net822));
 sg13g2_tiehi \board_state[439]$_DFFE_PP__823  (.L_HI(net823));
 sg13g2_tiehi \board_state[43]$_DFFE_PP__824  (.L_HI(net824));
 sg13g2_tiehi \board_state[440]$_DFFE_PP__825  (.L_HI(net825));
 sg13g2_tiehi \board_state[441]$_DFFE_PP__826  (.L_HI(net826));
 sg13g2_tiehi \board_state[442]$_DFFE_PP__827  (.L_HI(net827));
 sg13g2_tiehi \board_state[443]$_DFFE_PP__828  (.L_HI(net828));
 sg13g2_tiehi \board_state[444]$_DFFE_PP__829  (.L_HI(net829));
 sg13g2_tiehi \board_state[445]$_DFFE_PP__830  (.L_HI(net830));
 sg13g2_tiehi \board_state[446]$_DFFE_PP__831  (.L_HI(net831));
 sg13g2_tiehi \board_state[447]$_DFFE_PP__832  (.L_HI(net832));
 sg13g2_tiehi \board_state[448]$_DFFE_PP__833  (.L_HI(net833));
 sg13g2_tiehi \board_state[449]$_DFFE_PP__834  (.L_HI(net834));
 sg13g2_tiehi \board_state[44]$_DFFE_PP__835  (.L_HI(net835));
 sg13g2_tiehi \board_state[450]$_DFFE_PP__836  (.L_HI(net836));
 sg13g2_tiehi \board_state[451]$_DFFE_PP__837  (.L_HI(net837));
 sg13g2_tiehi \board_state[452]$_DFFE_PP__838  (.L_HI(net838));
 sg13g2_tiehi \board_state[453]$_DFFE_PP__839  (.L_HI(net839));
 sg13g2_tiehi \board_state[454]$_DFFE_PP__840  (.L_HI(net840));
 sg13g2_tiehi \board_state[455]$_DFFE_PP__841  (.L_HI(net841));
 sg13g2_tiehi \board_state[456]$_DFFE_PP__842  (.L_HI(net842));
 sg13g2_tiehi \board_state[457]$_DFFE_PP__843  (.L_HI(net843));
 sg13g2_tiehi \board_state[458]$_DFFE_PP__844  (.L_HI(net844));
 sg13g2_tiehi \board_state[459]$_DFFE_PP__845  (.L_HI(net845));
 sg13g2_tiehi \board_state[45]$_DFFE_PP__846  (.L_HI(net846));
 sg13g2_tiehi \board_state[460]$_DFFE_PP__847  (.L_HI(net847));
 sg13g2_tiehi \board_state[461]$_DFFE_PP__848  (.L_HI(net848));
 sg13g2_tiehi \board_state[462]$_DFFE_PP__849  (.L_HI(net849));
 sg13g2_tiehi \board_state[463]$_DFFE_PP__850  (.L_HI(net850));
 sg13g2_tiehi \board_state[464]$_DFFE_PP__851  (.L_HI(net851));
 sg13g2_tiehi \board_state[465]$_DFFE_PP__852  (.L_HI(net852));
 sg13g2_tiehi \board_state[466]$_DFFE_PP__853  (.L_HI(net853));
 sg13g2_tiehi \board_state[467]$_DFFE_PP__854  (.L_HI(net854));
 sg13g2_tiehi \board_state[468]$_DFFE_PP__855  (.L_HI(net855));
 sg13g2_tiehi \board_state[469]$_DFFE_PP__856  (.L_HI(net856));
 sg13g2_tiehi \board_state[46]$_DFFE_PP__857  (.L_HI(net857));
 sg13g2_tiehi \board_state[470]$_DFFE_PP__858  (.L_HI(net858));
 sg13g2_tiehi \board_state[471]$_DFFE_PP__859  (.L_HI(net859));
 sg13g2_tiehi \board_state[472]$_DFFE_PP__860  (.L_HI(net860));
 sg13g2_tiehi \board_state[473]$_DFFE_PP__861  (.L_HI(net861));
 sg13g2_tiehi \board_state[474]$_DFFE_PP__862  (.L_HI(net862));
 sg13g2_tiehi \board_state[475]$_DFFE_PP__863  (.L_HI(net863));
 sg13g2_tiehi \board_state[476]$_DFFE_PP__864  (.L_HI(net864));
 sg13g2_tiehi \board_state[477]$_DFFE_PP__865  (.L_HI(net865));
 sg13g2_tiehi \board_state[478]$_DFFE_PP__866  (.L_HI(net866));
 sg13g2_tiehi \board_state[479]$_DFFE_PP__867  (.L_HI(net867));
 sg13g2_tiehi \board_state[47]$_DFFE_PP__868  (.L_HI(net868));
 sg13g2_tiehi \board_state[480]$_DFFE_PP__869  (.L_HI(net869));
 sg13g2_tiehi \board_state[481]$_DFFE_PP__870  (.L_HI(net870));
 sg13g2_tiehi \board_state[482]$_DFFE_PP__871  (.L_HI(net871));
 sg13g2_tiehi \board_state[483]$_DFFE_PP__872  (.L_HI(net872));
 sg13g2_tiehi \board_state[484]$_DFFE_PP__873  (.L_HI(net873));
 sg13g2_tiehi \board_state[485]$_DFFE_PP__874  (.L_HI(net874));
 sg13g2_tiehi \board_state[486]$_DFFE_PP__875  (.L_HI(net875));
 sg13g2_tiehi \board_state[487]$_DFFE_PP__876  (.L_HI(net876));
 sg13g2_tiehi \board_state[488]$_DFFE_PP__877  (.L_HI(net877));
 sg13g2_tiehi \board_state[489]$_DFFE_PP__878  (.L_HI(net878));
 sg13g2_tiehi \board_state[48]$_DFFE_PP__879  (.L_HI(net879));
 sg13g2_tiehi \board_state[490]$_DFFE_PP__880  (.L_HI(net880));
 sg13g2_tiehi \board_state[491]$_DFFE_PP__881  (.L_HI(net881));
 sg13g2_tiehi \board_state[492]$_DFFE_PP__882  (.L_HI(net882));
 sg13g2_tiehi \board_state[493]$_DFFE_PP__883  (.L_HI(net883));
 sg13g2_tiehi \board_state[494]$_DFFE_PP__884  (.L_HI(net884));
 sg13g2_tiehi \board_state[495]$_DFFE_PP__885  (.L_HI(net885));
 sg13g2_tiehi \board_state[496]$_DFFE_PP__886  (.L_HI(net886));
 sg13g2_tiehi \board_state[497]$_DFFE_PP__887  (.L_HI(net887));
 sg13g2_tiehi \board_state[498]$_DFFE_PP__888  (.L_HI(net888));
 sg13g2_tiehi \board_state[499]$_DFFE_PP__889  (.L_HI(net889));
 sg13g2_tiehi \board_state[49]$_DFFE_PP__890  (.L_HI(net890));
 sg13g2_tiehi \board_state[4]$_DFFE_PP__891  (.L_HI(net891));
 sg13g2_tiehi \board_state[500]$_DFFE_PP__892  (.L_HI(net892));
 sg13g2_tiehi \board_state[501]$_DFFE_PP__893  (.L_HI(net893));
 sg13g2_tiehi \board_state[502]$_DFFE_PP__894  (.L_HI(net894));
 sg13g2_tiehi \board_state[503]$_DFFE_PP__895  (.L_HI(net895));
 sg13g2_tiehi \board_state[504]$_DFFE_PP__896  (.L_HI(net896));
 sg13g2_tiehi \board_state[505]$_DFFE_PP__897  (.L_HI(net897));
 sg13g2_tiehi \board_state[506]$_DFFE_PP__898  (.L_HI(net898));
 sg13g2_tiehi \board_state[507]$_DFFE_PP__899  (.L_HI(net899));
 sg13g2_tiehi \board_state[508]$_DFFE_PP__900  (.L_HI(net900));
 sg13g2_tiehi \board_state[509]$_DFFE_PP__901  (.L_HI(net901));
 sg13g2_tiehi \board_state[50]$_DFFE_PP__902  (.L_HI(net902));
 sg13g2_tiehi \board_state[510]$_DFFE_PP__903  (.L_HI(net903));
 sg13g2_tiehi \board_state[511]$_DFFE_PP__904  (.L_HI(net904));
 sg13g2_tiehi \board_state[51]$_DFFE_PP__905  (.L_HI(net905));
 sg13g2_tiehi \board_state[52]$_DFFE_PP__906  (.L_HI(net906));
 sg13g2_tiehi \board_state[53]$_DFFE_PP__907  (.L_HI(net907));
 sg13g2_tiehi \board_state[54]$_DFFE_PP__908  (.L_HI(net908));
 sg13g2_tiehi \board_state[55]$_DFFE_PP__909  (.L_HI(net909));
 sg13g2_tiehi \board_state[56]$_DFFE_PP__910  (.L_HI(net910));
 sg13g2_tiehi \board_state[57]$_DFFE_PP__911  (.L_HI(net911));
 sg13g2_tiehi \board_state[58]$_DFFE_PP__912  (.L_HI(net912));
 sg13g2_tiehi \board_state[59]$_DFFE_PP__913  (.L_HI(net913));
 sg13g2_tiehi \board_state[5]$_DFFE_PP__914  (.L_HI(net914));
 sg13g2_tiehi \board_state[60]$_DFFE_PP__915  (.L_HI(net915));
 sg13g2_tiehi \board_state[61]$_DFFE_PP__916  (.L_HI(net916));
 sg13g2_tiehi \board_state[62]$_DFFE_PP__917  (.L_HI(net917));
 sg13g2_tiehi \board_state[63]$_DFFE_PP__918  (.L_HI(net918));
 sg13g2_tiehi \board_state[64]$_DFFE_PP__919  (.L_HI(net919));
 sg13g2_tiehi \board_state[65]$_DFFE_PP__920  (.L_HI(net920));
 sg13g2_tiehi \board_state[66]$_DFFE_PP__921  (.L_HI(net921));
 sg13g2_tiehi \board_state[67]$_DFFE_PP__922  (.L_HI(net922));
 sg13g2_tiehi \board_state[68]$_DFFE_PP__923  (.L_HI(net923));
 sg13g2_tiehi \board_state[69]$_DFFE_PP__924  (.L_HI(net924));
 sg13g2_tiehi \board_state[6]$_DFFE_PP__925  (.L_HI(net925));
 sg13g2_tiehi \board_state[70]$_DFFE_PP__926  (.L_HI(net926));
 sg13g2_tiehi \board_state[71]$_DFFE_PP__927  (.L_HI(net927));
 sg13g2_tiehi \board_state[72]$_DFFE_PP__928  (.L_HI(net928));
 sg13g2_tiehi \board_state[73]$_DFFE_PP__929  (.L_HI(net929));
 sg13g2_tiehi \board_state[74]$_DFFE_PP__930  (.L_HI(net930));
 sg13g2_tiehi \board_state[75]$_DFFE_PP__931  (.L_HI(net931));
 sg13g2_tiehi \board_state[76]$_DFFE_PP__932  (.L_HI(net932));
 sg13g2_tiehi \board_state[77]$_DFFE_PP__933  (.L_HI(net933));
 sg13g2_tiehi \board_state[78]$_DFFE_PP__934  (.L_HI(net934));
 sg13g2_tiehi \board_state[79]$_DFFE_PP__935  (.L_HI(net935));
 sg13g2_tiehi \board_state[7]$_DFFE_PP__936  (.L_HI(net936));
 sg13g2_tiehi \board_state[80]$_DFFE_PP__937  (.L_HI(net937));
 sg13g2_tiehi \board_state[81]$_DFFE_PP__938  (.L_HI(net938));
 sg13g2_tiehi \board_state[82]$_DFFE_PP__939  (.L_HI(net939));
 sg13g2_tiehi \board_state[83]$_DFFE_PP__940  (.L_HI(net940));
 sg13g2_tiehi \board_state[84]$_DFFE_PP__941  (.L_HI(net941));
 sg13g2_tiehi \board_state[85]$_DFFE_PP__942  (.L_HI(net942));
 sg13g2_tiehi \board_state[86]$_DFFE_PP__943  (.L_HI(net943));
 sg13g2_tiehi \board_state[87]$_DFFE_PP__944  (.L_HI(net944));
 sg13g2_tiehi \board_state[88]$_DFFE_PP__945  (.L_HI(net945));
 sg13g2_tiehi \board_state[89]$_DFFE_PP__946  (.L_HI(net946));
 sg13g2_tiehi \board_state[8]$_DFFE_PP__947  (.L_HI(net947));
 sg13g2_tiehi \board_state[90]$_DFFE_PP__948  (.L_HI(net948));
 sg13g2_tiehi \board_state[91]$_DFFE_PP__949  (.L_HI(net949));
 sg13g2_tiehi \board_state[92]$_DFFE_PP__950  (.L_HI(net950));
 sg13g2_tiehi \board_state[93]$_DFFE_PP__951  (.L_HI(net951));
 sg13g2_tiehi \board_state[94]$_DFFE_PP__952  (.L_HI(net952));
 sg13g2_tiehi \board_state[95]$_DFFE_PP__953  (.L_HI(net953));
 sg13g2_tiehi \board_state[96]$_DFFE_PP__954  (.L_HI(net954));
 sg13g2_tiehi \board_state[97]$_DFFE_PP__955  (.L_HI(net955));
 sg13g2_tiehi \board_state[98]$_DFFE_PP__956  (.L_HI(net956));
 sg13g2_tiehi \board_state[99]$_DFFE_PP__957  (.L_HI(net957));
 sg13g2_tiehi \board_state[9]$_DFFE_PP__958  (.L_HI(net958));
 sg13g2_tiehi \board_state_next[0]$_SDFFCE_PP0P__959  (.L_HI(net959));
 sg13g2_tiehi \board_state_next[100]$_DFFE_PP__960  (.L_HI(net960));
 sg13g2_tiehi \board_state_next[101]$_DFFE_PP__961  (.L_HI(net961));
 sg13g2_tiehi \board_state_next[102]$_DFFE_PP__962  (.L_HI(net962));
 sg13g2_tiehi \board_state_next[103]$_DFFE_PP__963  (.L_HI(net963));
 sg13g2_tiehi \board_state_next[104]$_DFFE_PP__964  (.L_HI(net964));
 sg13g2_tiehi \board_state_next[105]$_DFFE_PP__965  (.L_HI(net965));
 sg13g2_tiehi \board_state_next[106]$_DFFE_PP__966  (.L_HI(net966));
 sg13g2_tiehi \board_state_next[107]$_DFFE_PP__967  (.L_HI(net967));
 sg13g2_tiehi \board_state_next[108]$_DFFE_PP__968  (.L_HI(net968));
 sg13g2_tiehi \board_state_next[109]$_DFFE_PP__969  (.L_HI(net969));
 sg13g2_tiehi \board_state_next[10]$_DFFE_PP__970  (.L_HI(net970));
 sg13g2_tiehi \board_state_next[110]$_DFFE_PP__971  (.L_HI(net971));
 sg13g2_tiehi \board_state_next[111]$_DFFE_PP__972  (.L_HI(net972));
 sg13g2_tiehi \board_state_next[112]$_DFFE_PP__973  (.L_HI(net973));
 sg13g2_tiehi \board_state_next[113]$_DFFE_PP__974  (.L_HI(net974));
 sg13g2_tiehi \board_state_next[114]$_DFFE_PP__975  (.L_HI(net975));
 sg13g2_tiehi \board_state_next[115]$_DFFE_PP__976  (.L_HI(net976));
 sg13g2_tiehi \board_state_next[116]$_DFFE_PP__977  (.L_HI(net977));
 sg13g2_tiehi \board_state_next[117]$_DFFE_PP__978  (.L_HI(net978));
 sg13g2_tiehi \board_state_next[118]$_DFFE_PP__979  (.L_HI(net979));
 sg13g2_tiehi \board_state_next[119]$_DFFE_PP__980  (.L_HI(net980));
 sg13g2_tiehi \board_state_next[11]$_DFFE_PP__981  (.L_HI(net981));
 sg13g2_tiehi \board_state_next[120]$_DFFE_PP__982  (.L_HI(net982));
 sg13g2_tiehi \board_state_next[121]$_DFFE_PP__983  (.L_HI(net983));
 sg13g2_tiehi \board_state_next[122]$_DFFE_PP__984  (.L_HI(net984));
 sg13g2_tiehi \board_state_next[123]$_DFFE_PP__985  (.L_HI(net985));
 sg13g2_tiehi \board_state_next[124]$_DFFE_PP__986  (.L_HI(net986));
 sg13g2_tiehi \board_state_next[125]$_DFFE_PP__987  (.L_HI(net987));
 sg13g2_tiehi \board_state_next[126]$_DFFE_PP__988  (.L_HI(net988));
 sg13g2_tiehi \board_state_next[127]$_DFFE_PP__989  (.L_HI(net989));
 sg13g2_tiehi \board_state_next[128]$_DFFE_PP__990  (.L_HI(net990));
 sg13g2_tiehi \board_state_next[129]$_DFFE_PP__991  (.L_HI(net991));
 sg13g2_tiehi \board_state_next[12]$_DFFE_PP__992  (.L_HI(net992));
 sg13g2_tiehi \board_state_next[130]$_DFFE_PP__993  (.L_HI(net993));
 sg13g2_tiehi \board_state_next[131]$_DFFE_PP__994  (.L_HI(net994));
 sg13g2_tiehi \board_state_next[132]$_DFFE_PP__995  (.L_HI(net995));
 sg13g2_tiehi \board_state_next[133]$_DFFE_PP__996  (.L_HI(net996));
 sg13g2_tiehi \board_state_next[134]$_DFFE_PP__997  (.L_HI(net997));
 sg13g2_tiehi \board_state_next[135]$_DFFE_PP__998  (.L_HI(net998));
 sg13g2_tiehi \board_state_next[136]$_DFFE_PP__999  (.L_HI(net999));
 sg13g2_tiehi \board_state_next[137]$_DFFE_PP__1000  (.L_HI(net1000));
 sg13g2_tiehi \board_state_next[138]$_DFFE_PP__1001  (.L_HI(net1001));
 sg13g2_tiehi \board_state_next[139]$_DFFE_PP__1002  (.L_HI(net1002));
 sg13g2_tiehi \board_state_next[13]$_DFFE_PP__1003  (.L_HI(net1003));
 sg13g2_tiehi \board_state_next[140]$_DFFE_PP__1004  (.L_HI(net1004));
 sg13g2_tiehi \board_state_next[141]$_DFFE_PP__1005  (.L_HI(net1005));
 sg13g2_tiehi \board_state_next[142]$_DFFE_PP__1006  (.L_HI(net1006));
 sg13g2_tiehi \board_state_next[143]$_DFFE_PP__1007  (.L_HI(net1007));
 sg13g2_tiehi \board_state_next[144]$_DFFE_PP__1008  (.L_HI(net1008));
 sg13g2_tiehi \board_state_next[145]$_DFFE_PP__1009  (.L_HI(net1009));
 sg13g2_tiehi \board_state_next[146]$_DFFE_PP__1010  (.L_HI(net1010));
 sg13g2_tiehi \board_state_next[147]$_DFFE_PP__1011  (.L_HI(net1011));
 sg13g2_tiehi \board_state_next[148]$_DFFE_PP__1012  (.L_HI(net1012));
 sg13g2_tiehi \board_state_next[149]$_DFFE_PP__1013  (.L_HI(net1013));
 sg13g2_tiehi \board_state_next[14]$_DFFE_PP__1014  (.L_HI(net1014));
 sg13g2_tiehi \board_state_next[150]$_DFFE_PP__1015  (.L_HI(net1015));
 sg13g2_tiehi \board_state_next[151]$_DFFE_PP__1016  (.L_HI(net1016));
 sg13g2_tiehi \board_state_next[152]$_DFFE_PP__1017  (.L_HI(net1017));
 sg13g2_tiehi \board_state_next[153]$_DFFE_PP__1018  (.L_HI(net1018));
 sg13g2_tiehi \board_state_next[154]$_DFFE_PP__1019  (.L_HI(net1019));
 sg13g2_tiehi \board_state_next[155]$_DFFE_PP__1020  (.L_HI(net1020));
 sg13g2_tiehi \board_state_next[156]$_DFFE_PP__1021  (.L_HI(net1021));
 sg13g2_tiehi \board_state_next[157]$_DFFE_PP__1022  (.L_HI(net1022));
 sg13g2_tiehi \board_state_next[158]$_DFFE_PP__1023  (.L_HI(net1023));
 sg13g2_tiehi \board_state_next[159]$_DFFE_PP__1024  (.L_HI(net1024));
 sg13g2_tiehi \board_state_next[15]$_DFFE_PP__1025  (.L_HI(net1025));
 sg13g2_tiehi \board_state_next[160]$_DFFE_PP__1026  (.L_HI(net1026));
 sg13g2_tiehi \board_state_next[161]$_DFFE_PP__1027  (.L_HI(net1027));
 sg13g2_tiehi \board_state_next[162]$_DFFE_PP__1028  (.L_HI(net1028));
 sg13g2_tiehi \board_state_next[163]$_DFFE_PP__1029  (.L_HI(net1029));
 sg13g2_tiehi \board_state_next[164]$_DFFE_PP__1030  (.L_HI(net1030));
 sg13g2_tiehi \board_state_next[165]$_DFFE_PP__1031  (.L_HI(net1031));
 sg13g2_tiehi \board_state_next[166]$_DFFE_PP__1032  (.L_HI(net1032));
 sg13g2_tiehi \board_state_next[167]$_DFFE_PP__1033  (.L_HI(net1033));
 sg13g2_tiehi \board_state_next[168]$_DFFE_PP__1034  (.L_HI(net1034));
 sg13g2_tiehi \board_state_next[169]$_DFFE_PP__1035  (.L_HI(net1035));
 sg13g2_tiehi \board_state_next[16]$_DFFE_PP__1036  (.L_HI(net1036));
 sg13g2_tiehi \board_state_next[170]$_DFFE_PP__1037  (.L_HI(net1037));
 sg13g2_tiehi \board_state_next[171]$_DFFE_PP__1038  (.L_HI(net1038));
 sg13g2_tiehi \board_state_next[172]$_DFFE_PP__1039  (.L_HI(net1039));
 sg13g2_tiehi \board_state_next[173]$_DFFE_PP__1040  (.L_HI(net1040));
 sg13g2_tiehi \board_state_next[174]$_DFFE_PP__1041  (.L_HI(net1041));
 sg13g2_tiehi \board_state_next[175]$_DFFE_PP__1042  (.L_HI(net1042));
 sg13g2_tiehi \board_state_next[176]$_DFFE_PP__1043  (.L_HI(net1043));
 sg13g2_tiehi \board_state_next[177]$_DFFE_PP__1044  (.L_HI(net1044));
 sg13g2_tiehi \board_state_next[178]$_DFFE_PP__1045  (.L_HI(net1045));
 sg13g2_tiehi \board_state_next[179]$_DFFE_PP__1046  (.L_HI(net1046));
 sg13g2_tiehi \board_state_next[17]$_DFFE_PP__1047  (.L_HI(net1047));
 sg13g2_tiehi \board_state_next[180]$_DFFE_PP__1048  (.L_HI(net1048));
 sg13g2_tiehi \board_state_next[181]$_DFFE_PP__1049  (.L_HI(net1049));
 sg13g2_tiehi \board_state_next[182]$_DFFE_PP__1050  (.L_HI(net1050));
 sg13g2_tiehi \board_state_next[183]$_DFFE_PP__1051  (.L_HI(net1051));
 sg13g2_tiehi \board_state_next[184]$_DFFE_PP__1052  (.L_HI(net1052));
 sg13g2_tiehi \board_state_next[185]$_DFFE_PP__1053  (.L_HI(net1053));
 sg13g2_tiehi \board_state_next[186]$_DFFE_PP__1054  (.L_HI(net1054));
 sg13g2_tiehi \board_state_next[187]$_DFFE_PP__1055  (.L_HI(net1055));
 sg13g2_tiehi \board_state_next[188]$_DFFE_PP__1056  (.L_HI(net1056));
 sg13g2_tiehi \board_state_next[189]$_DFFE_PP__1057  (.L_HI(net1057));
 sg13g2_tiehi \board_state_next[18]$_DFFE_PP__1058  (.L_HI(net1058));
 sg13g2_tiehi \board_state_next[190]$_DFFE_PP__1059  (.L_HI(net1059));
 sg13g2_tiehi \board_state_next[191]$_DFFE_PP__1060  (.L_HI(net1060));
 sg13g2_tiehi \board_state_next[192]$_DFFE_PP__1061  (.L_HI(net1061));
 sg13g2_tiehi \board_state_next[193]$_DFFE_PP__1062  (.L_HI(net1062));
 sg13g2_tiehi \board_state_next[194]$_DFFE_PP__1063  (.L_HI(net1063));
 sg13g2_tiehi \board_state_next[195]$_DFFE_PP__1064  (.L_HI(net1064));
 sg13g2_tiehi \board_state_next[196]$_DFFE_PP__1065  (.L_HI(net1065));
 sg13g2_tiehi \board_state_next[197]$_DFFE_PP__1066  (.L_HI(net1066));
 sg13g2_tiehi \board_state_next[198]$_DFFE_PP__1067  (.L_HI(net1067));
 sg13g2_tiehi \board_state_next[199]$_DFFE_PP__1068  (.L_HI(net1068));
 sg13g2_tiehi \board_state_next[19]$_DFFE_PP__1069  (.L_HI(net1069));
 sg13g2_tiehi \board_state_next[1]$_DFFE_PP__1070  (.L_HI(net1070));
 sg13g2_tiehi \board_state_next[200]$_DFFE_PP__1071  (.L_HI(net1071));
 sg13g2_tiehi \board_state_next[201]$_DFFE_PP__1072  (.L_HI(net1072));
 sg13g2_tiehi \board_state_next[202]$_DFFE_PP__1073  (.L_HI(net1073));
 sg13g2_tiehi \board_state_next[203]$_DFFE_PP__1074  (.L_HI(net1074));
 sg13g2_tiehi \board_state_next[204]$_DFFE_PP__1075  (.L_HI(net1075));
 sg13g2_tiehi \board_state_next[205]$_DFFE_PP__1076  (.L_HI(net1076));
 sg13g2_tiehi \board_state_next[206]$_DFFE_PP__1077  (.L_HI(net1077));
 sg13g2_tiehi \board_state_next[207]$_DFFE_PP__1078  (.L_HI(net1078));
 sg13g2_tiehi \board_state_next[208]$_DFFE_PP__1079  (.L_HI(net1079));
 sg13g2_tiehi \board_state_next[209]$_DFFE_PP__1080  (.L_HI(net1080));
 sg13g2_tiehi \board_state_next[20]$_DFFE_PP__1081  (.L_HI(net1081));
 sg13g2_tiehi \board_state_next[210]$_DFFE_PP__1082  (.L_HI(net1082));
 sg13g2_tiehi \board_state_next[211]$_DFFE_PP__1083  (.L_HI(net1083));
 sg13g2_tiehi \board_state_next[212]$_DFFE_PP__1084  (.L_HI(net1084));
 sg13g2_tiehi \board_state_next[213]$_DFFE_PP__1085  (.L_HI(net1085));
 sg13g2_tiehi \board_state_next[214]$_DFFE_PP__1086  (.L_HI(net1086));
 sg13g2_tiehi \board_state_next[215]$_DFFE_PP__1087  (.L_HI(net1087));
 sg13g2_tiehi \board_state_next[216]$_DFFE_PP__1088  (.L_HI(net1088));
 sg13g2_tiehi \board_state_next[217]$_DFFE_PP__1089  (.L_HI(net1089));
 sg13g2_tiehi \board_state_next[218]$_DFFE_PP__1090  (.L_HI(net1090));
 sg13g2_tiehi \board_state_next[219]$_DFFE_PP__1091  (.L_HI(net1091));
 sg13g2_tiehi \board_state_next[21]$_DFFE_PP__1092  (.L_HI(net1092));
 sg13g2_tiehi \board_state_next[220]$_DFFE_PP__1093  (.L_HI(net1093));
 sg13g2_tiehi \board_state_next[221]$_DFFE_PP__1094  (.L_HI(net1094));
 sg13g2_tiehi \board_state_next[222]$_DFFE_PP__1095  (.L_HI(net1095));
 sg13g2_tiehi \board_state_next[223]$_DFFE_PP__1096  (.L_HI(net1096));
 sg13g2_tiehi \board_state_next[224]$_DFFE_PP__1097  (.L_HI(net1097));
 sg13g2_tiehi \board_state_next[225]$_DFFE_PP__1098  (.L_HI(net1098));
 sg13g2_tiehi \board_state_next[226]$_DFFE_PP__1099  (.L_HI(net1099));
 sg13g2_tiehi \board_state_next[227]$_DFFE_PP__1100  (.L_HI(net1100));
 sg13g2_tiehi \board_state_next[228]$_DFFE_PP__1101  (.L_HI(net1101));
 sg13g2_tiehi \board_state_next[229]$_DFFE_PP__1102  (.L_HI(net1102));
 sg13g2_tiehi \board_state_next[22]$_DFFE_PP__1103  (.L_HI(net1103));
 sg13g2_tiehi \board_state_next[230]$_DFFE_PP__1104  (.L_HI(net1104));
 sg13g2_tiehi \board_state_next[231]$_DFFE_PP__1105  (.L_HI(net1105));
 sg13g2_tiehi \board_state_next[232]$_DFFE_PP__1106  (.L_HI(net1106));
 sg13g2_tiehi \board_state_next[233]$_DFFE_PP__1107  (.L_HI(net1107));
 sg13g2_tiehi \board_state_next[234]$_DFFE_PP__1108  (.L_HI(net1108));
 sg13g2_tiehi \board_state_next[235]$_DFFE_PP__1109  (.L_HI(net1109));
 sg13g2_tiehi \board_state_next[236]$_DFFE_PP__1110  (.L_HI(net1110));
 sg13g2_tiehi \board_state_next[237]$_DFFE_PP__1111  (.L_HI(net1111));
 sg13g2_tiehi \board_state_next[238]$_DFFE_PP__1112  (.L_HI(net1112));
 sg13g2_tiehi \board_state_next[239]$_DFFE_PP__1113  (.L_HI(net1113));
 sg13g2_tiehi \board_state_next[23]$_DFFE_PP__1114  (.L_HI(net1114));
 sg13g2_tiehi \board_state_next[240]$_DFFE_PP__1115  (.L_HI(net1115));
 sg13g2_tiehi \board_state_next[241]$_DFFE_PP__1116  (.L_HI(net1116));
 sg13g2_tiehi \board_state_next[242]$_DFFE_PP__1117  (.L_HI(net1117));
 sg13g2_tiehi \board_state_next[243]$_DFFE_PP__1118  (.L_HI(net1118));
 sg13g2_tiehi \board_state_next[244]$_DFFE_PP__1119  (.L_HI(net1119));
 sg13g2_tiehi \board_state_next[245]$_DFFE_PP__1120  (.L_HI(net1120));
 sg13g2_tiehi \board_state_next[246]$_DFFE_PP__1121  (.L_HI(net1121));
 sg13g2_tiehi \board_state_next[247]$_DFFE_PP__1122  (.L_HI(net1122));
 sg13g2_tiehi \board_state_next[248]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \board_state_next[249]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \board_state_next[24]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \board_state_next[250]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \board_state_next[251]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \board_state_next[252]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \board_state_next[253]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \board_state_next[254]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \board_state_next[255]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \board_state_next[256]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \board_state_next[257]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \board_state_next[258]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \board_state_next[259]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \board_state_next[25]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \board_state_next[260]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \board_state_next[261]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \board_state_next[262]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \board_state_next[263]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \board_state_next[264]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \board_state_next[265]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \board_state_next[266]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \board_state_next[267]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \board_state_next[268]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \board_state_next[269]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \board_state_next[26]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \board_state_next[270]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \board_state_next[271]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \board_state_next[272]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \board_state_next[273]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \board_state_next[274]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \board_state_next[275]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \board_state_next[276]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \board_state_next[277]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \board_state_next[278]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \board_state_next[279]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \board_state_next[27]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \board_state_next[280]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \board_state_next[281]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \board_state_next[282]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \board_state_next[283]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \board_state_next[284]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \board_state_next[285]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \board_state_next[286]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \board_state_next[287]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \board_state_next[288]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \board_state_next[289]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \board_state_next[28]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \board_state_next[290]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \board_state_next[291]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \board_state_next[292]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \board_state_next[293]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \board_state_next[294]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \board_state_next[295]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \board_state_next[296]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \board_state_next[297]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \board_state_next[298]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \board_state_next[299]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \board_state_next[29]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \board_state_next[2]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \board_state_next[300]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \board_state_next[301]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \board_state_next[302]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \board_state_next[303]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \board_state_next[304]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \board_state_next[305]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \board_state_next[306]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \board_state_next[307]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \board_state_next[308]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \board_state_next[309]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \board_state_next[30]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \board_state_next[310]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \board_state_next[311]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \board_state_next[312]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \board_state_next[313]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \board_state_next[314]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \board_state_next[315]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \board_state_next[316]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \board_state_next[317]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \board_state_next[318]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \board_state_next[319]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \board_state_next[31]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \board_state_next[320]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \board_state_next[321]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \board_state_next[322]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \board_state_next[323]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \board_state_next[324]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \board_state_next[325]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \board_state_next[326]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \board_state_next[327]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \board_state_next[328]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \board_state_next[329]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \board_state_next[32]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \board_state_next[330]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \board_state_next[331]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \board_state_next[332]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \board_state_next[333]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \board_state_next[334]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \board_state_next[335]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \board_state_next[336]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \board_state_next[337]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \board_state_next[338]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \board_state_next[339]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \board_state_next[33]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \board_state_next[340]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \board_state_next[341]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \board_state_next[342]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \board_state_next[343]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \board_state_next[344]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \board_state_next[345]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \board_state_next[346]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \board_state_next[347]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \board_state_next[348]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \board_state_next[349]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \board_state_next[34]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \board_state_next[350]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \board_state_next[351]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \board_state_next[352]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \board_state_next[353]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \board_state_next[354]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \board_state_next[355]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \board_state_next[356]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \board_state_next[357]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \board_state_next[358]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \board_state_next[359]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \board_state_next[35]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \board_state_next[360]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \board_state_next[361]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \board_state_next[362]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \board_state_next[363]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \board_state_next[364]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \board_state_next[365]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \board_state_next[366]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \board_state_next[367]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \board_state_next[368]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \board_state_next[369]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \board_state_next[36]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \board_state_next[370]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \board_state_next[371]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \board_state_next[372]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \board_state_next[373]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \board_state_next[374]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \board_state_next[375]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \board_state_next[376]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \board_state_next[377]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \board_state_next[378]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \board_state_next[379]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \board_state_next[37]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \board_state_next[380]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \board_state_next[381]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \board_state_next[382]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \board_state_next[383]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \board_state_next[384]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \board_state_next[385]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \board_state_next[386]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \board_state_next[387]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \board_state_next[388]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \board_state_next[389]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \board_state_next[38]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \board_state_next[390]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \board_state_next[391]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \board_state_next[392]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \board_state_next[393]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \board_state_next[394]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \board_state_next[395]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \board_state_next[396]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \board_state_next[397]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \board_state_next[398]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \board_state_next[399]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \board_state_next[39]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \board_state_next[3]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \board_state_next[400]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \board_state_next[401]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \board_state_next[402]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \board_state_next[403]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \board_state_next[404]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \board_state_next[405]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \board_state_next[406]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \board_state_next[407]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \board_state_next[408]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \board_state_next[409]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \board_state_next[40]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \board_state_next[410]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \board_state_next[411]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \board_state_next[412]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \board_state_next[413]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \board_state_next[414]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \board_state_next[415]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \board_state_next[416]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \board_state_next[417]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \board_state_next[418]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \board_state_next[419]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \board_state_next[41]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \board_state_next[420]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \board_state_next[421]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \board_state_next[422]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \board_state_next[423]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \board_state_next[424]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \board_state_next[425]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \board_state_next[426]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \board_state_next[427]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \board_state_next[428]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \board_state_next[429]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \board_state_next[42]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \board_state_next[430]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \board_state_next[431]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \board_state_next[432]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \board_state_next[433]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \board_state_next[434]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \board_state_next[435]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \board_state_next[436]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \board_state_next[437]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \board_state_next[438]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \board_state_next[439]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \board_state_next[43]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \board_state_next[440]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \board_state_next[441]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \board_state_next[442]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \board_state_next[443]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \board_state_next[444]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \board_state_next[445]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \board_state_next[446]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \board_state_next[447]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \board_state_next[448]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \board_state_next[449]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \board_state_next[44]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \board_state_next[450]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \board_state_next[451]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \board_state_next[452]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \board_state_next[453]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \board_state_next[454]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \board_state_next[455]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \board_state_next[456]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \board_state_next[457]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \board_state_next[458]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \board_state_next[459]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \board_state_next[45]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \board_state_next[460]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \board_state_next[461]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \board_state_next[462]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \board_state_next[463]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \board_state_next[464]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \board_state_next[465]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \board_state_next[466]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \board_state_next[467]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \board_state_next[468]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \board_state_next[469]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \board_state_next[46]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \board_state_next[470]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \board_state_next[471]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \board_state_next[472]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \board_state_next[473]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \board_state_next[474]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \board_state_next[475]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \board_state_next[476]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \board_state_next[477]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \board_state_next[478]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \board_state_next[479]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \board_state_next[47]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \board_state_next[480]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \board_state_next[481]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \board_state_next[482]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \board_state_next[483]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \board_state_next[484]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \board_state_next[485]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \board_state_next[486]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \board_state_next[487]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \board_state_next[488]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \board_state_next[489]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \board_state_next[48]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \board_state_next[490]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \board_state_next[491]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \board_state_next[492]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \board_state_next[493]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \board_state_next[494]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \board_state_next[495]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \board_state_next[496]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \board_state_next[497]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \board_state_next[498]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \board_state_next[499]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \board_state_next[49]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \board_state_next[4]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \board_state_next[500]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \board_state_next[501]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \board_state_next[502]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \board_state_next[503]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \board_state_next[504]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \board_state_next[505]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \board_state_next[506]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \board_state_next[507]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \board_state_next[508]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \board_state_next[509]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \board_state_next[50]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \board_state_next[510]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \board_state_next[511]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \board_state_next[51]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \board_state_next[52]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \board_state_next[53]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \board_state_next[54]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \board_state_next[55]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \board_state_next[56]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \board_state_next[57]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \board_state_next[58]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \board_state_next[59]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \board_state_next[5]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \board_state_next[60]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \board_state_next[61]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \board_state_next[62]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \board_state_next[63]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \board_state_next[64]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \board_state_next[65]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \board_state_next[66]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \board_state_next[67]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \board_state_next[68]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \board_state_next[69]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \board_state_next[6]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \board_state_next[70]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \board_state_next[71]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \board_state_next[72]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \board_state_next[73]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \board_state_next[74]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \board_state_next[75]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \board_state_next[76]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \board_state_next[77]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \board_state_next[78]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \board_state_next[79]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \board_state_next[7]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \board_state_next[80]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \board_state_next[81]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \board_state_next[82]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \board_state_next[83]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \board_state_next[84]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \board_state_next[85]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \board_state_next[86]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \board_state_next[87]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \board_state_next[88]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \board_state_next[89]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \board_state_next[8]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \board_state_next[90]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \board_state_next[91]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \board_state_next[92]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \board_state_next[93]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \board_state_next[94]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \board_state_next[95]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \board_state_next[96]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \board_state_next[97]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \board_state_next[98]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \board_state_next[99]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \board_state_next[9]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \colindex[0]$_SDFFE_PN0P__1471  (.L_HI(net1471));
 sg13g2_tiehi \colindex[1]$_SDFFE_PN0P__1472  (.L_HI(net1472));
 sg13g2_tiehi \colindex[2]$_SDFFE_PN0P__1473  (.L_HI(net1473));
 sg13g2_tiehi \colindex[3]$_SDFFE_PN0P__1474  (.L_HI(net1474));
 sg13g2_tiehi \colindex[4]$_SDFFE_PN0P__1475  (.L_HI(net1475));
 sg13g2_tiehi \colindex[5]$_SDFFE_PN0P__1476  (.L_HI(net1476));
 sg13g2_tiehi \hvsync_inst.hpos[0]$_SDFF_PN0__1477  (.L_HI(net1477));
 sg13g2_tiehi \hvsync_inst.hpos[1]$_SDFF_PN0__1478  (.L_HI(net1478));
 sg13g2_tiehi \hvsync_inst.hpos[2]$_SDFF_PN0__1479  (.L_HI(net1479));
 sg13g2_tiehi \hvsync_inst.hpos[3]$_SDFF_PN0__1480  (.L_HI(net1480));
 sg13g2_tiehi \hvsync_inst.hpos[4]$_SDFF_PN0__1481  (.L_HI(net1481));
 sg13g2_tiehi \hvsync_inst.hpos[5]$_SDFF_PN0__1482  (.L_HI(net1482));
 sg13g2_tiehi \hvsync_inst.hpos[6]$_SDFF_PN0__1483  (.L_HI(net1483));
 sg13g2_tiehi \hvsync_inst.hpos[7]$_SDFF_PN0__1484  (.L_HI(net1484));
 sg13g2_tiehi \hvsync_inst.hpos[8]$_SDFF_PN0__1485  (.L_HI(net1485));
 sg13g2_tiehi \hvsync_inst.hpos[9]$_SDFF_PN0__1486  (.L_HI(net1486));
 sg13g2_tiehi \hvsync_inst.hsync$_DFF_P__1487  (.L_HI(net1487));
 sg13g2_tiehi \hvsync_inst.vpos[0]$_SDFFCE_PP0N__1488  (.L_HI(net1488));
 sg13g2_tiehi \hvsync_inst.vpos[1]$_SDFFCE_PP0N__1489  (.L_HI(net1489));
 sg13g2_tiehi \hvsync_inst.vpos[2]$_SDFFCE_PP0N__1490  (.L_HI(net1490));
 sg13g2_tiehi \hvsync_inst.vpos[3]$_SDFFCE_PP0N__1491  (.L_HI(net1491));
 sg13g2_tiehi \hvsync_inst.vpos[4]$_SDFFCE_PP0N__1492  (.L_HI(net1492));
 sg13g2_tiehi \hvsync_inst.vpos[5]$_SDFFCE_PP0N__1493  (.L_HI(net1493));
 sg13g2_tiehi \hvsync_inst.vpos[6]$_SDFFCE_PP0N__1494  (.L_HI(net1494));
 sg13g2_tiehi \hvsync_inst.vpos[7]$_SDFFCE_PP0N__1495  (.L_HI(net1495));
 sg13g2_tiehi \hvsync_inst.vpos[8]$_SDFFCE_PP0N__1496  (.L_HI(net1496));
 sg13g2_tiehi \hvsync_inst.vpos[9]$_SDFFCE_PP0N__1497  (.L_HI(net1497));
 sg13g2_tiehi \hvsync_inst.vsync$_DFF_P__1498  (.L_HI(net1498));
 sg13g2_tiehi \index[0]$_SDFFE_PN0P__1499  (.L_HI(net1499));
 sg13g2_tiehi \index[1]$_SDFFE_PN0P__1500  (.L_HI(net1500));
 sg13g2_tiehi \index[2]$_SDFFE_PN0P__1501  (.L_HI(net1501));
 sg13g2_tiehi \index[3]$_SDFFE_PN0P__1502  (.L_HI(net1502));
 sg13g2_tiehi \index[4]$_SDFFE_PN0P__1503  (.L_HI(net1503));
 sg13g2_tiehi \index[5]$_SDFFE_PN0P__1504  (.L_HI(net1504));
 sg13g2_tiehi \index[6]$_SDFFE_PN0P__1505  (.L_HI(net1505));
 sg13g2_tiehi \index[7]$_SDFFE_PN0P__1506  (.L_HI(net1506));
 sg13g2_tiehi \index[8]$_SDFFE_PN0P__1507  (.L_HI(net1507));
 sg13g2_tiehi \lfsr.lfsr_reg[0]$_SDFF_PN1__1508  (.L_HI(net1508));
 sg13g2_tiehi \lfsr.lfsr_reg[10]$_SDFF_PN0__1509  (.L_HI(net1509));
 sg13g2_tiehi \lfsr.lfsr_reg[11]$_SDFF_PN0__1510  (.L_HI(net1510));
 sg13g2_tiehi \lfsr.lfsr_reg[12]$_SDFF_PN0__1511  (.L_HI(net1511));
 sg13g2_tiehi \lfsr.lfsr_reg[13]$_SDFF_PN0__1512  (.L_HI(net1512));
 sg13g2_tiehi \lfsr.lfsr_reg[14]$_SDFF_PN0__1513  (.L_HI(net1513));
 sg13g2_tiehi \lfsr.lfsr_reg[15]$_SDFF_PN0__1514  (.L_HI(net1514));
 sg13g2_tiehi \lfsr.lfsr_reg[1]$_SDFF_PN0__1515  (.L_HI(net1515));
 sg13g2_tiehi \lfsr.lfsr_reg[2]$_SDFF_PN0__1516  (.L_HI(net1516));
 sg13g2_tiehi \lfsr.lfsr_reg[3]$_SDFF_PN0__1517  (.L_HI(net1517));
 sg13g2_tiehi \lfsr.lfsr_reg[4]$_SDFF_PN0__1518  (.L_HI(net1518));
 sg13g2_tiehi \lfsr.lfsr_reg[5]$_SDFF_PN0__1519  (.L_HI(net1519));
 sg13g2_tiehi \lfsr.lfsr_reg[6]$_SDFF_PN0__1520  (.L_HI(net1520));
 sg13g2_tiehi \lfsr.lfsr_reg[7]$_SDFF_PN0__1521  (.L_HI(net1521));
 sg13g2_tiehi \lfsr.lfsr_reg[8]$_SDFF_PN0__1522  (.L_HI(net1522));
 sg13g2_tiehi \lfsr.lfsr_reg[9]$_SDFF_PN0__1523  (.L_HI(net1523));
 sg13g2_tiehi \neigh_index[0]$_SDFFE_PN0P__1524  (.L_HI(net1524));
 sg13g2_tiehi \neigh_index[1]$_SDFFE_PN0P__1525  (.L_HI(net1525));
 sg13g2_tiehi \neigh_index[2]$_SDFFE_PN0P__1526  (.L_HI(net1526));
 sg13g2_tiehi \neigh_index[3]$_SDFFE_PN0P__1527  (.L_HI(net1527));
 sg13g2_tiehi \num_neighbors[0]$_SDFFE_PN0P__1528  (.L_HI(net1528));
 sg13g2_tiehi \num_neighbors[1]$_SDFFE_PN0P__1529  (.L_HI(net1529));
 sg13g2_tiehi \num_neighbors[2]$_SDFFE_PN0P__1530  (.L_HI(net1530));
 sg13g2_tiehi \num_neighbors[3]$_SDFFE_PN0P__1531  (.L_HI(net1531));
 sg13g2_tiehi \running$_SDFFE_PN0P__1532  (.L_HI(net1532));
 sg13g2_tiehi \timer[0]$_SDFFE_PN0P__1533  (.L_HI(net1533));
 sg13g2_tiehi \timer[10]$_SDFFE_PN0P__1534  (.L_HI(net1534));
 sg13g2_tiehi \timer[11]$_SDFFE_PN0P__1535  (.L_HI(net1535));
 sg13g2_tiehi \timer[12]$_SDFFE_PN0P__1536  (.L_HI(net1536));
 sg13g2_tiehi \timer[13]$_SDFFE_PN0P__1537  (.L_HI(net1537));
 sg13g2_tiehi \timer[14]$_SDFFE_PN0P__1538  (.L_HI(net1538));
 sg13g2_tiehi \timer[15]$_SDFFE_PN0P__1539  (.L_HI(net1539));
 sg13g2_tiehi \timer[16]$_SDFFE_PN0P__1540  (.L_HI(net1540));
 sg13g2_tiehi \timer[17]$_SDFFE_PN0P__1541  (.L_HI(net1541));
 sg13g2_tiehi \timer[18]$_SDFFE_PN0P__1542  (.L_HI(net1542));
 sg13g2_tiehi \timer[19]$_SDFFE_PN0P__1543  (.L_HI(net1543));
 sg13g2_tiehi \timer[1]$_SDFFE_PN0P__1544  (.L_HI(net1544));
 sg13g2_tiehi \timer[20]$_SDFFE_PN0P__1545  (.L_HI(net1545));
 sg13g2_tiehi \timer[21]$_SDFFE_PN0P__1546  (.L_HI(net1546));
 sg13g2_tiehi \timer[22]$_SDFFE_PN0P__1547  (.L_HI(net1547));
 sg13g2_tiehi \timer[23]$_SDFFE_PN0P__1548  (.L_HI(net1548));
 sg13g2_tiehi \timer[24]$_SDFFE_PN0P__1549  (.L_HI(net1549));
 sg13g2_tiehi \timer[25]$_SDFFE_PN0P__1550  (.L_HI(net1550));
 sg13g2_tiehi \timer[26]$_SDFFE_PN0P__1551  (.L_HI(net1551));
 sg13g2_tiehi \timer[27]$_SDFFE_PN0P__1552  (.L_HI(net1552));
 sg13g2_tiehi \timer[28]$_SDFFE_PN0P__1553  (.L_HI(net1553));
 sg13g2_tiehi \timer[29]$_SDFFE_PN0P__1554  (.L_HI(net1554));
 sg13g2_tiehi \timer[2]$_SDFFE_PN0P__1555  (.L_HI(net1555));
 sg13g2_tiehi \timer[30]$_SDFFE_PN0P__1556  (.L_HI(net1556));
 sg13g2_tiehi \timer[31]$_SDFFE_PN0P__1557  (.L_HI(net1557));
 sg13g2_tiehi \timer[3]$_SDFFE_PN0P__1558  (.L_HI(net1558));
 sg13g2_tiehi \timer[4]$_SDFFE_PN0P__1559  (.L_HI(net1559));
 sg13g2_tiehi \timer[5]$_SDFFE_PN0P__1560  (.L_HI(net1560));
 sg13g2_tiehi \timer[6]$_SDFFE_PN0P__1561  (.L_HI(net1561));
 sg13g2_tiehi \timer[7]$_SDFFE_PN0P__1562  (.L_HI(net1562));
 sg13g2_tiehi \timer[8]$_SDFFE_PN0P__1563  (.L_HI(net1563));
 sg13g2_tiehi \timer[9]$_SDFFE_PN0P__1564  (.L_HI(net1564));
 sg13g2_tiehi \txindex[0]$_SDFFE_PN0P__1565  (.L_HI(net1565));
 sg13g2_tiehi \txindex[1]$_SDFFE_PN0P__1566  (.L_HI(net1566));
 sg13g2_tiehi \txindex[2]$_SDFFE_PN0P__1567  (.L_HI(net1567));
 sg13g2_tiehi \txindex[3]$_SDFFE_PN0P__1568  (.L_HI(net1568));
 sg13g2_tiehi \txindex[4]$_SDFFE_PN0P__1569  (.L_HI(net1569));
 sg13g2_tiehi \txindex[5]$_SDFFE_PN0P__1570  (.L_HI(net1570));
 sg13g2_tiehi \txstate[0]$_DFF_P__1571  (.L_HI(net1571));
 sg13g2_tiehi \txstate[2]$_DFF_P__1572  (.L_HI(net1572));
 sg13g2_tiehi \txstate[3]$_DFF_P__1573  (.L_HI(net1573));
 sg13g2_tiehi \txstate[4]$_DFF_P__1574  (.L_HI(net1574));
 sg13g2_tiehi \txstate[5]$_DFF_P__1575  (.L_HI(net1575));
 sg13g2_tiehi \txstate[6]$_DFF_P__1576  (.L_HI(net1576));
 sg13g2_tiehi \txstate[7]$_DFF_P__1577  (.L_HI(net1577));
 sg13g2_tiehi \txstate[8]$_DFF_P__1578  (.L_HI(net1578));
 sg13g2_tiehi \uart_rx_inst.bitIndex[0]$_SDFFE_PN0P__1579  (.L_HI(net1579));
 sg13g2_tiehi \uart_rx_inst.bitIndex[1]$_SDFFE_PN0P__1580  (.L_HI(net1580));
 sg13g2_tiehi \uart_rx_inst.bitIndex[2]$_SDFFE_PN0P__1581  (.L_HI(net1581));
 sg13g2_tiehi \uart_rx_inst.data[0]$_SDFFE_PN0P__1582  (.L_HI(net1582));
 sg13g2_tiehi \uart_rx_inst.data[1]$_SDFFE_PN0P__1583  (.L_HI(net1583));
 sg13g2_tiehi \uart_rx_inst.data[2]$_SDFFE_PN0P__1584  (.L_HI(net1584));
 sg13g2_tiehi \uart_rx_inst.data[3]$_SDFFE_PN0P__1585  (.L_HI(net1585));
 sg13g2_tiehi \uart_rx_inst.data[4]$_SDFFE_PN0P__1586  (.L_HI(net1586));
 sg13g2_tiehi \uart_rx_inst.data[5]$_SDFFE_PN0P__1587  (.L_HI(net1587));
 sg13g2_tiehi \uart_rx_inst.data[6]$_SDFFE_PN0P__1588  (.L_HI(net1588));
 sg13g2_tiehi \uart_rx_inst.data[7]$_SDFFE_PN0P__1589  (.L_HI(net1589));
 sg13g2_tiehi \uart_rx_inst.inputReg[0]$_SDFFE_PN1P__1590  (.L_HI(net1590));
 sg13g2_tiehi \uart_rx_inst.inputReg[1]$_SDFFE_PN1P__1591  (.L_HI(net1591));
 sg13g2_tiehi \uart_rx_inst.inputReg[2]$_SDFFE_PN1P__1592  (.L_HI(net1592));
 sg13g2_tiehi \uart_rx_inst.out[0]$_SDFFE_PN0P__1593  (.L_HI(net1593));
 sg13g2_tiehi \uart_rx_inst.out[1]$_SDFFE_PN0P__1594  (.L_HI(net1594));
 sg13g2_tiehi \uart_rx_inst.out[2]$_SDFFE_PN0P__1595  (.L_HI(net1595));
 sg13g2_tiehi \uart_rx_inst.out[3]$_SDFFE_PN0P__1596  (.L_HI(net1596));
 sg13g2_tiehi \uart_rx_inst.out[4]$_SDFFE_PN0P__1597  (.L_HI(net1597));
 sg13g2_tiehi \uart_rx_inst.out[5]$_SDFFE_PN0P__1598  (.L_HI(net1598));
 sg13g2_tiehi \uart_rx_inst.out[6]$_SDFFE_PN0P__1599  (.L_HI(net1599));
 sg13g2_tiehi \uart_rx_inst.out[7]$_SDFFE_PN0P__1600  (.L_HI(net1600));
 sg13g2_tiehi \uart_rx_inst.out_latched$_SDFFE_PP0P__1601  (.L_HI(net1601));
 sg13g2_tiehi \uart_rx_inst.rxCounter[0]$_SDFF_PN0__1602  (.L_HI(net1602));
 sg13g2_tiehi \uart_rx_inst.rxCounter[1]$_SDFF_PN0__1603  (.L_HI(net1603));
 sg13g2_tiehi \uart_rx_inst.rxCounter[2]$_SDFF_PN0__1604  (.L_HI(net1604));
 sg13g2_tiehi \uart_rx_inst.rxCounter[3]$_SDFF_PN0__1605  (.L_HI(net1605));
 sg13g2_tiehi \uart_rx_inst.sampleCount[0]$_SDFFE_PN0P__1606  (.L_HI(net1606));
 sg13g2_tiehi \uart_rx_inst.sampleCount[1]$_SDFFE_PN0P__1607  (.L_HI(net1607));
 sg13g2_tiehi \uart_rx_inst.sampleCount[2]$_SDFFE_PN0P__1608  (.L_HI(net1608));
 sg13g2_tiehi \uart_rx_inst.sampleCount[3]$_SDFFE_PN0P__1609  (.L_HI(net1609));
 sg13g2_tiehi \uart_rx_inst.state[0]$_DFF_P__1610  (.L_HI(net1610));
 sg13g2_tiehi \uart_rx_inst.state[1]$_DFF_P__1611  (.L_HI(net1611));
 sg13g2_tiehi \uart_rx_inst.state[2]$_DFF_P__1612  (.L_HI(net1612));
 sg13g2_tiehi \uart_rx_inst.state[3]$_DFF_P__1613  (.L_HI(net1613));
 sg13g2_tiehi \uart_rx_inst.valid$_SDFFE_PN0P__1614  (.L_HI(net1614));
 sg13g2_tiehi \uart_rx_ready$_SDFFE_PN0P__1615  (.L_HI(net1615));
 sg13g2_tiehi \uart_tx_data[0]$_SDFFE_PN0P__1616  (.L_HI(net1616));
 sg13g2_tiehi \uart_tx_data[1]$_SDFFE_PN0P__1617  (.L_HI(net1617));
 sg13g2_tiehi \uart_tx_data[2]$_SDFFE_PN0P__1618  (.L_HI(net1618));
 sg13g2_tiehi \uart_tx_data[3]$_SDFFE_PN0P__1619  (.L_HI(net1619));
 sg13g2_tiehi \uart_tx_data[4]$_SDFFE_PN0P__1620  (.L_HI(net1620));
 sg13g2_tiehi \uart_tx_data[5]$_SDFFE_PN0P__1621  (.L_HI(net1621));
 sg13g2_tiehi \uart_tx_data[6]$_SDFFE_PN0P__1622  (.L_HI(net1622));
 sg13g2_tiehi \uart_tx_inst.bitIndex[0]$_SDFFE_PN0P__1623  (.L_HI(net1623));
 sg13g2_tiehi \uart_tx_inst.bitIndex[1]$_SDFFE_PN0P__1624  (.L_HI(net1624));
 sg13g2_tiehi \uart_tx_inst.bitIndex[2]$_SDFFE_PN0P__1625  (.L_HI(net1625));
 sg13g2_tiehi \uart_tx_inst.data[0]$_SDFFE_PN0P__1626  (.L_HI(net1626));
 sg13g2_tiehi \uart_tx_inst.data[1]$_SDFFE_PN0P__1627  (.L_HI(net1627));
 sg13g2_tiehi \uart_tx_inst.data[2]$_SDFFE_PN0P__1628  (.L_HI(net1628));
 sg13g2_tiehi \uart_tx_inst.data[3]$_SDFFE_PN0P__1629  (.L_HI(net1629));
 sg13g2_tiehi \uart_tx_inst.data[4]$_SDFFE_PN0P__1630  (.L_HI(net1630));
 sg13g2_tiehi \uart_tx_inst.data[5]$_SDFFE_PN0P__1631  (.L_HI(net1631));
 sg13g2_tiehi \uart_tx_inst.data[6]$_SDFFE_PN0P__1632  (.L_HI(net1632));
 sg13g2_tiehi \uart_tx_inst.out$_SDFFE_PN1P__1633  (.L_HI(net1633));
 sg13g2_tiehi \uart_tx_inst.ready$_SDFFE_PP0P__1634  (.L_HI(net1634));
 sg13g2_tiehi \uart_tx_inst.state[0]$_DFF_P__1635  (.L_HI(net1635));
 sg13g2_tiehi \uart_tx_inst.state[1]$_DFF_P__1636  (.L_HI(net1636));
 sg13g2_tiehi \uart_tx_inst.state[2]$_DFF_P__1637  (.L_HI(net1637));
 sg13g2_tiehi \uart_tx_inst.state[3]$_DFF_P__1638  (.L_HI(net1638));
 sg13g2_tiehi \uart_tx_inst.txCounter[0]$_SDFFE_PN0N__1639  (.L_HI(net1639));
 sg13g2_tiehi \uart_tx_inst.txCounter[1]$_SDFFE_PN0N__1640  (.L_HI(net1640));
 sg13g2_tiehi \uart_tx_inst.txCounter[2]$_SDFFE_PN0N__1641  (.L_HI(net1641));
 sg13g2_tiehi \uart_tx_inst.txCounter[3]$_SDFFE_PN0N__1642  (.L_HI(net1642));
 sg13g2_tiehi \uart_tx_inst.txCounter[4]$_SDFFE_PN0N__1643  (.L_HI(net1643));
 sg13g2_tiehi \uart_tx_inst.txCounter[5]$_SDFFE_PN0N__1644  (.L_HI(net1644));
 sg13g2_tiehi \uart_tx_inst.txCounter[6]$_SDFFE_PN0N__1645  (.L_HI(net1645));
 sg13g2_tiehi \uart_tx_inst.txCounter[7]$_SDFFE_PN0N__1646  (.L_HI(net1646));
 sg13g2_tiehi \uart_tx_valid$_SDFFE_PN0P__1647  (.L_HI(net1647));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_62_clk (.X(clknet_leaf_62_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_63_clk (.X(clknet_leaf_63_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_64_clk (.X(clknet_leaf_64_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_65_clk (.X(clknet_leaf_65_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_66_clk (.X(clknet_leaf_66_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_67_clk (.X(clknet_leaf_67_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_68_clk (.X(clknet_leaf_68_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_69_clk (.X(clknet_leaf_69_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_70_clk (.X(clknet_leaf_70_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_71_clk (.X(clknet_leaf_71_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_72_clk (.X(clknet_leaf_72_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_73_clk (.X(clknet_leaf_73_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_74_clk (.X(clknet_leaf_74_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_75_clk (.X(clknet_leaf_75_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_76_clk (.X(clknet_leaf_76_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_77_clk (.X(clknet_leaf_77_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_78_clk (.X(clknet_leaf_78_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_79_clk (.X(clknet_leaf_79_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_80_clk (.X(clknet_leaf_80_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_81_clk (.X(clknet_leaf_81_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_82_clk (.X(clknet_leaf_82_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_83_clk (.X(clknet_leaf_83_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_84_clk (.X(clknet_leaf_84_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_85_clk (.X(clknet_leaf_85_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_86_clk (.X(clknet_leaf_86_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_87_clk (.X(clknet_leaf_87_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_88_clk (.X(clknet_leaf_88_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_89_clk (.X(clknet_leaf_89_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_90_clk (.X(clknet_leaf_90_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_91_clk (.X(clknet_leaf_91_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_92_clk (.X(clknet_leaf_92_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_93_clk (.X(clknet_leaf_93_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_94_clk (.X(clknet_leaf_94_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_95_clk (.X(clknet_leaf_95_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_96_clk (.X(clknet_leaf_96_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_97_clk (.X(clknet_leaf_97_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_98_clk (.X(clknet_leaf_98_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_99_clk (.X(clknet_leaf_99_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_100_clk (.X(clknet_leaf_100_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_101_clk (.X(clknet_leaf_101_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_102_clk (.X(clknet_leaf_102_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_103_clk (.X(clknet_leaf_103_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_104_clk (.X(clknet_leaf_104_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_105_clk (.X(clknet_leaf_105_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_106_clk (.X(clknet_leaf_106_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_107_clk (.X(clknet_leaf_107_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_108_clk (.X(clknet_leaf_108_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_109_clk (.X(clknet_leaf_109_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_110_clk (.X(clknet_leaf_110_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_111_clk (.X(clknet_leaf_111_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_112_clk (.X(clknet_leaf_112_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_113_clk (.X(clknet_leaf_113_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_114_clk (.X(clknet_leaf_114_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_115_clk (.X(clknet_leaf_115_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_116_clk (.X(clknet_leaf_116_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_117_clk (.X(clknet_leaf_117_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_118_clk (.X(clknet_leaf_118_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_119_clk (.X(clknet_leaf_119_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_120_clk (.X(clknet_leaf_120_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_121_clk (.X(clknet_leaf_121_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_122_clk (.X(clknet_leaf_122_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_123_clk (.X(clknet_leaf_123_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_124_clk (.X(clknet_leaf_124_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_125_clk (.X(clknet_leaf_125_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_126_clk (.X(clknet_leaf_126_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_127_clk (.X(clknet_leaf_127_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_128_clk (.X(clknet_leaf_128_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_129_clk (.X(clknet_leaf_129_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_130_clk (.X(clknet_leaf_130_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_131_clk (.X(clknet_leaf_131_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_132_clk (.X(clknet_leaf_132_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_133_clk (.X(clknet_leaf_133_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_134_clk (.X(clknet_leaf_134_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_135_clk (.X(clknet_leaf_135_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_136_clk (.X(clknet_leaf_136_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_137_clk (.X(clknet_leaf_137_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_138_clk (.X(clknet_leaf_138_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_139_clk (.X(clknet_leaf_139_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_140_clk (.X(clknet_leaf_140_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_141_clk (.X(clknet_leaf_141_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_142_clk (.X(clknet_leaf_142_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_143_clk (.X(clknet_leaf_143_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_144_clk (.X(clknet_leaf_144_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_145_clk (.X(clknet_leaf_145_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_146_clk (.X(clknet_leaf_146_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_147_clk (.X(clknet_leaf_147_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_148_clk (.X(clknet_leaf_148_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_149_clk (.X(clknet_leaf_149_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_150_clk (.X(clknet_leaf_150_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_151_clk (.X(clknet_leaf_151_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_152_clk (.X(clknet_leaf_152_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_153_clk (.X(clknet_leaf_153_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_154_clk (.X(clknet_leaf_154_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_155_clk (.X(clknet_leaf_155_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_156_clk (.X(clknet_leaf_156_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_157_clk (.X(clknet_leaf_157_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_153_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_leaf_157_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_11_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_leaf_140_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_25_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_36_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_45_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_46_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_49_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_50_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_38_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_44_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_124_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_51_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_52_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_83_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_86_clk));
 sg13g2_buf_8 clkload21 (.A(clknet_leaf_63_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0045_));
 sg13g2_antennanp ANTENNA_2 (.A(_3389_));
 sg13g2_antennanp ANTENNA_3 (.A(_4150_));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(net11));
 sg13g2_antennanp ANTENNA_6 (.A(net11));
 sg13g2_antennanp ANTENNA_7 (.A(_0045_));
 sg13g2_antennanp ANTENNA_8 (.A(_4150_));
 sg13g2_antennanp ANTENNA_9 (.A(clk));
 sg13g2_antennanp ANTENNA_10 (.A(net11));
 sg13g2_antennanp ANTENNA_11 (.A(net11));
 sg13g2_antennanp ANTENNA_12 (.A(_0045_));
 sg13g2_antennanp ANTENNA_13 (.A(_4150_));
 sg13g2_antennanp ANTENNA_14 (.A(clk));
 sg13g2_antennanp ANTENNA_15 (.A(net11));
 sg13g2_antennanp ANTENNA_16 (.A(net11));
 sg13g2_antennanp ANTENNA_17 (.A(_4150_));
 sg13g2_antennanp ANTENNA_18 (.A(clk));
 sg13g2_antennanp ANTENNA_19 (.A(net11));
 sg13g2_antennanp ANTENNA_20 (.A(net11));
 sg13g2_antennanp ANTENNA_21 (.A(_4150_));
 sg13g2_antennanp ANTENNA_22 (.A(clk));
 sg13g2_antennanp ANTENNA_23 (.A(net11));
 sg13g2_antennanp ANTENNA_24 (.A(net11));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_4 FILLER_0_182 ();
 sg13g2_fill_2 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_4 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_fill_1 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_decap_8 FILLER_0_240 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_4 FILLER_0_261 ();
 sg13g2_fill_2 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_fill_2 FILLER_0_313 ();
 sg13g2_fill_1 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_4 FILLER_0_348 ();
 sg13g2_fill_1 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_4 FILLER_0_378 ();
 sg13g2_fill_1 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_fill_2 FILLER_0_400 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_fill_1 FILLER_0_420 ();
 sg13g2_fill_1 FILLER_0_425 ();
 sg13g2_decap_8 FILLER_0_430 ();
 sg13g2_decap_8 FILLER_0_437 ();
 sg13g2_decap_8 FILLER_0_444 ();
 sg13g2_decap_4 FILLER_0_451 ();
 sg13g2_decap_8 FILLER_0_465 ();
 sg13g2_decap_8 FILLER_0_472 ();
 sg13g2_decap_4 FILLER_0_479 ();
 sg13g2_decap_8 FILLER_0_517 ();
 sg13g2_decap_8 FILLER_0_524 ();
 sg13g2_decap_8 FILLER_0_531 ();
 sg13g2_decap_8 FILLER_0_538 ();
 sg13g2_decap_8 FILLER_0_545 ();
 sg13g2_decap_4 FILLER_0_556 ();
 sg13g2_decap_8 FILLER_0_564 ();
 sg13g2_decap_8 FILLER_0_571 ();
 sg13g2_decap_8 FILLER_0_578 ();
 sg13g2_decap_8 FILLER_0_593 ();
 sg13g2_decap_8 FILLER_0_600 ();
 sg13g2_decap_8 FILLER_0_607 ();
 sg13g2_decap_8 FILLER_0_614 ();
 sg13g2_decap_8 FILLER_0_631 ();
 sg13g2_decap_8 FILLER_0_638 ();
 sg13g2_fill_2 FILLER_0_645 ();
 sg13g2_fill_1 FILLER_0_647 ();
 sg13g2_decap_8 FILLER_0_652 ();
 sg13g2_decap_8 FILLER_0_659 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_8 FILLER_0_673 ();
 sg13g2_decap_8 FILLER_0_680 ();
 sg13g2_decap_8 FILLER_0_687 ();
 sg13g2_decap_8 FILLER_0_694 ();
 sg13g2_decap_8 FILLER_0_701 ();
 sg13g2_decap_8 FILLER_0_708 ();
 sg13g2_decap_8 FILLER_0_715 ();
 sg13g2_decap_8 FILLER_0_722 ();
 sg13g2_decap_8 FILLER_0_729 ();
 sg13g2_decap_8 FILLER_0_736 ();
 sg13g2_decap_8 FILLER_0_743 ();
 sg13g2_decap_8 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_757 ();
 sg13g2_decap_8 FILLER_0_764 ();
 sg13g2_decap_8 FILLER_0_771 ();
 sg13g2_decap_8 FILLER_0_778 ();
 sg13g2_decap_8 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_decap_8 FILLER_0_799 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_8 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_820 ();
 sg13g2_decap_8 FILLER_0_827 ();
 sg13g2_decap_8 FILLER_0_834 ();
 sg13g2_decap_8 FILLER_0_841 ();
 sg13g2_decap_8 FILLER_0_848 ();
 sg13g2_decap_8 FILLER_0_855 ();
 sg13g2_decap_8 FILLER_0_862 ();
 sg13g2_decap_8 FILLER_0_869 ();
 sg13g2_decap_8 FILLER_0_876 ();
 sg13g2_decap_8 FILLER_0_883 ();
 sg13g2_decap_8 FILLER_0_890 ();
 sg13g2_decap_8 FILLER_0_897 ();
 sg13g2_decap_8 FILLER_0_904 ();
 sg13g2_decap_8 FILLER_0_911 ();
 sg13g2_decap_8 FILLER_0_918 ();
 sg13g2_decap_8 FILLER_0_925 ();
 sg13g2_decap_8 FILLER_0_932 ();
 sg13g2_decap_8 FILLER_0_939 ();
 sg13g2_decap_4 FILLER_0_946 ();
 sg13g2_fill_2 FILLER_0_950 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_986 ();
 sg13g2_decap_8 FILLER_0_993 ();
 sg13g2_decap_8 FILLER_0_1000 ();
 sg13g2_decap_8 FILLER_0_1007 ();
 sg13g2_decap_8 FILLER_0_1014 ();
 sg13g2_decap_8 FILLER_0_1021 ();
 sg13g2_decap_8 FILLER_0_1028 ();
 sg13g2_decap_8 FILLER_0_1035 ();
 sg13g2_decap_8 FILLER_0_1042 ();
 sg13g2_decap_8 FILLER_0_1049 ();
 sg13g2_decap_4 FILLER_0_1056 ();
 sg13g2_fill_2 FILLER_0_1060 ();
 sg13g2_decap_8 FILLER_0_1066 ();
 sg13g2_decap_8 FILLER_0_1073 ();
 sg13g2_fill_1 FILLER_0_1080 ();
 sg13g2_decap_8 FILLER_0_1111 ();
 sg13g2_decap_8 FILLER_0_1118 ();
 sg13g2_decap_8 FILLER_0_1125 ();
 sg13g2_decap_8 FILLER_0_1132 ();
 sg13g2_fill_1 FILLER_0_1139 ();
 sg13g2_decap_4 FILLER_0_1144 ();
 sg13g2_fill_2 FILLER_0_1148 ();
 sg13g2_decap_8 FILLER_0_1160 ();
 sg13g2_fill_1 FILLER_0_1167 ();
 sg13g2_decap_8 FILLER_0_1198 ();
 sg13g2_decap_8 FILLER_0_1205 ();
 sg13g2_decap_8 FILLER_0_1212 ();
 sg13g2_decap_8 FILLER_0_1219 ();
 sg13g2_decap_8 FILLER_0_1226 ();
 sg13g2_decap_8 FILLER_0_1233 ();
 sg13g2_decap_8 FILLER_0_1240 ();
 sg13g2_decap_8 FILLER_0_1247 ();
 sg13g2_decap_8 FILLER_0_1254 ();
 sg13g2_decap_8 FILLER_0_1261 ();
 sg13g2_decap_8 FILLER_0_1268 ();
 sg13g2_decap_8 FILLER_0_1275 ();
 sg13g2_decap_8 FILLER_0_1282 ();
 sg13g2_decap_8 FILLER_0_1289 ();
 sg13g2_decap_8 FILLER_0_1296 ();
 sg13g2_decap_8 FILLER_0_1303 ();
 sg13g2_decap_8 FILLER_0_1310 ();
 sg13g2_decap_8 FILLER_0_1317 ();
 sg13g2_fill_2 FILLER_0_1324 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_fill_2 FILLER_1_56 ();
 sg13g2_fill_1 FILLER_1_58 ();
 sg13g2_decap_8 FILLER_1_85 ();
 sg13g2_decap_8 FILLER_1_92 ();
 sg13g2_decap_8 FILLER_1_99 ();
 sg13g2_decap_4 FILLER_1_106 ();
 sg13g2_fill_1 FILLER_1_110 ();
 sg13g2_decap_8 FILLER_1_157 ();
 sg13g2_decap_8 FILLER_1_164 ();
 sg13g2_decap_8 FILLER_1_171 ();
 sg13g2_fill_1 FILLER_1_178 ();
 sg13g2_fill_2 FILLER_1_205 ();
 sg13g2_fill_1 FILLER_1_207 ();
 sg13g2_decap_8 FILLER_1_248 ();
 sg13g2_fill_1 FILLER_1_255 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_fill_2 FILLER_1_420 ();
 sg13g2_fill_1 FILLER_1_422 ();
 sg13g2_fill_1 FILLER_1_457 ();
 sg13g2_fill_2 FILLER_1_462 ();
 sg13g2_fill_2 FILLER_1_526 ();
 sg13g2_fill_1 FILLER_1_528 ();
 sg13g2_decap_4 FILLER_1_533 ();
 sg13g2_fill_2 FILLER_1_537 ();
 sg13g2_fill_2 FILLER_1_543 ();
 sg13g2_fill_1 FILLER_1_571 ();
 sg13g2_fill_2 FILLER_1_576 ();
 sg13g2_fill_1 FILLER_1_578 ();
 sg13g2_fill_1 FILLER_1_605 ();
 sg13g2_fill_1 FILLER_1_620 ();
 sg13g2_decap_8 FILLER_1_625 ();
 sg13g2_fill_1 FILLER_1_632 ();
 sg13g2_decap_8 FILLER_1_669 ();
 sg13g2_decap_8 FILLER_1_676 ();
 sg13g2_decap_8 FILLER_1_683 ();
 sg13g2_decap_8 FILLER_1_690 ();
 sg13g2_decap_8 FILLER_1_697 ();
 sg13g2_decap_8 FILLER_1_704 ();
 sg13g2_decap_8 FILLER_1_711 ();
 sg13g2_decap_8 FILLER_1_718 ();
 sg13g2_decap_8 FILLER_1_725 ();
 sg13g2_decap_8 FILLER_1_732 ();
 sg13g2_decap_8 FILLER_1_739 ();
 sg13g2_decap_8 FILLER_1_746 ();
 sg13g2_decap_8 FILLER_1_753 ();
 sg13g2_decap_8 FILLER_1_760 ();
 sg13g2_decap_8 FILLER_1_767 ();
 sg13g2_decap_8 FILLER_1_774 ();
 sg13g2_decap_8 FILLER_1_781 ();
 sg13g2_decap_8 FILLER_1_788 ();
 sg13g2_decap_8 FILLER_1_795 ();
 sg13g2_decap_8 FILLER_1_802 ();
 sg13g2_decap_8 FILLER_1_809 ();
 sg13g2_decap_8 FILLER_1_816 ();
 sg13g2_fill_2 FILLER_1_823 ();
 sg13g2_fill_1 FILLER_1_855 ();
 sg13g2_decap_8 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_1_867 ();
 sg13g2_decap_8 FILLER_1_874 ();
 sg13g2_decap_8 FILLER_1_881 ();
 sg13g2_decap_8 FILLER_1_888 ();
 sg13g2_decap_8 FILLER_1_895 ();
 sg13g2_decap_8 FILLER_1_902 ();
 sg13g2_decap_8 FILLER_1_909 ();
 sg13g2_decap_8 FILLER_1_916 ();
 sg13g2_decap_8 FILLER_1_923 ();
 sg13g2_fill_2 FILLER_1_930 ();
 sg13g2_fill_1 FILLER_1_932 ();
 sg13g2_fill_1 FILLER_1_967 ();
 sg13g2_decap_8 FILLER_1_998 ();
 sg13g2_decap_8 FILLER_1_1005 ();
 sg13g2_decap_8 FILLER_1_1012 ();
 sg13g2_decap_8 FILLER_1_1019 ();
 sg13g2_decap_8 FILLER_1_1026 ();
 sg13g2_decap_8 FILLER_1_1033 ();
 sg13g2_fill_1 FILLER_1_1040 ();
 sg13g2_decap_4 FILLER_1_1085 ();
 sg13g2_fill_1 FILLER_1_1089 ();
 sg13g2_decap_8 FILLER_1_1104 ();
 sg13g2_fill_2 FILLER_1_1111 ();
 sg13g2_decap_4 FILLER_1_1123 ();
 sg13g2_fill_2 FILLER_1_1127 ();
 sg13g2_decap_4 FILLER_1_1159 ();
 sg13g2_fill_2 FILLER_1_1163 ();
 sg13g2_decap_8 FILLER_1_1191 ();
 sg13g2_decap_8 FILLER_1_1208 ();
 sg13g2_decap_8 FILLER_1_1215 ();
 sg13g2_decap_8 FILLER_1_1222 ();
 sg13g2_decap_8 FILLER_1_1229 ();
 sg13g2_decap_8 FILLER_1_1236 ();
 sg13g2_decap_8 FILLER_1_1243 ();
 sg13g2_decap_8 FILLER_1_1250 ();
 sg13g2_decap_8 FILLER_1_1257 ();
 sg13g2_decap_8 FILLER_1_1264 ();
 sg13g2_decap_8 FILLER_1_1271 ();
 sg13g2_decap_8 FILLER_1_1278 ();
 sg13g2_decap_8 FILLER_1_1285 ();
 sg13g2_decap_8 FILLER_1_1292 ();
 sg13g2_decap_8 FILLER_1_1299 ();
 sg13g2_decap_8 FILLER_1_1306 ();
 sg13g2_decap_8 FILLER_1_1313 ();
 sg13g2_decap_4 FILLER_1_1320 ();
 sg13g2_fill_2 FILLER_1_1324 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_fill_2 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_92 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_4 FILLER_2_172 ();
 sg13g2_fill_2 FILLER_2_176 ();
 sg13g2_fill_2 FILLER_2_250 ();
 sg13g2_fill_2 FILLER_2_256 ();
 sg13g2_fill_1 FILLER_2_294 ();
 sg13g2_fill_1 FILLER_2_335 ();
 sg13g2_fill_2 FILLER_2_372 ();
 sg13g2_fill_1 FILLER_2_374 ();
 sg13g2_fill_1 FILLER_2_421 ();
 sg13g2_fill_1 FILLER_2_458 ();
 sg13g2_decap_4 FILLER_2_495 ();
 sg13g2_fill_1 FILLER_2_499 ();
 sg13g2_decap_4 FILLER_2_504 ();
 sg13g2_fill_1 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_513 ();
 sg13g2_decap_4 FILLER_2_520 ();
 sg13g2_fill_2 FILLER_2_570 ();
 sg13g2_fill_2 FILLER_2_608 ();
 sg13g2_fill_1 FILLER_2_610 ();
 sg13g2_decap_8 FILLER_2_675 ();
 sg13g2_decap_8 FILLER_2_682 ();
 sg13g2_decap_8 FILLER_2_689 ();
 sg13g2_decap_8 FILLER_2_696 ();
 sg13g2_decap_8 FILLER_2_703 ();
 sg13g2_decap_8 FILLER_2_710 ();
 sg13g2_decap_8 FILLER_2_717 ();
 sg13g2_decap_8 FILLER_2_724 ();
 sg13g2_decap_8 FILLER_2_731 ();
 sg13g2_decap_8 FILLER_2_738 ();
 sg13g2_decap_8 FILLER_2_745 ();
 sg13g2_decap_8 FILLER_2_752 ();
 sg13g2_decap_8 FILLER_2_759 ();
 sg13g2_decap_8 FILLER_2_766 ();
 sg13g2_decap_8 FILLER_2_773 ();
 sg13g2_decap_8 FILLER_2_780 ();
 sg13g2_decap_8 FILLER_2_787 ();
 sg13g2_decap_8 FILLER_2_794 ();
 sg13g2_decap_8 FILLER_2_801 ();
 sg13g2_decap_8 FILLER_2_808 ();
 sg13g2_decap_8 FILLER_2_815 ();
 sg13g2_decap_8 FILLER_2_822 ();
 sg13g2_fill_2 FILLER_2_829 ();
 sg13g2_fill_1 FILLER_2_831 ();
 sg13g2_decap_8 FILLER_2_842 ();
 sg13g2_fill_1 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_880 ();
 sg13g2_decap_8 FILLER_2_887 ();
 sg13g2_decap_8 FILLER_2_894 ();
 sg13g2_decap_8 FILLER_2_901 ();
 sg13g2_decap_8 FILLER_2_908 ();
 sg13g2_decap_8 FILLER_2_915 ();
 sg13g2_decap_4 FILLER_2_922 ();
 sg13g2_decap_8 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1015 ();
 sg13g2_decap_8 FILLER_2_1022 ();
 sg13g2_decap_8 FILLER_2_1029 ();
 sg13g2_decap_8 FILLER_2_1036 ();
 sg13g2_fill_2 FILLER_2_1043 ();
 sg13g2_fill_2 FILLER_2_1179 ();
 sg13g2_decap_8 FILLER_2_1233 ();
 sg13g2_decap_8 FILLER_2_1240 ();
 sg13g2_decap_8 FILLER_2_1247 ();
 sg13g2_decap_8 FILLER_2_1254 ();
 sg13g2_decap_8 FILLER_2_1261 ();
 sg13g2_decap_8 FILLER_2_1268 ();
 sg13g2_decap_8 FILLER_2_1275 ();
 sg13g2_decap_8 FILLER_2_1282 ();
 sg13g2_decap_8 FILLER_2_1289 ();
 sg13g2_decap_8 FILLER_2_1296 ();
 sg13g2_decap_8 FILLER_2_1303 ();
 sg13g2_decap_8 FILLER_2_1310 ();
 sg13g2_decap_8 FILLER_2_1317 ();
 sg13g2_fill_2 FILLER_2_1324 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_4 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_fill_2 FILLER_3_91 ();
 sg13g2_fill_2 FILLER_3_101 ();
 sg13g2_fill_1 FILLER_3_103 ();
 sg13g2_fill_1 FILLER_3_138 ();
 sg13g2_decap_8 FILLER_3_164 ();
 sg13g2_decap_4 FILLER_3_171 ();
 sg13g2_fill_1 FILLER_3_175 ();
 sg13g2_decap_4 FILLER_3_190 ();
 sg13g2_fill_1 FILLER_3_194 ();
 sg13g2_fill_2 FILLER_3_256 ();
 sg13g2_fill_1 FILLER_3_258 ();
 sg13g2_fill_2 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_325 ();
 sg13g2_decap_4 FILLER_3_332 ();
 sg13g2_fill_1 FILLER_3_370 ();
 sg13g2_fill_1 FILLER_3_375 ();
 sg13g2_fill_1 FILLER_3_397 ();
 sg13g2_fill_1 FILLER_3_402 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_fill_1 FILLER_3_469 ();
 sg13g2_fill_2 FILLER_3_474 ();
 sg13g2_fill_2 FILLER_3_480 ();
 sg13g2_fill_2 FILLER_3_492 ();
 sg13g2_decap_8 FILLER_3_515 ();
 sg13g2_fill_1 FILLER_3_522 ();
 sg13g2_fill_2 FILLER_3_569 ();
 sg13g2_fill_1 FILLER_3_585 ();
 sg13g2_fill_2 FILLER_3_607 ();
 sg13g2_fill_1 FILLER_3_609 ();
 sg13g2_fill_2 FILLER_3_618 ();
 sg13g2_fill_1 FILLER_3_620 ();
 sg13g2_decap_8 FILLER_3_668 ();
 sg13g2_decap_8 FILLER_3_675 ();
 sg13g2_decap_8 FILLER_3_682 ();
 sg13g2_decap_8 FILLER_3_689 ();
 sg13g2_decap_8 FILLER_3_696 ();
 sg13g2_decap_8 FILLER_3_703 ();
 sg13g2_decap_8 FILLER_3_710 ();
 sg13g2_decap_8 FILLER_3_717 ();
 sg13g2_decap_8 FILLER_3_724 ();
 sg13g2_decap_8 FILLER_3_731 ();
 sg13g2_decap_8 FILLER_3_738 ();
 sg13g2_decap_8 FILLER_3_745 ();
 sg13g2_decap_8 FILLER_3_752 ();
 sg13g2_decap_8 FILLER_3_759 ();
 sg13g2_decap_8 FILLER_3_766 ();
 sg13g2_decap_8 FILLER_3_773 ();
 sg13g2_decap_8 FILLER_3_780 ();
 sg13g2_decap_8 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_794 ();
 sg13g2_decap_8 FILLER_3_801 ();
 sg13g2_decap_4 FILLER_3_808 ();
 sg13g2_fill_1 FILLER_3_812 ();
 sg13g2_fill_2 FILLER_3_863 ();
 sg13g2_fill_1 FILLER_3_865 ();
 sg13g2_decap_8 FILLER_3_892 ();
 sg13g2_decap_8 FILLER_3_899 ();
 sg13g2_decap_8 FILLER_3_906 ();
 sg13g2_decap_4 FILLER_3_913 ();
 sg13g2_fill_1 FILLER_3_917 ();
 sg13g2_fill_2 FILLER_3_967 ();
 sg13g2_decap_8 FILLER_3_1005 ();
 sg13g2_decap_8 FILLER_3_1012 ();
 sg13g2_decap_8 FILLER_3_1019 ();
 sg13g2_decap_8 FILLER_3_1026 ();
 sg13g2_decap_8 FILLER_3_1033 ();
 sg13g2_fill_1 FILLER_3_1086 ();
 sg13g2_fill_2 FILLER_3_1175 ();
 sg13g2_fill_2 FILLER_3_1187 ();
 sg13g2_fill_1 FILLER_3_1189 ();
 sg13g2_fill_2 FILLER_3_1194 ();
 sg13g2_fill_1 FILLER_3_1196 ();
 sg13g2_decap_8 FILLER_3_1219 ();
 sg13g2_decap_8 FILLER_3_1226 ();
 sg13g2_decap_8 FILLER_3_1233 ();
 sg13g2_decap_8 FILLER_3_1240 ();
 sg13g2_decap_8 FILLER_3_1247 ();
 sg13g2_decap_8 FILLER_3_1254 ();
 sg13g2_decap_8 FILLER_3_1261 ();
 sg13g2_decap_8 FILLER_3_1268 ();
 sg13g2_decap_8 FILLER_3_1275 ();
 sg13g2_decap_8 FILLER_3_1282 ();
 sg13g2_decap_8 FILLER_3_1289 ();
 sg13g2_decap_8 FILLER_3_1296 ();
 sg13g2_decap_8 FILLER_3_1303 ();
 sg13g2_decap_8 FILLER_3_1310 ();
 sg13g2_decap_8 FILLER_3_1317 ();
 sg13g2_fill_2 FILLER_3_1324 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_4 FILLER_4_35 ();
 sg13g2_fill_2 FILLER_4_39 ();
 sg13g2_decap_4 FILLER_4_55 ();
 sg13g2_fill_2 FILLER_4_59 ();
 sg13g2_fill_2 FILLER_4_65 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_decap_4 FILLER_4_95 ();
 sg13g2_fill_2 FILLER_4_103 ();
 sg13g2_fill_1 FILLER_4_105 ();
 sg13g2_decap_4 FILLER_4_128 ();
 sg13g2_fill_2 FILLER_4_132 ();
 sg13g2_decap_8 FILLER_4_155 ();
 sg13g2_decap_8 FILLER_4_162 ();
 sg13g2_fill_2 FILLER_4_169 ();
 sg13g2_fill_1 FILLER_4_171 ();
 sg13g2_fill_2 FILLER_4_184 ();
 sg13g2_decap_8 FILLER_4_190 ();
 sg13g2_fill_2 FILLER_4_197 ();
 sg13g2_fill_1 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_4_204 ();
 sg13g2_decap_4 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_219 ();
 sg13g2_decap_8 FILLER_4_247 ();
 sg13g2_fill_2 FILLER_4_254 ();
 sg13g2_fill_1 FILLER_4_256 ();
 sg13g2_fill_1 FILLER_4_261 ();
 sg13g2_fill_1 FILLER_4_266 ();
 sg13g2_fill_1 FILLER_4_271 ();
 sg13g2_fill_1 FILLER_4_276 ();
 sg13g2_fill_2 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_328 ();
 sg13g2_fill_2 FILLER_4_335 ();
 sg13g2_fill_1 FILLER_4_381 ();
 sg13g2_decap_4 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_415 ();
 sg13g2_decap_8 FILLER_4_422 ();
 sg13g2_decap_8 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_4_436 ();
 sg13g2_decap_8 FILLER_4_443 ();
 sg13g2_decap_4 FILLER_4_450 ();
 sg13g2_fill_1 FILLER_4_454 ();
 sg13g2_decap_8 FILLER_4_459 ();
 sg13g2_decap_8 FILLER_4_466 ();
 sg13g2_fill_2 FILLER_4_515 ();
 sg13g2_fill_2 FILLER_4_529 ();
 sg13g2_fill_2 FILLER_4_582 ();
 sg13g2_fill_1 FILLER_4_584 ();
 sg13g2_decap_8 FILLER_4_606 ();
 sg13g2_decap_8 FILLER_4_613 ();
 sg13g2_fill_2 FILLER_4_620 ();
 sg13g2_fill_1 FILLER_4_622 ();
 sg13g2_decap_8 FILLER_4_641 ();
 sg13g2_decap_8 FILLER_4_648 ();
 sg13g2_fill_2 FILLER_4_655 ();
 sg13g2_decap_8 FILLER_4_678 ();
 sg13g2_decap_8 FILLER_4_685 ();
 sg13g2_decap_8 FILLER_4_692 ();
 sg13g2_decap_8 FILLER_4_699 ();
 sg13g2_decap_8 FILLER_4_706 ();
 sg13g2_decap_8 FILLER_4_713 ();
 sg13g2_decap_8 FILLER_4_720 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_decap_8 FILLER_4_734 ();
 sg13g2_decap_8 FILLER_4_741 ();
 sg13g2_decap_8 FILLER_4_748 ();
 sg13g2_decap_8 FILLER_4_755 ();
 sg13g2_decap_8 FILLER_4_762 ();
 sg13g2_decap_8 FILLER_4_769 ();
 sg13g2_decap_8 FILLER_4_776 ();
 sg13g2_decap_8 FILLER_4_783 ();
 sg13g2_decap_8 FILLER_4_790 ();
 sg13g2_decap_8 FILLER_4_797 ();
 sg13g2_decap_8 FILLER_4_804 ();
 sg13g2_decap_8 FILLER_4_811 ();
 sg13g2_decap_4 FILLER_4_818 ();
 sg13g2_fill_2 FILLER_4_858 ();
 sg13g2_fill_1 FILLER_4_860 ();
 sg13g2_fill_2 FILLER_4_875 ();
 sg13g2_decap_4 FILLER_4_881 ();
 sg13g2_decap_8 FILLER_4_895 ();
 sg13g2_decap_8 FILLER_4_902 ();
 sg13g2_decap_4 FILLER_4_945 ();
 sg13g2_decap_8 FILLER_4_961 ();
 sg13g2_fill_2 FILLER_4_968 ();
 sg13g2_fill_1 FILLER_4_970 ();
 sg13g2_decap_8 FILLER_4_999 ();
 sg13g2_decap_8 FILLER_4_1006 ();
 sg13g2_decap_8 FILLER_4_1013 ();
 sg13g2_decap_8 FILLER_4_1020 ();
 sg13g2_decap_8 FILLER_4_1027 ();
 sg13g2_decap_8 FILLER_4_1034 ();
 sg13g2_decap_4 FILLER_4_1041 ();
 sg13g2_fill_2 FILLER_4_1045 ();
 sg13g2_fill_2 FILLER_4_1059 ();
 sg13g2_fill_1 FILLER_4_1061 ();
 sg13g2_decap_8 FILLER_4_1072 ();
 sg13g2_decap_4 FILLER_4_1079 ();
 sg13g2_fill_1 FILLER_4_1083 ();
 sg13g2_decap_8 FILLER_4_1120 ();
 sg13g2_decap_8 FILLER_4_1157 ();
 sg13g2_decap_4 FILLER_4_1164 ();
 sg13g2_fill_1 FILLER_4_1168 ();
 sg13g2_decap_8 FILLER_4_1173 ();
 sg13g2_decap_8 FILLER_4_1180 ();
 sg13g2_decap_8 FILLER_4_1187 ();
 sg13g2_decap_8 FILLER_4_1194 ();
 sg13g2_fill_1 FILLER_4_1201 ();
 sg13g2_decap_8 FILLER_4_1242 ();
 sg13g2_decap_8 FILLER_4_1249 ();
 sg13g2_decap_8 FILLER_4_1256 ();
 sg13g2_decap_8 FILLER_4_1263 ();
 sg13g2_decap_8 FILLER_4_1270 ();
 sg13g2_decap_8 FILLER_4_1277 ();
 sg13g2_decap_8 FILLER_4_1284 ();
 sg13g2_decap_8 FILLER_4_1291 ();
 sg13g2_decap_8 FILLER_4_1298 ();
 sg13g2_decap_8 FILLER_4_1305 ();
 sg13g2_decap_8 FILLER_4_1312 ();
 sg13g2_decap_8 FILLER_4_1319 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_94 ();
 sg13g2_decap_8 FILLER_5_101 ();
 sg13g2_decap_8 FILLER_5_108 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_decap_8 FILLER_5_163 ();
 sg13g2_decap_4 FILLER_5_220 ();
 sg13g2_fill_2 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_247 ();
 sg13g2_fill_2 FILLER_5_254 ();
 sg13g2_fill_1 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_decap_8 FILLER_5_268 ();
 sg13g2_decap_8 FILLER_5_275 ();
 sg13g2_decap_4 FILLER_5_282 ();
 sg13g2_fill_2 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_fill_2 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_4 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_412 ();
 sg13g2_decap_8 FILLER_5_419 ();
 sg13g2_fill_1 FILLER_5_426 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_fill_1 FILLER_5_476 ();
 sg13g2_fill_1 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_519 ();
 sg13g2_decap_8 FILLER_5_526 ();
 sg13g2_decap_8 FILLER_5_533 ();
 sg13g2_fill_1 FILLER_5_540 ();
 sg13g2_decap_4 FILLER_5_545 ();
 sg13g2_fill_1 FILLER_5_549 ();
 sg13g2_fill_1 FILLER_5_554 ();
 sg13g2_fill_1 FILLER_5_576 ();
 sg13g2_decap_8 FILLER_5_610 ();
 sg13g2_decap_4 FILLER_5_617 ();
 sg13g2_decap_8 FILLER_5_625 ();
 sg13g2_decap_4 FILLER_5_632 ();
 sg13g2_fill_2 FILLER_5_636 ();
 sg13g2_decap_8 FILLER_5_694 ();
 sg13g2_decap_8 FILLER_5_701 ();
 sg13g2_decap_8 FILLER_5_708 ();
 sg13g2_decap_8 FILLER_5_715 ();
 sg13g2_decap_8 FILLER_5_722 ();
 sg13g2_decap_8 FILLER_5_729 ();
 sg13g2_decap_4 FILLER_5_736 ();
 sg13g2_fill_1 FILLER_5_740 ();
 sg13g2_fill_1 FILLER_5_745 ();
 sg13g2_decap_8 FILLER_5_750 ();
 sg13g2_decap_8 FILLER_5_757 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_fill_2 FILLER_5_781 ();
 sg13g2_fill_1 FILLER_5_783 ();
 sg13g2_fill_2 FILLER_5_794 ();
 sg13g2_fill_1 FILLER_5_796 ();
 sg13g2_decap_8 FILLER_5_815 ();
 sg13g2_decap_8 FILLER_5_822 ();
 sg13g2_fill_2 FILLER_5_829 ();
 sg13g2_fill_2 FILLER_5_879 ();
 sg13g2_decap_8 FILLER_5_907 ();
 sg13g2_fill_2 FILLER_5_914 ();
 sg13g2_fill_1 FILLER_5_916 ();
 sg13g2_decap_8 FILLER_5_921 ();
 sg13g2_fill_1 FILLER_5_928 ();
 sg13g2_decap_8 FILLER_5_933 ();
 sg13g2_decap_8 FILLER_5_950 ();
 sg13g2_fill_1 FILLER_5_957 ();
 sg13g2_decap_8 FILLER_5_966 ();
 sg13g2_fill_2 FILLER_5_973 ();
 sg13g2_decap_4 FILLER_5_1001 ();
 sg13g2_fill_2 FILLER_5_1005 ();
 sg13g2_decap_8 FILLER_5_1017 ();
 sg13g2_decap_8 FILLER_5_1024 ();
 sg13g2_decap_8 FILLER_5_1031 ();
 sg13g2_decap_8 FILLER_5_1078 ();
 sg13g2_decap_8 FILLER_5_1085 ();
 sg13g2_fill_2 FILLER_5_1096 ();
 sg13g2_fill_1 FILLER_5_1098 ();
 sg13g2_decap_8 FILLER_5_1109 ();
 sg13g2_fill_2 FILLER_5_1126 ();
 sg13g2_decap_8 FILLER_5_1154 ();
 sg13g2_decap_4 FILLER_5_1161 ();
 sg13g2_decap_4 FILLER_5_1195 ();
 sg13g2_fill_2 FILLER_5_1199 ();
 sg13g2_decap_8 FILLER_5_1241 ();
 sg13g2_decap_8 FILLER_5_1248 ();
 sg13g2_decap_8 FILLER_5_1255 ();
 sg13g2_decap_8 FILLER_5_1262 ();
 sg13g2_decap_8 FILLER_5_1269 ();
 sg13g2_decap_8 FILLER_5_1276 ();
 sg13g2_decap_8 FILLER_5_1283 ();
 sg13g2_decap_8 FILLER_5_1290 ();
 sg13g2_decap_8 FILLER_5_1297 ();
 sg13g2_decap_8 FILLER_5_1304 ();
 sg13g2_decap_8 FILLER_5_1311 ();
 sg13g2_decap_8 FILLER_5_1318 ();
 sg13g2_fill_1 FILLER_5_1325 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_fill_2 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_16 ();
 sg13g2_fill_2 FILLER_6_47 ();
 sg13g2_decap_4 FILLER_6_96 ();
 sg13g2_fill_2 FILLER_6_136 ();
 sg13g2_decap_8 FILLER_6_159 ();
 sg13g2_decap_8 FILLER_6_166 ();
 sg13g2_decap_4 FILLER_6_173 ();
 sg13g2_fill_1 FILLER_6_177 ();
 sg13g2_fill_2 FILLER_6_204 ();
 sg13g2_fill_1 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_233 ();
 sg13g2_fill_2 FILLER_6_255 ();
 sg13g2_fill_1 FILLER_6_257 ();
 sg13g2_fill_1 FILLER_6_279 ();
 sg13g2_decap_4 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_fill_2 FILLER_6_390 ();
 sg13g2_fill_1 FILLER_6_392 ();
 sg13g2_decap_4 FILLER_6_414 ();
 sg13g2_fill_1 FILLER_6_422 ();
 sg13g2_fill_2 FILLER_6_449 ();
 sg13g2_fill_2 FILLER_6_461 ();
 sg13g2_fill_2 FILLER_6_467 ();
 sg13g2_decap_8 FILLER_6_495 ();
 sg13g2_fill_2 FILLER_6_502 ();
 sg13g2_fill_1 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_526 ();
 sg13g2_decap_4 FILLER_6_533 ();
 sg13g2_fill_2 FILLER_6_537 ();
 sg13g2_decap_4 FILLER_6_544 ();
 sg13g2_decap_4 FILLER_6_561 ();
 sg13g2_decap_4 FILLER_6_601 ();
 sg13g2_fill_1 FILLER_6_605 ();
 sg13g2_fill_2 FILLER_6_822 ();
 sg13g2_decap_4 FILLER_6_828 ();
 sg13g2_fill_2 FILLER_6_832 ();
 sg13g2_decap_4 FILLER_6_914 ();
 sg13g2_fill_1 FILLER_6_918 ();
 sg13g2_decap_8 FILLER_6_955 ();
 sg13g2_fill_2 FILLER_6_962 ();
 sg13g2_fill_1 FILLER_6_964 ();
 sg13g2_decap_4 FILLER_6_979 ();
 sg13g2_decap_8 FILLER_6_987 ();
 sg13g2_fill_2 FILLER_6_994 ();
 sg13g2_fill_1 FILLER_6_996 ();
 sg13g2_decap_8 FILLER_6_1023 ();
 sg13g2_decap_8 FILLER_6_1030 ();
 sg13g2_decap_4 FILLER_6_1037 ();
 sg13g2_fill_2 FILLER_6_1041 ();
 sg13g2_decap_8 FILLER_6_1079 ();
 sg13g2_decap_8 FILLER_6_1086 ();
 sg13g2_fill_2 FILLER_6_1093 ();
 sg13g2_fill_1 FILLER_6_1095 ();
 sg13g2_fill_2 FILLER_6_1162 ();
 sg13g2_fill_1 FILLER_6_1164 ();
 sg13g2_decap_8 FILLER_6_1195 ();
 sg13g2_fill_1 FILLER_6_1202 ();
 sg13g2_decap_8 FILLER_6_1239 ();
 sg13g2_decap_8 FILLER_6_1246 ();
 sg13g2_decap_8 FILLER_6_1253 ();
 sg13g2_decap_8 FILLER_6_1260 ();
 sg13g2_decap_8 FILLER_6_1267 ();
 sg13g2_decap_8 FILLER_6_1274 ();
 sg13g2_decap_8 FILLER_6_1281 ();
 sg13g2_decap_8 FILLER_6_1288 ();
 sg13g2_decap_8 FILLER_6_1295 ();
 sg13g2_decap_8 FILLER_6_1302 ();
 sg13g2_decap_8 FILLER_6_1309 ();
 sg13g2_decap_8 FILLER_6_1316 ();
 sg13g2_fill_2 FILLER_6_1323 ();
 sg13g2_fill_1 FILLER_6_1325 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_4 FILLER_7_14 ();
 sg13g2_fill_2 FILLER_7_18 ();
 sg13g2_decap_8 FILLER_7_34 ();
 sg13g2_fill_2 FILLER_7_41 ();
 sg13g2_fill_1 FILLER_7_43 ();
 sg13g2_fill_1 FILLER_7_48 ();
 sg13g2_fill_1 FILLER_7_63 ();
 sg13g2_decap_4 FILLER_7_68 ();
 sg13g2_fill_1 FILLER_7_72 ();
 sg13g2_fill_2 FILLER_7_122 ();
 sg13g2_decap_8 FILLER_7_128 ();
 sg13g2_fill_2 FILLER_7_135 ();
 sg13g2_fill_1 FILLER_7_137 ();
 sg13g2_decap_8 FILLER_7_159 ();
 sg13g2_decap_8 FILLER_7_166 ();
 sg13g2_fill_1 FILLER_7_173 ();
 sg13g2_fill_2 FILLER_7_184 ();
 sg13g2_fill_1 FILLER_7_186 ();
 sg13g2_decap_8 FILLER_7_191 ();
 sg13g2_decap_4 FILLER_7_223 ();
 sg13g2_fill_1 FILLER_7_227 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_fill_2 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_decap_4 FILLER_7_295 ();
 sg13g2_decap_4 FILLER_7_339 ();
 sg13g2_fill_2 FILLER_7_343 ();
 sg13g2_fill_1 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_fill_2 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_fill_2 FILLER_7_409 ();
 sg13g2_fill_1 FILLER_7_411 ();
 sg13g2_fill_1 FILLER_7_430 ();
 sg13g2_fill_1 FILLER_7_457 ();
 sg13g2_fill_1 FILLER_7_479 ();
 sg13g2_fill_2 FILLER_7_484 ();
 sg13g2_decap_8 FILLER_7_512 ();
 sg13g2_decap_8 FILLER_7_519 ();
 sg13g2_decap_8 FILLER_7_526 ();
 sg13g2_fill_1 FILLER_7_537 ();
 sg13g2_fill_2 FILLER_7_548 ();
 sg13g2_fill_1 FILLER_7_550 ();
 sg13g2_fill_1 FILLER_7_568 ();
 sg13g2_fill_2 FILLER_7_583 ();
 sg13g2_fill_1 FILLER_7_585 ();
 sg13g2_fill_2 FILLER_7_607 ();
 sg13g2_fill_1 FILLER_7_609 ();
 sg13g2_fill_2 FILLER_7_654 ();
 sg13g2_fill_2 FILLER_7_666 ();
 sg13g2_fill_1 FILLER_7_668 ();
 sg13g2_fill_2 FILLER_7_699 ();
 sg13g2_fill_2 FILLER_7_723 ();
 sg13g2_fill_1 FILLER_7_725 ();
 sg13g2_fill_2 FILLER_7_736 ();
 sg13g2_fill_1 FILLER_7_738 ();
 sg13g2_fill_2 FILLER_7_805 ();
 sg13g2_fill_1 FILLER_7_807 ();
 sg13g2_decap_8 FILLER_7_834 ();
 sg13g2_fill_1 FILLER_7_841 ();
 sg13g2_decap_8 FILLER_7_852 ();
 sg13g2_decap_8 FILLER_7_859 ();
 sg13g2_decap_8 FILLER_7_866 ();
 sg13g2_decap_8 FILLER_7_873 ();
 sg13g2_decap_4 FILLER_7_880 ();
 sg13g2_fill_2 FILLER_7_884 ();
 sg13g2_decap_4 FILLER_7_894 ();
 sg13g2_fill_2 FILLER_7_898 ();
 sg13g2_decap_8 FILLER_7_910 ();
 sg13g2_fill_1 FILLER_7_917 ();
 sg13g2_fill_1 FILLER_7_932 ();
 sg13g2_fill_1 FILLER_7_959 ();
 sg13g2_fill_1 FILLER_7_1012 ();
 sg13g2_decap_4 FILLER_7_1039 ();
 sg13g2_fill_2 FILLER_7_1043 ();
 sg13g2_decap_4 FILLER_7_1097 ();
 sg13g2_decap_8 FILLER_7_1105 ();
 sg13g2_decap_8 FILLER_7_1112 ();
 sg13g2_decap_8 FILLER_7_1119 ();
 sg13g2_decap_8 FILLER_7_1126 ();
 sg13g2_decap_8 FILLER_7_1133 ();
 sg13g2_fill_2 FILLER_7_1140 ();
 sg13g2_decap_4 FILLER_7_1146 ();
 sg13g2_fill_1 FILLER_7_1150 ();
 sg13g2_decap_4 FILLER_7_1199 ();
 sg13g2_decap_8 FILLER_7_1213 ();
 sg13g2_decap_8 FILLER_7_1224 ();
 sg13g2_decap_8 FILLER_7_1231 ();
 sg13g2_decap_8 FILLER_7_1238 ();
 sg13g2_decap_8 FILLER_7_1245 ();
 sg13g2_decap_8 FILLER_7_1252 ();
 sg13g2_decap_8 FILLER_7_1259 ();
 sg13g2_decap_8 FILLER_7_1266 ();
 sg13g2_decap_8 FILLER_7_1273 ();
 sg13g2_decap_8 FILLER_7_1280 ();
 sg13g2_decap_8 FILLER_7_1287 ();
 sg13g2_decap_8 FILLER_7_1294 ();
 sg13g2_decap_8 FILLER_7_1301 ();
 sg13g2_decap_8 FILLER_7_1308 ();
 sg13g2_decap_8 FILLER_7_1315 ();
 sg13g2_decap_4 FILLER_7_1322 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_4 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_62 ();
 sg13g2_fill_1 FILLER_8_69 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_98 ();
 sg13g2_decap_4 FILLER_8_103 ();
 sg13g2_fill_1 FILLER_8_107 ();
 sg13g2_fill_2 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_167 ();
 sg13g2_fill_1 FILLER_8_173 ();
 sg13g2_decap_8 FILLER_8_178 ();
 sg13g2_fill_1 FILLER_8_185 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_4 FILLER_8_203 ();
 sg13g2_fill_2 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_fill_2 FILLER_8_270 ();
 sg13g2_fill_2 FILLER_8_280 ();
 sg13g2_fill_1 FILLER_8_282 ();
 sg13g2_fill_2 FILLER_8_293 ();
 sg13g2_decap_4 FILLER_8_316 ();
 sg13g2_fill_2 FILLER_8_330 ();
 sg13g2_fill_2 FILLER_8_341 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_fill_1 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_366 ();
 sg13g2_decap_8 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_decap_4 FILLER_8_408 ();
 sg13g2_fill_1 FILLER_8_463 ();
 sg13g2_decap_8 FILLER_8_500 ();
 sg13g2_decap_4 FILLER_8_507 ();
 sg13g2_fill_1 FILLER_8_511 ();
 sg13g2_decap_4 FILLER_8_517 ();
 sg13g2_fill_1 FILLER_8_521 ();
 sg13g2_decap_4 FILLER_8_562 ();
 sg13g2_fill_2 FILLER_8_571 ();
 sg13g2_fill_1 FILLER_8_573 ();
 sg13g2_decap_8 FILLER_8_614 ();
 sg13g2_fill_1 FILLER_8_621 ();
 sg13g2_fill_1 FILLER_8_653 ();
 sg13g2_decap_8 FILLER_8_664 ();
 sg13g2_decap_8 FILLER_8_671 ();
 sg13g2_decap_8 FILLER_8_682 ();
 sg13g2_decap_8 FILLER_8_689 ();
 sg13g2_decap_4 FILLER_8_696 ();
 sg13g2_fill_2 FILLER_8_700 ();
 sg13g2_fill_2 FILLER_8_738 ();
 sg13g2_fill_1 FILLER_8_788 ();
 sg13g2_fill_1 FILLER_8_829 ();
 sg13g2_decap_4 FILLER_8_840 ();
 sg13g2_fill_1 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_875 ();
 sg13g2_fill_1 FILLER_8_882 ();
 sg13g2_fill_2 FILLER_8_909 ();
 sg13g2_fill_1 FILLER_8_911 ();
 sg13g2_fill_2 FILLER_8_922 ();
 sg13g2_decap_4 FILLER_8_959 ();
 sg13g2_fill_1 FILLER_8_963 ();
 sg13g2_fill_2 FILLER_8_1010 ();
 sg13g2_fill_2 FILLER_8_1054 ();
 sg13g2_fill_1 FILLER_8_1056 ();
 sg13g2_decap_8 FILLER_8_1067 ();
 sg13g2_fill_2 FILLER_8_1104 ();
 sg13g2_fill_1 FILLER_8_1106 ();
 sg13g2_decap_8 FILLER_8_1111 ();
 sg13g2_fill_1 FILLER_8_1118 ();
 sg13g2_decap_8 FILLER_8_1123 ();
 sg13g2_fill_1 FILLER_8_1130 ();
 sg13g2_fill_2 FILLER_8_1157 ();
 sg13g2_fill_1 FILLER_8_1159 ();
 sg13g2_decap_4 FILLER_8_1200 ();
 sg13g2_decap_8 FILLER_8_1234 ();
 sg13g2_decap_8 FILLER_8_1241 ();
 sg13g2_decap_8 FILLER_8_1248 ();
 sg13g2_decap_8 FILLER_8_1255 ();
 sg13g2_decap_8 FILLER_8_1262 ();
 sg13g2_decap_8 FILLER_8_1269 ();
 sg13g2_decap_8 FILLER_8_1276 ();
 sg13g2_decap_8 FILLER_8_1283 ();
 sg13g2_decap_8 FILLER_8_1290 ();
 sg13g2_decap_8 FILLER_8_1297 ();
 sg13g2_decap_8 FILLER_8_1304 ();
 sg13g2_decap_8 FILLER_8_1311 ();
 sg13g2_decap_8 FILLER_8_1318 ();
 sg13g2_fill_1 FILLER_8_1325 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_18 ();
 sg13g2_decap_4 FILLER_9_40 ();
 sg13g2_fill_2 FILLER_9_44 ();
 sg13g2_decap_8 FILLER_9_67 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_4 FILLER_9_95 ();
 sg13g2_decap_4 FILLER_9_109 ();
 sg13g2_fill_2 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_145 ();
 sg13g2_decap_8 FILLER_9_152 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_fill_2 FILLER_9_166 ();
 sg13g2_decap_4 FILLER_9_181 ();
 sg13g2_fill_1 FILLER_9_185 ();
 sg13g2_fill_2 FILLER_9_194 ();
 sg13g2_decap_8 FILLER_9_226 ();
 sg13g2_decap_8 FILLER_9_233 ();
 sg13g2_decap_4 FILLER_9_240 ();
 sg13g2_fill_2 FILLER_9_259 ();
 sg13g2_fill_1 FILLER_9_261 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_fill_2 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_fill_2 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_367 ();
 sg13g2_decap_4 FILLER_9_411 ();
 sg13g2_decap_4 FILLER_9_451 ();
 sg13g2_fill_1 FILLER_9_455 ();
 sg13g2_fill_1 FILLER_9_464 ();
 sg13g2_fill_1 FILLER_9_474 ();
 sg13g2_fill_1 FILLER_9_479 ();
 sg13g2_decap_8 FILLER_9_484 ();
 sg13g2_decap_8 FILLER_9_491 ();
 sg13g2_decap_8 FILLER_9_498 ();
 sg13g2_decap_8 FILLER_9_505 ();
 sg13g2_decap_8 FILLER_9_516 ();
 sg13g2_decap_8 FILLER_9_523 ();
 sg13g2_decap_8 FILLER_9_530 ();
 sg13g2_fill_1 FILLER_9_537 ();
 sg13g2_decap_8 FILLER_9_580 ();
 sg13g2_decap_8 FILLER_9_587 ();
 sg13g2_fill_1 FILLER_9_594 ();
 sg13g2_decap_8 FILLER_9_599 ();
 sg13g2_decap_8 FILLER_9_606 ();
 sg13g2_decap_8 FILLER_9_613 ();
 sg13g2_decap_8 FILLER_9_620 ();
 sg13g2_decap_8 FILLER_9_627 ();
 sg13g2_fill_2 FILLER_9_634 ();
 sg13g2_decap_8 FILLER_9_645 ();
 sg13g2_fill_1 FILLER_9_652 ();
 sg13g2_decap_8 FILLER_9_661 ();
 sg13g2_decap_8 FILLER_9_668 ();
 sg13g2_decap_8 FILLER_9_675 ();
 sg13g2_decap_8 FILLER_9_682 ();
 sg13g2_decap_8 FILLER_9_689 ();
 sg13g2_fill_2 FILLER_9_696 ();
 sg13g2_decap_8 FILLER_9_738 ();
 sg13g2_decap_8 FILLER_9_745 ();
 sg13g2_decap_4 FILLER_9_752 ();
 sg13g2_fill_1 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_761 ();
 sg13g2_decap_8 FILLER_9_768 ();
 sg13g2_decap_8 FILLER_9_775 ();
 sg13g2_decap_8 FILLER_9_782 ();
 sg13g2_decap_8 FILLER_9_789 ();
 sg13g2_fill_2 FILLER_9_796 ();
 sg13g2_fill_1 FILLER_9_798 ();
 sg13g2_decap_4 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_815 ();
 sg13g2_decap_4 FILLER_9_852 ();
 sg13g2_decap_8 FILLER_9_864 ();
 sg13g2_decap_8 FILLER_9_871 ();
 sg13g2_decap_8 FILLER_9_878 ();
 sg13g2_fill_2 FILLER_9_967 ();
 sg13g2_fill_1 FILLER_9_969 ();
 sg13g2_decap_8 FILLER_9_984 ();
 sg13g2_decap_4 FILLER_9_995 ();
 sg13g2_fill_2 FILLER_9_999 ();
 sg13g2_fill_2 FILLER_9_1051 ();
 sg13g2_decap_8 FILLER_9_1057 ();
 sg13g2_fill_2 FILLER_9_1064 ();
 sg13g2_fill_1 FILLER_9_1084 ();
 sg13g2_fill_1 FILLER_9_1098 ();
 sg13g2_fill_2 FILLER_9_1147 ();
 sg13g2_fill_2 FILLER_9_1159 ();
 sg13g2_fill_2 FILLER_9_1197 ();
 sg13g2_fill_1 FILLER_9_1199 ();
 sg13g2_decap_8 FILLER_9_1240 ();
 sg13g2_decap_8 FILLER_9_1247 ();
 sg13g2_decap_8 FILLER_9_1254 ();
 sg13g2_decap_8 FILLER_9_1261 ();
 sg13g2_decap_8 FILLER_9_1268 ();
 sg13g2_decap_8 FILLER_9_1275 ();
 sg13g2_decap_8 FILLER_9_1282 ();
 sg13g2_decap_8 FILLER_9_1289 ();
 sg13g2_decap_8 FILLER_9_1296 ();
 sg13g2_decap_8 FILLER_9_1303 ();
 sg13g2_decap_8 FILLER_9_1310 ();
 sg13g2_decap_8 FILLER_9_1317 ();
 sg13g2_fill_2 FILLER_9_1324 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_90 ();
 sg13g2_decap_4 FILLER_10_101 ();
 sg13g2_fill_1 FILLER_10_109 ();
 sg13g2_fill_2 FILLER_10_120 ();
 sg13g2_fill_2 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_fill_2 FILLER_10_261 ();
 sg13g2_fill_2 FILLER_10_299 ();
 sg13g2_fill_1 FILLER_10_301 ();
 sg13g2_decap_4 FILLER_10_333 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_353 ();
 sg13g2_fill_1 FILLER_10_355 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_fill_1 FILLER_10_409 ();
 sg13g2_fill_1 FILLER_10_418 ();
 sg13g2_decap_8 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_10_430 ();
 sg13g2_fill_2 FILLER_10_437 ();
 sg13g2_fill_2 FILLER_10_453 ();
 sg13g2_fill_1 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_481 ();
 sg13g2_fill_2 FILLER_10_488 ();
 sg13g2_fill_2 FILLER_10_498 ();
 sg13g2_decap_8 FILLER_10_530 ();
 sg13g2_decap_8 FILLER_10_537 ();
 sg13g2_decap_4 FILLER_10_581 ();
 sg13g2_fill_2 FILLER_10_585 ();
 sg13g2_decap_8 FILLER_10_591 ();
 sg13g2_fill_1 FILLER_10_598 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_fill_1 FILLER_10_646 ();
 sg13g2_decap_8 FILLER_10_691 ();
 sg13g2_decap_8 FILLER_10_698 ();
 sg13g2_decap_4 FILLER_10_705 ();
 sg13g2_decap_8 FILLER_10_745 ();
 sg13g2_decap_8 FILLER_10_752 ();
 sg13g2_decap_8 FILLER_10_759 ();
 sg13g2_decap_8 FILLER_10_766 ();
 sg13g2_fill_2 FILLER_10_773 ();
 sg13g2_decap_8 FILLER_10_785 ();
 sg13g2_decap_4 FILLER_10_800 ();
 sg13g2_fill_2 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_878 ();
 sg13g2_decap_8 FILLER_10_885 ();
 sg13g2_fill_1 FILLER_10_892 ();
 sg13g2_decap_4 FILLER_10_949 ();
 sg13g2_decap_8 FILLER_10_957 ();
 sg13g2_decap_4 FILLER_10_968 ();
 sg13g2_fill_2 FILLER_10_972 ();
 sg13g2_decap_4 FILLER_10_984 ();
 sg13g2_fill_2 FILLER_10_988 ();
 sg13g2_decap_8 FILLER_10_1000 ();
 sg13g2_decap_4 FILLER_10_1007 ();
 sg13g2_fill_1 FILLER_10_1011 ();
 sg13g2_decap_4 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1030 ();
 sg13g2_decap_8 FILLER_10_1035 ();
 sg13g2_decap_8 FILLER_10_1042 ();
 sg13g2_decap_4 FILLER_10_1049 ();
 sg13g2_fill_1 FILLER_10_1053 ();
 sg13g2_fill_2 FILLER_10_1064 ();
 sg13g2_decap_4 FILLER_10_1070 ();
 sg13g2_fill_2 FILLER_10_1074 ();
 sg13g2_fill_2 FILLER_10_1096 ();
 sg13g2_decap_4 FILLER_10_1124 ();
 sg13g2_fill_1 FILLER_10_1128 ();
 sg13g2_decap_4 FILLER_10_1133 ();
 sg13g2_decap_8 FILLER_10_1141 ();
 sg13g2_decap_8 FILLER_10_1148 ();
 sg13g2_fill_1 FILLER_10_1155 ();
 sg13g2_fill_2 FILLER_10_1182 ();
 sg13g2_fill_1 FILLER_10_1184 ();
 sg13g2_fill_2 FILLER_10_1203 ();
 sg13g2_decap_8 FILLER_10_1241 ();
 sg13g2_decap_8 FILLER_10_1248 ();
 sg13g2_decap_8 FILLER_10_1255 ();
 sg13g2_decap_8 FILLER_10_1262 ();
 sg13g2_decap_8 FILLER_10_1269 ();
 sg13g2_decap_8 FILLER_10_1276 ();
 sg13g2_decap_8 FILLER_10_1283 ();
 sg13g2_decap_8 FILLER_10_1290 ();
 sg13g2_decap_8 FILLER_10_1297 ();
 sg13g2_decap_8 FILLER_10_1304 ();
 sg13g2_decap_8 FILLER_10_1311 ();
 sg13g2_decap_8 FILLER_10_1318 ();
 sg13g2_fill_1 FILLER_10_1325 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_5 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_60 ();
 sg13g2_decap_8 FILLER_11_83 ();
 sg13g2_decap_8 FILLER_11_90 ();
 sg13g2_fill_2 FILLER_11_97 ();
 sg13g2_decap_4 FILLER_11_113 ();
 sg13g2_fill_2 FILLER_11_117 ();
 sg13g2_fill_2 FILLER_11_123 ();
 sg13g2_fill_1 FILLER_11_125 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_fill_1 FILLER_11_179 ();
 sg13g2_decap_4 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_192 ();
 sg13g2_fill_2 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_264 ();
 sg13g2_fill_2 FILLER_11_274 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_309 ();
 sg13g2_decap_8 FILLER_11_316 ();
 sg13g2_fill_2 FILLER_11_323 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_fill_1 FILLER_11_336 ();
 sg13g2_fill_2 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_415 ();
 sg13g2_decap_4 FILLER_11_422 ();
 sg13g2_fill_1 FILLER_11_430 ();
 sg13g2_fill_1 FILLER_11_452 ();
 sg13g2_fill_2 FILLER_11_457 ();
 sg13g2_decap_4 FILLER_11_485 ();
 sg13g2_fill_2 FILLER_11_489 ();
 sg13g2_fill_2 FILLER_11_541 ();
 sg13g2_fill_1 FILLER_11_543 ();
 sg13g2_fill_1 FILLER_11_558 ();
 sg13g2_decap_4 FILLER_11_595 ();
 sg13g2_fill_1 FILLER_11_599 ();
 sg13g2_fill_2 FILLER_11_621 ();
 sg13g2_fill_2 FILLER_11_664 ();
 sg13g2_fill_1 FILLER_11_666 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_fill_2 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_720 ();
 sg13g2_decap_4 FILLER_11_727 ();
 sg13g2_decap_8 FILLER_11_741 ();
 sg13g2_fill_2 FILLER_11_822 ();
 sg13g2_fill_1 FILLER_11_824 ();
 sg13g2_decap_8 FILLER_11_829 ();
 sg13g2_decap_4 FILLER_11_836 ();
 sg13g2_decap_4 FILLER_11_906 ();
 sg13g2_fill_2 FILLER_11_910 ();
 sg13g2_decap_8 FILLER_11_916 ();
 sg13g2_decap_4 FILLER_11_923 ();
 sg13g2_fill_1 FILLER_11_927 ();
 sg13g2_decap_8 FILLER_11_932 ();
 sg13g2_decap_4 FILLER_11_939 ();
 sg13g2_fill_2 FILLER_11_943 ();
 sg13g2_decap_4 FILLER_11_971 ();
 sg13g2_fill_2 FILLER_11_975 ();
 sg13g2_decap_4 FILLER_11_1003 ();
 sg13g2_fill_1 FILLER_11_1021 ();
 sg13g2_decap_8 FILLER_11_1048 ();
 sg13g2_decap_8 FILLER_11_1115 ();
 sg13g2_decap_8 FILLER_11_1122 ();
 sg13g2_decap_8 FILLER_11_1129 ();
 sg13g2_fill_2 FILLER_11_1136 ();
 sg13g2_fill_1 FILLER_11_1138 ();
 sg13g2_decap_4 FILLER_11_1161 ();
 sg13g2_decap_8 FILLER_11_1179 ();
 sg13g2_decap_8 FILLER_11_1186 ();
 sg13g2_decap_8 FILLER_11_1193 ();
 sg13g2_decap_8 FILLER_11_1200 ();
 sg13g2_fill_2 FILLER_11_1207 ();
 sg13g2_fill_1 FILLER_11_1209 ();
 sg13g2_decap_8 FILLER_11_1231 ();
 sg13g2_decap_8 FILLER_11_1238 ();
 sg13g2_decap_8 FILLER_11_1245 ();
 sg13g2_decap_8 FILLER_11_1252 ();
 sg13g2_decap_8 FILLER_11_1259 ();
 sg13g2_decap_8 FILLER_11_1266 ();
 sg13g2_decap_8 FILLER_11_1273 ();
 sg13g2_decap_8 FILLER_11_1280 ();
 sg13g2_decap_8 FILLER_11_1287 ();
 sg13g2_decap_8 FILLER_11_1294 ();
 sg13g2_decap_8 FILLER_11_1301 ();
 sg13g2_decap_8 FILLER_11_1308 ();
 sg13g2_decap_8 FILLER_11_1315 ();
 sg13g2_decap_4 FILLER_11_1322 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_fill_2 FILLER_12_20 ();
 sg13g2_fill_1 FILLER_12_22 ();
 sg13g2_fill_1 FILLER_12_67 ();
 sg13g2_fill_1 FILLER_12_73 ();
 sg13g2_fill_1 FILLER_12_138 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_decap_8 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_178 ();
 sg13g2_decap_8 FILLER_12_185 ();
 sg13g2_fill_2 FILLER_12_192 ();
 sg13g2_fill_1 FILLER_12_194 ();
 sg13g2_decap_4 FILLER_12_209 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_4 FILLER_12_224 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_decap_4 FILLER_12_250 ();
 sg13g2_fill_2 FILLER_12_254 ();
 sg13g2_fill_2 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_342 ();
 sg13g2_fill_2 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_4 FILLER_12_413 ();
 sg13g2_fill_2 FILLER_12_417 ();
 sg13g2_fill_2 FILLER_12_455 ();
 sg13g2_fill_1 FILLER_12_457 ();
 sg13g2_decap_8 FILLER_12_488 ();
 sg13g2_decap_8 FILLER_12_531 ();
 sg13g2_decap_4 FILLER_12_538 ();
 sg13g2_fill_2 FILLER_12_542 ();
 sg13g2_fill_1 FILLER_12_570 ();
 sg13g2_decap_4 FILLER_12_581 ();
 sg13g2_fill_1 FILLER_12_585 ();
 sg13g2_decap_8 FILLER_12_620 ();
 sg13g2_fill_1 FILLER_12_627 ();
 sg13g2_decap_4 FILLER_12_632 ();
 sg13g2_fill_1 FILLER_12_636 ();
 sg13g2_fill_2 FILLER_12_684 ();
 sg13g2_fill_1 FILLER_12_686 ();
 sg13g2_fill_2 FILLER_12_712 ();
 sg13g2_fill_2 FILLER_12_740 ();
 sg13g2_fill_2 FILLER_12_772 ();
 sg13g2_fill_1 FILLER_12_774 ();
 sg13g2_decap_8 FILLER_12_815 ();
 sg13g2_decap_4 FILLER_12_822 ();
 sg13g2_fill_2 FILLER_12_856 ();
 sg13g2_decap_4 FILLER_12_872 ();
 sg13g2_fill_2 FILLER_12_876 ();
 sg13g2_decap_8 FILLER_12_900 ();
 sg13g2_fill_1 FILLER_12_907 ();
 sg13g2_decap_4 FILLER_12_916 ();
 sg13g2_fill_1 FILLER_12_920 ();
 sg13g2_decap_8 FILLER_12_925 ();
 sg13g2_fill_1 FILLER_12_932 ();
 sg13g2_decap_8 FILLER_12_943 ();
 sg13g2_fill_2 FILLER_12_950 ();
 sg13g2_decap_4 FILLER_12_1072 ();
 sg13g2_fill_2 FILLER_12_1076 ();
 sg13g2_fill_1 FILLER_12_1170 ();
 sg13g2_decap_8 FILLER_12_1197 ();
 sg13g2_fill_2 FILLER_12_1204 ();
 sg13g2_fill_1 FILLER_12_1206 ();
 sg13g2_decap_8 FILLER_12_1259 ();
 sg13g2_decap_8 FILLER_12_1266 ();
 sg13g2_decap_8 FILLER_12_1273 ();
 sg13g2_decap_8 FILLER_12_1280 ();
 sg13g2_decap_8 FILLER_12_1287 ();
 sg13g2_decap_8 FILLER_12_1294 ();
 sg13g2_decap_8 FILLER_12_1301 ();
 sg13g2_decap_8 FILLER_12_1308 ();
 sg13g2_decap_8 FILLER_12_1315 ();
 sg13g2_decap_4 FILLER_12_1322 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_decap_4 FILLER_13_15 ();
 sg13g2_fill_1 FILLER_13_19 ();
 sg13g2_decap_4 FILLER_13_33 ();
 sg13g2_decap_4 FILLER_13_55 ();
 sg13g2_fill_2 FILLER_13_59 ();
 sg13g2_decap_8 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_94 ();
 sg13g2_fill_1 FILLER_13_100 ();
 sg13g2_fill_2 FILLER_13_111 ();
 sg13g2_fill_1 FILLER_13_139 ();
 sg13g2_fill_2 FILLER_13_150 ();
 sg13g2_decap_8 FILLER_13_178 ();
 sg13g2_decap_4 FILLER_13_189 ();
 sg13g2_fill_1 FILLER_13_197 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_decap_8 FILLER_13_209 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_2 FILLER_13_259 ();
 sg13g2_fill_1 FILLER_13_279 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_fill_2 FILLER_13_294 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_fill_2 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_fill_2 FILLER_13_417 ();
 sg13g2_fill_1 FILLER_13_419 ();
 sg13g2_decap_4 FILLER_13_475 ();
 sg13g2_decap_4 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_4 FILLER_13_504 ();
 sg13g2_fill_1 FILLER_13_508 ();
 sg13g2_decap_8 FILLER_13_513 ();
 sg13g2_decap_8 FILLER_13_520 ();
 sg13g2_decap_8 FILLER_13_527 ();
 sg13g2_decap_8 FILLER_13_534 ();
 sg13g2_decap_4 FILLER_13_541 ();
 sg13g2_fill_2 FILLER_13_545 ();
 sg13g2_decap_4 FILLER_13_556 ();
 sg13g2_decap_4 FILLER_13_581 ();
 sg13g2_fill_1 FILLER_13_585 ();
 sg13g2_fill_2 FILLER_13_616 ();
 sg13g2_decap_4 FILLER_13_630 ();
 sg13g2_fill_1 FILLER_13_670 ();
 sg13g2_decap_8 FILLER_13_675 ();
 sg13g2_fill_2 FILLER_13_682 ();
 sg13g2_fill_1 FILLER_13_684 ();
 sg13g2_decap_8 FILLER_13_706 ();
 sg13g2_fill_2 FILLER_13_713 ();
 sg13g2_fill_1 FILLER_13_715 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_fill_1 FILLER_13_749 ();
 sg13g2_decap_4 FILLER_13_754 ();
 sg13g2_fill_2 FILLER_13_794 ();
 sg13g2_fill_1 FILLER_13_796 ();
 sg13g2_decap_8 FILLER_13_815 ();
 sg13g2_decap_4 FILLER_13_822 ();
 sg13g2_fill_1 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_867 ();
 sg13g2_fill_2 FILLER_13_874 ();
 sg13g2_fill_1 FILLER_13_876 ();
 sg13g2_fill_1 FILLER_13_913 ();
 sg13g2_decap_4 FILLER_13_940 ();
 sg13g2_fill_1 FILLER_13_944 ();
 sg13g2_fill_1 FILLER_13_971 ();
 sg13g2_fill_1 FILLER_13_982 ();
 sg13g2_fill_1 FILLER_13_997 ();
 sg13g2_fill_1 FILLER_13_1042 ();
 sg13g2_fill_1 FILLER_13_1047 ();
 sg13g2_fill_2 FILLER_13_1052 ();
 sg13g2_fill_2 FILLER_13_1062 ();
 sg13g2_fill_1 FILLER_13_1064 ();
 sg13g2_fill_2 FILLER_13_1091 ();
 sg13g2_fill_2 FILLER_13_1119 ();
 sg13g2_fill_1 FILLER_13_1121 ();
 sg13g2_decap_4 FILLER_13_1148 ();
 sg13g2_fill_2 FILLER_13_1152 ();
 sg13g2_fill_2 FILLER_13_1180 ();
 sg13g2_fill_1 FILLER_13_1182 ();
 sg13g2_decap_4 FILLER_13_1187 ();
 sg13g2_fill_2 FILLER_13_1191 ();
 sg13g2_decap_8 FILLER_13_1285 ();
 sg13g2_decap_8 FILLER_13_1292 ();
 sg13g2_decap_8 FILLER_13_1299 ();
 sg13g2_decap_8 FILLER_13_1306 ();
 sg13g2_decap_8 FILLER_13_1313 ();
 sg13g2_decap_4 FILLER_13_1320 ();
 sg13g2_fill_2 FILLER_13_1324 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_34 ();
 sg13g2_decap_8 FILLER_14_41 ();
 sg13g2_decap_8 FILLER_14_48 ();
 sg13g2_fill_1 FILLER_14_55 ();
 sg13g2_fill_2 FILLER_14_74 ();
 sg13g2_decap_8 FILLER_14_80 ();
 sg13g2_decap_8 FILLER_14_87 ();
 sg13g2_decap_8 FILLER_14_94 ();
 sg13g2_decap_8 FILLER_14_101 ();
 sg13g2_decap_8 FILLER_14_108 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_decap_8 FILLER_14_125 ();
 sg13g2_decap_4 FILLER_14_132 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_157 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_4 FILLER_14_292 ();
 sg13g2_fill_2 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_fill_2 FILLER_14_334 ();
 sg13g2_fill_1 FILLER_14_336 ();
 sg13g2_fill_2 FILLER_14_341 ();
 sg13g2_fill_1 FILLER_14_343 ();
 sg13g2_decap_4 FILLER_14_362 ();
 sg13g2_fill_1 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_fill_2 FILLER_14_395 ();
 sg13g2_fill_1 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_419 ();
 sg13g2_fill_2 FILLER_14_423 ();
 sg13g2_decap_8 FILLER_14_456 ();
 sg13g2_fill_1 FILLER_14_467 ();
 sg13g2_fill_2 FILLER_14_478 ();
 sg13g2_decap_4 FILLER_14_553 ();
 sg13g2_fill_2 FILLER_14_557 ();
 sg13g2_decap_8 FILLER_14_580 ();
 sg13g2_decap_4 FILLER_14_605 ();
 sg13g2_fill_2 FILLER_14_622 ();
 sg13g2_fill_1 FILLER_14_624 ();
 sg13g2_decap_8 FILLER_14_629 ();
 sg13g2_decap_8 FILLER_14_636 ();
 sg13g2_decap_8 FILLER_14_643 ();
 sg13g2_fill_1 FILLER_14_650 ();
 sg13g2_decap_8 FILLER_14_655 ();
 sg13g2_decap_8 FILLER_14_662 ();
 sg13g2_fill_2 FILLER_14_669 ();
 sg13g2_fill_1 FILLER_14_671 ();
 sg13g2_decap_8 FILLER_14_698 ();
 sg13g2_decap_8 FILLER_14_705 ();
 sg13g2_decap_8 FILLER_14_712 ();
 sg13g2_fill_2 FILLER_14_719 ();
 sg13g2_fill_1 FILLER_14_721 ();
 sg13g2_decap_4 FILLER_14_726 ();
 sg13g2_decap_8 FILLER_14_740 ();
 sg13g2_fill_1 FILLER_14_747 ();
 sg13g2_decap_4 FILLER_14_756 ();
 sg13g2_decap_4 FILLER_14_786 ();
 sg13g2_fill_2 FILLER_14_790 ();
 sg13g2_decap_8 FILLER_14_823 ();
 sg13g2_fill_1 FILLER_14_830 ();
 sg13g2_decap_8 FILLER_14_867 ();
 sg13g2_decap_8 FILLER_14_874 ();
 sg13g2_decap_8 FILLER_14_881 ();
 sg13g2_fill_1 FILLER_14_888 ();
 sg13g2_fill_2 FILLER_14_893 ();
 sg13g2_fill_1 FILLER_14_895 ();
 sg13g2_decap_8 FILLER_14_900 ();
 sg13g2_decap_4 FILLER_14_907 ();
 sg13g2_fill_1 FILLER_14_911 ();
 sg13g2_decap_4 FILLER_14_948 ();
 sg13g2_fill_2 FILLER_14_952 ();
 sg13g2_decap_8 FILLER_14_976 ();
 sg13g2_fill_1 FILLER_14_983 ();
 sg13g2_decap_8 FILLER_14_988 ();
 sg13g2_decap_4 FILLER_14_995 ();
 sg13g2_fill_1 FILLER_14_999 ();
 sg13g2_decap_8 FILLER_14_1012 ();
 sg13g2_decap_4 FILLER_14_1019 ();
 sg13g2_fill_1 FILLER_14_1023 ();
 sg13g2_decap_8 FILLER_14_1032 ();
 sg13g2_decap_4 FILLER_14_1039 ();
 sg13g2_fill_2 FILLER_14_1043 ();
 sg13g2_decap_8 FILLER_14_1109 ();
 sg13g2_decap_8 FILLER_14_1116 ();
 sg13g2_fill_2 FILLER_14_1123 ();
 sg13g2_decap_4 FILLER_14_1159 ();
 sg13g2_decap_8 FILLER_14_1167 ();
 sg13g2_fill_2 FILLER_14_1274 ();
 sg13g2_decap_8 FILLER_14_1280 ();
 sg13g2_decap_8 FILLER_14_1287 ();
 sg13g2_decap_8 FILLER_14_1294 ();
 sg13g2_decap_8 FILLER_14_1301 ();
 sg13g2_decap_8 FILLER_14_1308 ();
 sg13g2_decap_8 FILLER_14_1315 ();
 sg13g2_decap_4 FILLER_14_1322 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_30 ();
 sg13g2_decap_8 FILLER_15_52 ();
 sg13g2_fill_2 FILLER_15_59 ();
 sg13g2_decap_8 FILLER_15_82 ();
 sg13g2_decap_4 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_108 ();
 sg13g2_decap_4 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_121 ();
 sg13g2_decap_4 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_250 ();
 sg13g2_decap_8 FILLER_15_257 ();
 sg13g2_decap_8 FILLER_15_264 ();
 sg13g2_decap_8 FILLER_15_271 ();
 sg13g2_fill_2 FILLER_15_278 ();
 sg13g2_fill_1 FILLER_15_280 ();
 sg13g2_decap_4 FILLER_15_289 ();
 sg13g2_fill_1 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_fill_2 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_4 FILLER_15_431 ();
 sg13g2_fill_2 FILLER_15_493 ();
 sg13g2_fill_2 FILLER_15_516 ();
 sg13g2_fill_1 FILLER_15_552 ();
 sg13g2_fill_1 FILLER_15_563 ();
 sg13g2_fill_1 FILLER_15_574 ();
 sg13g2_fill_1 FILLER_15_596 ();
 sg13g2_fill_2 FILLER_15_652 ();
 sg13g2_fill_2 FILLER_15_664 ();
 sg13g2_fill_1 FILLER_15_666 ();
 sg13g2_decap_8 FILLER_15_709 ();
 sg13g2_decap_8 FILLER_15_716 ();
 sg13g2_decap_8 FILLER_15_723 ();
 sg13g2_decap_8 FILLER_15_730 ();
 sg13g2_fill_1 FILLER_15_737 ();
 sg13g2_decap_4 FILLER_15_748 ();
 sg13g2_fill_1 FILLER_15_752 ();
 sg13g2_fill_2 FILLER_15_779 ();
 sg13g2_fill_1 FILLER_15_781 ();
 sg13g2_decap_8 FILLER_15_820 ();
 sg13g2_decap_8 FILLER_15_827 ();
 sg13g2_fill_2 FILLER_15_834 ();
 sg13g2_fill_2 FILLER_15_840 ();
 sg13g2_decap_4 FILLER_15_846 ();
 sg13g2_fill_1 FILLER_15_850 ();
 sg13g2_decap_8 FILLER_15_861 ();
 sg13g2_fill_2 FILLER_15_868 ();
 sg13g2_fill_1 FILLER_15_870 ();
 sg13g2_decap_8 FILLER_15_907 ();
 sg13g2_decap_4 FILLER_15_914 ();
 sg13g2_fill_1 FILLER_15_918 ();
 sg13g2_fill_2 FILLER_15_959 ();
 sg13g2_fill_2 FILLER_15_973 ();
 sg13g2_fill_1 FILLER_15_975 ();
 sg13g2_decap_8 FILLER_15_980 ();
 sg13g2_decap_8 FILLER_15_987 ();
 sg13g2_decap_8 FILLER_15_994 ();
 sg13g2_decap_4 FILLER_15_1001 ();
 sg13g2_fill_2 FILLER_15_1005 ();
 sg13g2_decap_8 FILLER_15_1037 ();
 sg13g2_decap_4 FILLER_15_1044 ();
 sg13g2_decap_8 FILLER_15_1066 ();
 sg13g2_fill_2 FILLER_15_1077 ();
 sg13g2_fill_1 FILLER_15_1079 ();
 sg13g2_decap_8 FILLER_15_1110 ();
 sg13g2_fill_1 FILLER_15_1117 ();
 sg13g2_decap_4 FILLER_15_1130 ();
 sg13g2_decap_8 FILLER_15_1152 ();
 sg13g2_decap_8 FILLER_15_1159 ();
 sg13g2_decap_4 FILLER_15_1166 ();
 sg13g2_fill_1 FILLER_15_1182 ();
 sg13g2_decap_4 FILLER_15_1191 ();
 sg13g2_decap_8 FILLER_15_1209 ();
 sg13g2_decap_8 FILLER_15_1216 ();
 sg13g2_decap_8 FILLER_15_1223 ();
 sg13g2_decap_8 FILLER_15_1230 ();
 sg13g2_fill_1 FILLER_15_1237 ();
 sg13g2_decap_8 FILLER_15_1284 ();
 sg13g2_decap_8 FILLER_15_1291 ();
 sg13g2_decap_8 FILLER_15_1298 ();
 sg13g2_decap_8 FILLER_15_1305 ();
 sg13g2_decap_8 FILLER_15_1312 ();
 sg13g2_decap_8 FILLER_15_1319 ();
 sg13g2_decap_8 FILLER_16_54 ();
 sg13g2_decap_4 FILLER_16_61 ();
 sg13g2_fill_1 FILLER_16_65 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_decap_4 FILLER_16_174 ();
 sg13g2_fill_2 FILLER_16_178 ();
 sg13g2_fill_2 FILLER_16_184 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_234 ();
 sg13g2_decap_4 FILLER_16_241 ();
 sg13g2_fill_2 FILLER_16_245 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_2 FILLER_16_298 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_decap_4 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_340 ();
 sg13g2_fill_2 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_405 ();
 sg13g2_decap_4 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_fill_2 FILLER_16_441 ();
 sg13g2_fill_1 FILLER_16_443 ();
 sg13g2_fill_2 FILLER_16_517 ();
 sg13g2_fill_2 FILLER_16_571 ();
 sg13g2_decap_4 FILLER_16_583 ();
 sg13g2_fill_2 FILLER_16_587 ();
 sg13g2_fill_2 FILLER_16_625 ();
 sg13g2_fill_2 FILLER_16_671 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_fill_1 FILLER_16_714 ();
 sg13g2_fill_1 FILLER_16_741 ();
 sg13g2_fill_1 FILLER_16_768 ();
 sg13g2_fill_1 FILLER_16_779 ();
 sg13g2_fill_2 FILLER_16_790 ();
 sg13g2_fill_2 FILLER_16_802 ();
 sg13g2_decap_8 FILLER_16_808 ();
 sg13g2_decap_8 FILLER_16_815 ();
 sg13g2_decap_8 FILLER_16_822 ();
 sg13g2_decap_4 FILLER_16_829 ();
 sg13g2_fill_2 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_897 ();
 sg13g2_decap_8 FILLER_16_904 ();
 sg13g2_decap_8 FILLER_16_911 ();
 sg13g2_decap_8 FILLER_16_918 ();
 sg13g2_decap_8 FILLER_16_925 ();
 sg13g2_fill_2 FILLER_16_932 ();
 sg13g2_fill_2 FILLER_16_938 ();
 sg13g2_fill_2 FILLER_16_966 ();
 sg13g2_fill_1 FILLER_16_968 ();
 sg13g2_fill_2 FILLER_16_995 ();
 sg13g2_decap_8 FILLER_16_1033 ();
 sg13g2_decap_8 FILLER_16_1040 ();
 sg13g2_decap_8 FILLER_16_1047 ();
 sg13g2_fill_2 FILLER_16_1054 ();
 sg13g2_fill_1 FILLER_16_1056 ();
 sg13g2_fill_2 FILLER_16_1083 ();
 sg13g2_decap_8 FILLER_16_1095 ();
 sg13g2_decap_8 FILLER_16_1102 ();
 sg13g2_decap_8 FILLER_16_1109 ();
 sg13g2_decap_4 FILLER_16_1142 ();
 sg13g2_fill_2 FILLER_16_1146 ();
 sg13g2_fill_2 FILLER_16_1174 ();
 sg13g2_decap_4 FILLER_16_1212 ();
 sg13g2_fill_2 FILLER_16_1216 ();
 sg13g2_fill_1 FILLER_16_1258 ();
 sg13g2_decap_4 FILLER_16_1263 ();
 sg13g2_decap_8 FILLER_16_1271 ();
 sg13g2_decap_8 FILLER_16_1278 ();
 sg13g2_decap_8 FILLER_16_1285 ();
 sg13g2_decap_8 FILLER_16_1292 ();
 sg13g2_decap_8 FILLER_16_1299 ();
 sg13g2_decap_8 FILLER_16_1306 ();
 sg13g2_decap_8 FILLER_16_1313 ();
 sg13g2_decap_4 FILLER_16_1320 ();
 sg13g2_fill_2 FILLER_16_1324 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_62 ();
 sg13g2_decap_8 FILLER_17_85 ();
 sg13g2_fill_2 FILLER_17_92 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_fill_2 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_decap_8 FILLER_17_241 ();
 sg13g2_decap_8 FILLER_17_248 ();
 sg13g2_decap_4 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_4 FILLER_17_340 ();
 sg13g2_fill_1 FILLER_17_344 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_fill_1 FILLER_17_393 ();
 sg13g2_fill_1 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_419 ();
 sg13g2_fill_2 FILLER_17_431 ();
 sg13g2_fill_1 FILLER_17_433 ();
 sg13g2_decap_8 FILLER_17_444 ();
 sg13g2_fill_2 FILLER_17_451 ();
 sg13g2_decap_4 FILLER_17_514 ();
 sg13g2_fill_1 FILLER_17_518 ();
 sg13g2_fill_2 FILLER_17_540 ();
 sg13g2_decap_8 FILLER_17_547 ();
 sg13g2_decap_8 FILLER_17_554 ();
 sg13g2_fill_2 FILLER_17_569 ();
 sg13g2_decap_8 FILLER_17_592 ();
 sg13g2_fill_1 FILLER_17_599 ();
 sg13g2_decap_8 FILLER_17_618 ();
 sg13g2_fill_2 FILLER_17_634 ();
 sg13g2_fill_2 FILLER_17_646 ();
 sg13g2_fill_1 FILLER_17_648 ();
 sg13g2_fill_1 FILLER_17_675 ();
 sg13g2_decap_8 FILLER_17_684 ();
 sg13g2_decap_8 FILLER_17_691 ();
 sg13g2_fill_2 FILLER_17_698 ();
 sg13g2_decap_8 FILLER_17_710 ();
 sg13g2_decap_4 FILLER_17_717 ();
 sg13g2_fill_1 FILLER_17_725 ();
 sg13g2_fill_1 FILLER_17_736 ();
 sg13g2_fill_2 FILLER_17_747 ();
 sg13g2_fill_1 FILLER_17_753 ();
 sg13g2_fill_2 FILLER_17_764 ();
 sg13g2_fill_2 FILLER_17_770 ();
 sg13g2_fill_1 FILLER_17_772 ();
 sg13g2_decap_4 FILLER_17_777 ();
 sg13g2_fill_2 FILLER_17_781 ();
 sg13g2_decap_8 FILLER_17_787 ();
 sg13g2_decap_8 FILLER_17_794 ();
 sg13g2_decap_8 FILLER_17_801 ();
 sg13g2_decap_8 FILLER_17_808 ();
 sg13g2_decap_8 FILLER_17_815 ();
 sg13g2_decap_8 FILLER_17_822 ();
 sg13g2_decap_8 FILLER_17_829 ();
 sg13g2_fill_2 FILLER_17_836 ();
 sg13g2_fill_1 FILLER_17_838 ();
 sg13g2_fill_1 FILLER_17_864 ();
 sg13g2_decap_8 FILLER_17_909 ();
 sg13g2_decap_8 FILLER_17_916 ();
 sg13g2_decap_8 FILLER_17_923 ();
 sg13g2_decap_8 FILLER_17_930 ();
 sg13g2_fill_2 FILLER_17_937 ();
 sg13g2_decap_4 FILLER_17_953 ();
 sg13g2_fill_1 FILLER_17_957 ();
 sg13g2_fill_2 FILLER_17_1044 ();
 sg13g2_fill_2 FILLER_17_1184 ();
 sg13g2_fill_2 FILLER_17_1226 ();
 sg13g2_decap_8 FILLER_17_1272 ();
 sg13g2_decap_8 FILLER_17_1279 ();
 sg13g2_decap_8 FILLER_17_1286 ();
 sg13g2_decap_8 FILLER_17_1293 ();
 sg13g2_decap_8 FILLER_17_1300 ();
 sg13g2_decap_8 FILLER_17_1307 ();
 sg13g2_decap_8 FILLER_17_1314 ();
 sg13g2_decap_4 FILLER_17_1321 ();
 sg13g2_fill_1 FILLER_17_1325 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_17 ();
 sg13g2_fill_2 FILLER_18_24 ();
 sg13g2_decap_4 FILLER_18_31 ();
 sg13g2_fill_1 FILLER_18_45 ();
 sg13g2_fill_2 FILLER_18_79 ();
 sg13g2_fill_1 FILLER_18_81 ();
 sg13g2_decap_4 FILLER_18_92 ();
 sg13g2_fill_2 FILLER_18_96 ();
 sg13g2_decap_8 FILLER_18_128 ();
 sg13g2_fill_1 FILLER_18_135 ();
 sg13g2_decap_4 FILLER_18_157 ();
 sg13g2_decap_8 FILLER_18_171 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_fill_1 FILLER_18_185 ();
 sg13g2_fill_2 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_197 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_209 ();
 sg13g2_decap_8 FILLER_18_250 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_317 ();
 sg13g2_fill_2 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_fill_2 FILLER_18_356 ();
 sg13g2_decap_4 FILLER_18_366 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_fill_1 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_446 ();
 sg13g2_fill_2 FILLER_18_453 ();
 sg13g2_fill_1 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_460 ();
 sg13g2_decap_8 FILLER_18_467 ();
 sg13g2_decap_8 FILLER_18_474 ();
 sg13g2_fill_2 FILLER_18_481 ();
 sg13g2_decap_8 FILLER_18_487 ();
 sg13g2_fill_2 FILLER_18_494 ();
 sg13g2_fill_1 FILLER_18_496 ();
 sg13g2_decap_4 FILLER_18_518 ();
 sg13g2_fill_2 FILLER_18_522 ();
 sg13g2_decap_8 FILLER_18_537 ();
 sg13g2_decap_8 FILLER_18_544 ();
 sg13g2_decap_8 FILLER_18_551 ();
 sg13g2_fill_2 FILLER_18_558 ();
 sg13g2_fill_1 FILLER_18_570 ();
 sg13g2_decap_8 FILLER_18_579 ();
 sg13g2_decap_8 FILLER_18_594 ();
 sg13g2_fill_2 FILLER_18_601 ();
 sg13g2_fill_1 FILLER_18_603 ();
 sg13g2_decap_4 FILLER_18_608 ();
 sg13g2_fill_2 FILLER_18_612 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_4 FILLER_18_637 ();
 sg13g2_fill_2 FILLER_18_651 ();
 sg13g2_fill_1 FILLER_18_653 ();
 sg13g2_decap_4 FILLER_18_667 ();
 sg13g2_decap_8 FILLER_18_681 ();
 sg13g2_decap_8 FILLER_18_688 ();
 sg13g2_fill_2 FILLER_18_695 ();
 sg13g2_fill_1 FILLER_18_697 ();
 sg13g2_decap_8 FILLER_18_702 ();
 sg13g2_decap_8 FILLER_18_709 ();
 sg13g2_decap_8 FILLER_18_746 ();
 sg13g2_decap_8 FILLER_18_753 ();
 sg13g2_decap_4 FILLER_18_760 ();
 sg13g2_fill_1 FILLER_18_764 ();
 sg13g2_fill_2 FILLER_18_773 ();
 sg13g2_fill_2 FILLER_18_835 ();
 sg13g2_fill_1 FILLER_18_837 ();
 sg13g2_fill_1 FILLER_18_852 ();
 sg13g2_fill_1 FILLER_18_889 ();
 sg13g2_decap_8 FILLER_18_920 ();
 sg13g2_decap_8 FILLER_18_927 ();
 sg13g2_fill_2 FILLER_18_934 ();
 sg13g2_fill_1 FILLER_18_936 ();
 sg13g2_decap_8 FILLER_18_947 ();
 sg13g2_fill_2 FILLER_18_954 ();
 sg13g2_fill_1 FILLER_18_956 ();
 sg13g2_fill_1 FILLER_18_991 ();
 sg13g2_fill_2 FILLER_18_996 ();
 sg13g2_fill_1 FILLER_18_998 ();
 sg13g2_fill_1 FILLER_18_1009 ();
 sg13g2_fill_2 FILLER_18_1020 ();
 sg13g2_fill_1 FILLER_18_1052 ();
 sg13g2_fill_1 FILLER_18_1057 ();
 sg13g2_fill_2 FILLER_18_1068 ();
 sg13g2_decap_4 FILLER_18_1082 ();
 sg13g2_fill_1 FILLER_18_1096 ();
 sg13g2_decap_8 FILLER_18_1101 ();
 sg13g2_decap_8 FILLER_18_1108 ();
 sg13g2_fill_2 FILLER_18_1115 ();
 sg13g2_fill_1 FILLER_18_1117 ();
 sg13g2_fill_1 FILLER_18_1122 ();
 sg13g2_fill_1 FILLER_18_1133 ();
 sg13g2_fill_1 FILLER_18_1144 ();
 sg13g2_fill_1 FILLER_18_1149 ();
 sg13g2_decap_8 FILLER_18_1228 ();
 sg13g2_decap_4 FILLER_18_1235 ();
 sg13g2_fill_1 FILLER_18_1239 ();
 sg13g2_decap_8 FILLER_18_1254 ();
 sg13g2_decap_8 FILLER_18_1261 ();
 sg13g2_fill_1 FILLER_18_1268 ();
 sg13g2_decap_8 FILLER_18_1295 ();
 sg13g2_decap_8 FILLER_18_1302 ();
 sg13g2_decap_8 FILLER_18_1309 ();
 sg13g2_decap_8 FILLER_18_1316 ();
 sg13g2_fill_2 FILLER_18_1323 ();
 sg13g2_fill_1 FILLER_18_1325 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_4 FILLER_19_63 ();
 sg13g2_fill_1 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_72 ();
 sg13g2_decap_8 FILLER_19_79 ();
 sg13g2_decap_4 FILLER_19_86 ();
 sg13g2_decap_8 FILLER_19_94 ();
 sg13g2_decap_8 FILLER_19_101 ();
 sg13g2_decap_4 FILLER_19_108 ();
 sg13g2_decap_8 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_4 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_fill_2 FILLER_19_279 ();
 sg13g2_decap_8 FILLER_19_285 ();
 sg13g2_fill_1 FILLER_19_292 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_decap_4 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_350 ();
 sg13g2_decap_4 FILLER_19_364 ();
 sg13g2_fill_1 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_457 ();
 sg13g2_decap_8 FILLER_19_464 ();
 sg13g2_decap_8 FILLER_19_471 ();
 sg13g2_decap_8 FILLER_19_478 ();
 sg13g2_fill_2 FILLER_19_485 ();
 sg13g2_fill_1 FILLER_19_487 ();
 sg13g2_decap_4 FILLER_19_492 ();
 sg13g2_decap_8 FILLER_19_557 ();
 sg13g2_decap_8 FILLER_19_568 ();
 sg13g2_decap_8 FILLER_19_575 ();
 sg13g2_decap_8 FILLER_19_582 ();
 sg13g2_decap_8 FILLER_19_597 ();
 sg13g2_decap_8 FILLER_19_604 ();
 sg13g2_fill_2 FILLER_19_611 ();
 sg13g2_fill_1 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_628 ();
 sg13g2_decap_8 FILLER_19_635 ();
 sg13g2_decap_4 FILLER_19_642 ();
 sg13g2_fill_2 FILLER_19_646 ();
 sg13g2_fill_1 FILLER_19_661 ();
 sg13g2_fill_1 FILLER_19_666 ();
 sg13g2_decap_4 FILLER_19_721 ();
 sg13g2_fill_2 FILLER_19_725 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_fill_1 FILLER_19_796 ();
 sg13g2_decap_4 FILLER_19_807 ();
 sg13g2_fill_1 FILLER_19_811 ();
 sg13g2_fill_2 FILLER_19_876 ();
 sg13g2_decap_8 FILLER_19_882 ();
 sg13g2_fill_2 FILLER_19_889 ();
 sg13g2_fill_2 FILLER_19_911 ();
 sg13g2_decap_4 FILLER_19_947 ();
 sg13g2_fill_1 FILLER_19_951 ();
 sg13g2_fill_2 FILLER_19_962 ();
 sg13g2_fill_1 FILLER_19_964 ();
 sg13g2_decap_8 FILLER_19_969 ();
 sg13g2_decap_8 FILLER_19_976 ();
 sg13g2_decap_8 FILLER_19_983 ();
 sg13g2_fill_2 FILLER_19_990 ();
 sg13g2_fill_1 FILLER_19_992 ();
 sg13g2_decap_8 FILLER_19_997 ();
 sg13g2_decap_4 FILLER_19_1004 ();
 sg13g2_fill_2 FILLER_19_1008 ();
 sg13g2_fill_1 FILLER_19_1020 ();
 sg13g2_decap_4 FILLER_19_1031 ();
 sg13g2_decap_8 FILLER_19_1039 ();
 sg13g2_decap_8 FILLER_19_1046 ();
 sg13g2_decap_8 FILLER_19_1053 ();
 sg13g2_fill_2 FILLER_19_1060 ();
 sg13g2_fill_1 FILLER_19_1062 ();
 sg13g2_decap_8 FILLER_19_1099 ();
 sg13g2_decap_8 FILLER_19_1106 ();
 sg13g2_decap_4 FILLER_19_1113 ();
 sg13g2_fill_2 FILLER_19_1117 ();
 sg13g2_decap_8 FILLER_19_1133 ();
 sg13g2_decap_8 FILLER_19_1140 ();
 sg13g2_decap_8 FILLER_19_1147 ();
 sg13g2_decap_8 FILLER_19_1154 ();
 sg13g2_decap_8 FILLER_19_1165 ();
 sg13g2_fill_2 FILLER_19_1172 ();
 sg13g2_fill_2 FILLER_19_1186 ();
 sg13g2_decap_4 FILLER_19_1214 ();
 sg13g2_fill_2 FILLER_19_1218 ();
 sg13g2_decap_4 FILLER_19_1250 ();
 sg13g2_decap_8 FILLER_19_1290 ();
 sg13g2_decap_8 FILLER_19_1297 ();
 sg13g2_decap_8 FILLER_19_1304 ();
 sg13g2_decap_8 FILLER_19_1311 ();
 sg13g2_decap_8 FILLER_19_1318 ();
 sg13g2_fill_1 FILLER_19_1325 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_20 ();
 sg13g2_fill_2 FILLER_20_51 ();
 sg13g2_fill_1 FILLER_20_53 ();
 sg13g2_fill_2 FILLER_20_64 ();
 sg13g2_fill_1 FILLER_20_66 ();
 sg13g2_fill_2 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_fill_2 FILLER_20_106 ();
 sg13g2_decap_8 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_136 ();
 sg13g2_fill_1 FILLER_20_141 ();
 sg13g2_decap_8 FILLER_20_146 ();
 sg13g2_decap_8 FILLER_20_153 ();
 sg13g2_decap_8 FILLER_20_160 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_decap_4 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_293 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_decap_8 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_314 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_4 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_fill_2 FILLER_20_449 ();
 sg13g2_fill_1 FILLER_20_451 ();
 sg13g2_fill_2 FILLER_20_462 ();
 sg13g2_fill_2 FILLER_20_485 ();
 sg13g2_fill_2 FILLER_20_523 ();
 sg13g2_fill_1 FILLER_20_525 ();
 sg13g2_fill_1 FILLER_20_530 ();
 sg13g2_decap_4 FILLER_20_540 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_fill_1 FILLER_20_611 ();
 sg13g2_fill_1 FILLER_20_622 ();
 sg13g2_decap_4 FILLER_20_631 ();
 sg13g2_fill_1 FILLER_20_635 ();
 sg13g2_decap_4 FILLER_20_657 ();
 sg13g2_decap_4 FILLER_20_665 ();
 sg13g2_fill_2 FILLER_20_669 ();
 sg13g2_fill_2 FILLER_20_681 ();
 sg13g2_fill_2 FILLER_20_709 ();
 sg13g2_fill_1 FILLER_20_737 ();
 sg13g2_fill_2 FILLER_20_764 ();
 sg13g2_fill_2 FILLER_20_792 ();
 sg13g2_fill_2 FILLER_20_820 ();
 sg13g2_decap_4 FILLER_20_846 ();
 sg13g2_fill_2 FILLER_20_912 ();
 sg13g2_decap_4 FILLER_20_950 ();
 sg13g2_decap_4 FILLER_20_980 ();
 sg13g2_fill_2 FILLER_20_984 ();
 sg13g2_decap_4 FILLER_20_1022 ();
 sg13g2_fill_2 FILLER_20_1026 ();
 sg13g2_fill_2 FILLER_20_1072 ();
 sg13g2_fill_2 FILLER_20_1078 ();
 sg13g2_decap_8 FILLER_20_1084 ();
 sg13g2_decap_8 FILLER_20_1091 ();
 sg13g2_decap_4 FILLER_20_1098 ();
 sg13g2_fill_1 FILLER_20_1102 ();
 sg13g2_decap_8 FILLER_20_1133 ();
 sg13g2_decap_8 FILLER_20_1140 ();
 sg13g2_decap_8 FILLER_20_1147 ();
 sg13g2_fill_1 FILLER_20_1154 ();
 sg13g2_decap_4 FILLER_20_1159 ();
 sg13g2_decap_8 FILLER_20_1173 ();
 sg13g2_fill_1 FILLER_20_1180 ();
 sg13g2_fill_2 FILLER_20_1201 ();
 sg13g2_fill_1 FILLER_20_1203 ();
 sg13g2_decap_8 FILLER_20_1208 ();
 sg13g2_decap_8 FILLER_20_1215 ();
 sg13g2_decap_8 FILLER_20_1222 ();
 sg13g2_fill_2 FILLER_20_1229 ();
 sg13g2_fill_1 FILLER_20_1231 ();
 sg13g2_fill_2 FILLER_20_1236 ();
 sg13g2_fill_1 FILLER_20_1238 ();
 sg13g2_fill_2 FILLER_20_1249 ();
 sg13g2_fill_1 FILLER_20_1251 ();
 sg13g2_fill_1 FILLER_20_1276 ();
 sg13g2_decap_4 FILLER_20_1281 ();
 sg13g2_fill_2 FILLER_20_1285 ();
 sg13g2_decap_8 FILLER_20_1313 ();
 sg13g2_decap_4 FILLER_20_1320 ();
 sg13g2_fill_2 FILLER_20_1324 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_fill_2 FILLER_21_20 ();
 sg13g2_fill_2 FILLER_21_26 ();
 sg13g2_fill_1 FILLER_21_90 ();
 sg13g2_fill_2 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_182 ();
 sg13g2_decap_4 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_decap_4 FILLER_21_225 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_4 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_363 ();
 sg13g2_fill_2 FILLER_21_370 ();
 sg13g2_fill_1 FILLER_21_393 ();
 sg13g2_fill_1 FILLER_21_407 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_1 FILLER_21_438 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_fill_1 FILLER_21_504 ();
 sg13g2_decap_4 FILLER_21_509 ();
 sg13g2_decap_4 FILLER_21_544 ();
 sg13g2_fill_2 FILLER_21_578 ();
 sg13g2_fill_2 FILLER_21_584 ();
 sg13g2_fill_1 FILLER_21_586 ();
 sg13g2_decap_8 FILLER_21_643 ();
 sg13g2_fill_1 FILLER_21_650 ();
 sg13g2_fill_1 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_720 ();
 sg13g2_decap_8 FILLER_21_727 ();
 sg13g2_decap_8 FILLER_21_734 ();
 sg13g2_decap_4 FILLER_21_759 ();
 sg13g2_fill_1 FILLER_21_773 ();
 sg13g2_decap_4 FILLER_21_784 ();
 sg13g2_decap_4 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_806 ();
 sg13g2_decap_8 FILLER_21_813 ();
 sg13g2_decap_4 FILLER_21_820 ();
 sg13g2_fill_2 FILLER_21_824 ();
 sg13g2_decap_4 FILLER_21_856 ();
 sg13g2_fill_1 FILLER_21_860 ();
 sg13g2_decap_8 FILLER_21_875 ();
 sg13g2_decap_8 FILLER_21_882 ();
 sg13g2_decap_4 FILLER_21_889 ();
 sg13g2_fill_1 FILLER_21_893 ();
 sg13g2_decap_4 FILLER_21_898 ();
 sg13g2_fill_2 FILLER_21_912 ();
 sg13g2_fill_1 FILLER_21_914 ();
 sg13g2_fill_2 FILLER_21_919 ();
 sg13g2_fill_1 FILLER_21_957 ();
 sg13g2_fill_2 FILLER_21_984 ();
 sg13g2_fill_1 FILLER_21_986 ();
 sg13g2_fill_1 FILLER_21_1013 ();
 sg13g2_fill_2 FILLER_21_1024 ();
 sg13g2_fill_1 FILLER_21_1026 ();
 sg13g2_fill_2 FILLER_21_1063 ();
 sg13g2_fill_1 FILLER_21_1065 ();
 sg13g2_decap_8 FILLER_21_1092 ();
 sg13g2_fill_2 FILLER_21_1099 ();
 sg13g2_decap_8 FILLER_21_1141 ();
 sg13g2_fill_2 FILLER_21_1174 ();
 sg13g2_fill_2 FILLER_21_1180 ();
 sg13g2_fill_1 FILLER_21_1182 ();
 sg13g2_fill_2 FILLER_21_1193 ();
 sg13g2_fill_1 FILLER_21_1195 ();
 sg13g2_fill_2 FILLER_21_1222 ();
 sg13g2_fill_1 FILLER_21_1224 ();
 sg13g2_decap_8 FILLER_21_1251 ();
 sg13g2_decap_8 FILLER_21_1258 ();
 sg13g2_decap_8 FILLER_21_1265 ();
 sg13g2_fill_2 FILLER_21_1272 ();
 sg13g2_decap_4 FILLER_21_1284 ();
 sg13g2_decap_8 FILLER_21_1292 ();
 sg13g2_decap_8 FILLER_21_1299 ();
 sg13g2_decap_8 FILLER_21_1306 ();
 sg13g2_decap_8 FILLER_21_1313 ();
 sg13g2_decap_4 FILLER_21_1320 ();
 sg13g2_fill_2 FILLER_21_1324 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_58 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_1 FILLER_22_101 ();
 sg13g2_decap_4 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_131 ();
 sg13g2_decap_4 FILLER_22_138 ();
 sg13g2_fill_2 FILLER_22_142 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_4 FILLER_22_334 ();
 sg13g2_decap_4 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_414 ();
 sg13g2_decap_8 FILLER_22_437 ();
 sg13g2_fill_1 FILLER_22_444 ();
 sg13g2_decap_8 FILLER_22_496 ();
 sg13g2_decap_8 FILLER_22_503 ();
 sg13g2_decap_8 FILLER_22_510 ();
 sg13g2_decap_8 FILLER_22_517 ();
 sg13g2_decap_8 FILLER_22_524 ();
 sg13g2_fill_1 FILLER_22_566 ();
 sg13g2_fill_1 FILLER_22_571 ();
 sg13g2_fill_1 FILLER_22_602 ();
 sg13g2_fill_2 FILLER_22_642 ();
 sg13g2_fill_1 FILLER_22_644 ();
 sg13g2_fill_2 FILLER_22_649 ();
 sg13g2_fill_2 FILLER_22_661 ();
 sg13g2_decap_8 FILLER_22_689 ();
 sg13g2_fill_2 FILLER_22_696 ();
 sg13g2_fill_1 FILLER_22_698 ();
 sg13g2_fill_1 FILLER_22_703 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_decap_8 FILLER_22_754 ();
 sg13g2_decap_4 FILLER_22_761 ();
 sg13g2_fill_1 FILLER_22_765 ();
 sg13g2_fill_2 FILLER_22_774 ();
 sg13g2_fill_2 FILLER_22_780 ();
 sg13g2_fill_1 FILLER_22_782 ();
 sg13g2_fill_1 FILLER_22_787 ();
 sg13g2_decap_4 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_820 ();
 sg13g2_fill_2 FILLER_22_827 ();
 sg13g2_fill_1 FILLER_22_829 ();
 sg13g2_fill_1 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_897 ();
 sg13g2_fill_2 FILLER_22_904 ();
 sg13g2_fill_1 FILLER_22_906 ();
 sg13g2_decap_4 FILLER_22_949 ();
 sg13g2_decap_8 FILLER_22_977 ();
 sg13g2_fill_2 FILLER_22_984 ();
 sg13g2_decap_4 FILLER_22_991 ();
 sg13g2_fill_1 FILLER_22_995 ();
 sg13g2_decap_8 FILLER_22_1056 ();
 sg13g2_fill_2 FILLER_22_1063 ();
 sg13g2_fill_2 FILLER_22_1109 ();
 sg13g2_fill_1 FILLER_22_1111 ();
 sg13g2_fill_1 FILLER_22_1138 ();
 sg13g2_decap_8 FILLER_22_1217 ();
 sg13g2_decap_8 FILLER_22_1224 ();
 sg13g2_decap_8 FILLER_22_1231 ();
 sg13g2_decap_8 FILLER_22_1238 ();
 sg13g2_fill_1 FILLER_22_1245 ();
 sg13g2_decap_8 FILLER_22_1260 ();
 sg13g2_decap_8 FILLER_22_1267 ();
 sg13g2_fill_1 FILLER_22_1274 ();
 sg13g2_decap_8 FILLER_22_1301 ();
 sg13g2_decap_8 FILLER_22_1308 ();
 sg13g2_decap_8 FILLER_22_1315 ();
 sg13g2_decap_4 FILLER_22_1322 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_34 ();
 sg13g2_fill_2 FILLER_23_57 ();
 sg13g2_fill_1 FILLER_23_59 ();
 sg13g2_fill_2 FILLER_23_64 ();
 sg13g2_fill_1 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_71 ();
 sg13g2_decap_8 FILLER_23_94 ();
 sg13g2_decap_8 FILLER_23_101 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_fill_2 FILLER_23_115 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_fill_2 FILLER_23_139 ();
 sg13g2_fill_1 FILLER_23_141 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_decap_4 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_317 ();
 sg13g2_decap_8 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_331 ();
 sg13g2_fill_1 FILLER_23_333 ();
 sg13g2_fill_2 FILLER_23_369 ();
 sg13g2_decap_4 FILLER_23_433 ();
 sg13g2_decap_4 FILLER_23_503 ();
 sg13g2_fill_1 FILLER_23_507 ();
 sg13g2_decap_4 FILLER_23_512 ();
 sg13g2_decap_4 FILLER_23_524 ();
 sg13g2_fill_2 FILLER_23_542 ();
 sg13g2_decap_8 FILLER_23_548 ();
 sg13g2_decap_8 FILLER_23_555 ();
 sg13g2_decap_8 FILLER_23_562 ();
 sg13g2_decap_8 FILLER_23_569 ();
 sg13g2_decap_4 FILLER_23_576 ();
 sg13g2_decap_4 FILLER_23_598 ();
 sg13g2_fill_2 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_612 ();
 sg13g2_decap_8 FILLER_23_619 ();
 sg13g2_decap_4 FILLER_23_630 ();
 sg13g2_fill_2 FILLER_23_634 ();
 sg13g2_fill_1 FILLER_23_640 ();
 sg13g2_fill_2 FILLER_23_662 ();
 sg13g2_fill_1 FILLER_23_664 ();
 sg13g2_decap_8 FILLER_23_675 ();
 sg13g2_decap_8 FILLER_23_729 ();
 sg13g2_decap_4 FILLER_23_736 ();
 sg13g2_fill_2 FILLER_23_740 ();
 sg13g2_decap_4 FILLER_23_766 ();
 sg13g2_decap_8 FILLER_23_822 ();
 sg13g2_fill_2 FILLER_23_829 ();
 sg13g2_decap_4 FILLER_23_861 ();
 sg13g2_fill_1 FILLER_23_865 ();
 sg13g2_decap_8 FILLER_23_922 ();
 sg13g2_fill_2 FILLER_23_929 ();
 sg13g2_fill_1 FILLER_23_931 ();
 sg13g2_decap_8 FILLER_23_940 ();
 sg13g2_decap_8 FILLER_23_973 ();
 sg13g2_decap_8 FILLER_23_980 ();
 sg13g2_fill_2 FILLER_23_987 ();
 sg13g2_fill_1 FILLER_23_989 ();
 sg13g2_decap_8 FILLER_23_994 ();
 sg13g2_fill_2 FILLER_23_1001 ();
 sg13g2_fill_1 FILLER_23_1003 ();
 sg13g2_decap_8 FILLER_23_1008 ();
 sg13g2_fill_2 FILLER_23_1015 ();
 sg13g2_fill_1 FILLER_23_1017 ();
 sg13g2_decap_8 FILLER_23_1046 ();
 sg13g2_decap_8 FILLER_23_1053 ();
 sg13g2_decap_8 FILLER_23_1060 ();
 sg13g2_fill_2 FILLER_23_1067 ();
 sg13g2_fill_1 FILLER_23_1069 ();
 sg13g2_decap_8 FILLER_23_1100 ();
 sg13g2_fill_1 FILLER_23_1107 ();
 sg13g2_decap_4 FILLER_23_1112 ();
 sg13g2_decap_4 FILLER_23_1130 ();
 sg13g2_fill_1 FILLER_23_1134 ();
 sg13g2_decap_8 FILLER_23_1149 ();
 sg13g2_decap_8 FILLER_23_1156 ();
 sg13g2_decap_4 FILLER_23_1173 ();
 sg13g2_fill_2 FILLER_23_1187 ();
 sg13g2_fill_1 FILLER_23_1189 ();
 sg13g2_fill_1 FILLER_23_1194 ();
 sg13g2_fill_1 FILLER_23_1229 ();
 sg13g2_decap_4 FILLER_23_1256 ();
 sg13g2_fill_2 FILLER_23_1260 ();
 sg13g2_decap_8 FILLER_23_1298 ();
 sg13g2_decap_8 FILLER_23_1305 ();
 sg13g2_decap_8 FILLER_23_1312 ();
 sg13g2_decap_8 FILLER_23_1319 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_16 ();
 sg13g2_decap_4 FILLER_24_23 ();
 sg13g2_fill_2 FILLER_24_31 ();
 sg13g2_fill_1 FILLER_24_41 ();
 sg13g2_decap_4 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_55 ();
 sg13g2_decap_8 FILLER_24_62 ();
 sg13g2_decap_8 FILLER_24_90 ();
 sg13g2_decap_8 FILLER_24_97 ();
 sg13g2_decap_8 FILLER_24_104 ();
 sg13g2_decap_8 FILLER_24_111 ();
 sg13g2_decap_4 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_decap_8 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_187 ();
 sg13g2_fill_2 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_4 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_4 FILLER_24_268 ();
 sg13g2_decap_4 FILLER_24_276 ();
 sg13g2_decap_4 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_339 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_fill_2 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_407 ();
 sg13g2_fill_2 FILLER_24_415 ();
 sg13g2_fill_2 FILLER_24_421 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_4 FILLER_24_434 ();
 sg13g2_fill_2 FILLER_24_438 ();
 sg13g2_decap_4 FILLER_24_454 ();
 sg13g2_fill_2 FILLER_24_494 ();
 sg13g2_decap_8 FILLER_24_501 ();
 sg13g2_decap_8 FILLER_24_508 ();
 sg13g2_decap_4 FILLER_24_515 ();
 sg13g2_decap_8 FILLER_24_563 ();
 sg13g2_decap_8 FILLER_24_570 ();
 sg13g2_decap_8 FILLER_24_577 ();
 sg13g2_decap_8 FILLER_24_613 ();
 sg13g2_fill_1 FILLER_24_624 ();
 sg13g2_decap_4 FILLER_24_635 ();
 sg13g2_decap_4 FILLER_24_644 ();
 sg13g2_fill_1 FILLER_24_648 ();
 sg13g2_fill_1 FILLER_24_653 ();
 sg13g2_fill_1 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_720 ();
 sg13g2_decap_8 FILLER_24_727 ();
 sg13g2_fill_2 FILLER_24_734 ();
 sg13g2_fill_1 FILLER_24_798 ();
 sg13g2_decap_4 FILLER_24_835 ();
 sg13g2_fill_1 FILLER_24_839 ();
 sg13g2_fill_1 FILLER_24_844 ();
 sg13g2_fill_1 FILLER_24_855 ();
 sg13g2_fill_1 FILLER_24_866 ();
 sg13g2_fill_2 FILLER_24_877 ();
 sg13g2_decap_8 FILLER_24_891 ();
 sg13g2_decap_4 FILLER_24_898 ();
 sg13g2_fill_1 FILLER_24_902 ();
 sg13g2_decap_4 FILLER_24_907 ();
 sg13g2_fill_2 FILLER_24_911 ();
 sg13g2_decap_4 FILLER_24_923 ();
 sg13g2_fill_2 FILLER_24_927 ();
 sg13g2_fill_2 FILLER_24_937 ();
 sg13g2_fill_1 FILLER_24_939 ();
 sg13g2_decap_4 FILLER_24_950 ();
 sg13g2_fill_1 FILLER_24_954 ();
 sg13g2_fill_2 FILLER_24_969 ();
 sg13g2_decap_4 FILLER_24_1007 ();
 sg13g2_fill_1 FILLER_24_1011 ();
 sg13g2_decap_8 FILLER_24_1020 ();
 sg13g2_fill_2 FILLER_24_1027 ();
 sg13g2_fill_2 FILLER_24_1049 ();
 sg13g2_decap_4 FILLER_24_1061 ();
 sg13g2_decap_8 FILLER_24_1091 ();
 sg13g2_decap_8 FILLER_24_1098 ();
 sg13g2_decap_8 FILLER_24_1105 ();
 sg13g2_decap_8 FILLER_24_1116 ();
 sg13g2_fill_2 FILLER_24_1123 ();
 sg13g2_fill_1 FILLER_24_1125 ();
 sg13g2_decap_4 FILLER_24_1136 ();
 sg13g2_fill_1 FILLER_24_1140 ();
 sg13g2_decap_8 FILLER_24_1145 ();
 sg13g2_decap_8 FILLER_24_1152 ();
 sg13g2_fill_2 FILLER_24_1159 ();
 sg13g2_decap_8 FILLER_24_1187 ();
 sg13g2_fill_2 FILLER_24_1194 ();
 sg13g2_fill_1 FILLER_24_1200 ();
 sg13g2_fill_1 FILLER_24_1237 ();
 sg13g2_decap_8 FILLER_24_1294 ();
 sg13g2_decap_8 FILLER_24_1301 ();
 sg13g2_decap_8 FILLER_24_1308 ();
 sg13g2_decap_8 FILLER_24_1315 ();
 sg13g2_decap_4 FILLER_24_1322 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_20 ();
 sg13g2_fill_1 FILLER_25_27 ();
 sg13g2_fill_2 FILLER_25_59 ();
 sg13g2_fill_1 FILLER_25_61 ();
 sg13g2_decap_4 FILLER_25_66 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_92 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_fill_2 FILLER_25_125 ();
 sg13g2_decap_8 FILLER_25_132 ();
 sg13g2_decap_8 FILLER_25_139 ();
 sg13g2_decap_8 FILLER_25_146 ();
 sg13g2_decap_8 FILLER_25_153 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_fill_1 FILLER_25_182 ();
 sg13g2_decap_4 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_221 ();
 sg13g2_decap_4 FILLER_25_228 ();
 sg13g2_fill_1 FILLER_25_232 ();
 sg13g2_decap_4 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_275 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_363 ();
 sg13g2_fill_1 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_fill_1 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_414 ();
 sg13g2_fill_1 FILLER_25_425 ();
 sg13g2_fill_1 FILLER_25_430 ();
 sg13g2_fill_2 FILLER_25_435 ();
 sg13g2_fill_1 FILLER_25_447 ();
 sg13g2_decap_8 FILLER_25_452 ();
 sg13g2_fill_2 FILLER_25_459 ();
 sg13g2_fill_1 FILLER_25_461 ();
 sg13g2_fill_1 FILLER_25_466 ();
 sg13g2_fill_2 FILLER_25_488 ();
 sg13g2_fill_2 FILLER_25_498 ();
 sg13g2_fill_1 FILLER_25_500 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_fill_2 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_590 ();
 sg13g2_fill_1 FILLER_25_597 ();
 sg13g2_fill_1 FILLER_25_628 ();
 sg13g2_decap_8 FILLER_25_655 ();
 sg13g2_fill_1 FILLER_25_662 ();
 sg13g2_fill_1 FILLER_25_673 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_4 FILLER_25_728 ();
 sg13g2_fill_2 FILLER_25_732 ();
 sg13g2_fill_2 FILLER_25_764 ();
 sg13g2_fill_1 FILLER_25_766 ();
 sg13g2_fill_2 FILLER_25_823 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_8 FILLER_25_856 ();
 sg13g2_fill_1 FILLER_25_863 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_decap_8 FILLER_25_875 ();
 sg13g2_decap_8 FILLER_25_882 ();
 sg13g2_fill_1 FILLER_25_889 ();
 sg13g2_decap_4 FILLER_25_900 ();
 sg13g2_decap_8 FILLER_25_908 ();
 sg13g2_decap_8 FILLER_25_915 ();
 sg13g2_fill_1 FILLER_25_922 ();
 sg13g2_fill_1 FILLER_25_953 ();
 sg13g2_fill_1 FILLER_25_980 ();
 sg13g2_fill_1 FILLER_25_991 ();
 sg13g2_fill_2 FILLER_25_1018 ();
 sg13g2_decap_4 FILLER_25_1050 ();
 sg13g2_decap_8 FILLER_25_1090 ();
 sg13g2_decap_4 FILLER_25_1097 ();
 sg13g2_fill_1 FILLER_25_1101 ();
 sg13g2_decap_4 FILLER_25_1158 ();
 sg13g2_fill_1 FILLER_25_1170 ();
 sg13g2_decap_8 FILLER_25_1175 ();
 sg13g2_decap_8 FILLER_25_1182 ();
 sg13g2_decap_8 FILLER_25_1189 ();
 sg13g2_decap_8 FILLER_25_1196 ();
 sg13g2_fill_2 FILLER_25_1203 ();
 sg13g2_decap_8 FILLER_25_1229 ();
 sg13g2_fill_1 FILLER_25_1236 ();
 sg13g2_decap_4 FILLER_25_1241 ();
 sg13g2_decap_4 FILLER_25_1253 ();
 sg13g2_fill_1 FILLER_25_1281 ();
 sg13g2_decap_8 FILLER_25_1286 ();
 sg13g2_fill_2 FILLER_25_1293 ();
 sg13g2_fill_1 FILLER_25_1295 ();
 sg13g2_decap_8 FILLER_25_1304 ();
 sg13g2_decap_8 FILLER_25_1311 ();
 sg13g2_decap_8 FILLER_25_1318 ();
 sg13g2_fill_1 FILLER_25_1325 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_31 ();
 sg13g2_decap_4 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_fill_1 FILLER_26_78 ();
 sg13g2_fill_2 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_128 ();
 sg13g2_decap_4 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_fill_2 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_205 ();
 sg13g2_decap_8 FILLER_26_212 ();
 sg13g2_decap_4 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_fill_1 FILLER_26_261 ();
 sg13g2_decap_4 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_4 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_403 ();
 sg13g2_fill_1 FILLER_26_413 ();
 sg13g2_fill_1 FILLER_26_418 ();
 sg13g2_fill_2 FILLER_26_445 ();
 sg13g2_fill_2 FILLER_26_457 ();
 sg13g2_fill_1 FILLER_26_459 ();
 sg13g2_decap_4 FILLER_26_470 ();
 sg13g2_decap_4 FILLER_26_545 ();
 sg13g2_decap_8 FILLER_26_570 ();
 sg13g2_fill_1 FILLER_26_577 ();
 sg13g2_fill_1 FILLER_26_590 ();
 sg13g2_decap_8 FILLER_26_664 ();
 sg13g2_fill_1 FILLER_26_671 ();
 sg13g2_decap_4 FILLER_26_676 ();
 sg13g2_decap_8 FILLER_26_688 ();
 sg13g2_decap_4 FILLER_26_695 ();
 sg13g2_fill_2 FILLER_26_703 ();
 sg13g2_decap_8 FILLER_26_715 ();
 sg13g2_decap_8 FILLER_26_722 ();
 sg13g2_decap_8 FILLER_26_729 ();
 sg13g2_decap_4 FILLER_26_736 ();
 sg13g2_fill_2 FILLER_26_740 ();
 sg13g2_fill_2 FILLER_26_750 ();
 sg13g2_fill_1 FILLER_26_752 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_4 FILLER_26_770 ();
 sg13g2_fill_1 FILLER_26_774 ();
 sg13g2_decap_8 FILLER_26_779 ();
 sg13g2_decap_8 FILLER_26_786 ();
 sg13g2_decap_4 FILLER_26_793 ();
 sg13g2_fill_1 FILLER_26_797 ();
 sg13g2_fill_1 FILLER_26_810 ();
 sg13g2_fill_1 FILLER_26_821 ();
 sg13g2_fill_2 FILLER_26_894 ();
 sg13g2_fill_1 FILLER_26_896 ();
 sg13g2_fill_2 FILLER_26_923 ();
 sg13g2_fill_1 FILLER_26_925 ();
 sg13g2_fill_1 FILLER_26_930 ();
 sg13g2_fill_2 FILLER_26_957 ();
 sg13g2_fill_1 FILLER_26_959 ();
 sg13g2_decap_8 FILLER_26_964 ();
 sg13g2_fill_2 FILLER_26_971 ();
 sg13g2_fill_1 FILLER_26_973 ();
 sg13g2_fill_2 FILLER_26_1014 ();
 sg13g2_fill_1 FILLER_26_1016 ();
 sg13g2_decap_4 FILLER_26_1021 ();
 sg13g2_fill_2 FILLER_26_1025 ();
 sg13g2_decap_4 FILLER_26_1057 ();
 sg13g2_fill_2 FILLER_26_1061 ();
 sg13g2_decap_8 FILLER_26_1081 ();
 sg13g2_decap_8 FILLER_26_1088 ();
 sg13g2_fill_2 FILLER_26_1095 ();
 sg13g2_fill_1 FILLER_26_1097 ();
 sg13g2_decap_4 FILLER_26_1134 ();
 sg13g2_fill_2 FILLER_26_1208 ();
 sg13g2_fill_1 FILLER_26_1214 ();
 sg13g2_fill_2 FILLER_26_1255 ();
 sg13g2_decap_8 FILLER_26_1261 ();
 sg13g2_decap_8 FILLER_26_1268 ();
 sg13g2_decap_8 FILLER_26_1275 ();
 sg13g2_fill_1 FILLER_26_1282 ();
 sg13g2_fill_2 FILLER_26_1323 ();
 sg13g2_fill_1 FILLER_26_1325 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_5 ();
 sg13g2_fill_1 FILLER_27_10 ();
 sg13g2_decap_4 FILLER_27_37 ();
 sg13g2_fill_2 FILLER_27_41 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_165 ();
 sg13g2_fill_2 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_287 ();
 sg13g2_decap_4 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_318 ();
 sg13g2_fill_2 FILLER_27_325 ();
 sg13g2_fill_1 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_fill_1 FILLER_27_405 ();
 sg13g2_fill_1 FILLER_27_416 ();
 sg13g2_fill_1 FILLER_27_469 ();
 sg13g2_fill_1 FILLER_27_540 ();
 sg13g2_fill_1 FILLER_27_562 ();
 sg13g2_fill_2 FILLER_27_583 ();
 sg13g2_fill_2 FILLER_27_606 ();
 sg13g2_fill_2 FILLER_27_612 ();
 sg13g2_fill_1 FILLER_27_618 ();
 sg13g2_fill_2 FILLER_27_629 ();
 sg13g2_fill_1 FILLER_27_631 ();
 sg13g2_decap_8 FILLER_27_657 ();
 sg13g2_decap_8 FILLER_27_664 ();
 sg13g2_decap_8 FILLER_27_671 ();
 sg13g2_decap_8 FILLER_27_678 ();
 sg13g2_decap_8 FILLER_27_685 ();
 sg13g2_decap_8 FILLER_27_692 ();
 sg13g2_fill_2 FILLER_27_699 ();
 sg13g2_fill_1 FILLER_27_701 ();
 sg13g2_decap_8 FILLER_27_771 ();
 sg13g2_decap_8 FILLER_27_778 ();
 sg13g2_decap_8 FILLER_27_785 ();
 sg13g2_decap_4 FILLER_27_792 ();
 sg13g2_fill_2 FILLER_27_796 ();
 sg13g2_fill_1 FILLER_27_808 ();
 sg13g2_fill_2 FILLER_27_887 ();
 sg13g2_decap_8 FILLER_27_929 ();
 sg13g2_fill_1 FILLER_27_936 ();
 sg13g2_decap_8 FILLER_27_947 ();
 sg13g2_decap_4 FILLER_27_954 ();
 sg13g2_decap_4 FILLER_27_970 ();
 sg13g2_fill_2 FILLER_27_974 ();
 sg13g2_decap_8 FILLER_27_1020 ();
 sg13g2_decap_8 FILLER_27_1027 ();
 sg13g2_decap_8 FILLER_27_1034 ();
 sg13g2_fill_1 FILLER_27_1041 ();
 sg13g2_decap_8 FILLER_27_1050 ();
 sg13g2_decap_4 FILLER_27_1057 ();
 sg13g2_fill_2 FILLER_27_1061 ();
 sg13g2_fill_2 FILLER_27_1099 ();
 sg13g2_fill_1 FILLER_27_1101 ();
 sg13g2_fill_2 FILLER_27_1148 ();
 sg13g2_fill_1 FILLER_27_1150 ();
 sg13g2_fill_1 FILLER_27_1177 ();
 sg13g2_fill_1 FILLER_27_1204 ();
 sg13g2_fill_1 FILLER_27_1225 ();
 sg13g2_decap_8 FILLER_27_1252 ();
 sg13g2_decap_8 FILLER_27_1259 ();
 sg13g2_fill_1 FILLER_27_1266 ();
 sg13g2_fill_1 FILLER_27_1281 ();
 sg13g2_decap_4 FILLER_27_1322 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_8 ();
 sg13g2_fill_2 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_55 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_decap_4 FILLER_28_65 ();
 sg13g2_fill_2 FILLER_28_69 ();
 sg13g2_fill_2 FILLER_28_94 ();
 sg13g2_fill_1 FILLER_28_117 ();
 sg13g2_fill_2 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_171 ();
 sg13g2_fill_2 FILLER_28_181 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_248 ();
 sg13g2_decap_4 FILLER_28_337 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_decap_4 FILLER_28_356 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_fill_2 FILLER_28_374 ();
 sg13g2_fill_1 FILLER_28_397 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_28_414 ();
 sg13g2_fill_1 FILLER_28_421 ();
 sg13g2_fill_1 FILLER_28_432 ();
 sg13g2_fill_1 FILLER_28_454 ();
 sg13g2_fill_1 FILLER_28_485 ();
 sg13g2_fill_2 FILLER_28_496 ();
 sg13g2_fill_1 FILLER_28_524 ();
 sg13g2_fill_1 FILLER_28_551 ();
 sg13g2_decap_4 FILLER_28_573 ();
 sg13g2_fill_1 FILLER_28_577 ();
 sg13g2_fill_2 FILLER_28_609 ();
 sg13g2_fill_2 FILLER_28_624 ();
 sg13g2_decap_8 FILLER_28_640 ();
 sg13g2_decap_8 FILLER_28_647 ();
 sg13g2_decap_4 FILLER_28_654 ();
 sg13g2_fill_2 FILLER_28_658 ();
 sg13g2_fill_1 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_675 ();
 sg13g2_fill_1 FILLER_28_682 ();
 sg13g2_decap_8 FILLER_28_687 ();
 sg13g2_decap_8 FILLER_28_694 ();
 sg13g2_decap_4 FILLER_28_701 ();
 sg13g2_fill_1 FILLER_28_705 ();
 sg13g2_decap_4 FILLER_28_732 ();
 sg13g2_fill_2 FILLER_28_736 ();
 sg13g2_decap_8 FILLER_28_768 ();
 sg13g2_fill_1 FILLER_28_775 ();
 sg13g2_fill_2 FILLER_28_812 ();
 sg13g2_fill_1 FILLER_28_814 ();
 sg13g2_decap_8 FILLER_28_853 ();
 sg13g2_decap_8 FILLER_28_860 ();
 sg13g2_fill_1 FILLER_28_867 ();
 sg13g2_decap_4 FILLER_28_872 ();
 sg13g2_fill_2 FILLER_28_876 ();
 sg13g2_decap_4 FILLER_28_896 ();
 sg13g2_fill_2 FILLER_28_910 ();
 sg13g2_fill_1 FILLER_28_912 ();
 sg13g2_decap_4 FILLER_28_939 ();
 sg13g2_fill_1 FILLER_28_943 ();
 sg13g2_fill_1 FILLER_28_948 ();
 sg13g2_fill_1 FILLER_28_975 ();
 sg13g2_fill_2 FILLER_28_986 ();
 sg13g2_fill_1 FILLER_28_998 ();
 sg13g2_fill_2 FILLER_28_1003 ();
 sg13g2_decap_8 FILLER_28_1009 ();
 sg13g2_decap_8 FILLER_28_1016 ();
 sg13g2_fill_2 FILLER_28_1023 ();
 sg13g2_fill_1 FILLER_28_1025 ();
 sg13g2_decap_8 FILLER_28_1052 ();
 sg13g2_decap_4 FILLER_28_1059 ();
 sg13g2_fill_2 FILLER_28_1063 ();
 sg13g2_decap_8 FILLER_28_1095 ();
 sg13g2_decap_8 FILLER_28_1102 ();
 sg13g2_fill_2 FILLER_28_1109 ();
 sg13g2_fill_1 FILLER_28_1111 ();
 sg13g2_decap_8 FILLER_28_1116 ();
 sg13g2_fill_2 FILLER_28_1123 ();
 sg13g2_fill_1 FILLER_28_1125 ();
 sg13g2_decap_4 FILLER_28_1136 ();
 sg13g2_fill_2 FILLER_28_1140 ();
 sg13g2_fill_1 FILLER_28_1146 ();
 sg13g2_fill_1 FILLER_28_1157 ();
 sg13g2_fill_1 FILLER_28_1172 ();
 sg13g2_fill_1 FILLER_28_1177 ();
 sg13g2_decap_8 FILLER_28_1248 ();
 sg13g2_decap_8 FILLER_28_1255 ();
 sg13g2_fill_2 FILLER_28_1266 ();
 sg13g2_fill_1 FILLER_28_1268 ();
 sg13g2_decap_8 FILLER_28_1295 ();
 sg13g2_decap_4 FILLER_28_1302 ();
 sg13g2_fill_1 FILLER_28_1306 ();
 sg13g2_decap_8 FILLER_28_1311 ();
 sg13g2_decap_8 FILLER_28_1318 ();
 sg13g2_fill_1 FILLER_28_1325 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_11 ();
 sg13g2_fill_1 FILLER_29_16 ();
 sg13g2_decap_8 FILLER_29_31 ();
 sg13g2_fill_2 FILLER_29_38 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_decap_8 FILLER_29_90 ();
 sg13g2_decap_8 FILLER_29_97 ();
 sg13g2_decap_8 FILLER_29_104 ();
 sg13g2_decap_4 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_195 ();
 sg13g2_decap_4 FILLER_29_201 ();
 sg13g2_fill_2 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_275 ();
 sg13g2_decap_8 FILLER_29_282 ();
 sg13g2_decap_8 FILLER_29_289 ();
 sg13g2_decap_4 FILLER_29_296 ();
 sg13g2_decap_4 FILLER_29_333 ();
 sg13g2_fill_1 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_4 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_359 ();
 sg13g2_decap_8 FILLER_29_366 ();
 sg13g2_fill_2 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_29_409 ();
 sg13g2_decap_4 FILLER_29_416 ();
 sg13g2_fill_2 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_430 ();
 sg13g2_fill_1 FILLER_29_432 ();
 sg13g2_decap_8 FILLER_29_446 ();
 sg13g2_fill_2 FILLER_29_457 ();
 sg13g2_fill_2 FILLER_29_467 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_490 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_decap_4 FILLER_29_508 ();
 sg13g2_fill_1 FILLER_29_512 ();
 sg13g2_fill_2 FILLER_29_517 ();
 sg13g2_fill_1 FILLER_29_519 ();
 sg13g2_decap_4 FILLER_29_539 ();
 sg13g2_decap_4 FILLER_29_564 ();
 sg13g2_fill_1 FILLER_29_568 ();
 sg13g2_decap_4 FILLER_29_590 ();
 sg13g2_decap_4 FILLER_29_615 ();
 sg13g2_fill_1 FILLER_29_619 ();
 sg13g2_decap_8 FILLER_29_624 ();
 sg13g2_decap_4 FILLER_29_631 ();
 sg13g2_fill_1 FILLER_29_635 ();
 sg13g2_fill_1 FILLER_29_665 ();
 sg13g2_fill_2 FILLER_29_707 ();
 sg13g2_decap_4 FILLER_29_730 ();
 sg13g2_fill_1 FILLER_29_734 ();
 sg13g2_fill_2 FILLER_29_805 ();
 sg13g2_fill_1 FILLER_29_807 ();
 sg13g2_decap_8 FILLER_29_834 ();
 sg13g2_decap_8 FILLER_29_841 ();
 sg13g2_decap_8 FILLER_29_848 ();
 sg13g2_decap_8 FILLER_29_855 ();
 sg13g2_fill_1 FILLER_29_888 ();
 sg13g2_fill_1 FILLER_29_925 ();
 sg13g2_fill_2 FILLER_29_962 ();
 sg13g2_fill_2 FILLER_29_990 ();
 sg13g2_fill_2 FILLER_29_1018 ();
 sg13g2_fill_1 FILLER_29_1060 ();
 sg13g2_decap_8 FILLER_29_1096 ();
 sg13g2_decap_8 FILLER_29_1103 ();
 sg13g2_fill_2 FILLER_29_1110 ();
 sg13g2_fill_1 FILLER_29_1112 ();
 sg13g2_decap_4 FILLER_29_1139 ();
 sg13g2_fill_2 FILLER_29_1143 ();
 sg13g2_fill_2 FILLER_29_1149 ();
 sg13g2_fill_1 FILLER_29_1151 ();
 sg13g2_decap_8 FILLER_29_1160 ();
 sg13g2_decap_8 FILLER_29_1167 ();
 sg13g2_decap_8 FILLER_29_1174 ();
 sg13g2_fill_1 FILLER_29_1181 ();
 sg13g2_fill_2 FILLER_29_1194 ();
 sg13g2_fill_1 FILLER_29_1196 ();
 sg13g2_fill_2 FILLER_29_1233 ();
 sg13g2_fill_1 FILLER_29_1235 ();
 sg13g2_decap_4 FILLER_29_1284 ();
 sg13g2_fill_2 FILLER_29_1298 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_32 ();
 sg13g2_decap_4 FILLER_30_37 ();
 sg13g2_decap_8 FILLER_30_45 ();
 sg13g2_fill_2 FILLER_30_52 ();
 sg13g2_decap_8 FILLER_30_58 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_4 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_127 ();
 sg13g2_decap_8 FILLER_30_134 ();
 sg13g2_fill_1 FILLER_30_141 ();
 sg13g2_decap_8 FILLER_30_146 ();
 sg13g2_decap_8 FILLER_30_153 ();
 sg13g2_decap_8 FILLER_30_160 ();
 sg13g2_decap_8 FILLER_30_167 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_decap_4 FILLER_30_211 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_fill_2 FILLER_30_246 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_4 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_329 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_decap_4 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_362 ();
 sg13g2_fill_2 FILLER_30_384 ();
 sg13g2_fill_2 FILLER_30_412 ();
 sg13g2_decap_4 FILLER_30_418 ();
 sg13g2_fill_1 FILLER_30_422 ();
 sg13g2_fill_2 FILLER_30_440 ();
 sg13g2_fill_1 FILLER_30_447 ();
 sg13g2_fill_2 FILLER_30_452 ();
 sg13g2_fill_1 FILLER_30_454 ();
 sg13g2_decap_4 FILLER_30_459 ();
 sg13g2_fill_2 FILLER_30_463 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_fill_2 FILLER_30_511 ();
 sg13g2_fill_1 FILLER_30_513 ();
 sg13g2_fill_2 FILLER_30_519 ();
 sg13g2_fill_2 FILLER_30_525 ();
 sg13g2_fill_1 FILLER_30_527 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_fill_2 FILLER_30_539 ();
 sg13g2_fill_1 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_573 ();
 sg13g2_decap_8 FILLER_30_580 ();
 sg13g2_decap_8 FILLER_30_587 ();
 sg13g2_fill_1 FILLER_30_594 ();
 sg13g2_decap_8 FILLER_30_603 ();
 sg13g2_decap_8 FILLER_30_614 ();
 sg13g2_fill_1 FILLER_30_621 ();
 sg13g2_fill_2 FILLER_30_626 ();
 sg13g2_fill_2 FILLER_30_636 ();
 sg13g2_fill_1 FILLER_30_638 ();
 sg13g2_fill_1 FILLER_30_649 ();
 sg13g2_fill_2 FILLER_30_671 ();
 sg13g2_fill_1 FILLER_30_673 ();
 sg13g2_fill_1 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_743 ();
 sg13g2_decap_4 FILLER_30_750 ();
 sg13g2_fill_1 FILLER_30_754 ();
 sg13g2_fill_1 FILLER_30_765 ();
 sg13g2_decap_4 FILLER_30_806 ();
 sg13g2_fill_1 FILLER_30_810 ();
 sg13g2_fill_2 FILLER_30_825 ();
 sg13g2_fill_1 FILLER_30_827 ();
 sg13g2_fill_2 FILLER_30_838 ();
 sg13g2_fill_2 FILLER_30_907 ();
 sg13g2_fill_2 FILLER_30_923 ();
 sg13g2_fill_1 FILLER_30_925 ();
 sg13g2_fill_2 FILLER_30_942 ();
 sg13g2_decap_8 FILLER_30_968 ();
 sg13g2_fill_1 FILLER_30_975 ();
 sg13g2_fill_1 FILLER_30_980 ();
 sg13g2_decap_8 FILLER_30_1007 ();
 sg13g2_decap_4 FILLER_30_1014 ();
 sg13g2_decap_8 FILLER_30_1082 ();
 sg13g2_decap_8 FILLER_30_1089 ();
 sg13g2_decap_8 FILLER_30_1096 ();
 sg13g2_decap_4 FILLER_30_1113 ();
 sg13g2_fill_2 FILLER_30_1117 ();
 sg13g2_decap_4 FILLER_30_1123 ();
 sg13g2_decap_8 FILLER_30_1141 ();
 sg13g2_decap_8 FILLER_30_1148 ();
 sg13g2_decap_8 FILLER_30_1155 ();
 sg13g2_fill_2 FILLER_30_1162 ();
 sg13g2_fill_1 FILLER_30_1164 ();
 sg13g2_decap_8 FILLER_30_1183 ();
 sg13g2_decap_8 FILLER_30_1190 ();
 sg13g2_decap_4 FILLER_30_1197 ();
 sg13g2_fill_2 FILLER_30_1201 ();
 sg13g2_decap_8 FILLER_30_1207 ();
 sg13g2_decap_8 FILLER_30_1214 ();
 sg13g2_fill_1 FILLER_30_1221 ();
 sg13g2_decap_8 FILLER_30_1227 ();
 sg13g2_fill_2 FILLER_30_1234 ();
 sg13g2_fill_1 FILLER_30_1236 ();
 sg13g2_fill_2 FILLER_30_1241 ();
 sg13g2_decap_8 FILLER_30_1279 ();
 sg13g2_fill_1 FILLER_30_1286 ();
 sg13g2_fill_2 FILLER_30_1297 ();
 sg13g2_fill_1 FILLER_30_1299 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_38 ();
 sg13g2_decap_8 FILLER_31_106 ();
 sg13g2_decap_4 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_117 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_8 FILLER_31_167 ();
 sg13g2_decap_8 FILLER_31_174 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_fill_2 FILLER_31_220 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_254 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_4 FILLER_31_406 ();
 sg13g2_fill_2 FILLER_31_410 ();
 sg13g2_decap_4 FILLER_31_422 ();
 sg13g2_decap_4 FILLER_31_452 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_4 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_508 ();
 sg13g2_decap_8 FILLER_31_515 ();
 sg13g2_fill_1 FILLER_31_522 ();
 sg13g2_decap_8 FILLER_31_527 ();
 sg13g2_decap_8 FILLER_31_534 ();
 sg13g2_decap_4 FILLER_31_541 ();
 sg13g2_fill_1 FILLER_31_545 ();
 sg13g2_decap_8 FILLER_31_550 ();
 sg13g2_decap_8 FILLER_31_557 ();
 sg13g2_decap_8 FILLER_31_564 ();
 sg13g2_decap_8 FILLER_31_571 ();
 sg13g2_fill_1 FILLER_31_578 ();
 sg13g2_fill_1 FILLER_31_583 ();
 sg13g2_fill_1 FILLER_31_588 ();
 sg13g2_fill_1 FILLER_31_607 ();
 sg13g2_fill_1 FILLER_31_652 ();
 sg13g2_fill_2 FILLER_31_692 ();
 sg13g2_fill_1 FILLER_31_694 ();
 sg13g2_fill_2 FILLER_31_705 ();
 sg13g2_decap_8 FILLER_31_738 ();
 sg13g2_decap_8 FILLER_31_745 ();
 sg13g2_decap_8 FILLER_31_752 ();
 sg13g2_decap_8 FILLER_31_759 ();
 sg13g2_decap_8 FILLER_31_766 ();
 sg13g2_decap_8 FILLER_31_773 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_fill_2 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_832 ();
 sg13g2_decap_8 FILLER_31_839 ();
 sg13g2_fill_1 FILLER_31_846 ();
 sg13g2_decap_8 FILLER_31_851 ();
 sg13g2_decap_8 FILLER_31_858 ();
 sg13g2_decap_4 FILLER_31_865 ();
 sg13g2_fill_1 FILLER_31_869 ();
 sg13g2_fill_1 FILLER_31_874 ();
 sg13g2_fill_2 FILLER_31_901 ();
 sg13g2_fill_1 FILLER_31_903 ();
 sg13g2_fill_2 FILLER_31_930 ();
 sg13g2_fill_1 FILLER_31_932 ();
 sg13g2_decap_8 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_966 ();
 sg13g2_decap_8 FILLER_31_973 ();
 sg13g2_decap_8 FILLER_31_980 ();
 sg13g2_fill_2 FILLER_31_987 ();
 sg13g2_fill_1 FILLER_31_989 ();
 sg13g2_decap_8 FILLER_31_994 ();
 sg13g2_decap_8 FILLER_31_1001 ();
 sg13g2_decap_8 FILLER_31_1008 ();
 sg13g2_decap_8 FILLER_31_1015 ();
 sg13g2_fill_2 FILLER_31_1022 ();
 sg13g2_decap_4 FILLER_31_1028 ();
 sg13g2_decap_8 FILLER_31_1052 ();
 sg13g2_decap_8 FILLER_31_1059 ();
 sg13g2_decap_4 FILLER_31_1096 ();
 sg13g2_fill_1 FILLER_31_1100 ();
 sg13g2_fill_2 FILLER_31_1163 ();
 sg13g2_fill_1 FILLER_31_1165 ();
 sg13g2_decap_8 FILLER_31_1192 ();
 sg13g2_fill_1 FILLER_31_1199 ();
 sg13g2_fill_1 FILLER_31_1210 ();
 sg13g2_fill_1 FILLER_31_1215 ();
 sg13g2_fill_1 FILLER_31_1242 ();
 sg13g2_fill_1 FILLER_31_1269 ();
 sg13g2_decap_8 FILLER_31_1278 ();
 sg13g2_fill_2 FILLER_31_1285 ();
 sg13g2_fill_1 FILLER_31_1287 ();
 sg13g2_decap_8 FILLER_31_1298 ();
 sg13g2_fill_1 FILLER_31_1305 ();
 sg13g2_decap_8 FILLER_31_1310 ();
 sg13g2_decap_8 FILLER_31_1317 ();
 sg13g2_fill_2 FILLER_31_1324 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_37 ();
 sg13g2_fill_1 FILLER_32_52 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_1 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_113 ();
 sg13g2_fill_2 FILLER_32_117 ();
 sg13g2_fill_2 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_decap_8 FILLER_32_310 ();
 sg13g2_fill_2 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_decap_4 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_4 FILLER_32_393 ();
 sg13g2_fill_1 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_406 ();
 sg13g2_fill_2 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_417 ();
 sg13g2_fill_2 FILLER_32_424 ();
 sg13g2_fill_1 FILLER_32_426 ();
 sg13g2_fill_2 FILLER_32_514 ();
 sg13g2_fill_2 FILLER_32_557 ();
 sg13g2_decap_4 FILLER_32_620 ();
 sg13g2_fill_2 FILLER_32_624 ();
 sg13g2_decap_8 FILLER_32_647 ();
 sg13g2_fill_2 FILLER_32_654 ();
 sg13g2_fill_1 FILLER_32_656 ();
 sg13g2_fill_2 FILLER_32_674 ();
 sg13g2_decap_8 FILLER_32_694 ();
 sg13g2_decap_8 FILLER_32_727 ();
 sg13g2_decap_8 FILLER_32_734 ();
 sg13g2_decap_8 FILLER_32_741 ();
 sg13g2_decap_8 FILLER_32_748 ();
 sg13g2_fill_2 FILLER_32_755 ();
 sg13g2_decap_8 FILLER_32_765 ();
 sg13g2_decap_4 FILLER_32_772 ();
 sg13g2_fill_1 FILLER_32_776 ();
 sg13g2_decap_4 FILLER_32_803 ();
 sg13g2_fill_1 FILLER_32_807 ();
 sg13g2_decap_8 FILLER_32_844 ();
 sg13g2_decap_8 FILLER_32_851 ();
 sg13g2_decap_8 FILLER_32_858 ();
 sg13g2_decap_8 FILLER_32_865 ();
 sg13g2_decap_8 FILLER_32_872 ();
 sg13g2_fill_1 FILLER_32_879 ();
 sg13g2_decap_4 FILLER_32_894 ();
 sg13g2_decap_8 FILLER_32_928 ();
 sg13g2_decap_4 FILLER_32_935 ();
 sg13g2_fill_1 FILLER_32_939 ();
 sg13g2_decap_4 FILLER_32_954 ();
 sg13g2_fill_1 FILLER_32_958 ();
 sg13g2_decap_4 FILLER_32_969 ();
 sg13g2_decap_8 FILLER_32_1059 ();
 sg13g2_decap_4 FILLER_32_1066 ();
 sg13g2_fill_1 FILLER_32_1070 ();
 sg13g2_fill_2 FILLER_32_1081 ();
 sg13g2_decap_8 FILLER_32_1087 ();
 sg13g2_fill_1 FILLER_32_1114 ();
 sg13g2_fill_1 FILLER_32_1141 ();
 sg13g2_fill_2 FILLER_32_1168 ();
 sg13g2_fill_1 FILLER_32_1232 ();
 sg13g2_fill_2 FILLER_32_1253 ();
 sg13g2_decap_4 FILLER_32_1271 ();
 sg13g2_fill_2 FILLER_32_1285 ();
 sg13g2_fill_1 FILLER_32_1287 ();
 sg13g2_fill_2 FILLER_32_1292 ();
 sg13g2_fill_2 FILLER_32_1324 ();
 sg13g2_fill_2 FILLER_33_44 ();
 sg13g2_decap_8 FILLER_33_101 ();
 sg13g2_decap_8 FILLER_33_108 ();
 sg13g2_decap_8 FILLER_33_115 ();
 sg13g2_decap_4 FILLER_33_122 ();
 sg13g2_decap_4 FILLER_33_130 ();
 sg13g2_fill_2 FILLER_33_138 ();
 sg13g2_decap_4 FILLER_33_144 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_181 ();
 sg13g2_fill_1 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_4 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_decap_4 FILLER_33_321 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_4 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_428 ();
 sg13g2_decap_4 FILLER_33_434 ();
 sg13g2_fill_2 FILLER_33_443 ();
 sg13g2_fill_1 FILLER_33_466 ();
 sg13g2_fill_1 FILLER_33_578 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_fill_1 FILLER_33_616 ();
 sg13g2_fill_2 FILLER_33_684 ();
 sg13g2_decap_4 FILLER_33_712 ();
 sg13g2_decap_8 FILLER_33_724 ();
 sg13g2_decap_8 FILLER_33_731 ();
 sg13g2_decap_4 FILLER_33_738 ();
 sg13g2_decap_8 FILLER_33_746 ();
 sg13g2_decap_8 FILLER_33_753 ();
 sg13g2_decap_4 FILLER_33_760 ();
 sg13g2_fill_1 FILLER_33_820 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_decap_8 FILLER_33_859 ();
 sg13g2_decap_8 FILLER_33_866 ();
 sg13g2_decap_8 FILLER_33_873 ();
 sg13g2_decap_8 FILLER_33_890 ();
 sg13g2_fill_2 FILLER_33_897 ();
 sg13g2_fill_2 FILLER_33_903 ();
 sg13g2_fill_2 FILLER_33_915 ();
 sg13g2_fill_1 FILLER_33_917 ();
 sg13g2_decap_8 FILLER_33_928 ();
 sg13g2_fill_2 FILLER_33_935 ();
 sg13g2_fill_1 FILLER_33_937 ();
 sg13g2_fill_1 FILLER_33_942 ();
 sg13g2_decap_8 FILLER_33_989 ();
 sg13g2_decap_8 FILLER_33_996 ();
 sg13g2_decap_4 FILLER_33_1003 ();
 sg13g2_decap_4 FILLER_33_1021 ();
 sg13g2_fill_1 FILLER_33_1025 ();
 sg13g2_decap_8 FILLER_33_1036 ();
 sg13g2_fill_1 FILLER_33_1047 ();
 sg13g2_decap_4 FILLER_33_1056 ();
 sg13g2_fill_2 FILLER_33_1064 ();
 sg13g2_decap_8 FILLER_33_1102 ();
 sg13g2_decap_4 FILLER_33_1109 ();
 sg13g2_decap_8 FILLER_33_1127 ();
 sg13g2_decap_8 FILLER_33_1134 ();
 sg13g2_fill_2 FILLER_33_1189 ();
 sg13g2_fill_2 FILLER_33_1195 ();
 sg13g2_fill_1 FILLER_33_1197 ();
 sg13g2_fill_1 FILLER_33_1224 ();
 sg13g2_decap_4 FILLER_33_1229 ();
 sg13g2_fill_1 FILLER_33_1233 ();
 sg13g2_fill_2 FILLER_33_1244 ();
 sg13g2_fill_1 FILLER_33_1246 ();
 sg13g2_fill_2 FILLER_33_1277 ();
 sg13g2_fill_1 FILLER_33_1279 ();
 sg13g2_decap_8 FILLER_33_1314 ();
 sg13g2_decap_4 FILLER_33_1321 ();
 sg13g2_fill_1 FILLER_33_1325 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_12 ();
 sg13g2_fill_1 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_19 ();
 sg13g2_fill_2 FILLER_34_24 ();
 sg13g2_fill_1 FILLER_34_26 ();
 sg13g2_fill_1 FILLER_34_40 ();
 sg13g2_fill_1 FILLER_34_51 ();
 sg13g2_fill_1 FILLER_34_61 ();
 sg13g2_decap_4 FILLER_34_66 ();
 sg13g2_fill_2 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_124 ();
 sg13g2_decap_4 FILLER_34_131 ();
 sg13g2_decap_8 FILLER_34_139 ();
 sg13g2_decap_8 FILLER_34_146 ();
 sg13g2_decap_4 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_fill_2 FILLER_34_210 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_decap_4 FILLER_34_268 ();
 sg13g2_fill_1 FILLER_34_272 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_decap_8 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_324 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_fill_2 FILLER_34_338 ();
 sg13g2_fill_1 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_356 ();
 sg13g2_fill_2 FILLER_34_363 ();
 sg13g2_fill_1 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_370 ();
 sg13g2_fill_1 FILLER_34_383 ();
 sg13g2_fill_1 FILLER_34_388 ();
 sg13g2_decap_4 FILLER_34_419 ();
 sg13g2_fill_1 FILLER_34_423 ();
 sg13g2_fill_1 FILLER_34_428 ();
 sg13g2_decap_4 FILLER_34_443 ();
 sg13g2_fill_1 FILLER_34_447 ();
 sg13g2_decap_8 FILLER_34_452 ();
 sg13g2_fill_2 FILLER_34_464 ();
 sg13g2_decap_4 FILLER_34_474 ();
 sg13g2_fill_1 FILLER_34_478 ();
 sg13g2_fill_1 FILLER_34_522 ();
 sg13g2_fill_1 FILLER_34_533 ();
 sg13g2_fill_1 FILLER_34_538 ();
 sg13g2_fill_1 FILLER_34_544 ();
 sg13g2_decap_8 FILLER_34_574 ();
 sg13g2_fill_1 FILLER_34_585 ();
 sg13g2_decap_4 FILLER_34_590 ();
 sg13g2_fill_1 FILLER_34_594 ();
 sg13g2_fill_2 FILLER_34_599 ();
 sg13g2_fill_2 FILLER_34_605 ();
 sg13g2_fill_1 FILLER_34_607 ();
 sg13g2_fill_2 FILLER_34_663 ();
 sg13g2_fill_1 FILLER_34_665 ();
 sg13g2_fill_2 FILLER_34_670 ();
 sg13g2_fill_1 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_728 ();
 sg13g2_decap_8 FILLER_34_735 ();
 sg13g2_decap_8 FILLER_34_742 ();
 sg13g2_fill_2 FILLER_34_775 ();
 sg13g2_fill_1 FILLER_34_777 ();
 sg13g2_fill_2 FILLER_34_782 ();
 sg13g2_fill_1 FILLER_34_784 ();
 sg13g2_fill_2 FILLER_34_790 ();
 sg13g2_fill_1 FILLER_34_792 ();
 sg13g2_fill_2 FILLER_34_798 ();
 sg13g2_fill_1 FILLER_34_800 ();
 sg13g2_decap_4 FILLER_34_810 ();
 sg13g2_fill_1 FILLER_34_814 ();
 sg13g2_decap_4 FILLER_34_853 ();
 sg13g2_fill_1 FILLER_34_919 ();
 sg13g2_fill_2 FILLER_34_924 ();
 sg13g2_fill_1 FILLER_34_926 ();
 sg13g2_decap_8 FILLER_34_969 ();
 sg13g2_decap_8 FILLER_34_976 ();
 sg13g2_fill_1 FILLER_34_983 ();
 sg13g2_decap_8 FILLER_34_988 ();
 sg13g2_decap_8 FILLER_34_995 ();
 sg13g2_decap_8 FILLER_34_1002 ();
 sg13g2_decap_8 FILLER_34_1009 ();
 sg13g2_decap_4 FILLER_34_1016 ();
 sg13g2_fill_2 FILLER_34_1060 ();
 sg13g2_decap_8 FILLER_34_1098 ();
 sg13g2_decap_8 FILLER_34_1105 ();
 sg13g2_decap_8 FILLER_34_1112 ();
 sg13g2_decap_8 FILLER_34_1119 ();
 sg13g2_decap_8 FILLER_34_1126 ();
 sg13g2_decap_4 FILLER_34_1133 ();
 sg13g2_decap_8 FILLER_34_1185 ();
 sg13g2_decap_8 FILLER_34_1192 ();
 sg13g2_decap_8 FILLER_34_1199 ();
 sg13g2_decap_4 FILLER_34_1210 ();
 sg13g2_fill_2 FILLER_34_1240 ();
 sg13g2_fill_1 FILLER_34_1242 ();
 sg13g2_fill_1 FILLER_34_1257 ();
 sg13g2_decap_8 FILLER_34_1262 ();
 sg13g2_decap_8 FILLER_34_1269 ();
 sg13g2_decap_8 FILLER_34_1276 ();
 sg13g2_fill_2 FILLER_34_1283 ();
 sg13g2_decap_4 FILLER_34_1295 ();
 sg13g2_fill_1 FILLER_34_1325 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_decap_8 FILLER_35_58 ();
 sg13g2_decap_8 FILLER_35_65 ();
 sg13g2_fill_1 FILLER_35_72 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_decap_4 FILLER_35_101 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_177 ();
 sg13g2_fill_1 FILLER_35_179 ();
 sg13g2_decap_4 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_241 ();
 sg13g2_fill_2 FILLER_35_248 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_decap_4 FILLER_35_261 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_decap_4 FILLER_35_307 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_fill_2 FILLER_35_336 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_decap_4 FILLER_35_422 ();
 sg13g2_fill_2 FILLER_35_426 ();
 sg13g2_fill_2 FILLER_35_443 ();
 sg13g2_fill_1 FILLER_35_445 ();
 sg13g2_decap_4 FILLER_35_463 ();
 sg13g2_fill_2 FILLER_35_467 ();
 sg13g2_fill_1 FILLER_35_487 ();
 sg13g2_fill_2 FILLER_35_501 ();
 sg13g2_fill_1 FILLER_35_503 ();
 sg13g2_decap_8 FILLER_35_508 ();
 sg13g2_decap_8 FILLER_35_515 ();
 sg13g2_decap_8 FILLER_35_522 ();
 sg13g2_decap_8 FILLER_35_529 ();
 sg13g2_decap_8 FILLER_35_536 ();
 sg13g2_decap_8 FILLER_35_543 ();
 sg13g2_fill_2 FILLER_35_554 ();
 sg13g2_fill_1 FILLER_35_556 ();
 sg13g2_fill_2 FILLER_35_562 ();
 sg13g2_decap_4 FILLER_35_570 ();
 sg13g2_fill_1 FILLER_35_574 ();
 sg13g2_decap_8 FILLER_35_593 ();
 sg13g2_fill_1 FILLER_35_600 ();
 sg13g2_fill_1 FILLER_35_615 ();
 sg13g2_fill_2 FILLER_35_663 ();
 sg13g2_fill_2 FILLER_35_673 ();
 sg13g2_fill_1 FILLER_35_690 ();
 sg13g2_decap_8 FILLER_35_717 ();
 sg13g2_fill_1 FILLER_35_724 ();
 sg13g2_decap_8 FILLER_35_729 ();
 sg13g2_decap_8 FILLER_35_741 ();
 sg13g2_decap_8 FILLER_35_748 ();
 sg13g2_fill_1 FILLER_35_755 ();
 sg13g2_fill_2 FILLER_35_765 ();
 sg13g2_decap_8 FILLER_35_776 ();
 sg13g2_decap_4 FILLER_35_783 ();
 sg13g2_decap_8 FILLER_35_796 ();
 sg13g2_fill_2 FILLER_35_803 ();
 sg13g2_fill_1 FILLER_35_805 ();
 sg13g2_fill_1 FILLER_35_810 ();
 sg13g2_fill_2 FILLER_35_819 ();
 sg13g2_fill_1 FILLER_35_825 ();
 sg13g2_fill_2 FILLER_35_898 ();
 sg13g2_decap_8 FILLER_35_904 ();
 sg13g2_fill_2 FILLER_35_911 ();
 sg13g2_fill_1 FILLER_35_913 ();
 sg13g2_decap_8 FILLER_35_918 ();
 sg13g2_decap_8 FILLER_35_925 ();
 sg13g2_fill_2 FILLER_35_932 ();
 sg13g2_fill_1 FILLER_35_934 ();
 sg13g2_fill_2 FILLER_35_963 ();
 sg13g2_decap_4 FILLER_35_1001 ();
 sg13g2_fill_2 FILLER_35_1005 ();
 sg13g2_decap_8 FILLER_35_1039 ();
 sg13g2_fill_2 FILLER_35_1046 ();
 sg13g2_fill_1 FILLER_35_1048 ();
 sg13g2_fill_1 FILLER_35_1105 ();
 sg13g2_decap_8 FILLER_35_1110 ();
 sg13g2_fill_2 FILLER_35_1117 ();
 sg13g2_fill_1 FILLER_35_1119 ();
 sg13g2_decap_8 FILLER_35_1160 ();
 sg13g2_decap_8 FILLER_35_1203 ();
 sg13g2_fill_2 FILLER_35_1220 ();
 sg13g2_decap_4 FILLER_35_1274 ();
 sg13g2_fill_2 FILLER_35_1278 ();
 sg13g2_fill_2 FILLER_35_1324 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_fill_1 FILLER_36_6 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_decap_8 FILLER_36_38 ();
 sg13g2_fill_1 FILLER_36_45 ();
 sg13g2_fill_2 FILLER_36_61 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_4 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_fill_2 FILLER_36_115 ();
 sg13g2_fill_2 FILLER_36_247 ();
 sg13g2_fill_1 FILLER_36_249 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_decap_4 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_330 ();
 sg13g2_fill_2 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_415 ();
 sg13g2_decap_8 FILLER_36_422 ();
 sg13g2_decap_4 FILLER_36_429 ();
 sg13g2_fill_1 FILLER_36_433 ();
 sg13g2_fill_1 FILLER_36_460 ();
 sg13g2_fill_1 FILLER_36_497 ();
 sg13g2_fill_2 FILLER_36_506 ();
 sg13g2_decap_4 FILLER_36_516 ();
 sg13g2_fill_1 FILLER_36_520 ();
 sg13g2_decap_8 FILLER_36_535 ();
 sg13g2_fill_1 FILLER_36_542 ();
 sg13g2_decap_4 FILLER_36_547 ();
 sg13g2_fill_1 FILLER_36_551 ();
 sg13g2_decap_4 FILLER_36_560 ();
 sg13g2_decap_8 FILLER_36_568 ();
 sg13g2_fill_1 FILLER_36_575 ();
 sg13g2_decap_4 FILLER_36_580 ();
 sg13g2_fill_1 FILLER_36_584 ();
 sg13g2_decap_8 FILLER_36_589 ();
 sg13g2_fill_2 FILLER_36_596 ();
 sg13g2_decap_4 FILLER_36_620 ();
 sg13g2_fill_2 FILLER_36_628 ();
 sg13g2_decap_8 FILLER_36_634 ();
 sg13g2_fill_2 FILLER_36_641 ();
 sg13g2_decap_4 FILLER_36_674 ();
 sg13g2_fill_1 FILLER_36_697 ();
 sg13g2_fill_1 FILLER_36_702 ();
 sg13g2_decap_8 FILLER_36_711 ();
 sg13g2_fill_1 FILLER_36_718 ();
 sg13g2_decap_8 FILLER_36_771 ();
 sg13g2_decap_4 FILLER_36_778 ();
 sg13g2_fill_1 FILLER_36_782 ();
 sg13g2_fill_1 FILLER_36_817 ();
 sg13g2_fill_2 FILLER_36_823 ();
 sg13g2_fill_1 FILLER_36_825 ();
 sg13g2_fill_2 FILLER_36_852 ();
 sg13g2_fill_1 FILLER_36_854 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_decap_4 FILLER_36_891 ();
 sg13g2_fill_2 FILLER_36_895 ();
 sg13g2_fill_1 FILLER_36_907 ();
 sg13g2_fill_2 FILLER_36_934 ();
 sg13g2_fill_2 FILLER_36_940 ();
 sg13g2_fill_2 FILLER_36_968 ();
 sg13g2_decap_4 FILLER_36_996 ();
 sg13g2_decap_8 FILLER_36_1038 ();
 sg13g2_decap_8 FILLER_36_1045 ();
 sg13g2_fill_2 FILLER_36_1052 ();
 sg13g2_fill_1 FILLER_36_1062 ();
 sg13g2_decap_4 FILLER_36_1067 ();
 sg13g2_fill_1 FILLER_36_1071 ();
 sg13g2_fill_2 FILLER_36_1118 ();
 sg13g2_fill_2 FILLER_36_1150 ();
 sg13g2_fill_1 FILLER_36_1152 ();
 sg13g2_fill_2 FILLER_36_1163 ();
 sg13g2_fill_1 FILLER_36_1165 ();
 sg13g2_fill_1 FILLER_36_1176 ();
 sg13g2_fill_2 FILLER_36_1207 ();
 sg13g2_decap_8 FILLER_36_1245 ();
 sg13g2_decap_8 FILLER_36_1252 ();
 sg13g2_decap_8 FILLER_36_1259 ();
 sg13g2_decap_8 FILLER_36_1266 ();
 sg13g2_decap_8 FILLER_36_1273 ();
 sg13g2_decap_4 FILLER_36_1280 ();
 sg13g2_fill_1 FILLER_36_1284 ();
 sg13g2_fill_1 FILLER_36_1325 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_22 ();
 sg13g2_decap_8 FILLER_37_29 ();
 sg13g2_decap_8 FILLER_37_36 ();
 sg13g2_fill_1 FILLER_37_43 ();
 sg13g2_fill_2 FILLER_37_48 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_decap_8 FILLER_37_114 ();
 sg13g2_decap_8 FILLER_37_121 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_fill_2 FILLER_37_180 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_187 ();
 sg13g2_decap_8 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_201 ();
 sg13g2_decap_4 FILLER_37_208 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_4 FILLER_37_245 ();
 sg13g2_fill_1 FILLER_37_249 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_fill_1 FILLER_37_296 ();
 sg13g2_fill_1 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_decap_4 FILLER_37_353 ();
 sg13g2_fill_1 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_37_409 ();
 sg13g2_decap_4 FILLER_37_416 ();
 sg13g2_fill_1 FILLER_37_507 ();
 sg13g2_decap_8 FILLER_37_512 ();
 sg13g2_fill_2 FILLER_37_519 ();
 sg13g2_fill_1 FILLER_37_561 ();
 sg13g2_fill_2 FILLER_37_566 ();
 sg13g2_fill_2 FILLER_37_572 ();
 sg13g2_fill_2 FILLER_37_578 ();
 sg13g2_fill_1 FILLER_37_580 ();
 sg13g2_decap_8 FILLER_37_590 ();
 sg13g2_fill_1 FILLER_37_597 ();
 sg13g2_fill_2 FILLER_37_603 ();
 sg13g2_fill_1 FILLER_37_605 ();
 sg13g2_fill_2 FILLER_37_610 ();
 sg13g2_fill_1 FILLER_37_625 ();
 sg13g2_decap_8 FILLER_37_634 ();
 sg13g2_decap_8 FILLER_37_666 ();
 sg13g2_decap_4 FILLER_37_673 ();
 sg13g2_decap_8 FILLER_37_682 ();
 sg13g2_decap_4 FILLER_37_689 ();
 sg13g2_fill_2 FILLER_37_693 ();
 sg13g2_decap_4 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_708 ();
 sg13g2_decap_8 FILLER_37_715 ();
 sg13g2_decap_4 FILLER_37_722 ();
 sg13g2_decap_4 FILLER_37_730 ();
 sg13g2_fill_1 FILLER_37_734 ();
 sg13g2_fill_1 FILLER_37_761 ();
 sg13g2_decap_8 FILLER_37_850 ();
 sg13g2_decap_8 FILLER_37_857 ();
 sg13g2_decap_8 FILLER_37_864 ();
 sg13g2_fill_1 FILLER_37_871 ();
 sg13g2_decap_8 FILLER_37_876 ();
 sg13g2_decap_8 FILLER_37_883 ();
 sg13g2_decap_4 FILLER_37_890 ();
 sg13g2_fill_2 FILLER_37_894 ();
 sg13g2_fill_2 FILLER_37_942 ();
 sg13g2_fill_2 FILLER_37_970 ();
 sg13g2_fill_1 FILLER_37_972 ();
 sg13g2_fill_1 FILLER_37_977 ();
 sg13g2_fill_2 FILLER_37_1004 ();
 sg13g2_fill_1 FILLER_37_1006 ();
 sg13g2_decap_8 FILLER_37_1037 ();
 sg13g2_fill_1 FILLER_37_1044 ();
 sg13g2_decap_4 FILLER_37_1121 ();
 sg13g2_fill_2 FILLER_37_1133 ();
 sg13g2_fill_1 FILLER_37_1135 ();
 sg13g2_decap_4 FILLER_37_1196 ();
 sg13g2_fill_1 FILLER_37_1200 ();
 sg13g2_decap_4 FILLER_37_1231 ();
 sg13g2_fill_2 FILLER_37_1235 ();
 sg13g2_decap_8 FILLER_37_1277 ();
 sg13g2_decap_4 FILLER_37_1294 ();
 sg13g2_fill_2 FILLER_37_1298 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_37 ();
 sg13g2_fill_2 FILLER_38_52 ();
 sg13g2_fill_1 FILLER_38_54 ();
 sg13g2_fill_2 FILLER_38_59 ();
 sg13g2_fill_1 FILLER_38_61 ();
 sg13g2_decap_8 FILLER_38_129 ();
 sg13g2_decap_4 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_149 ();
 sg13g2_decap_8 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_163 ();
 sg13g2_decap_4 FILLER_38_170 ();
 sg13g2_fill_1 FILLER_38_174 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_249 ();
 sg13g2_decap_4 FILLER_38_256 ();
 sg13g2_fill_2 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_266 ();
 sg13g2_decap_4 FILLER_38_290 ();
 sg13g2_decap_8 FILLER_38_298 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_decap_4 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_316 ();
 sg13g2_fill_2 FILLER_38_329 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_decap_4 FILLER_38_346 ();
 sg13g2_fill_1 FILLER_38_350 ();
 sg13g2_fill_2 FILLER_38_355 ();
 sg13g2_decap_4 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_fill_1 FILLER_38_400 ();
 sg13g2_decap_8 FILLER_38_422 ();
 sg13g2_decap_4 FILLER_38_429 ();
 sg13g2_fill_1 FILLER_38_433 ();
 sg13g2_decap_8 FILLER_38_489 ();
 sg13g2_decap_4 FILLER_38_496 ();
 sg13g2_fill_1 FILLER_38_500 ();
 sg13g2_decap_4 FILLER_38_574 ();
 sg13g2_decap_8 FILLER_38_597 ();
 sg13g2_decap_8 FILLER_38_604 ();
 sg13g2_fill_2 FILLER_38_625 ();
 sg13g2_decap_8 FILLER_38_641 ();
 sg13g2_fill_2 FILLER_38_648 ();
 sg13g2_decap_8 FILLER_38_676 ();
 sg13g2_decap_8 FILLER_38_683 ();
 sg13g2_decap_4 FILLER_38_690 ();
 sg13g2_fill_2 FILLER_38_694 ();
 sg13g2_decap_8 FILLER_38_701 ();
 sg13g2_decap_8 FILLER_38_712 ();
 sg13g2_fill_2 FILLER_38_749 ();
 sg13g2_fill_1 FILLER_38_751 ();
 sg13g2_decap_8 FILLER_38_761 ();
 sg13g2_decap_4 FILLER_38_768 ();
 sg13g2_fill_2 FILLER_38_772 ();
 sg13g2_decap_4 FILLER_38_778 ();
 sg13g2_fill_1 FILLER_38_782 ();
 sg13g2_fill_1 FILLER_38_788 ();
 sg13g2_fill_1 FILLER_38_793 ();
 sg13g2_fill_2 FILLER_38_799 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_4 FILLER_38_847 ();
 sg13g2_fill_2 FILLER_38_851 ();
 sg13g2_decap_8 FILLER_38_882 ();
 sg13g2_decap_8 FILLER_38_889 ();
 sg13g2_decap_4 FILLER_38_896 ();
 sg13g2_fill_1 FILLER_38_968 ();
 sg13g2_fill_1 FILLER_38_989 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_decap_8 FILLER_38_1001 ();
 sg13g2_decap_4 FILLER_38_1008 ();
 sg13g2_fill_2 FILLER_38_1012 ();
 sg13g2_decap_8 FILLER_38_1050 ();
 sg13g2_decap_4 FILLER_38_1057 ();
 sg13g2_fill_1 FILLER_38_1061 ();
 sg13g2_decap_8 FILLER_38_1110 ();
 sg13g2_decap_8 FILLER_38_1117 ();
 sg13g2_decap_8 FILLER_38_1124 ();
 sg13g2_fill_1 FILLER_38_1131 ();
 sg13g2_decap_4 FILLER_38_1136 ();
 sg13g2_decap_8 FILLER_38_1164 ();
 sg13g2_decap_8 FILLER_38_1233 ();
 sg13g2_decap_4 FILLER_38_1240 ();
 sg13g2_decap_8 FILLER_38_1310 ();
 sg13g2_decap_8 FILLER_38_1317 ();
 sg13g2_fill_2 FILLER_38_1324 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_4 FILLER_39_94 ();
 sg13g2_fill_1 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_120 ();
 sg13g2_decap_8 FILLER_39_127 ();
 sg13g2_decap_8 FILLER_39_134 ();
 sg13g2_fill_2 FILLER_39_141 ();
 sg13g2_decap_4 FILLER_39_155 ();
 sg13g2_fill_2 FILLER_39_159 ();
 sg13g2_decap_8 FILLER_39_173 ();
 sg13g2_decap_8 FILLER_39_180 ();
 sg13g2_decap_8 FILLER_39_187 ();
 sg13g2_decap_8 FILLER_39_194 ();
 sg13g2_fill_2 FILLER_39_201 ();
 sg13g2_fill_1 FILLER_39_203 ();
 sg13g2_fill_2 FILLER_39_208 ();
 sg13g2_decap_4 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_232 ();
 sg13g2_decap_8 FILLER_39_239 ();
 sg13g2_decap_4 FILLER_39_246 ();
 sg13g2_fill_1 FILLER_39_259 ();
 sg13g2_fill_2 FILLER_39_274 ();
 sg13g2_decap_8 FILLER_39_323 ();
 sg13g2_decap_8 FILLER_39_330 ();
 sg13g2_fill_1 FILLER_39_337 ();
 sg13g2_fill_2 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_357 ();
 sg13g2_fill_1 FILLER_39_362 ();
 sg13g2_fill_1 FILLER_39_373 ();
 sg13g2_fill_1 FILLER_39_395 ();
 sg13g2_fill_2 FILLER_39_417 ();
 sg13g2_fill_1 FILLER_39_419 ();
 sg13g2_fill_1 FILLER_39_473 ();
 sg13g2_fill_1 FILLER_39_535 ();
 sg13g2_fill_1 FILLER_39_562 ();
 sg13g2_decap_4 FILLER_39_567 ();
 sg13g2_fill_1 FILLER_39_571 ();
 sg13g2_decap_8 FILLER_39_602 ();
 sg13g2_decap_4 FILLER_39_609 ();
 sg13g2_fill_2 FILLER_39_613 ();
 sg13g2_decap_4 FILLER_39_620 ();
 sg13g2_decap_8 FILLER_39_650 ();
 sg13g2_fill_2 FILLER_39_657 ();
 sg13g2_fill_2 FILLER_39_674 ();
 sg13g2_fill_2 FILLER_39_702 ();
 sg13g2_fill_1 FILLER_39_704 ();
 sg13g2_decap_8 FILLER_39_709 ();
 sg13g2_decap_8 FILLER_39_716 ();
 sg13g2_decap_8 FILLER_39_723 ();
 sg13g2_decap_8 FILLER_39_730 ();
 sg13g2_fill_2 FILLER_39_737 ();
 sg13g2_fill_1 FILLER_39_739 ();
 sg13g2_decap_4 FILLER_39_748 ();
 sg13g2_fill_2 FILLER_39_752 ();
 sg13g2_decap_4 FILLER_39_758 ();
 sg13g2_fill_1 FILLER_39_762 ();
 sg13g2_decap_8 FILLER_39_789 ();
 sg13g2_fill_1 FILLER_39_796 ();
 sg13g2_fill_2 FILLER_39_809 ();
 sg13g2_decap_8 FILLER_39_819 ();
 sg13g2_decap_8 FILLER_39_826 ();
 sg13g2_decap_8 FILLER_39_833 ();
 sg13g2_decap_8 FILLER_39_840 ();
 sg13g2_decap_4 FILLER_39_847 ();
 sg13g2_fill_1 FILLER_39_851 ();
 sg13g2_decap_4 FILLER_39_904 ();
 sg13g2_fill_1 FILLER_39_908 ();
 sg13g2_decap_8 FILLER_39_917 ();
 sg13g2_decap_8 FILLER_39_924 ();
 sg13g2_decap_4 FILLER_39_931 ();
 sg13g2_fill_2 FILLER_39_935 ();
 sg13g2_decap_4 FILLER_39_941 ();
 sg13g2_fill_1 FILLER_39_945 ();
 sg13g2_decap_8 FILLER_39_960 ();
 sg13g2_decap_8 FILLER_39_967 ();
 sg13g2_decap_8 FILLER_39_974 ();
 sg13g2_fill_2 FILLER_39_981 ();
 sg13g2_decap_4 FILLER_39_1023 ();
 sg13g2_decap_8 FILLER_39_1041 ();
 sg13g2_decap_4 FILLER_39_1048 ();
 sg13g2_fill_1 FILLER_39_1052 ();
 sg13g2_fill_2 FILLER_39_1061 ();
 sg13g2_fill_1 FILLER_39_1063 ();
 sg13g2_fill_1 FILLER_39_1068 ();
 sg13g2_decap_4 FILLER_39_1089 ();
 sg13g2_fill_1 FILLER_39_1093 ();
 sg13g2_decap_8 FILLER_39_1124 ();
 sg13g2_decap_8 FILLER_39_1131 ();
 sg13g2_fill_2 FILLER_39_1138 ();
 sg13g2_fill_1 FILLER_39_1140 ();
 sg13g2_decap_8 FILLER_39_1145 ();
 sg13g2_decap_8 FILLER_39_1152 ();
 sg13g2_decap_8 FILLER_39_1159 ();
 sg13g2_decap_8 FILLER_39_1166 ();
 sg13g2_decap_8 FILLER_39_1173 ();
 sg13g2_decap_4 FILLER_39_1180 ();
 sg13g2_fill_1 FILLER_39_1184 ();
 sg13g2_decap_8 FILLER_39_1231 ();
 sg13g2_decap_8 FILLER_39_1238 ();
 sg13g2_decap_4 FILLER_39_1245 ();
 sg13g2_decap_8 FILLER_39_1269 ();
 sg13g2_decap_4 FILLER_39_1276 ();
 sg13g2_fill_1 FILLER_39_1280 ();
 sg13g2_decap_4 FILLER_39_1295 ();
 sg13g2_fill_1 FILLER_39_1299 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_1 FILLER_40_66 ();
 sg13g2_fill_2 FILLER_40_71 ();
 sg13g2_fill_1 FILLER_40_73 ();
 sg13g2_decap_8 FILLER_40_78 ();
 sg13g2_decap_8 FILLER_40_114 ();
 sg13g2_decap_4 FILLER_40_121 ();
 sg13g2_fill_2 FILLER_40_125 ();
 sg13g2_decap_4 FILLER_40_200 ();
 sg13g2_fill_1 FILLER_40_204 ();
 sg13g2_fill_2 FILLER_40_270 ();
 sg13g2_decap_4 FILLER_40_302 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_decap_8 FILLER_40_328 ();
 sg13g2_fill_1 FILLER_40_335 ();
 sg13g2_fill_1 FILLER_40_387 ();
 sg13g2_decap_4 FILLER_40_430 ();
 sg13g2_fill_2 FILLER_40_434 ();
 sg13g2_fill_1 FILLER_40_440 ();
 sg13g2_decap_8 FILLER_40_445 ();
 sg13g2_decap_4 FILLER_40_452 ();
 sg13g2_fill_2 FILLER_40_460 ();
 sg13g2_fill_1 FILLER_40_509 ();
 sg13g2_decap_4 FILLER_40_518 ();
 sg13g2_fill_2 FILLER_40_522 ();
 sg13g2_decap_4 FILLER_40_529 ();
 sg13g2_fill_1 FILLER_40_533 ();
 sg13g2_fill_2 FILLER_40_538 ();
 sg13g2_fill_1 FILLER_40_540 ();
 sg13g2_decap_4 FILLER_40_562 ();
 sg13g2_fill_1 FILLER_40_566 ();
 sg13g2_fill_1 FILLER_40_599 ();
 sg13g2_decap_8 FILLER_40_604 ();
 sg13g2_decap_8 FILLER_40_611 ();
 sg13g2_fill_1 FILLER_40_618 ();
 sg13g2_decap_8 FILLER_40_674 ();
 sg13g2_decap_4 FILLER_40_681 ();
 sg13g2_decap_4 FILLER_40_694 ();
 sg13g2_fill_1 FILLER_40_698 ();
 sg13g2_decap_4 FILLER_40_729 ();
 sg13g2_fill_1 FILLER_40_733 ();
 sg13g2_decap_4 FILLER_40_742 ();
 sg13g2_fill_1 FILLER_40_746 ();
 sg13g2_fill_1 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_782 ();
 sg13g2_decap_8 FILLER_40_789 ();
 sg13g2_decap_8 FILLER_40_796 ();
 sg13g2_decap_8 FILLER_40_803 ();
 sg13g2_decap_8 FILLER_40_810 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_decap_8 FILLER_40_824 ();
 sg13g2_fill_1 FILLER_40_831 ();
 sg13g2_fill_2 FILLER_40_862 ();
 sg13g2_fill_1 FILLER_40_880 ();
 sg13g2_decap_8 FILLER_40_907 ();
 sg13g2_decap_8 FILLER_40_914 ();
 sg13g2_decap_8 FILLER_40_921 ();
 sg13g2_decap_8 FILLER_40_928 ();
 sg13g2_fill_2 FILLER_40_935 ();
 sg13g2_fill_1 FILLER_40_937 ();
 sg13g2_decap_8 FILLER_40_945 ();
 sg13g2_decap_8 FILLER_40_978 ();
 sg13g2_fill_1 FILLER_40_985 ();
 sg13g2_decap_4 FILLER_40_1026 ();
 sg13g2_fill_1 FILLER_40_1030 ();
 sg13g2_decap_4 FILLER_40_1057 ();
 sg13g2_fill_1 FILLER_40_1061 ();
 sg13g2_fill_2 FILLER_40_1088 ();
 sg13g2_fill_1 FILLER_40_1090 ();
 sg13g2_fill_2 FILLER_40_1095 ();
 sg13g2_fill_1 FILLER_40_1097 ();
 sg13g2_decap_4 FILLER_40_1124 ();
 sg13g2_fill_2 FILLER_40_1128 ();
 sg13g2_decap_8 FILLER_40_1160 ();
 sg13g2_decap_8 FILLER_40_1167 ();
 sg13g2_decap_8 FILLER_40_1178 ();
 sg13g2_decap_8 FILLER_40_1185 ();
 sg13g2_decap_8 FILLER_40_1192 ();
 sg13g2_fill_2 FILLER_40_1199 ();
 sg13g2_fill_1 FILLER_40_1201 ();
 sg13g2_decap_8 FILLER_40_1232 ();
 sg13g2_decap_8 FILLER_40_1239 ();
 sg13g2_decap_8 FILLER_40_1246 ();
 sg13g2_decap_8 FILLER_40_1253 ();
 sg13g2_decap_4 FILLER_40_1260 ();
 sg13g2_fill_1 FILLER_40_1264 ();
 sg13g2_decap_8 FILLER_40_1299 ();
 sg13g2_decap_8 FILLER_40_1314 ();
 sg13g2_decap_4 FILLER_40_1321 ();
 sg13g2_fill_1 FILLER_40_1325 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_11 ();
 sg13g2_decap_8 FILLER_41_74 ();
 sg13g2_decap_8 FILLER_41_81 ();
 sg13g2_decap_8 FILLER_41_88 ();
 sg13g2_decap_8 FILLER_41_95 ();
 sg13g2_decap_8 FILLER_41_102 ();
 sg13g2_decap_8 FILLER_41_109 ();
 sg13g2_decap_8 FILLER_41_116 ();
 sg13g2_decap_4 FILLER_41_123 ();
 sg13g2_fill_1 FILLER_41_152 ();
 sg13g2_fill_1 FILLER_41_179 ();
 sg13g2_fill_2 FILLER_41_237 ();
 sg13g2_fill_2 FILLER_41_260 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_fill_2 FILLER_41_272 ();
 sg13g2_fill_1 FILLER_41_274 ();
 sg13g2_fill_2 FILLER_41_301 ();
 sg13g2_fill_1 FILLER_41_303 ();
 sg13g2_fill_2 FILLER_41_325 ();
 sg13g2_fill_1 FILLER_41_327 ();
 sg13g2_fill_2 FILLER_41_338 ();
 sg13g2_fill_2 FILLER_41_372 ();
 sg13g2_fill_2 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_4 FILLER_41_413 ();
 sg13g2_fill_2 FILLER_41_417 ();
 sg13g2_decap_8 FILLER_41_423 ();
 sg13g2_fill_2 FILLER_41_430 ();
 sg13g2_fill_1 FILLER_41_432 ();
 sg13g2_fill_1 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_499 ();
 sg13g2_fill_2 FILLER_41_506 ();
 sg13g2_fill_1 FILLER_41_508 ();
 sg13g2_decap_8 FILLER_41_513 ();
 sg13g2_decap_8 FILLER_41_520 ();
 sg13g2_decap_4 FILLER_41_527 ();
 sg13g2_fill_2 FILLER_41_531 ();
 sg13g2_decap_8 FILLER_41_538 ();
 sg13g2_fill_2 FILLER_41_545 ();
 sg13g2_decap_4 FILLER_41_573 ();
 sg13g2_fill_2 FILLER_41_577 ();
 sg13g2_decap_4 FILLER_41_653 ();
 sg13g2_fill_1 FILLER_41_657 ();
 sg13g2_decap_4 FILLER_41_666 ();
 sg13g2_fill_1 FILLER_41_670 ();
 sg13g2_decap_4 FILLER_41_675 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_fill_2 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_706 ();
 sg13g2_fill_2 FILLER_41_713 ();
 sg13g2_fill_1 FILLER_41_715 ();
 sg13g2_fill_2 FILLER_41_719 ();
 sg13g2_fill_2 FILLER_41_734 ();
 sg13g2_fill_1 FILLER_41_736 ();
 sg13g2_fill_2 FILLER_41_745 ();
 sg13g2_fill_1 FILLER_41_747 ();
 sg13g2_fill_1 FILLER_41_752 ();
 sg13g2_fill_1 FILLER_41_766 ();
 sg13g2_decap_8 FILLER_41_801 ();
 sg13g2_fill_1 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_846 ();
 sg13g2_fill_1 FILLER_41_853 ();
 sg13g2_fill_2 FILLER_41_863 ();
 sg13g2_decap_4 FILLER_41_895 ();
 sg13g2_fill_2 FILLER_41_899 ();
 sg13g2_fill_2 FILLER_41_968 ();
 sg13g2_decap_8 FILLER_41_974 ();
 sg13g2_decap_8 FILLER_41_981 ();
 sg13g2_decap_4 FILLER_41_988 ();
 sg13g2_decap_4 FILLER_41_1018 ();
 sg13g2_fill_2 FILLER_41_1022 ();
 sg13g2_fill_2 FILLER_41_1050 ();
 sg13g2_fill_1 FILLER_41_1078 ();
 sg13g2_fill_2 FILLER_41_1083 ();
 sg13g2_fill_1 FILLER_41_1085 ();
 sg13g2_decap_8 FILLER_41_1116 ();
 sg13g2_fill_2 FILLER_41_1123 ();
 sg13g2_fill_1 FILLER_41_1125 ();
 sg13g2_fill_1 FILLER_41_1152 ();
 sg13g2_decap_4 FILLER_41_1209 ();
 sg13g2_fill_2 FILLER_41_1213 ();
 sg13g2_decap_8 FILLER_41_1219 ();
 sg13g2_fill_2 FILLER_41_1226 ();
 sg13g2_fill_1 FILLER_41_1228 ();
 sg13g2_decap_4 FILLER_41_1269 ();
 sg13g2_decap_8 FILLER_41_1277 ();
 sg13g2_decap_8 FILLER_41_1284 ();
 sg13g2_decap_8 FILLER_41_1291 ();
 sg13g2_decap_8 FILLER_41_1298 ();
 sg13g2_decap_8 FILLER_41_1305 ();
 sg13g2_decap_8 FILLER_41_1312 ();
 sg13g2_decap_8 FILLER_41_1319 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_12 ();
 sg13g2_fill_1 FILLER_42_23 ();
 sg13g2_fill_2 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_40 ();
 sg13g2_decap_8 FILLER_42_51 ();
 sg13g2_decap_8 FILLER_42_58 ();
 sg13g2_decap_8 FILLER_42_65 ();
 sg13g2_decap_8 FILLER_42_72 ();
 sg13g2_decap_8 FILLER_42_79 ();
 sg13g2_fill_2 FILLER_42_86 ();
 sg13g2_fill_1 FILLER_42_88 ();
 sg13g2_decap_8 FILLER_42_115 ();
 sg13g2_decap_8 FILLER_42_122 ();
 sg13g2_decap_8 FILLER_42_129 ();
 sg13g2_decap_4 FILLER_42_136 ();
 sg13g2_fill_2 FILLER_42_166 ();
 sg13g2_decap_8 FILLER_42_197 ();
 sg13g2_fill_2 FILLER_42_307 ();
 sg13g2_fill_1 FILLER_42_338 ();
 sg13g2_decap_4 FILLER_42_344 ();
 sg13g2_decap_8 FILLER_42_352 ();
 sg13g2_fill_2 FILLER_42_363 ();
 sg13g2_fill_1 FILLER_42_365 ();
 sg13g2_fill_1 FILLER_42_370 ();
 sg13g2_fill_2 FILLER_42_385 ();
 sg13g2_fill_2 FILLER_42_391 ();
 sg13g2_fill_2 FILLER_42_403 ();
 sg13g2_fill_1 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_fill_1 FILLER_42_490 ();
 sg13g2_decap_4 FILLER_42_495 ();
 sg13g2_fill_2 FILLER_42_533 ();
 sg13g2_fill_2 FILLER_42_540 ();
 sg13g2_fill_1 FILLER_42_542 ();
 sg13g2_decap_4 FILLER_42_564 ();
 sg13g2_fill_2 FILLER_42_568 ();
 sg13g2_decap_8 FILLER_42_580 ();
 sg13g2_fill_2 FILLER_42_587 ();
 sg13g2_decap_8 FILLER_42_619 ();
 sg13g2_decap_4 FILLER_42_626 ();
 sg13g2_fill_1 FILLER_42_630 ();
 sg13g2_decap_8 FILLER_42_635 ();
 sg13g2_decap_8 FILLER_42_642 ();
 sg13g2_decap_8 FILLER_42_649 ();
 sg13g2_decap_4 FILLER_42_669 ();
 sg13g2_fill_2 FILLER_42_697 ();
 sg13g2_fill_2 FILLER_42_709 ();
 sg13g2_fill_2 FILLER_42_728 ();
 sg13g2_fill_1 FILLER_42_733 ();
 sg13g2_fill_1 FILLER_42_759 ();
 sg13g2_fill_1 FILLER_42_765 ();
 sg13g2_fill_1 FILLER_42_775 ();
 sg13g2_decap_8 FILLER_42_785 ();
 sg13g2_decap_4 FILLER_42_792 ();
 sg13g2_fill_1 FILLER_42_838 ();
 sg13g2_decap_8 FILLER_42_843 ();
 sg13g2_decap_8 FILLER_42_850 ();
 sg13g2_fill_1 FILLER_42_857 ();
 sg13g2_decap_8 FILLER_42_888 ();
 sg13g2_decap_8 FILLER_42_895 ();
 sg13g2_decap_4 FILLER_42_902 ();
 sg13g2_fill_1 FILLER_42_911 ();
 sg13g2_fill_1 FILLER_42_938 ();
 sg13g2_fill_1 FILLER_42_943 ();
 sg13g2_decap_8 FILLER_42_991 ();
 sg13g2_fill_2 FILLER_42_998 ();
 sg13g2_fill_1 FILLER_42_1000 ();
 sg13g2_decap_8 FILLER_42_1015 ();
 sg13g2_fill_2 FILLER_42_1022 ();
 sg13g2_fill_1 FILLER_42_1038 ();
 sg13g2_decap_8 FILLER_42_1043 ();
 sg13g2_decap_8 FILLER_42_1050 ();
 sg13g2_fill_2 FILLER_42_1057 ();
 sg13g2_decap_4 FILLER_42_1063 ();
 sg13g2_fill_2 FILLER_42_1067 ();
 sg13g2_fill_2 FILLER_42_1079 ();
 sg13g2_fill_1 FILLER_42_1081 ();
 sg13g2_decap_8 FILLER_42_1092 ();
 sg13g2_decap_8 FILLER_42_1109 ();
 sg13g2_fill_1 FILLER_42_1116 ();
 sg13g2_fill_2 FILLER_42_1173 ();
 sg13g2_decap_4 FILLER_42_1203 ();
 sg13g2_fill_2 FILLER_42_1207 ();
 sg13g2_fill_2 FILLER_42_1217 ();
 sg13g2_fill_1 FILLER_42_1219 ();
 sg13g2_decap_4 FILLER_42_1261 ();
 sg13g2_fill_2 FILLER_42_1275 ();
 sg13g2_decap_8 FILLER_42_1303 ();
 sg13g2_decap_8 FILLER_42_1310 ();
 sg13g2_decap_8 FILLER_42_1317 ();
 sg13g2_fill_2 FILLER_42_1324 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_fill_2 FILLER_43_42 ();
 sg13g2_fill_2 FILLER_43_62 ();
 sg13g2_fill_1 FILLER_43_64 ();
 sg13g2_decap_8 FILLER_43_69 ();
 sg13g2_fill_2 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_78 ();
 sg13g2_fill_1 FILLER_43_89 ();
 sg13g2_decap_4 FILLER_43_139 ();
 sg13g2_fill_1 FILLER_43_143 ();
 sg13g2_decap_8 FILLER_43_148 ();
 sg13g2_fill_1 FILLER_43_155 ();
 sg13g2_decap_4 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_176 ();
 sg13g2_decap_8 FILLER_43_183 ();
 sg13g2_decap_8 FILLER_43_190 ();
 sg13g2_decap_8 FILLER_43_197 ();
 sg13g2_fill_2 FILLER_43_239 ();
 sg13g2_fill_2 FILLER_43_245 ();
 sg13g2_fill_1 FILLER_43_247 ();
 sg13g2_fill_1 FILLER_43_258 ();
 sg13g2_fill_2 FILLER_43_264 ();
 sg13g2_fill_2 FILLER_43_270 ();
 sg13g2_fill_2 FILLER_43_280 ();
 sg13g2_fill_1 FILLER_43_282 ();
 sg13g2_decap_8 FILLER_43_312 ();
 sg13g2_fill_1 FILLER_43_319 ();
 sg13g2_fill_1 FILLER_43_324 ();
 sg13g2_decap_4 FILLER_43_329 ();
 sg13g2_fill_2 FILLER_43_333 ();
 sg13g2_decap_8 FILLER_43_339 ();
 sg13g2_decap_8 FILLER_43_346 ();
 sg13g2_fill_1 FILLER_43_353 ();
 sg13g2_decap_8 FILLER_43_358 ();
 sg13g2_decap_4 FILLER_43_365 ();
 sg13g2_fill_2 FILLER_43_369 ();
 sg13g2_fill_1 FILLER_43_457 ();
 sg13g2_fill_1 FILLER_43_493 ();
 sg13g2_fill_2 FILLER_43_504 ();
 sg13g2_fill_1 FILLER_43_510 ();
 sg13g2_fill_1 FILLER_43_537 ();
 sg13g2_fill_1 FILLER_43_543 ();
 sg13g2_fill_2 FILLER_43_565 ();
 sg13g2_fill_2 FILLER_43_571 ();
 sg13g2_fill_1 FILLER_43_573 ();
 sg13g2_fill_2 FILLER_43_600 ();
 sg13g2_fill_1 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_607 ();
 sg13g2_decap_8 FILLER_43_614 ();
 sg13g2_decap_4 FILLER_43_621 ();
 sg13g2_decap_8 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_644 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_fill_2 FILLER_43_688 ();
 sg13g2_fill_1 FILLER_43_690 ();
 sg13g2_fill_1 FILLER_43_735 ();
 sg13g2_decap_4 FILLER_43_745 ();
 sg13g2_fill_1 FILLER_43_767 ();
 sg13g2_decap_4 FILLER_43_772 ();
 sg13g2_fill_2 FILLER_43_781 ();
 sg13g2_decap_4 FILLER_43_786 ();
 sg13g2_fill_1 FILLER_43_790 ();
 sg13g2_decap_8 FILLER_43_842 ();
 sg13g2_decap_8 FILLER_43_849 ();
 sg13g2_decap_4 FILLER_43_856 ();
 sg13g2_fill_2 FILLER_43_860 ();
 sg13g2_fill_1 FILLER_43_871 ();
 sg13g2_decap_8 FILLER_43_898 ();
 sg13g2_fill_2 FILLER_43_905 ();
 sg13g2_fill_2 FILLER_43_912 ();
 sg13g2_decap_8 FILLER_43_982 ();
 sg13g2_decap_8 FILLER_43_989 ();
 sg13g2_decap_8 FILLER_43_996 ();
 sg13g2_decap_8 FILLER_43_1003 ();
 sg13g2_decap_8 FILLER_43_1010 ();
 sg13g2_decap_8 FILLER_43_1017 ();
 sg13g2_decap_8 FILLER_43_1024 ();
 sg13g2_fill_2 FILLER_43_1031 ();
 sg13g2_fill_1 FILLER_43_1033 ();
 sg13g2_decap_4 FILLER_43_1037 ();
 sg13g2_fill_1 FILLER_43_1041 ();
 sg13g2_decap_8 FILLER_43_1068 ();
 sg13g2_decap_8 FILLER_43_1075 ();
 sg13g2_decap_8 FILLER_43_1082 ();
 sg13g2_decap_8 FILLER_43_1089 ();
 sg13g2_decap_4 FILLER_43_1096 ();
 sg13g2_fill_2 FILLER_43_1108 ();
 sg13g2_fill_1 FILLER_43_1110 ();
 sg13g2_decap_8 FILLER_43_1116 ();
 sg13g2_fill_1 FILLER_43_1123 ();
 sg13g2_decap_4 FILLER_43_1132 ();
 sg13g2_fill_2 FILLER_43_1136 ();
 sg13g2_decap_8 FILLER_43_1148 ();
 sg13g2_decap_8 FILLER_43_1155 ();
 sg13g2_fill_2 FILLER_43_1162 ();
 sg13g2_fill_1 FILLER_43_1164 ();
 sg13g2_fill_2 FILLER_43_1217 ();
 sg13g2_fill_1 FILLER_43_1219 ();
 sg13g2_decap_8 FILLER_43_1300 ();
 sg13g2_decap_8 FILLER_43_1307 ();
 sg13g2_decap_8 FILLER_43_1314 ();
 sg13g2_decap_4 FILLER_43_1321 ();
 sg13g2_fill_1 FILLER_43_1325 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_fill_1 FILLER_44_35 ();
 sg13g2_decap_4 FILLER_44_50 ();
 sg13g2_fill_1 FILLER_44_80 ();
 sg13g2_fill_1 FILLER_44_107 ();
 sg13g2_fill_2 FILLER_44_160 ();
 sg13g2_decap_8 FILLER_44_170 ();
 sg13g2_decap_8 FILLER_44_208 ();
 sg13g2_decap_8 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_222 ();
 sg13g2_decap_8 FILLER_44_229 ();
 sg13g2_decap_8 FILLER_44_236 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_decap_8 FILLER_44_271 ();
 sg13g2_decap_8 FILLER_44_278 ();
 sg13g2_decap_4 FILLER_44_285 ();
 sg13g2_fill_2 FILLER_44_289 ();
 sg13g2_decap_8 FILLER_44_296 ();
 sg13g2_decap_8 FILLER_44_303 ();
 sg13g2_fill_2 FILLER_44_310 ();
 sg13g2_fill_1 FILLER_44_312 ();
 sg13g2_decap_8 FILLER_44_318 ();
 sg13g2_fill_2 FILLER_44_325 ();
 sg13g2_decap_8 FILLER_44_340 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_decap_8 FILLER_44_356 ();
 sg13g2_decap_4 FILLER_44_363 ();
 sg13g2_decap_8 FILLER_44_372 ();
 sg13g2_decap_4 FILLER_44_379 ();
 sg13g2_fill_1 FILLER_44_383 ();
 sg13g2_fill_2 FILLER_44_410 ();
 sg13g2_fill_2 FILLER_44_425 ();
 sg13g2_fill_1 FILLER_44_432 ();
 sg13g2_fill_2 FILLER_44_437 ();
 sg13g2_fill_1 FILLER_44_443 ();
 sg13g2_fill_2 FILLER_44_454 ();
 sg13g2_fill_2 FILLER_44_466 ();
 sg13g2_decap_8 FILLER_44_472 ();
 sg13g2_decap_8 FILLER_44_479 ();
 sg13g2_fill_2 FILLER_44_486 ();
 sg13g2_fill_1 FILLER_44_488 ();
 sg13g2_fill_2 FILLER_44_612 ();
 sg13g2_fill_1 FILLER_44_614 ();
 sg13g2_fill_2 FILLER_44_619 ();
 sg13g2_fill_1 FILLER_44_621 ();
 sg13g2_decap_8 FILLER_44_648 ();
 sg13g2_decap_8 FILLER_44_655 ();
 sg13g2_fill_2 FILLER_44_662 ();
 sg13g2_fill_2 FILLER_44_668 ();
 sg13g2_fill_1 FILLER_44_674 ();
 sg13g2_fill_1 FILLER_44_679 ();
 sg13g2_fill_1 FILLER_44_690 ();
 sg13g2_decap_4 FILLER_44_697 ();
 sg13g2_fill_1 FILLER_44_701 ();
 sg13g2_fill_1 FILLER_44_707 ();
 sg13g2_fill_1 FILLER_44_728 ();
 sg13g2_fill_2 FILLER_44_733 ();
 sg13g2_decap_4 FILLER_44_739 ();
 sg13g2_fill_2 FILLER_44_765 ();
 sg13g2_fill_1 FILLER_44_771 ();
 sg13g2_fill_2 FILLER_44_777 ();
 sg13g2_fill_2 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_820 ();
 sg13g2_fill_2 FILLER_44_827 ();
 sg13g2_fill_1 FILLER_44_829 ();
 sg13g2_decap_8 FILLER_44_834 ();
 sg13g2_decap_8 FILLER_44_896 ();
 sg13g2_decap_8 FILLER_44_903 ();
 sg13g2_fill_2 FILLER_44_920 ();
 sg13g2_fill_1 FILLER_44_922 ();
 sg13g2_decap_8 FILLER_44_931 ();
 sg13g2_decap_4 FILLER_44_938 ();
 sg13g2_fill_2 FILLER_44_942 ();
 sg13g2_fill_1 FILLER_44_950 ();
 sg13g2_fill_2 FILLER_44_971 ();
 sg13g2_decap_4 FILLER_44_1003 ();
 sg13g2_fill_2 FILLER_44_1033 ();
 sg13g2_decap_4 FILLER_44_1065 ();
 sg13g2_decap_8 FILLER_44_1099 ();
 sg13g2_decap_8 FILLER_44_1106 ();
 sg13g2_decap_8 FILLER_44_1113 ();
 sg13g2_decap_8 FILLER_44_1146 ();
 sg13g2_decap_8 FILLER_44_1153 ();
 sg13g2_decap_8 FILLER_44_1160 ();
 sg13g2_decap_8 FILLER_44_1167 ();
 sg13g2_fill_1 FILLER_44_1174 ();
 sg13g2_fill_2 FILLER_44_1225 ();
 sg13g2_fill_1 FILLER_44_1227 ();
 sg13g2_fill_2 FILLER_44_1258 ();
 sg13g2_fill_2 FILLER_44_1286 ();
 sg13g2_decap_8 FILLER_44_1292 ();
 sg13g2_decap_8 FILLER_44_1299 ();
 sg13g2_decap_8 FILLER_44_1306 ();
 sg13g2_decap_8 FILLER_44_1313 ();
 sg13g2_decap_4 FILLER_44_1320 ();
 sg13g2_fill_2 FILLER_44_1324 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_77 ();
 sg13g2_fill_1 FILLER_45_82 ();
 sg13g2_decap_4 FILLER_45_118 ();
 sg13g2_fill_1 FILLER_45_122 ();
 sg13g2_fill_2 FILLER_45_144 ();
 sg13g2_decap_4 FILLER_45_150 ();
 sg13g2_fill_2 FILLER_45_154 ();
 sg13g2_decap_4 FILLER_45_174 ();
 sg13g2_fill_1 FILLER_45_178 ();
 sg13g2_decap_8 FILLER_45_200 ();
 sg13g2_decap_8 FILLER_45_207 ();
 sg13g2_decap_4 FILLER_45_214 ();
 sg13g2_fill_2 FILLER_45_218 ();
 sg13g2_decap_8 FILLER_45_225 ();
 sg13g2_decap_8 FILLER_45_232 ();
 sg13g2_decap_4 FILLER_45_239 ();
 sg13g2_fill_1 FILLER_45_243 ();
 sg13g2_fill_2 FILLER_45_258 ();
 sg13g2_decap_8 FILLER_45_286 ();
 sg13g2_decap_4 FILLER_45_293 ();
 sg13g2_fill_2 FILLER_45_297 ();
 sg13g2_decap_8 FILLER_45_303 ();
 sg13g2_decap_8 FILLER_45_310 ();
 sg13g2_decap_4 FILLER_45_321 ();
 sg13g2_fill_1 FILLER_45_325 ();
 sg13g2_decap_8 FILLER_45_335 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_decap_8 FILLER_45_349 ();
 sg13g2_decap_4 FILLER_45_356 ();
 sg13g2_fill_1 FILLER_45_379 ();
 sg13g2_fill_2 FILLER_45_388 ();
 sg13g2_fill_1 FILLER_45_390 ();
 sg13g2_fill_2 FILLER_45_395 ();
 sg13g2_fill_1 FILLER_45_397 ();
 sg13g2_fill_2 FILLER_45_442 ();
 sg13g2_fill_1 FILLER_45_444 ();
 sg13g2_decap_8 FILLER_45_452 ();
 sg13g2_fill_2 FILLER_45_459 ();
 sg13g2_fill_1 FILLER_45_461 ();
 sg13g2_decap_8 FILLER_45_466 ();
 sg13g2_decap_8 FILLER_45_473 ();
 sg13g2_decap_8 FILLER_45_480 ();
 sg13g2_decap_4 FILLER_45_487 ();
 sg13g2_fill_2 FILLER_45_491 ();
 sg13g2_fill_1 FILLER_45_516 ();
 sg13g2_decap_4 FILLER_45_553 ();
 sg13g2_fill_1 FILLER_45_557 ();
 sg13g2_decap_8 FILLER_45_562 ();
 sg13g2_decap_8 FILLER_45_569 ();
 sg13g2_fill_1 FILLER_45_576 ();
 sg13g2_decap_4 FILLER_45_658 ();
 sg13g2_fill_1 FILLER_45_662 ();
 sg13g2_decap_4 FILLER_45_668 ();
 sg13g2_fill_1 FILLER_45_672 ();
 sg13g2_fill_2 FILLER_45_682 ();
 sg13g2_fill_1 FILLER_45_684 ();
 sg13g2_fill_1 FILLER_45_694 ();
 sg13g2_fill_2 FILLER_45_700 ();
 sg13g2_fill_1 FILLER_45_716 ();
 sg13g2_fill_2 FILLER_45_734 ();
 sg13g2_fill_1 FILLER_45_744 ();
 sg13g2_fill_1 FILLER_45_761 ();
 sg13g2_fill_1 FILLER_45_797 ();
 sg13g2_fill_1 FILLER_45_807 ();
 sg13g2_fill_2 FILLER_45_818 ();
 sg13g2_decap_8 FILLER_45_825 ();
 sg13g2_decap_8 FILLER_45_832 ();
 sg13g2_fill_1 FILLER_45_876 ();
 sg13g2_fill_2 FILLER_45_881 ();
 sg13g2_decap_4 FILLER_45_887 ();
 sg13g2_fill_1 FILLER_45_891 ();
 sg13g2_decap_8 FILLER_45_896 ();
 sg13g2_fill_2 FILLER_45_903 ();
 sg13g2_decap_8 FILLER_45_939 ();
 sg13g2_decap_4 FILLER_45_946 ();
 sg13g2_decap_4 FILLER_45_956 ();
 sg13g2_decap_4 FILLER_45_992 ();
 sg13g2_fill_2 FILLER_45_1053 ();
 sg13g2_decap_4 FILLER_45_1068 ();
 sg13g2_fill_2 FILLER_45_1072 ();
 sg13g2_decap_4 FILLER_45_1098 ();
 sg13g2_decap_8 FILLER_45_1106 ();
 sg13g2_decap_4 FILLER_45_1113 ();
 sg13g2_fill_2 FILLER_45_1157 ();
 sg13g2_fill_1 FILLER_45_1159 ();
 sg13g2_fill_2 FILLER_45_1190 ();
 sg13g2_fill_1 FILLER_45_1192 ();
 sg13g2_decap_4 FILLER_45_1233 ();
 sg13g2_fill_2 FILLER_45_1241 ();
 sg13g2_fill_2 FILLER_45_1253 ();
 sg13g2_fill_1 FILLER_45_1255 ();
 sg13g2_fill_1 FILLER_45_1266 ();
 sg13g2_fill_2 FILLER_45_1271 ();
 sg13g2_fill_1 FILLER_45_1273 ();
 sg13g2_decap_8 FILLER_45_1288 ();
 sg13g2_decap_8 FILLER_45_1295 ();
 sg13g2_decap_8 FILLER_45_1302 ();
 sg13g2_decap_8 FILLER_45_1309 ();
 sg13g2_decap_8 FILLER_45_1316 ();
 sg13g2_fill_2 FILLER_45_1323 ();
 sg13g2_fill_1 FILLER_45_1325 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_15 ();
 sg13g2_fill_2 FILLER_46_22 ();
 sg13g2_fill_1 FILLER_46_42 ();
 sg13g2_decap_4 FILLER_46_47 ();
 sg13g2_fill_2 FILLER_46_55 ();
 sg13g2_fill_1 FILLER_46_78 ();
 sg13g2_fill_2 FILLER_46_89 ();
 sg13g2_fill_2 FILLER_46_95 ();
 sg13g2_decap_4 FILLER_46_101 ();
 sg13g2_decap_8 FILLER_46_114 ();
 sg13g2_fill_1 FILLER_46_121 ();
 sg13g2_decap_4 FILLER_46_143 ();
 sg13g2_fill_1 FILLER_46_214 ();
 sg13g2_fill_2 FILLER_46_241 ();
 sg13g2_fill_1 FILLER_46_243 ();
 sg13g2_fill_2 FILLER_46_265 ();
 sg13g2_decap_8 FILLER_46_307 ();
 sg13g2_decap_4 FILLER_46_314 ();
 sg13g2_fill_2 FILLER_46_333 ();
 sg13g2_fill_1 FILLER_46_335 ();
 sg13g2_fill_1 FILLER_46_378 ();
 sg13g2_decap_4 FILLER_46_389 ();
 sg13g2_fill_2 FILLER_46_393 ();
 sg13g2_decap_4 FILLER_46_400 ();
 sg13g2_fill_1 FILLER_46_404 ();
 sg13g2_fill_2 FILLER_46_414 ();
 sg13g2_decap_8 FILLER_46_435 ();
 sg13g2_fill_1 FILLER_46_442 ();
 sg13g2_fill_1 FILLER_46_454 ();
 sg13g2_decap_4 FILLER_46_466 ();
 sg13g2_fill_2 FILLER_46_474 ();
 sg13g2_fill_1 FILLER_46_528 ();
 sg13g2_fill_1 FILLER_46_539 ();
 sg13g2_fill_2 FILLER_46_544 ();
 sg13g2_fill_2 FILLER_46_554 ();
 sg13g2_fill_2 FILLER_46_566 ();
 sg13g2_decap_8 FILLER_46_572 ();
 sg13g2_decap_8 FILLER_46_579 ();
 sg13g2_decap_4 FILLER_46_586 ();
 sg13g2_fill_2 FILLER_46_590 ();
 sg13g2_fill_1 FILLER_46_596 ();
 sg13g2_fill_2 FILLER_46_605 ();
 sg13g2_fill_2 FILLER_46_615 ();
 sg13g2_fill_2 FILLER_46_623 ();
 sg13g2_fill_1 FILLER_46_635 ();
 sg13g2_fill_1 FILLER_46_641 ();
 sg13g2_fill_1 FILLER_46_646 ();
 sg13g2_decap_8 FILLER_46_657 ();
 sg13g2_decap_8 FILLER_46_664 ();
 sg13g2_decap_4 FILLER_46_675 ();
 sg13g2_fill_1 FILLER_46_679 ();
 sg13g2_fill_2 FILLER_46_712 ();
 sg13g2_fill_2 FILLER_46_718 ();
 sg13g2_fill_1 FILLER_46_720 ();
 sg13g2_fill_2 FILLER_46_744 ();
 sg13g2_fill_1 FILLER_46_746 ();
 sg13g2_fill_2 FILLER_46_757 ();
 sg13g2_fill_1 FILLER_46_764 ();
 sg13g2_decap_8 FILLER_46_774 ();
 sg13g2_fill_2 FILLER_46_781 ();
 sg13g2_fill_1 FILLER_46_783 ();
 sg13g2_decap_4 FILLER_46_790 ();
 sg13g2_fill_1 FILLER_46_794 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_fill_1 FILLER_46_819 ();
 sg13g2_decap_4 FILLER_46_837 ();
 sg13g2_fill_2 FILLER_46_841 ();
 sg13g2_decap_4 FILLER_46_851 ();
 sg13g2_fill_1 FILLER_46_855 ();
 sg13g2_fill_1 FILLER_46_859 ();
 sg13g2_fill_2 FILLER_46_864 ();
 sg13g2_decap_4 FILLER_46_877 ();
 sg13g2_decap_8 FILLER_46_886 ();
 sg13g2_decap_4 FILLER_46_893 ();
 sg13g2_decap_8 FILLER_46_905 ();
 sg13g2_fill_2 FILLER_46_912 ();
 sg13g2_fill_1 FILLER_46_914 ();
 sg13g2_decap_4 FILLER_46_927 ();
 sg13g2_fill_1 FILLER_46_931 ();
 sg13g2_decap_4 FILLER_46_1004 ();
 sg13g2_fill_1 FILLER_46_1008 ();
 sg13g2_decap_8 FILLER_46_1017 ();
 sg13g2_decap_4 FILLER_46_1024 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_fill_1 FILLER_46_1050 ();
 sg13g2_decap_8 FILLER_46_1059 ();
 sg13g2_fill_1 FILLER_46_1066 ();
 sg13g2_decap_4 FILLER_46_1119 ();
 sg13g2_decap_8 FILLER_46_1127 ();
 sg13g2_fill_2 FILLER_46_1134 ();
 sg13g2_decap_8 FILLER_46_1188 ();
 sg13g2_decap_8 FILLER_46_1195 ();
 sg13g2_decap_4 FILLER_46_1202 ();
 sg13g2_decap_8 FILLER_46_1210 ();
 sg13g2_decap_4 FILLER_46_1217 ();
 sg13g2_fill_1 FILLER_46_1221 ();
 sg13g2_decap_8 FILLER_46_1232 ();
 sg13g2_decap_8 FILLER_46_1239 ();
 sg13g2_decap_8 FILLER_46_1246 ();
 sg13g2_decap_4 FILLER_46_1253 ();
 sg13g2_fill_2 FILLER_46_1257 ();
 sg13g2_decap_8 FILLER_46_1301 ();
 sg13g2_decap_8 FILLER_46_1308 ();
 sg13g2_decap_8 FILLER_46_1315 ();
 sg13g2_decap_4 FILLER_46_1322 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_75 ();
 sg13g2_fill_2 FILLER_47_86 ();
 sg13g2_fill_1 FILLER_47_88 ();
 sg13g2_fill_1 FILLER_47_93 ();
 sg13g2_decap_8 FILLER_47_120 ();
 sg13g2_decap_8 FILLER_47_127 ();
 sg13g2_decap_8 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_141 ();
 sg13g2_fill_1 FILLER_47_182 ();
 sg13g2_fill_2 FILLER_47_187 ();
 sg13g2_fill_2 FILLER_47_193 ();
 sg13g2_fill_2 FILLER_47_262 ();
 sg13g2_fill_1 FILLER_47_264 ();
 sg13g2_decap_4 FILLER_47_281 ();
 sg13g2_fill_1 FILLER_47_285 ();
 sg13g2_fill_1 FILLER_47_296 ();
 sg13g2_decap_4 FILLER_47_342 ();
 sg13g2_fill_2 FILLER_47_352 ();
 sg13g2_fill_1 FILLER_47_354 ();
 sg13g2_decap_4 FILLER_47_385 ();
 sg13g2_fill_2 FILLER_47_389 ();
 sg13g2_fill_2 FILLER_47_395 ();
 sg13g2_decap_8 FILLER_47_412 ();
 sg13g2_decap_8 FILLER_47_419 ();
 sg13g2_fill_2 FILLER_47_426 ();
 sg13g2_fill_1 FILLER_47_428 ();
 sg13g2_decap_8 FILLER_47_433 ();
 sg13g2_decap_4 FILLER_47_440 ();
 sg13g2_fill_1 FILLER_47_444 ();
 sg13g2_decap_8 FILLER_47_450 ();
 sg13g2_decap_4 FILLER_47_457 ();
 sg13g2_fill_1 FILLER_47_461 ();
 sg13g2_fill_1 FILLER_47_466 ();
 sg13g2_fill_2 FILLER_47_507 ();
 sg13g2_fill_2 FILLER_47_513 ();
 sg13g2_fill_1 FILLER_47_515 ();
 sg13g2_fill_1 FILLER_47_537 ();
 sg13g2_fill_2 FILLER_47_559 ();
 sg13g2_fill_1 FILLER_47_561 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_fill_2 FILLER_47_616 ();
 sg13g2_fill_2 FILLER_47_631 ();
 sg13g2_fill_1 FILLER_47_633 ();
 sg13g2_decap_8 FILLER_47_642 ();
 sg13g2_fill_2 FILLER_47_649 ();
 sg13g2_fill_2 FILLER_47_656 ();
 sg13g2_fill_1 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_663 ();
 sg13g2_fill_2 FILLER_47_670 ();
 sg13g2_fill_2 FILLER_47_680 ();
 sg13g2_fill_2 FILLER_47_708 ();
 sg13g2_fill_1 FILLER_47_710 ();
 sg13g2_fill_2 FILLER_47_773 ();
 sg13g2_decap_4 FILLER_47_780 ();
 sg13g2_decap_4 FILLER_47_789 ();
 sg13g2_decap_8 FILLER_47_811 ();
 sg13g2_decap_8 FILLER_47_818 ();
 sg13g2_decap_8 FILLER_47_858 ();
 sg13g2_fill_2 FILLER_47_869 ();
 sg13g2_fill_2 FILLER_47_880 ();
 sg13g2_fill_1 FILLER_47_882 ();
 sg13g2_fill_2 FILLER_47_887 ();
 sg13g2_decap_4 FILLER_47_923 ();
 sg13g2_fill_1 FILLER_47_960 ();
 sg13g2_fill_1 FILLER_47_967 ();
 sg13g2_fill_1 FILLER_47_971 ();
 sg13g2_fill_1 FILLER_47_976 ();
 sg13g2_decap_8 FILLER_47_981 ();
 sg13g2_decap_4 FILLER_47_988 ();
 sg13g2_decap_8 FILLER_47_997 ();
 sg13g2_decap_8 FILLER_47_1004 ();
 sg13g2_decap_4 FILLER_47_1011 ();
 sg13g2_fill_2 FILLER_47_1015 ();
 sg13g2_fill_2 FILLER_47_1047 ();
 sg13g2_decap_8 FILLER_47_1075 ();
 sg13g2_fill_2 FILLER_47_1082 ();
 sg13g2_fill_1 FILLER_47_1094 ();
 sg13g2_fill_1 FILLER_47_1099 ();
 sg13g2_decap_4 FILLER_47_1126 ();
 sg13g2_fill_2 FILLER_47_1130 ();
 sg13g2_fill_1 FILLER_47_1140 ();
 sg13g2_fill_2 FILLER_47_1197 ();
 sg13g2_decap_4 FILLER_47_1229 ();
 sg13g2_decap_8 FILLER_47_1241 ();
 sg13g2_fill_1 FILLER_47_1248 ();
 sg13g2_decap_8 FILLER_47_1267 ();
 sg13g2_fill_2 FILLER_47_1274 ();
 sg13g2_decap_8 FILLER_47_1286 ();
 sg13g2_decap_4 FILLER_47_1293 ();
 sg13g2_fill_1 FILLER_47_1297 ();
 sg13g2_fill_2 FILLER_47_1324 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_4 ();
 sg13g2_fill_1 FILLER_48_26 ();
 sg13g2_decap_4 FILLER_48_82 ();
 sg13g2_fill_1 FILLER_48_86 ();
 sg13g2_decap_8 FILLER_48_134 ();
 sg13g2_fill_1 FILLER_48_141 ();
 sg13g2_decap_8 FILLER_48_176 ();
 sg13g2_decap_8 FILLER_48_183 ();
 sg13g2_decap_8 FILLER_48_190 ();
 sg13g2_fill_1 FILLER_48_218 ();
 sg13g2_decap_8 FILLER_48_223 ();
 sg13g2_fill_2 FILLER_48_230 ();
 sg13g2_fill_1 FILLER_48_232 ();
 sg13g2_fill_1 FILLER_48_237 ();
 sg13g2_decap_8 FILLER_48_309 ();
 sg13g2_decap_8 FILLER_48_316 ();
 sg13g2_decap_8 FILLER_48_323 ();
 sg13g2_decap_8 FILLER_48_330 ();
 sg13g2_decap_4 FILLER_48_337 ();
 sg13g2_fill_2 FILLER_48_341 ();
 sg13g2_decap_8 FILLER_48_353 ();
 sg13g2_fill_1 FILLER_48_360 ();
 sg13g2_decap_8 FILLER_48_365 ();
 sg13g2_fill_1 FILLER_48_372 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_fill_2 FILLER_48_434 ();
 sg13g2_fill_2 FILLER_48_445 ();
 sg13g2_decap_4 FILLER_48_452 ();
 sg13g2_fill_1 FILLER_48_456 ();
 sg13g2_decap_4 FILLER_48_465 ();
 sg13g2_fill_2 FILLER_48_481 ();
 sg13g2_fill_2 FILLER_48_496 ();
 sg13g2_fill_2 FILLER_48_524 ();
 sg13g2_fill_1 FILLER_48_547 ();
 sg13g2_fill_1 FILLER_48_564 ();
 sg13g2_fill_2 FILLER_48_572 ();
 sg13g2_decap_4 FILLER_48_578 ();
 sg13g2_fill_1 FILLER_48_582 ();
 sg13g2_fill_1 FILLER_48_629 ();
 sg13g2_decap_4 FILLER_48_645 ();
 sg13g2_fill_2 FILLER_48_658 ();
 sg13g2_fill_1 FILLER_48_660 ();
 sg13g2_decap_4 FILLER_48_665 ();
 sg13g2_fill_1 FILLER_48_676 ();
 sg13g2_decap_4 FILLER_48_681 ();
 sg13g2_fill_1 FILLER_48_685 ();
 sg13g2_decap_4 FILLER_48_690 ();
 sg13g2_fill_2 FILLER_48_694 ();
 sg13g2_fill_2 FILLER_48_730 ();
 sg13g2_decap_4 FILLER_48_736 ();
 sg13g2_fill_1 FILLER_48_745 ();
 sg13g2_fill_1 FILLER_48_753 ();
 sg13g2_fill_1 FILLER_48_758 ();
 sg13g2_fill_1 FILLER_48_764 ();
 sg13g2_fill_1 FILLER_48_791 ();
 sg13g2_fill_1 FILLER_48_818 ();
 sg13g2_decap_4 FILLER_48_865 ();
 sg13g2_fill_2 FILLER_48_874 ();
 sg13g2_decap_4 FILLER_48_880 ();
 sg13g2_fill_1 FILLER_48_884 ();
 sg13g2_fill_2 FILLER_48_931 ();
 sg13g2_fill_2 FILLER_48_942 ();
 sg13g2_decap_8 FILLER_48_965 ();
 sg13g2_decap_8 FILLER_48_972 ();
 sg13g2_decap_4 FILLER_48_979 ();
 sg13g2_fill_2 FILLER_48_983 ();
 sg13g2_decap_8 FILLER_48_989 ();
 sg13g2_fill_1 FILLER_48_996 ();
 sg13g2_decap_4 FILLER_48_1001 ();
 sg13g2_fill_2 FILLER_48_1016 ();
 sg13g2_fill_1 FILLER_48_1018 ();
 sg13g2_fill_2 FILLER_48_1034 ();
 sg13g2_fill_2 FILLER_48_1044 ();
 sg13g2_fill_1 FILLER_48_1046 ();
 sg13g2_fill_2 FILLER_48_1053 ();
 sg13g2_decap_8 FILLER_48_1081 ();
 sg13g2_decap_4 FILLER_48_1088 ();
 sg13g2_fill_1 FILLER_48_1092 ();
 sg13g2_decap_8 FILLER_48_1107 ();
 sg13g2_decap_8 FILLER_48_1114 ();
 sg13g2_decap_8 FILLER_48_1121 ();
 sg13g2_fill_1 FILLER_48_1128 ();
 sg13g2_decap_8 FILLER_48_1191 ();
 sg13g2_decap_4 FILLER_48_1198 ();
 sg13g2_fill_1 FILLER_48_1202 ();
 sg13g2_fill_2 FILLER_48_1239 ();
 sg13g2_fill_2 FILLER_48_1267 ();
 sg13g2_fill_1 FILLER_48_1295 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_7 ();
 sg13g2_decap_4 FILLER_49_12 ();
 sg13g2_fill_1 FILLER_49_76 ();
 sg13g2_decap_4 FILLER_49_91 ();
 sg13g2_fill_1 FILLER_49_95 ();
 sg13g2_fill_2 FILLER_49_100 ();
 sg13g2_fill_1 FILLER_49_102 ();
 sg13g2_fill_2 FILLER_49_155 ();
 sg13g2_fill_1 FILLER_49_157 ();
 sg13g2_fill_2 FILLER_49_174 ();
 sg13g2_fill_1 FILLER_49_176 ();
 sg13g2_decap_4 FILLER_49_187 ();
 sg13g2_fill_1 FILLER_49_191 ();
 sg13g2_decap_4 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_228 ();
 sg13g2_decap_4 FILLER_49_235 ();
 sg13g2_fill_1 FILLER_49_239 ();
 sg13g2_decap_4 FILLER_49_244 ();
 sg13g2_fill_2 FILLER_49_248 ();
 sg13g2_decap_4 FILLER_49_254 ();
 sg13g2_decap_8 FILLER_49_268 ();
 sg13g2_decap_8 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_282 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_4 FILLER_49_347 ();
 sg13g2_fill_1 FILLER_49_387 ();
 sg13g2_decap_4 FILLER_49_414 ();
 sg13g2_decap_8 FILLER_49_422 ();
 sg13g2_fill_2 FILLER_49_429 ();
 sg13g2_fill_1 FILLER_49_431 ();
 sg13g2_decap_4 FILLER_49_436 ();
 sg13g2_fill_2 FILLER_49_440 ();
 sg13g2_fill_2 FILLER_49_523 ();
 sg13g2_decap_8 FILLER_49_559 ();
 sg13g2_fill_2 FILLER_49_566 ();
 sg13g2_fill_1 FILLER_49_568 ();
 sg13g2_fill_1 FILLER_49_590 ();
 sg13g2_fill_1 FILLER_49_640 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_fill_2 FILLER_49_700 ();
 sg13g2_decap_4 FILLER_49_719 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_759 ();
 sg13g2_decap_4 FILLER_49_766 ();
 sg13g2_fill_1 FILLER_49_770 ();
 sg13g2_fill_1 FILLER_49_775 ();
 sg13g2_decap_8 FILLER_49_785 ();
 sg13g2_decap_4 FILLER_49_792 ();
 sg13g2_decap_8 FILLER_49_807 ();
 sg13g2_decap_8 FILLER_49_814 ();
 sg13g2_decap_4 FILLER_49_821 ();
 sg13g2_fill_1 FILLER_49_825 ();
 sg13g2_fill_2 FILLER_49_829 ();
 sg13g2_fill_1 FILLER_49_835 ();
 sg13g2_fill_1 FILLER_49_850 ();
 sg13g2_fill_2 FILLER_49_899 ();
 sg13g2_fill_1 FILLER_49_901 ();
 sg13g2_decap_4 FILLER_49_906 ();
 sg13g2_fill_1 FILLER_49_910 ();
 sg13g2_fill_2 FILLER_49_915 ();
 sg13g2_fill_1 FILLER_49_917 ();
 sg13g2_fill_1 FILLER_49_944 ();
 sg13g2_decap_8 FILLER_49_950 ();
 sg13g2_decap_8 FILLER_49_957 ();
 sg13g2_decap_4 FILLER_49_964 ();
 sg13g2_fill_1 FILLER_49_968 ();
 sg13g2_fill_2 FILLER_49_1042 ();
 sg13g2_fill_1 FILLER_49_1063 ();
 sg13g2_decap_8 FILLER_49_1068 ();
 sg13g2_decap_8 FILLER_49_1075 ();
 sg13g2_fill_2 FILLER_49_1082 ();
 sg13g2_decap_4 FILLER_49_1120 ();
 sg13g2_decap_8 FILLER_49_1128 ();
 sg13g2_decap_8 FILLER_49_1135 ();
 sg13g2_fill_2 FILLER_49_1152 ();
 sg13g2_decap_8 FILLER_49_1190 ();
 sg13g2_decap_4 FILLER_49_1197 ();
 sg13g2_fill_1 FILLER_49_1215 ();
 sg13g2_fill_1 FILLER_49_1220 ();
 sg13g2_fill_2 FILLER_49_1251 ();
 sg13g2_fill_1 FILLER_49_1253 ();
 sg13g2_decap_8 FILLER_49_1264 ();
 sg13g2_decap_8 FILLER_49_1271 ();
 sg13g2_fill_2 FILLER_49_1282 ();
 sg13g2_fill_1 FILLER_49_1284 ();
 sg13g2_decap_8 FILLER_49_1319 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_4 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_95 ();
 sg13g2_decap_4 FILLER_50_156 ();
 sg13g2_fill_1 FILLER_50_174 ();
 sg13g2_decap_8 FILLER_50_211 ();
 sg13g2_decap_4 FILLER_50_218 ();
 sg13g2_fill_1 FILLER_50_222 ();
 sg13g2_fill_1 FILLER_50_228 ();
 sg13g2_fill_2 FILLER_50_255 ();
 sg13g2_fill_1 FILLER_50_261 ();
 sg13g2_fill_2 FILLER_50_272 ();
 sg13g2_decap_8 FILLER_50_300 ();
 sg13g2_decap_8 FILLER_50_307 ();
 sg13g2_fill_1 FILLER_50_314 ();
 sg13g2_decap_4 FILLER_50_336 ();
 sg13g2_fill_1 FILLER_50_340 ();
 sg13g2_decap_8 FILLER_50_380 ();
 sg13g2_decap_8 FILLER_50_387 ();
 sg13g2_decap_8 FILLER_50_398 ();
 sg13g2_decap_8 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_50_412 ();
 sg13g2_decap_8 FILLER_50_419 ();
 sg13g2_decap_8 FILLER_50_467 ();
 sg13g2_decap_8 FILLER_50_474 ();
 sg13g2_decap_8 FILLER_50_481 ();
 sg13g2_fill_1 FILLER_50_488 ();
 sg13g2_decap_8 FILLER_50_493 ();
 sg13g2_fill_2 FILLER_50_500 ();
 sg13g2_fill_1 FILLER_50_502 ();
 sg13g2_fill_1 FILLER_50_507 ();
 sg13g2_decap_8 FILLER_50_512 ();
 sg13g2_decap_4 FILLER_50_540 ();
 sg13g2_decap_4 FILLER_50_565 ();
 sg13g2_fill_1 FILLER_50_569 ();
 sg13g2_fill_1 FILLER_50_629 ();
 sg13g2_fill_2 FILLER_50_674 ();
 sg13g2_fill_2 FILLER_50_682 ();
 sg13g2_fill_1 FILLER_50_684 ();
 sg13g2_fill_2 FILLER_50_698 ();
 sg13g2_fill_1 FILLER_50_700 ();
 sg13g2_fill_2 FILLER_50_709 ();
 sg13g2_fill_1 FILLER_50_711 ();
 sg13g2_decap_8 FILLER_50_717 ();
 sg13g2_fill_2 FILLER_50_724 ();
 sg13g2_fill_1 FILLER_50_726 ();
 sg13g2_decap_8 FILLER_50_732 ();
 sg13g2_decap_8 FILLER_50_739 ();
 sg13g2_decap_8 FILLER_50_746 ();
 sg13g2_decap_8 FILLER_50_753 ();
 sg13g2_fill_2 FILLER_50_760 ();
 sg13g2_fill_1 FILLER_50_762 ();
 sg13g2_decap_8 FILLER_50_767 ();
 sg13g2_decap_8 FILLER_50_774 ();
 sg13g2_decap_8 FILLER_50_781 ();
 sg13g2_decap_8 FILLER_50_788 ();
 sg13g2_fill_1 FILLER_50_795 ();
 sg13g2_decap_4 FILLER_50_843 ();
 sg13g2_fill_1 FILLER_50_847 ();
 sg13g2_fill_1 FILLER_50_853 ();
 sg13g2_fill_1 FILLER_50_860 ();
 sg13g2_fill_2 FILLER_50_866 ();
 sg13g2_fill_1 FILLER_50_868 ();
 sg13g2_fill_2 FILLER_50_878 ();
 sg13g2_fill_1 FILLER_50_880 ();
 sg13g2_decap_4 FILLER_50_886 ();
 sg13g2_fill_1 FILLER_50_890 ();
 sg13g2_fill_1 FILLER_50_924 ();
 sg13g2_fill_1 FILLER_50_930 ();
 sg13g2_fill_1 FILLER_50_935 ();
 sg13g2_fill_1 FILLER_50_948 ();
 sg13g2_fill_2 FILLER_50_954 ();
 sg13g2_fill_2 FILLER_50_960 ();
 sg13g2_decap_8 FILLER_50_971 ();
 sg13g2_fill_1 FILLER_50_978 ();
 sg13g2_decap_8 FILLER_50_983 ();
 sg13g2_decap_8 FILLER_50_1023 ();
 sg13g2_fill_2 FILLER_50_1048 ();
 sg13g2_fill_1 FILLER_50_1054 ();
 sg13g2_decap_4 FILLER_50_1060 ();
 sg13g2_decap_8 FILLER_50_1068 ();
 sg13g2_decap_4 FILLER_50_1075 ();
 sg13g2_fill_1 FILLER_50_1079 ();
 sg13g2_fill_2 FILLER_50_1124 ();
 sg13g2_fill_1 FILLER_50_1126 ();
 sg13g2_decap_4 FILLER_50_1163 ();
 sg13g2_fill_2 FILLER_50_1167 ();
 sg13g2_fill_2 FILLER_50_1173 ();
 sg13g2_fill_2 FILLER_50_1179 ();
 sg13g2_fill_2 FILLER_50_1237 ();
 sg13g2_decap_8 FILLER_50_1265 ();
 sg13g2_decap_8 FILLER_50_1272 ();
 sg13g2_decap_8 FILLER_50_1279 ();
 sg13g2_decap_8 FILLER_50_1286 ();
 sg13g2_fill_1 FILLER_50_1293 ();
 sg13g2_fill_2 FILLER_50_1324 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_fill_1 FILLER_51_11 ();
 sg13g2_fill_2 FILLER_51_22 ();
 sg13g2_decap_4 FILLER_51_32 ();
 sg13g2_fill_1 FILLER_51_36 ();
 sg13g2_fill_2 FILLER_51_55 ();
 sg13g2_fill_1 FILLER_51_57 ();
 sg13g2_fill_2 FILLER_51_72 ();
 sg13g2_decap_4 FILLER_51_78 ();
 sg13g2_fill_2 FILLER_51_82 ();
 sg13g2_fill_2 FILLER_51_94 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_4 FILLER_51_217 ();
 sg13g2_fill_1 FILLER_51_221 ();
 sg13g2_fill_2 FILLER_51_244 ();
 sg13g2_fill_1 FILLER_51_275 ();
 sg13g2_decap_8 FILLER_51_302 ();
 sg13g2_decap_8 FILLER_51_309 ();
 sg13g2_fill_1 FILLER_51_316 ();
 sg13g2_fill_1 FILLER_51_327 ();
 sg13g2_decap_4 FILLER_51_332 ();
 sg13g2_decap_8 FILLER_51_370 ();
 sg13g2_decap_8 FILLER_51_377 ();
 sg13g2_decap_8 FILLER_51_384 ();
 sg13g2_decap_8 FILLER_51_391 ();
 sg13g2_fill_2 FILLER_51_398 ();
 sg13g2_fill_1 FILLER_51_400 ();
 sg13g2_decap_4 FILLER_51_405 ();
 sg13g2_fill_2 FILLER_51_409 ();
 sg13g2_fill_2 FILLER_51_437 ();
 sg13g2_decap_8 FILLER_51_470 ();
 sg13g2_decap_8 FILLER_51_477 ();
 sg13g2_decap_8 FILLER_51_484 ();
 sg13g2_decap_8 FILLER_51_491 ();
 sg13g2_decap_8 FILLER_51_498 ();
 sg13g2_decap_8 FILLER_51_505 ();
 sg13g2_decap_8 FILLER_51_512 ();
 sg13g2_decap_8 FILLER_51_540 ();
 sg13g2_fill_2 FILLER_51_547 ();
 sg13g2_decap_4 FILLER_51_575 ();
 sg13g2_fill_1 FILLER_51_579 ();
 sg13g2_fill_2 FILLER_51_585 ();
 sg13g2_fill_1 FILLER_51_587 ();
 sg13g2_fill_1 FILLER_51_592 ();
 sg13g2_decap_8 FILLER_51_598 ();
 sg13g2_decap_4 FILLER_51_605 ();
 sg13g2_decap_4 FILLER_51_622 ();
 sg13g2_fill_1 FILLER_51_626 ();
 sg13g2_fill_2 FILLER_51_632 ();
 sg13g2_decap_4 FILLER_51_647 ();
 sg13g2_fill_1 FILLER_51_651 ();
 sg13g2_decap_4 FILLER_51_664 ();
 sg13g2_fill_2 FILLER_51_725 ();
 sg13g2_fill_1 FILLER_51_741 ();
 sg13g2_decap_4 FILLER_51_773 ();
 sg13g2_fill_1 FILLER_51_777 ();
 sg13g2_fill_1 FILLER_51_782 ();
 sg13g2_decap_8 FILLER_51_793 ();
 sg13g2_decap_8 FILLER_51_800 ();
 sg13g2_decap_8 FILLER_51_807 ();
 sg13g2_fill_2 FILLER_51_814 ();
 sg13g2_fill_1 FILLER_51_816 ();
 sg13g2_fill_1 FILLER_51_840 ();
 sg13g2_fill_1 FILLER_51_847 ();
 sg13g2_fill_1 FILLER_51_867 ();
 sg13g2_decap_8 FILLER_51_874 ();
 sg13g2_decap_8 FILLER_51_881 ();
 sg13g2_decap_8 FILLER_51_888 ();
 sg13g2_decap_8 FILLER_51_895 ();
 sg13g2_fill_2 FILLER_51_902 ();
 sg13g2_fill_1 FILLER_51_904 ();
 sg13g2_fill_2 FILLER_51_909 ();
 sg13g2_fill_1 FILLER_51_934 ();
 sg13g2_fill_2 FILLER_51_985 ();
 sg13g2_fill_1 FILLER_51_987 ();
 sg13g2_fill_1 FILLER_51_994 ();
 sg13g2_fill_2 FILLER_51_1004 ();
 sg13g2_fill_1 FILLER_51_1006 ();
 sg13g2_fill_2 FILLER_51_1032 ();
 sg13g2_fill_1 FILLER_51_1034 ();
 sg13g2_decap_8 FILLER_51_1065 ();
 sg13g2_fill_2 FILLER_51_1072 ();
 sg13g2_fill_1 FILLER_51_1074 ();
 sg13g2_fill_1 FILLER_51_1109 ();
 sg13g2_fill_1 FILLER_51_1140 ();
 sg13g2_fill_2 FILLER_51_1167 ();
 sg13g2_decap_8 FILLER_51_1179 ();
 sg13g2_decap_8 FILLER_51_1186 ();
 sg13g2_decap_4 FILLER_51_1193 ();
 sg13g2_fill_2 FILLER_51_1237 ();
 sg13g2_decap_8 FILLER_51_1277 ();
 sg13g2_fill_2 FILLER_51_1294 ();
 sg13g2_decap_8 FILLER_51_1310 ();
 sg13g2_decap_8 FILLER_51_1317 ();
 sg13g2_fill_2 FILLER_51_1324 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_fill_2 FILLER_52_46 ();
 sg13g2_fill_1 FILLER_52_48 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_2 FILLER_52_89 ();
 sg13g2_decap_8 FILLER_52_113 ();
 sg13g2_decap_8 FILLER_52_120 ();
 sg13g2_decap_8 FILLER_52_127 ();
 sg13g2_decap_8 FILLER_52_134 ();
 sg13g2_decap_8 FILLER_52_141 ();
 sg13g2_decap_4 FILLER_52_188 ();
 sg13g2_fill_1 FILLER_52_192 ();
 sg13g2_decap_4 FILLER_52_214 ();
 sg13g2_fill_2 FILLER_52_218 ();
 sg13g2_fill_2 FILLER_52_224 ();
 sg13g2_fill_1 FILLER_52_234 ();
 sg13g2_decap_8 FILLER_52_239 ();
 sg13g2_fill_2 FILLER_52_246 ();
 sg13g2_fill_2 FILLER_52_297 ();
 sg13g2_fill_1 FILLER_52_299 ();
 sg13g2_fill_1 FILLER_52_347 ();
 sg13g2_decap_4 FILLER_52_390 ();
 sg13g2_fill_2 FILLER_52_402 ();
 sg13g2_fill_1 FILLER_52_404 ();
 sg13g2_fill_1 FILLER_52_415 ();
 sg13g2_fill_1 FILLER_52_468 ();
 sg13g2_decap_4 FILLER_52_513 ();
 sg13g2_decap_4 FILLER_52_546 ();
 sg13g2_fill_1 FILLER_52_550 ();
 sg13g2_fill_1 FILLER_52_572 ();
 sg13g2_fill_2 FILLER_52_633 ();
 sg13g2_decap_8 FILLER_52_642 ();
 sg13g2_decap_4 FILLER_52_649 ();
 sg13g2_fill_1 FILLER_52_653 ();
 sg13g2_decap_8 FILLER_52_662 ();
 sg13g2_decap_4 FILLER_52_669 ();
 sg13g2_decap_8 FILLER_52_677 ();
 sg13g2_decap_4 FILLER_52_684 ();
 sg13g2_fill_2 FILLER_52_688 ();
 sg13g2_fill_1 FILLER_52_694 ();
 sg13g2_fill_1 FILLER_52_701 ();
 sg13g2_fill_1 FILLER_52_728 ();
 sg13g2_fill_2 FILLER_52_759 ();
 sg13g2_fill_1 FILLER_52_788 ();
 sg13g2_fill_2 FILLER_52_794 ();
 sg13g2_decap_8 FILLER_52_807 ();
 sg13g2_fill_2 FILLER_52_814 ();
 sg13g2_fill_1 FILLER_52_825 ();
 sg13g2_fill_1 FILLER_52_837 ();
 sg13g2_decap_8 FILLER_52_879 ();
 sg13g2_fill_1 FILLER_52_886 ();
 sg13g2_decap_4 FILLER_52_892 ();
 sg13g2_fill_1 FILLER_52_896 ();
 sg13g2_fill_1 FILLER_52_901 ();
 sg13g2_fill_2 FILLER_52_907 ();
 sg13g2_fill_1 FILLER_52_909 ();
 sg13g2_fill_2 FILLER_52_914 ();
 sg13g2_decap_4 FILLER_52_937 ();
 sg13g2_fill_2 FILLER_52_941 ();
 sg13g2_fill_2 FILLER_52_947 ();
 sg13g2_fill_1 FILLER_52_954 ();
 sg13g2_decap_4 FILLER_52_962 ();
 sg13g2_fill_2 FILLER_52_966 ();
 sg13g2_fill_1 FILLER_52_978 ();
 sg13g2_fill_2 FILLER_52_1012 ();
 sg13g2_fill_1 FILLER_52_1040 ();
 sg13g2_fill_2 FILLER_52_1067 ();
 sg13g2_decap_4 FILLER_52_1129 ();
 sg13g2_fill_1 FILLER_52_1133 ();
 sg13g2_fill_2 FILLER_52_1156 ();
 sg13g2_fill_2 FILLER_52_1166 ();
 sg13g2_fill_1 FILLER_52_1194 ();
 sg13g2_fill_1 FILLER_52_1203 ();
 sg13g2_fill_2 FILLER_52_1214 ();
 sg13g2_fill_2 FILLER_52_1220 ();
 sg13g2_fill_2 FILLER_52_1232 ();
 sg13g2_decap_8 FILLER_52_1290 ();
 sg13g2_fill_1 FILLER_52_1297 ();
 sg13g2_fill_2 FILLER_52_1324 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_14 ();
 sg13g2_fill_1 FILLER_53_16 ();
 sg13g2_decap_4 FILLER_53_25 ();
 sg13g2_decap_4 FILLER_53_43 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_fill_2 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_76 ();
 sg13g2_fill_2 FILLER_53_83 ();
 sg13g2_decap_4 FILLER_53_89 ();
 sg13g2_decap_4 FILLER_53_97 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_8 FILLER_53_161 ();
 sg13g2_fill_2 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_183 ();
 sg13g2_decap_8 FILLER_53_190 ();
 sg13g2_decap_8 FILLER_53_197 ();
 sg13g2_decap_8 FILLER_53_204 ();
 sg13g2_decap_4 FILLER_53_211 ();
 sg13g2_decap_8 FILLER_53_219 ();
 sg13g2_fill_2 FILLER_53_226 ();
 sg13g2_decap_8 FILLER_53_242 ();
 sg13g2_decap_8 FILLER_53_249 ();
 sg13g2_fill_2 FILLER_53_256 ();
 sg13g2_fill_1 FILLER_53_258 ();
 sg13g2_decap_8 FILLER_53_267 ();
 sg13g2_decap_4 FILLER_53_278 ();
 sg13g2_decap_4 FILLER_53_286 ();
 sg13g2_fill_2 FILLER_53_290 ();
 sg13g2_decap_8 FILLER_53_313 ();
 sg13g2_decap_8 FILLER_53_324 ();
 sg13g2_decap_8 FILLER_53_331 ();
 sg13g2_fill_2 FILLER_53_338 ();
 sg13g2_fill_1 FILLER_53_340 ();
 sg13g2_fill_1 FILLER_53_362 ();
 sg13g2_fill_1 FILLER_53_367 ();
 sg13g2_fill_1 FILLER_53_393 ();
 sg13g2_fill_2 FILLER_53_465 ();
 sg13g2_fill_1 FILLER_53_467 ();
 sg13g2_fill_1 FILLER_53_472 ();
 sg13g2_fill_1 FILLER_53_499 ();
 sg13g2_fill_1 FILLER_53_526 ();
 sg13g2_fill_1 FILLER_53_535 ();
 sg13g2_decap_4 FILLER_53_557 ();
 sg13g2_decap_8 FILLER_53_574 ();
 sg13g2_fill_1 FILLER_53_581 ();
 sg13g2_decap_8 FILLER_53_586 ();
 sg13g2_decap_8 FILLER_53_597 ();
 sg13g2_fill_1 FILLER_53_608 ();
 sg13g2_decap_8 FILLER_53_642 ();
 sg13g2_decap_8 FILLER_53_649 ();
 sg13g2_decap_4 FILLER_53_656 ();
 sg13g2_fill_1 FILLER_53_660 ();
 sg13g2_fill_2 FILLER_53_675 ();
 sg13g2_fill_1 FILLER_53_677 ();
 sg13g2_decap_8 FILLER_53_688 ();
 sg13g2_fill_1 FILLER_53_695 ();
 sg13g2_fill_1 FILLER_53_714 ();
 sg13g2_decap_8 FILLER_53_750 ();
 sg13g2_decap_4 FILLER_53_757 ();
 sg13g2_decap_8 FILLER_53_770 ();
 sg13g2_decap_8 FILLER_53_777 ();
 sg13g2_decap_8 FILLER_53_790 ();
 sg13g2_decap_4 FILLER_53_797 ();
 sg13g2_fill_1 FILLER_53_801 ();
 sg13g2_decap_8 FILLER_53_807 ();
 sg13g2_fill_1 FILLER_53_814 ();
 sg13g2_fill_2 FILLER_53_820 ();
 sg13g2_fill_1 FILLER_53_822 ();
 sg13g2_fill_1 FILLER_53_828 ();
 sg13g2_fill_1 FILLER_53_840 ();
 sg13g2_fill_2 FILLER_53_852 ();
 sg13g2_decap_4 FILLER_53_864 ();
 sg13g2_fill_2 FILLER_53_868 ();
 sg13g2_fill_2 FILLER_53_932 ();
 sg13g2_fill_1 FILLER_53_934 ();
 sg13g2_fill_2 FILLER_53_944 ();
 sg13g2_decap_4 FILLER_53_951 ();
 sg13g2_decap_8 FILLER_53_959 ();
 sg13g2_decap_8 FILLER_53_966 ();
 sg13g2_fill_1 FILLER_53_1002 ();
 sg13g2_decap_4 FILLER_53_1038 ();
 sg13g2_decap_8 FILLER_53_1058 ();
 sg13g2_decap_8 FILLER_53_1065 ();
 sg13g2_fill_2 FILLER_53_1072 ();
 sg13g2_fill_1 FILLER_53_1074 ();
 sg13g2_fill_1 FILLER_53_1079 ();
 sg13g2_fill_1 FILLER_53_1090 ();
 sg13g2_fill_1 FILLER_53_1101 ();
 sg13g2_fill_1 FILLER_53_1110 ();
 sg13g2_decap_4 FILLER_53_1121 ();
 sg13g2_fill_1 FILLER_53_1125 ();
 sg13g2_decap_8 FILLER_53_1136 ();
 sg13g2_fill_2 FILLER_53_1143 ();
 sg13g2_fill_1 FILLER_53_1145 ();
 sg13g2_fill_1 FILLER_53_1150 ();
 sg13g2_fill_2 FILLER_53_1161 ();
 sg13g2_fill_1 FILLER_53_1163 ();
 sg13g2_fill_2 FILLER_53_1186 ();
 sg13g2_decap_8 FILLER_53_1192 ();
 sg13g2_decap_8 FILLER_53_1199 ();
 sg13g2_fill_2 FILLER_53_1206 ();
 sg13g2_fill_1 FILLER_53_1208 ();
 sg13g2_fill_1 FILLER_53_1213 ();
 sg13g2_fill_1 FILLER_53_1240 ();
 sg13g2_fill_1 FILLER_53_1251 ();
 sg13g2_fill_2 FILLER_53_1262 ();
 sg13g2_fill_2 FILLER_53_1324 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_37 ();
 sg13g2_fill_1 FILLER_54_39 ();
 sg13g2_fill_1 FILLER_54_44 ();
 sg13g2_fill_1 FILLER_54_98 ();
 sg13g2_decap_4 FILLER_54_124 ();
 sg13g2_decap_8 FILLER_54_159 ();
 sg13g2_decap_8 FILLER_54_166 ();
 sg13g2_decap_8 FILLER_54_173 ();
 sg13g2_decap_4 FILLER_54_180 ();
 sg13g2_fill_2 FILLER_54_184 ();
 sg13g2_decap_4 FILLER_54_222 ();
 sg13g2_decap_8 FILLER_54_287 ();
 sg13g2_decap_8 FILLER_54_294 ();
 sg13g2_decap_8 FILLER_54_301 ();
 sg13g2_decap_8 FILLER_54_308 ();
 sg13g2_fill_2 FILLER_54_315 ();
 sg13g2_fill_1 FILLER_54_317 ();
 sg13g2_fill_2 FILLER_54_326 ();
 sg13g2_fill_1 FILLER_54_328 ();
 sg13g2_fill_2 FILLER_54_363 ();
 sg13g2_decap_8 FILLER_54_379 ();
 sg13g2_decap_8 FILLER_54_386 ();
 sg13g2_fill_2 FILLER_54_393 ();
 sg13g2_decap_4 FILLER_54_399 ();
 sg13g2_fill_1 FILLER_54_411 ();
 sg13g2_fill_2 FILLER_54_426 ();
 sg13g2_fill_1 FILLER_54_428 ();
 sg13g2_decap_4 FILLER_54_446 ();
 sg13g2_fill_1 FILLER_54_450 ();
 sg13g2_decap_4 FILLER_54_455 ();
 sg13g2_fill_1 FILLER_54_473 ();
 sg13g2_fill_1 FILLER_54_478 ();
 sg13g2_fill_1 FILLER_54_508 ();
 sg13g2_fill_1 FILLER_54_535 ();
 sg13g2_decap_8 FILLER_54_575 ();
 sg13g2_decap_4 FILLER_54_582 ();
 sg13g2_decap_8 FILLER_54_590 ();
 sg13g2_decap_8 FILLER_54_597 ();
 sg13g2_decap_4 FILLER_54_604 ();
 sg13g2_decap_8 FILLER_54_618 ();
 sg13g2_decap_8 FILLER_54_625 ();
 sg13g2_fill_2 FILLER_54_632 ();
 sg13g2_fill_1 FILLER_54_645 ();
 sg13g2_fill_2 FILLER_54_656 ();
 sg13g2_fill_1 FILLER_54_658 ();
 sg13g2_fill_2 FILLER_54_676 ();
 sg13g2_fill_1 FILLER_54_678 ();
 sg13g2_fill_2 FILLER_54_689 ();
 sg13g2_fill_1 FILLER_54_691 ();
 sg13g2_decap_4 FILLER_54_700 ();
 sg13g2_fill_1 FILLER_54_704 ();
 sg13g2_decap_8 FILLER_54_713 ();
 sg13g2_fill_2 FILLER_54_741 ();
 sg13g2_decap_4 FILLER_54_756 ();
 sg13g2_fill_1 FILLER_54_791 ();
 sg13g2_fill_1 FILLER_54_796 ();
 sg13g2_fill_1 FILLER_54_802 ();
 sg13g2_fill_2 FILLER_54_808 ();
 sg13g2_fill_1 FILLER_54_810 ();
 sg13g2_fill_1 FILLER_54_816 ();
 sg13g2_fill_1 FILLER_54_822 ();
 sg13g2_fill_1 FILLER_54_828 ();
 sg13g2_fill_2 FILLER_54_835 ();
 sg13g2_fill_1 FILLER_54_842 ();
 sg13g2_decap_8 FILLER_54_873 ();
 sg13g2_fill_2 FILLER_54_880 ();
 sg13g2_fill_1 FILLER_54_882 ();
 sg13g2_fill_2 FILLER_54_943 ();
 sg13g2_decap_4 FILLER_54_971 ();
 sg13g2_fill_2 FILLER_54_998 ();
 sg13g2_fill_2 FILLER_54_1004 ();
 sg13g2_decap_8 FILLER_54_1036 ();
 sg13g2_fill_2 FILLER_54_1079 ();
 sg13g2_fill_1 FILLER_54_1081 ();
 sg13g2_decap_8 FILLER_54_1086 ();
 sg13g2_decap_8 FILLER_54_1093 ();
 sg13g2_fill_1 FILLER_54_1100 ();
 sg13g2_decap_8 FILLER_54_1105 ();
 sg13g2_decap_8 FILLER_54_1112 ();
 sg13g2_fill_1 FILLER_54_1123 ();
 sg13g2_decap_8 FILLER_54_1134 ();
 sg13g2_decap_4 FILLER_54_1141 ();
 sg13g2_fill_2 FILLER_54_1145 ();
 sg13g2_decap_8 FILLER_54_1235 ();
 sg13g2_fill_2 FILLER_54_1242 ();
 sg13g2_fill_1 FILLER_54_1244 ();
 sg13g2_decap_8 FILLER_54_1249 ();
 sg13g2_decap_4 FILLER_54_1256 ();
 sg13g2_fill_1 FILLER_54_1260 ();
 sg13g2_decap_8 FILLER_54_1311 ();
 sg13g2_decap_8 FILLER_54_1318 ();
 sg13g2_fill_1 FILLER_54_1325 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_fill_2 FILLER_55_51 ();
 sg13g2_fill_2 FILLER_55_174 ();
 sg13g2_decap_8 FILLER_55_226 ();
 sg13g2_decap_8 FILLER_55_233 ();
 sg13g2_fill_1 FILLER_55_240 ();
 sg13g2_decap_8 FILLER_55_277 ();
 sg13g2_decap_8 FILLER_55_284 ();
 sg13g2_fill_2 FILLER_55_291 ();
 sg13g2_decap_4 FILLER_55_319 ();
 sg13g2_fill_2 FILLER_55_333 ();
 sg13g2_fill_1 FILLER_55_335 ();
 sg13g2_fill_1 FILLER_55_370 ();
 sg13g2_decap_4 FILLER_55_375 ();
 sg13g2_decap_4 FILLER_55_384 ();
 sg13g2_decap_8 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_decap_4 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_410 ();
 sg13g2_fill_2 FILLER_55_415 ();
 sg13g2_fill_1 FILLER_55_417 ();
 sg13g2_fill_2 FILLER_55_422 ();
 sg13g2_decap_4 FILLER_55_428 ();
 sg13g2_fill_1 FILLER_55_436 ();
 sg13g2_fill_2 FILLER_55_445 ();
 sg13g2_fill_2 FILLER_55_461 ();
 sg13g2_fill_1 FILLER_55_463 ();
 sg13g2_fill_2 FILLER_55_469 ();
 sg13g2_fill_1 FILLER_55_471 ();
 sg13g2_decap_4 FILLER_55_476 ();
 sg13g2_fill_1 FILLER_55_484 ();
 sg13g2_fill_1 FILLER_55_489 ();
 sg13g2_fill_2 FILLER_55_543 ();
 sg13g2_decap_8 FILLER_55_549 ();
 sg13g2_fill_2 FILLER_55_556 ();
 sg13g2_fill_1 FILLER_55_573 ();
 sg13g2_fill_2 FILLER_55_584 ();
 sg13g2_decap_8 FILLER_55_600 ();
 sg13g2_fill_2 FILLER_55_607 ();
 sg13g2_fill_2 FILLER_55_613 ();
 sg13g2_fill_2 FILLER_55_625 ();
 sg13g2_fill_1 FILLER_55_649 ();
 sg13g2_fill_1 FILLER_55_655 ();
 sg13g2_fill_1 FILLER_55_671 ();
 sg13g2_fill_1 FILLER_55_677 ();
 sg13g2_fill_1 FILLER_55_690 ();
 sg13g2_decap_8 FILLER_55_703 ();
 sg13g2_decap_8 FILLER_55_710 ();
 sg13g2_fill_1 FILLER_55_717 ();
 sg13g2_decap_4 FILLER_55_742 ();
 sg13g2_fill_2 FILLER_55_746 ();
 sg13g2_decap_4 FILLER_55_763 ();
 sg13g2_fill_1 FILLER_55_767 ();
 sg13g2_fill_1 FILLER_55_773 ();
 sg13g2_fill_1 FILLER_55_778 ();
 sg13g2_fill_1 FILLER_55_795 ();
 sg13g2_fill_1 FILLER_55_800 ();
 sg13g2_fill_1 FILLER_55_806 ();
 sg13g2_fill_1 FILLER_55_816 ();
 sg13g2_fill_2 FILLER_55_822 ();
 sg13g2_fill_1 FILLER_55_824 ();
 sg13g2_fill_1 FILLER_55_839 ();
 sg13g2_fill_1 FILLER_55_850 ();
 sg13g2_fill_1 FILLER_55_856 ();
 sg13g2_fill_1 FILLER_55_865 ();
 sg13g2_fill_1 FILLER_55_870 ();
 sg13g2_decap_8 FILLER_55_879 ();
 sg13g2_decap_8 FILLER_55_886 ();
 sg13g2_fill_1 FILLER_55_893 ();
 sg13g2_decap_8 FILLER_55_898 ();
 sg13g2_decap_4 FILLER_55_905 ();
 sg13g2_decap_4 FILLER_55_918 ();
 sg13g2_fill_1 FILLER_55_922 ();
 sg13g2_fill_1 FILLER_55_927 ();
 sg13g2_decap_8 FILLER_55_932 ();
 sg13g2_decap_8 FILLER_55_939 ();
 sg13g2_decap_4 FILLER_55_946 ();
 sg13g2_fill_2 FILLER_55_950 ();
 sg13g2_decap_4 FILLER_55_956 ();
 sg13g2_fill_1 FILLER_55_960 ();
 sg13g2_decap_8 FILLER_55_991 ();
 sg13g2_decap_8 FILLER_55_998 ();
 sg13g2_decap_8 FILLER_55_1005 ();
 sg13g2_decap_8 FILLER_55_1020 ();
 sg13g2_decap_8 FILLER_55_1027 ();
 sg13g2_decap_8 FILLER_55_1034 ();
 sg13g2_decap_8 FILLER_55_1041 ();
 sg13g2_decap_4 FILLER_55_1048 ();
 sg13g2_fill_2 FILLER_55_1062 ();
 sg13g2_fill_1 FILLER_55_1064 ();
 sg13g2_decap_4 FILLER_55_1075 ();
 sg13g2_fill_1 FILLER_55_1079 ();
 sg13g2_decap_8 FILLER_55_1084 ();
 sg13g2_decap_8 FILLER_55_1091 ();
 sg13g2_decap_8 FILLER_55_1098 ();
 sg13g2_decap_4 FILLER_55_1105 ();
 sg13g2_fill_2 FILLER_55_1109 ();
 sg13g2_decap_8 FILLER_55_1141 ();
 sg13g2_decap_4 FILLER_55_1148 ();
 sg13g2_fill_1 FILLER_55_1152 ();
 sg13g2_decap_8 FILLER_55_1157 ();
 sg13g2_fill_1 FILLER_55_1164 ();
 sg13g2_fill_2 FILLER_55_1175 ();
 sg13g2_fill_1 FILLER_55_1177 ();
 sg13g2_decap_8 FILLER_55_1186 ();
 sg13g2_decap_8 FILLER_55_1229 ();
 sg13g2_fill_1 FILLER_55_1246 ();
 sg13g2_fill_2 FILLER_55_1277 ();
 sg13g2_fill_1 FILLER_55_1279 ();
 sg13g2_fill_1 FILLER_55_1284 ();
 sg13g2_decap_4 FILLER_55_1295 ();
 sg13g2_decap_8 FILLER_55_1313 ();
 sg13g2_decap_4 FILLER_55_1320 ();
 sg13g2_fill_2 FILLER_55_1324 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_8 ();
 sg13g2_decap_8 FILLER_56_100 ();
 sg13g2_decap_8 FILLER_56_128 ();
 sg13g2_fill_2 FILLER_56_139 ();
 sg13g2_fill_1 FILLER_56_151 ();
 sg13g2_fill_2 FILLER_56_162 ();
 sg13g2_fill_2 FILLER_56_190 ();
 sg13g2_fill_1 FILLER_56_192 ();
 sg13g2_decap_8 FILLER_56_214 ();
 sg13g2_decap_8 FILLER_56_221 ();
 sg13g2_decap_8 FILLER_56_228 ();
 sg13g2_fill_1 FILLER_56_235 ();
 sg13g2_fill_2 FILLER_56_250 ();
 sg13g2_fill_2 FILLER_56_278 ();
 sg13g2_fill_1 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_323 ();
 sg13g2_fill_2 FILLER_56_330 ();
 sg13g2_fill_2 FILLER_56_344 ();
 sg13g2_fill_1 FILLER_56_346 ();
 sg13g2_fill_1 FILLER_56_377 ();
 sg13g2_decap_4 FILLER_56_482 ();
 sg13g2_fill_2 FILLER_56_486 ();
 sg13g2_fill_1 FILLER_56_496 ();
 sg13g2_fill_2 FILLER_56_551 ();
 sg13g2_fill_1 FILLER_56_553 ();
 sg13g2_fill_2 FILLER_56_567 ();
 sg13g2_fill_1 FILLER_56_569 ();
 sg13g2_decap_8 FILLER_56_574 ();
 sg13g2_fill_2 FILLER_56_581 ();
 sg13g2_decap_4 FILLER_56_591 ();
 sg13g2_fill_1 FILLER_56_599 ();
 sg13g2_decap_8 FILLER_56_604 ();
 sg13g2_decap_8 FILLER_56_611 ();
 sg13g2_decap_4 FILLER_56_618 ();
 sg13g2_fill_1 FILLER_56_639 ();
 sg13g2_fill_1 FILLER_56_645 ();
 sg13g2_fill_2 FILLER_56_653 ();
 sg13g2_fill_2 FILLER_56_663 ();
 sg13g2_decap_4 FILLER_56_702 ();
 sg13g2_fill_1 FILLER_56_706 ();
 sg13g2_fill_2 FILLER_56_724 ();
 sg13g2_fill_1 FILLER_56_726 ();
 sg13g2_decap_4 FILLER_56_737 ();
 sg13g2_decap_8 FILLER_56_754 ();
 sg13g2_fill_2 FILLER_56_761 ();
 sg13g2_decap_4 FILLER_56_767 ();
 sg13g2_fill_1 FILLER_56_776 ();
 sg13g2_fill_1 FILLER_56_782 ();
 sg13g2_decap_4 FILLER_56_787 ();
 sg13g2_fill_2 FILLER_56_797 ();
 sg13g2_fill_1 FILLER_56_799 ();
 sg13g2_fill_2 FILLER_56_806 ();
 sg13g2_fill_2 FILLER_56_813 ();
 sg13g2_fill_1 FILLER_56_815 ();
 sg13g2_decap_4 FILLER_56_825 ();
 sg13g2_fill_1 FILLER_56_829 ();
 sg13g2_fill_2 FILLER_56_835 ();
 sg13g2_fill_2 FILLER_56_843 ();
 sg13g2_fill_1 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_866 ();
 sg13g2_decap_4 FILLER_56_871 ();
 sg13g2_fill_1 FILLER_56_875 ();
 sg13g2_decap_8 FILLER_56_890 ();
 sg13g2_decap_8 FILLER_56_897 ();
 sg13g2_decap_8 FILLER_56_904 ();
 sg13g2_decap_4 FILLER_56_911 ();
 sg13g2_fill_1 FILLER_56_915 ();
 sg13g2_decap_8 FILLER_56_946 ();
 sg13g2_decap_8 FILLER_56_953 ();
 sg13g2_decap_8 FILLER_56_960 ();
 sg13g2_decap_8 FILLER_56_971 ();
 sg13g2_decap_8 FILLER_56_978 ();
 sg13g2_fill_2 FILLER_56_993 ();
 sg13g2_decap_8 FILLER_56_1021 ();
 sg13g2_decap_8 FILLER_56_1028 ();
 sg13g2_decap_4 FILLER_56_1035 ();
 sg13g2_fill_2 FILLER_56_1039 ();
 sg13g2_decap_4 FILLER_56_1045 ();
 sg13g2_fill_1 FILLER_56_1049 ();
 sg13g2_fill_2 FILLER_56_1086 ();
 sg13g2_fill_1 FILLER_56_1088 ();
 sg13g2_fill_1 FILLER_56_1099 ();
 sg13g2_decap_8 FILLER_56_1156 ();
 sg13g2_decap_8 FILLER_56_1163 ();
 sg13g2_fill_2 FILLER_56_1170 ();
 sg13g2_fill_2 FILLER_56_1198 ();
 sg13g2_fill_1 FILLER_56_1200 ();
 sg13g2_fill_2 FILLER_56_1205 ();
 sg13g2_decap_4 FILLER_56_1211 ();
 sg13g2_decap_4 FILLER_56_1225 ();
 sg13g2_fill_2 FILLER_56_1229 ();
 sg13g2_decap_8 FILLER_56_1265 ();
 sg13g2_decap_8 FILLER_56_1272 ();
 sg13g2_fill_1 FILLER_56_1279 ();
 sg13g2_decap_8 FILLER_56_1310 ();
 sg13g2_decap_8 FILLER_56_1317 ();
 sg13g2_fill_2 FILLER_56_1324 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_51 ();
 sg13g2_fill_1 FILLER_57_62 ();
 sg13g2_decap_8 FILLER_57_71 ();
 sg13g2_fill_2 FILLER_57_78 ();
 sg13g2_fill_1 FILLER_57_80 ();
 sg13g2_decap_4 FILLER_57_102 ();
 sg13g2_decap_8 FILLER_57_127 ();
 sg13g2_decap_8 FILLER_57_185 ();
 sg13g2_fill_1 FILLER_57_192 ();
 sg13g2_fill_2 FILLER_57_214 ();
 sg13g2_fill_1 FILLER_57_216 ();
 sg13g2_fill_2 FILLER_57_242 ();
 sg13g2_fill_1 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_307 ();
 sg13g2_fill_2 FILLER_57_314 ();
 sg13g2_fill_1 FILLER_57_316 ();
 sg13g2_fill_1 FILLER_57_361 ();
 sg13g2_decap_4 FILLER_57_366 ();
 sg13g2_fill_2 FILLER_57_370 ();
 sg13g2_decap_8 FILLER_57_376 ();
 sg13g2_decap_8 FILLER_57_383 ();
 sg13g2_decap_8 FILLER_57_390 ();
 sg13g2_fill_2 FILLER_57_397 ();
 sg13g2_fill_2 FILLER_57_404 ();
 sg13g2_fill_1 FILLER_57_406 ();
 sg13g2_decap_8 FILLER_57_464 ();
 sg13g2_fill_2 FILLER_57_471 ();
 sg13g2_fill_1 FILLER_57_473 ();
 sg13g2_fill_2 FILLER_57_505 ();
 sg13g2_decap_4 FILLER_57_523 ();
 sg13g2_fill_2 FILLER_57_553 ();
 sg13g2_fill_2 FILLER_57_564 ();
 sg13g2_fill_1 FILLER_57_566 ();
 sg13g2_fill_1 FILLER_57_576 ();
 sg13g2_fill_1 FILLER_57_582 ();
 sg13g2_fill_1 FILLER_57_588 ();
 sg13g2_fill_2 FILLER_57_594 ();
 sg13g2_decap_8 FILLER_57_600 ();
 sg13g2_decap_8 FILLER_57_607 ();
 sg13g2_decap_8 FILLER_57_614 ();
 sg13g2_fill_2 FILLER_57_621 ();
 sg13g2_fill_1 FILLER_57_623 ();
 sg13g2_fill_1 FILLER_57_646 ();
 sg13g2_fill_2 FILLER_57_652 ();
 sg13g2_fill_1 FILLER_57_654 ();
 sg13g2_fill_1 FILLER_57_680 ();
 sg13g2_fill_1 FILLER_57_686 ();
 sg13g2_fill_1 FILLER_57_703 ();
 sg13g2_decap_4 FILLER_57_714 ();
 sg13g2_decap_8 FILLER_57_723 ();
 sg13g2_decap_8 FILLER_57_730 ();
 sg13g2_decap_8 FILLER_57_737 ();
 sg13g2_decap_4 FILLER_57_744 ();
 sg13g2_fill_2 FILLER_57_748 ();
 sg13g2_decap_8 FILLER_57_755 ();
 sg13g2_decap_4 FILLER_57_762 ();
 sg13g2_fill_2 FILLER_57_770 ();
 sg13g2_fill_1 FILLER_57_791 ();
 sg13g2_fill_2 FILLER_57_804 ();
 sg13g2_fill_2 FILLER_57_812 ();
 sg13g2_fill_1 FILLER_57_814 ();
 sg13g2_fill_1 FILLER_57_841 ();
 sg13g2_fill_2 FILLER_57_845 ();
 sg13g2_fill_1 FILLER_57_847 ();
 sg13g2_decap_4 FILLER_57_852 ();
 sg13g2_fill_1 FILLER_57_866 ();
 sg13g2_fill_2 FILLER_57_886 ();
 sg13g2_fill_1 FILLER_57_898 ();
 sg13g2_decap_8 FILLER_57_925 ();
 sg13g2_decap_8 FILLER_57_932 ();
 sg13g2_decap_8 FILLER_57_939 ();
 sg13g2_decap_4 FILLER_57_946 ();
 sg13g2_fill_1 FILLER_57_950 ();
 sg13g2_decap_8 FILLER_57_954 ();
 sg13g2_decap_4 FILLER_57_961 ();
 sg13g2_fill_2 FILLER_57_965 ();
 sg13g2_decap_8 FILLER_57_977 ();
 sg13g2_decap_8 FILLER_57_1018 ();
 sg13g2_decap_8 FILLER_57_1025 ();
 sg13g2_fill_2 FILLER_57_1032 ();
 sg13g2_decap_8 FILLER_57_1146 ();
 sg13g2_decap_8 FILLER_57_1153 ();
 sg13g2_decap_4 FILLER_57_1160 ();
 sg13g2_decap_8 FILLER_57_1194 ();
 sg13g2_decap_8 FILLER_57_1201 ();
 sg13g2_decap_8 FILLER_57_1208 ();
 sg13g2_decap_8 FILLER_57_1215 ();
 sg13g2_decap_4 FILLER_57_1222 ();
 sg13g2_fill_2 FILLER_57_1236 ();
 sg13g2_decap_8 FILLER_57_1312 ();
 sg13g2_decap_8 FILLER_57_1319 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_9 ();
 sg13g2_decap_4 FILLER_58_24 ();
 sg13g2_fill_2 FILLER_58_32 ();
 sg13g2_fill_2 FILLER_58_38 ();
 sg13g2_decap_8 FILLER_58_44 ();
 sg13g2_decap_4 FILLER_58_51 ();
 sg13g2_decap_4 FILLER_58_68 ();
 sg13g2_fill_2 FILLER_58_72 ();
 sg13g2_decap_8 FILLER_58_82 ();
 sg13g2_decap_8 FILLER_58_89 ();
 sg13g2_decap_8 FILLER_58_96 ();
 sg13g2_fill_2 FILLER_58_103 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_fill_2 FILLER_58_133 ();
 sg13g2_fill_1 FILLER_58_135 ();
 sg13g2_decap_8 FILLER_58_150 ();
 sg13g2_fill_2 FILLER_58_161 ();
 sg13g2_decap_4 FILLER_58_184 ();
 sg13g2_fill_2 FILLER_58_188 ();
 sg13g2_decap_8 FILLER_58_216 ();
 sg13g2_fill_1 FILLER_58_223 ();
 sg13g2_decap_8 FILLER_58_232 ();
 sg13g2_decap_4 FILLER_58_239 ();
 sg13g2_fill_1 FILLER_58_243 ();
 sg13g2_fill_2 FILLER_58_257 ();
 sg13g2_fill_2 FILLER_58_289 ();
 sg13g2_fill_2 FILLER_58_295 ();
 sg13g2_decap_8 FILLER_58_318 ();
 sg13g2_decap_8 FILLER_58_325 ();
 sg13g2_fill_1 FILLER_58_346 ();
 sg13g2_fill_2 FILLER_58_351 ();
 sg13g2_fill_1 FILLER_58_353 ();
 sg13g2_decap_8 FILLER_58_358 ();
 sg13g2_decap_8 FILLER_58_365 ();
 sg13g2_decap_8 FILLER_58_372 ();
 sg13g2_fill_2 FILLER_58_379 ();
 sg13g2_fill_1 FILLER_58_381 ();
 sg13g2_decap_8 FILLER_58_411 ();
 sg13g2_decap_8 FILLER_58_474 ();
 sg13g2_fill_2 FILLER_58_481 ();
 sg13g2_decap_4 FILLER_58_491 ();
 sg13g2_decap_8 FILLER_58_557 ();
 sg13g2_decap_8 FILLER_58_564 ();
 sg13g2_decap_8 FILLER_58_571 ();
 sg13g2_fill_2 FILLER_58_587 ();
 sg13g2_fill_1 FILLER_58_589 ();
 sg13g2_decap_8 FILLER_58_599 ();
 sg13g2_decap_8 FILLER_58_606 ();
 sg13g2_decap_4 FILLER_58_652 ();
 sg13g2_fill_2 FILLER_58_656 ();
 sg13g2_fill_1 FILLER_58_664 ();
 sg13g2_fill_1 FILLER_58_683 ();
 sg13g2_fill_2 FILLER_58_709 ();
 sg13g2_fill_1 FILLER_58_711 ();
 sg13g2_fill_2 FILLER_58_720 ();
 sg13g2_fill_1 FILLER_58_722 ();
 sg13g2_fill_1 FILLER_58_727 ();
 sg13g2_decap_8 FILLER_58_737 ();
 sg13g2_decap_8 FILLER_58_744 ();
 sg13g2_decap_8 FILLER_58_751 ();
 sg13g2_decap_8 FILLER_58_758 ();
 sg13g2_decap_8 FILLER_58_765 ();
 sg13g2_decap_8 FILLER_58_772 ();
 sg13g2_fill_2 FILLER_58_779 ();
 sg13g2_fill_1 FILLER_58_781 ();
 sg13g2_decap_4 FILLER_58_791 ();
 sg13g2_fill_1 FILLER_58_795 ();
 sg13g2_fill_1 FILLER_58_800 ();
 sg13g2_fill_2 FILLER_58_827 ();
 sg13g2_decap_8 FILLER_58_859 ();
 sg13g2_fill_2 FILLER_58_866 ();
 sg13g2_fill_2 FILLER_58_879 ();
 sg13g2_fill_1 FILLER_58_881 ();
 sg13g2_fill_2 FILLER_58_887 ();
 sg13g2_fill_1 FILLER_58_897 ();
 sg13g2_fill_1 FILLER_58_910 ();
 sg13g2_fill_1 FILLER_58_916 ();
 sg13g2_decap_8 FILLER_58_921 ();
 sg13g2_fill_1 FILLER_58_933 ();
 sg13g2_fill_1 FILLER_58_939 ();
 sg13g2_fill_1 FILLER_58_950 ();
 sg13g2_fill_2 FILLER_58_990 ();
 sg13g2_fill_2 FILLER_58_996 ();
 sg13g2_decap_8 FILLER_58_1006 ();
 sg13g2_decap_8 FILLER_58_1013 ();
 sg13g2_decap_8 FILLER_58_1020 ();
 sg13g2_decap_8 FILLER_58_1027 ();
 sg13g2_decap_8 FILLER_58_1034 ();
 sg13g2_fill_2 FILLER_58_1041 ();
 sg13g2_decap_8 FILLER_58_1047 ();
 sg13g2_fill_1 FILLER_58_1054 ();
 sg13g2_decap_4 FILLER_58_1065 ();
 sg13g2_fill_1 FILLER_58_1069 ();
 sg13g2_fill_1 FILLER_58_1118 ();
 sg13g2_decap_8 FILLER_58_1139 ();
 sg13g2_decap_4 FILLER_58_1146 ();
 sg13g2_fill_1 FILLER_58_1150 ();
 sg13g2_decap_8 FILLER_58_1161 ();
 sg13g2_fill_1 FILLER_58_1168 ();
 sg13g2_decap_4 FILLER_58_1179 ();
 sg13g2_decap_8 FILLER_58_1187 ();
 sg13g2_decap_4 FILLER_58_1194 ();
 sg13g2_fill_2 FILLER_58_1210 ();
 sg13g2_fill_2 FILLER_58_1238 ();
 sg13g2_fill_1 FILLER_58_1240 ();
 sg13g2_fill_2 FILLER_58_1267 ();
 sg13g2_fill_1 FILLER_58_1269 ();
 sg13g2_fill_2 FILLER_58_1296 ();
 sg13g2_fill_1 FILLER_58_1298 ();
 sg13g2_fill_1 FILLER_58_1325 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_fill_2 FILLER_59_14 ();
 sg13g2_fill_1 FILLER_59_16 ();
 sg13g2_fill_1 FILLER_59_31 ();
 sg13g2_fill_2 FILLER_59_53 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_fill_2 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_128 ();
 sg13g2_decap_8 FILLER_59_135 ();
 sg13g2_fill_2 FILLER_59_142 ();
 sg13g2_fill_1 FILLER_59_144 ();
 sg13g2_fill_2 FILLER_59_171 ();
 sg13g2_fill_1 FILLER_59_173 ();
 sg13g2_decap_8 FILLER_59_179 ();
 sg13g2_fill_1 FILLER_59_186 ();
 sg13g2_decap_4 FILLER_59_205 ();
 sg13g2_fill_1 FILLER_59_214 ();
 sg13g2_decap_4 FILLER_59_219 ();
 sg13g2_decap_8 FILLER_59_227 ();
 sg13g2_decap_8 FILLER_59_234 ();
 sg13g2_decap_8 FILLER_59_241 ();
 sg13g2_decap_8 FILLER_59_248 ();
 sg13g2_decap_4 FILLER_59_255 ();
 sg13g2_fill_2 FILLER_59_259 ();
 sg13g2_fill_2 FILLER_59_291 ();
 sg13g2_decap_8 FILLER_59_314 ();
 sg13g2_decap_8 FILLER_59_321 ();
 sg13g2_fill_2 FILLER_59_328 ();
 sg13g2_decap_4 FILLER_59_344 ();
 sg13g2_fill_2 FILLER_59_348 ();
 sg13g2_fill_2 FILLER_59_354 ();
 sg13g2_decap_8 FILLER_59_400 ();
 sg13g2_decap_4 FILLER_59_407 ();
 sg13g2_fill_2 FILLER_59_422 ();
 sg13g2_fill_1 FILLER_59_424 ();
 sg13g2_decap_8 FILLER_59_438 ();
 sg13g2_decap_8 FILLER_59_445 ();
 sg13g2_decap_4 FILLER_59_452 ();
 sg13g2_fill_1 FILLER_59_456 ();
 sg13g2_decap_8 FILLER_59_461 ();
 sg13g2_decap_8 FILLER_59_468 ();
 sg13g2_decap_8 FILLER_59_475 ();
 sg13g2_decap_8 FILLER_59_482 ();
 sg13g2_decap_8 FILLER_59_489 ();
 sg13g2_decap_4 FILLER_59_496 ();
 sg13g2_decap_8 FILLER_59_514 ();
 sg13g2_fill_1 FILLER_59_521 ();
 sg13g2_fill_2 FILLER_59_527 ();
 sg13g2_fill_1 FILLER_59_529 ();
 sg13g2_fill_1 FILLER_59_534 ();
 sg13g2_fill_2 FILLER_59_539 ();
 sg13g2_fill_1 FILLER_59_541 ();
 sg13g2_decap_8 FILLER_59_546 ();
 sg13g2_fill_2 FILLER_59_553 ();
 sg13g2_fill_1 FILLER_59_555 ();
 sg13g2_decap_8 FILLER_59_561 ();
 sg13g2_decap_4 FILLER_59_568 ();
 sg13g2_fill_1 FILLER_59_577 ();
 sg13g2_fill_2 FILLER_59_586 ();
 sg13g2_decap_8 FILLER_59_593 ();
 sg13g2_decap_8 FILLER_59_600 ();
 sg13g2_decap_8 FILLER_59_607 ();
 sg13g2_fill_1 FILLER_59_624 ();
 sg13g2_fill_2 FILLER_59_647 ();
 sg13g2_fill_1 FILLER_59_649 ();
 sg13g2_decap_8 FILLER_59_665 ();
 sg13g2_fill_1 FILLER_59_672 ();
 sg13g2_decap_4 FILLER_59_678 ();
 sg13g2_fill_1 FILLER_59_682 ();
 sg13g2_fill_2 FILLER_59_701 ();
 sg13g2_fill_1 FILLER_59_708 ();
 sg13g2_fill_2 FILLER_59_727 ();
 sg13g2_fill_1 FILLER_59_729 ();
 sg13g2_fill_1 FILLER_59_737 ();
 sg13g2_decap_8 FILLER_59_742 ();
 sg13g2_decap_8 FILLER_59_749 ();
 sg13g2_decap_4 FILLER_59_756 ();
 sg13g2_fill_1 FILLER_59_760 ();
 sg13g2_fill_1 FILLER_59_787 ();
 sg13g2_fill_1 FILLER_59_792 ();
 sg13g2_fill_1 FILLER_59_798 ();
 sg13g2_fill_2 FILLER_59_815 ();
 sg13g2_fill_2 FILLER_59_826 ();
 sg13g2_decap_8 FILLER_59_844 ();
 sg13g2_decap_8 FILLER_59_851 ();
 sg13g2_decap_8 FILLER_59_858 ();
 sg13g2_fill_2 FILLER_59_901 ();
 sg13g2_fill_2 FILLER_59_911 ();
 sg13g2_fill_1 FILLER_59_918 ();
 sg13g2_fill_1 FILLER_59_973 ();
 sg13g2_fill_2 FILLER_59_993 ();
 sg13g2_decap_8 FILLER_59_1026 ();
 sg13g2_decap_4 FILLER_59_1033 ();
 sg13g2_decap_4 FILLER_59_1063 ();
 sg13g2_decap_8 FILLER_59_1093 ();
 sg13g2_decap_8 FILLER_59_1116 ();
 sg13g2_decap_4 FILLER_59_1123 ();
 sg13g2_fill_1 FILLER_59_1127 ();
 sg13g2_fill_2 FILLER_59_1132 ();
 sg13g2_fill_1 FILLER_59_1134 ();
 sg13g2_fill_1 FILLER_59_1165 ();
 sg13g2_fill_2 FILLER_59_1236 ();
 sg13g2_fill_1 FILLER_59_1238 ();
 sg13g2_fill_2 FILLER_59_1253 ();
 sg13g2_fill_1 FILLER_59_1255 ();
 sg13g2_decap_8 FILLER_59_1260 ();
 sg13g2_fill_1 FILLER_59_1267 ();
 sg13g2_fill_2 FILLER_59_1284 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_7 ();
 sg13g2_fill_2 FILLER_60_34 ();
 sg13g2_fill_1 FILLER_60_36 ();
 sg13g2_fill_2 FILLER_60_63 ();
 sg13g2_decap_4 FILLER_60_138 ();
 sg13g2_fill_1 FILLER_60_142 ();
 sg13g2_decap_4 FILLER_60_147 ();
 sg13g2_fill_2 FILLER_60_151 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_4 FILLER_60_238 ();
 sg13g2_fill_2 FILLER_60_242 ();
 sg13g2_decap_4 FILLER_60_262 ();
 sg13g2_fill_1 FILLER_60_266 ();
 sg13g2_decap_4 FILLER_60_271 ();
 sg13g2_fill_2 FILLER_60_275 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_60_329 ();
 sg13g2_decap_4 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_60_385 ();
 sg13g2_fill_2 FILLER_60_412 ();
 sg13g2_decap_8 FILLER_60_435 ();
 sg13g2_decap_8 FILLER_60_442 ();
 sg13g2_decap_8 FILLER_60_457 ();
 sg13g2_decap_8 FILLER_60_464 ();
 sg13g2_decap_4 FILLER_60_471 ();
 sg13g2_fill_2 FILLER_60_475 ();
 sg13g2_decap_8 FILLER_60_498 ();
 sg13g2_decap_8 FILLER_60_505 ();
 sg13g2_decap_8 FILLER_60_512 ();
 sg13g2_decap_8 FILLER_60_519 ();
 sg13g2_decap_8 FILLER_60_526 ();
 sg13g2_decap_8 FILLER_60_533 ();
 sg13g2_decap_8 FILLER_60_540 ();
 sg13g2_decap_4 FILLER_60_547 ();
 sg13g2_fill_2 FILLER_60_551 ();
 sg13g2_fill_2 FILLER_60_577 ();
 sg13g2_fill_1 FILLER_60_579 ();
 sg13g2_fill_1 FILLER_60_600 ();
 sg13g2_decap_8 FILLER_60_605 ();
 sg13g2_fill_2 FILLER_60_635 ();
 sg13g2_decap_8 FILLER_60_656 ();
 sg13g2_fill_1 FILLER_60_663 ();
 sg13g2_decap_4 FILLER_60_668 ();
 sg13g2_fill_2 FILLER_60_715 ();
 sg13g2_fill_2 FILLER_60_726 ();
 sg13g2_fill_1 FILLER_60_739 ();
 sg13g2_decap_8 FILLER_60_747 ();
 sg13g2_decap_4 FILLER_60_754 ();
 sg13g2_fill_2 FILLER_60_758 ();
 sg13g2_fill_2 FILLER_60_799 ();
 sg13g2_decap_8 FILLER_60_805 ();
 sg13g2_decap_4 FILLER_60_812 ();
 sg13g2_fill_1 FILLER_60_816 ();
 sg13g2_fill_1 FILLER_60_829 ();
 sg13g2_decap_8 FILLER_60_834 ();
 sg13g2_decap_8 FILLER_60_841 ();
 sg13g2_decap_4 FILLER_60_848 ();
 sg13g2_fill_2 FILLER_60_883 ();
 sg13g2_decap_4 FILLER_60_922 ();
 sg13g2_fill_1 FILLER_60_940 ();
 sg13g2_fill_1 FILLER_60_975 ();
 sg13g2_fill_1 FILLER_60_984 ();
 sg13g2_fill_2 FILLER_60_1004 ();
 sg13g2_fill_1 FILLER_60_1006 ();
 sg13g2_fill_2 FILLER_60_1011 ();
 sg13g2_decap_8 FILLER_60_1049 ();
 sg13g2_decap_8 FILLER_60_1056 ();
 sg13g2_decap_8 FILLER_60_1063 ();
 sg13g2_decap_4 FILLER_60_1070 ();
 sg13g2_decap_8 FILLER_60_1078 ();
 sg13g2_fill_2 FILLER_60_1095 ();
 sg13g2_fill_1 FILLER_60_1097 ();
 sg13g2_decap_8 FILLER_60_1102 ();
 sg13g2_decap_8 FILLER_60_1109 ();
 sg13g2_fill_2 FILLER_60_1116 ();
 sg13g2_fill_1 FILLER_60_1118 ();
 sg13g2_decap_4 FILLER_60_1161 ();
 sg13g2_fill_2 FILLER_60_1165 ();
 sg13g2_decap_8 FILLER_60_1203 ();
 sg13g2_fill_1 FILLER_60_1210 ();
 sg13g2_fill_2 FILLER_60_1215 ();
 sg13g2_fill_2 FILLER_60_1237 ();
 sg13g2_decap_8 FILLER_60_1249 ();
 sg13g2_decap_8 FILLER_60_1256 ();
 sg13g2_fill_2 FILLER_60_1263 ();
 sg13g2_decap_8 FILLER_60_1269 ();
 sg13g2_decap_4 FILLER_60_1289 ();
 sg13g2_decap_8 FILLER_60_1317 ();
 sg13g2_fill_2 FILLER_60_1324 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_27 ();
 sg13g2_fill_1 FILLER_61_48 ();
 sg13g2_decap_8 FILLER_61_116 ();
 sg13g2_decap_8 FILLER_61_123 ();
 sg13g2_decap_8 FILLER_61_130 ();
 sg13g2_decap_8 FILLER_61_137 ();
 sg13g2_decap_8 FILLER_61_144 ();
 sg13g2_decap_4 FILLER_61_151 ();
 sg13g2_fill_2 FILLER_61_155 ();
 sg13g2_decap_4 FILLER_61_222 ();
 sg13g2_decap_4 FILLER_61_231 ();
 sg13g2_fill_1 FILLER_61_235 ();
 sg13g2_fill_2 FILLER_61_240 ();
 sg13g2_decap_8 FILLER_61_263 ();
 sg13g2_decap_8 FILLER_61_270 ();
 sg13g2_decap_8 FILLER_61_277 ();
 sg13g2_decap_8 FILLER_61_314 ();
 sg13g2_decap_8 FILLER_61_321 ();
 sg13g2_decap_4 FILLER_61_328 ();
 sg13g2_fill_1 FILLER_61_336 ();
 sg13g2_decap_8 FILLER_61_341 ();
 sg13g2_fill_2 FILLER_61_374 ();
 sg13g2_fill_1 FILLER_61_376 ();
 sg13g2_fill_2 FILLER_61_392 ();
 sg13g2_fill_1 FILLER_61_394 ();
 sg13g2_decap_4 FILLER_61_399 ();
 sg13g2_fill_1 FILLER_61_403 ();
 sg13g2_decap_8 FILLER_61_414 ();
 sg13g2_decap_4 FILLER_61_421 ();
 sg13g2_fill_1 FILLER_61_425 ();
 sg13g2_decap_8 FILLER_61_440 ();
 sg13g2_decap_4 FILLER_61_447 ();
 sg13g2_fill_1 FILLER_61_451 ();
 sg13g2_decap_8 FILLER_61_488 ();
 sg13g2_decap_4 FILLER_61_495 ();
 sg13g2_fill_2 FILLER_61_499 ();
 sg13g2_decap_8 FILLER_61_522 ();
 sg13g2_decap_4 FILLER_61_529 ();
 sg13g2_fill_1 FILLER_61_600 ();
 sg13g2_fill_2 FILLER_61_606 ();
 sg13g2_fill_2 FILLER_61_625 ();
 sg13g2_fill_2 FILLER_61_636 ();
 sg13g2_fill_2 FILLER_61_692 ();
 sg13g2_decap_4 FILLER_61_699 ();
 sg13g2_fill_2 FILLER_61_709 ();
 sg13g2_fill_2 FILLER_61_715 ();
 sg13g2_fill_2 FILLER_61_722 ();
 sg13g2_fill_2 FILLER_61_728 ();
 sg13g2_fill_1 FILLER_61_730 ();
 sg13g2_fill_1 FILLER_61_767 ();
 sg13g2_fill_1 FILLER_61_772 ();
 sg13g2_fill_1 FILLER_61_799 ();
 sg13g2_fill_1 FILLER_61_806 ();
 sg13g2_fill_1 FILLER_61_821 ();
 sg13g2_decap_4 FILLER_61_827 ();
 sg13g2_fill_1 FILLER_61_835 ();
 sg13g2_fill_2 FILLER_61_845 ();
 sg13g2_fill_2 FILLER_61_855 ();
 sg13g2_fill_1 FILLER_61_857 ();
 sg13g2_decap_8 FILLER_61_862 ();
 sg13g2_decap_8 FILLER_61_892 ();
 sg13g2_fill_1 FILLER_61_903 ();
 sg13g2_decap_8 FILLER_61_908 ();
 sg13g2_decap_8 FILLER_61_915 ();
 sg13g2_fill_2 FILLER_61_922 ();
 sg13g2_fill_2 FILLER_61_942 ();
 sg13g2_fill_2 FILLER_61_950 ();
 sg13g2_fill_1 FILLER_61_952 ();
 sg13g2_fill_1 FILLER_61_962 ();
 sg13g2_fill_1 FILLER_61_967 ();
 sg13g2_fill_1 FILLER_61_974 ();
 sg13g2_fill_1 FILLER_61_980 ();
 sg13g2_decap_8 FILLER_61_999 ();
 sg13g2_decap_8 FILLER_61_1006 ();
 sg13g2_decap_4 FILLER_61_1017 ();
 sg13g2_fill_1 FILLER_61_1021 ();
 sg13g2_decap_8 FILLER_61_1026 ();
 sg13g2_decap_8 FILLER_61_1047 ();
 sg13g2_decap_8 FILLER_61_1064 ();
 sg13g2_decap_8 FILLER_61_1071 ();
 sg13g2_decap_4 FILLER_61_1078 ();
 sg13g2_fill_1 FILLER_61_1082 ();
 sg13g2_fill_2 FILLER_61_1145 ();
 sg13g2_fill_1 FILLER_61_1147 ();
 sg13g2_decap_8 FILLER_61_1188 ();
 sg13g2_fill_2 FILLER_61_1195 ();
 sg13g2_fill_2 FILLER_61_1241 ();
 sg13g2_decap_8 FILLER_61_1247 ();
 sg13g2_fill_2 FILLER_61_1280 ();
 sg13g2_fill_1 FILLER_61_1282 ();
 sg13g2_decap_4 FILLER_61_1287 ();
 sg13g2_decap_8 FILLER_61_1317 ();
 sg13g2_fill_2 FILLER_61_1324 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_6 ();
 sg13g2_decap_8 FILLER_62_17 ();
 sg13g2_decap_8 FILLER_62_24 ();
 sg13g2_fill_1 FILLER_62_31 ();
 sg13g2_decap_8 FILLER_62_48 ();
 sg13g2_decap_8 FILLER_62_55 ();
 sg13g2_decap_4 FILLER_62_66 ();
 sg13g2_decap_4 FILLER_62_92 ();
 sg13g2_fill_1 FILLER_62_104 ();
 sg13g2_decap_8 FILLER_62_110 ();
 sg13g2_decap_8 FILLER_62_117 ();
 sg13g2_fill_1 FILLER_62_124 ();
 sg13g2_decap_8 FILLER_62_155 ();
 sg13g2_decap_8 FILLER_62_162 ();
 sg13g2_decap_8 FILLER_62_169 ();
 sg13g2_decap_8 FILLER_62_184 ();
 sg13g2_fill_2 FILLER_62_201 ();
 sg13g2_fill_2 FILLER_62_207 ();
 sg13g2_fill_2 FILLER_62_213 ();
 sg13g2_fill_1 FILLER_62_215 ();
 sg13g2_fill_1 FILLER_62_221 ();
 sg13g2_fill_2 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_244 ();
 sg13g2_fill_1 FILLER_62_246 ();
 sg13g2_fill_2 FILLER_62_257 ();
 sg13g2_fill_2 FILLER_62_285 ();
 sg13g2_fill_1 FILLER_62_297 ();
 sg13g2_decap_8 FILLER_62_302 ();
 sg13g2_decap_4 FILLER_62_309 ();
 sg13g2_decap_4 FILLER_62_322 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_decap_8 FILLER_62_331 ();
 sg13g2_fill_2 FILLER_62_338 ();
 sg13g2_decap_8 FILLER_62_344 ();
 sg13g2_decap_8 FILLER_62_398 ();
 sg13g2_decap_8 FILLER_62_405 ();
 sg13g2_decap_4 FILLER_62_412 ();
 sg13g2_fill_2 FILLER_62_416 ();
 sg13g2_decap_8 FILLER_62_479 ();
 sg13g2_decap_4 FILLER_62_528 ();
 sg13g2_fill_2 FILLER_62_532 ();
 sg13g2_fill_2 FILLER_62_538 ();
 sg13g2_fill_1 FILLER_62_540 ();
 sg13g2_fill_2 FILLER_62_545 ();
 sg13g2_fill_1 FILLER_62_547 ();
 sg13g2_decap_4 FILLER_62_558 ();
 sg13g2_fill_1 FILLER_62_562 ();
 sg13g2_fill_1 FILLER_62_573 ();
 sg13g2_decap_4 FILLER_62_604 ();
 sg13g2_decap_4 FILLER_62_639 ();
 sg13g2_fill_1 FILLER_62_648 ();
 sg13g2_fill_1 FILLER_62_654 ();
 sg13g2_fill_2 FILLER_62_663 ();
 sg13g2_fill_1 FILLER_62_665 ();
 sg13g2_fill_2 FILLER_62_704 ();
 sg13g2_fill_2 FILLER_62_717 ();
 sg13g2_decap_8 FILLER_62_724 ();
 sg13g2_fill_1 FILLER_62_731 ();
 sg13g2_decap_8 FILLER_62_741 ();
 sg13g2_decap_8 FILLER_62_748 ();
 sg13g2_fill_2 FILLER_62_755 ();
 sg13g2_fill_1 FILLER_62_757 ();
 sg13g2_decap_4 FILLER_62_766 ();
 sg13g2_decap_4 FILLER_62_774 ();
 sg13g2_fill_2 FILLER_62_778 ();
 sg13g2_decap_8 FILLER_62_784 ();
 sg13g2_fill_1 FILLER_62_800 ();
 sg13g2_fill_2 FILLER_62_853 ();
 sg13g2_fill_1 FILLER_62_864 ();
 sg13g2_fill_1 FILLER_62_870 ();
 sg13g2_fill_1 FILLER_62_885 ();
 sg13g2_decap_8 FILLER_62_915 ();
 sg13g2_decap_8 FILLER_62_922 ();
 sg13g2_fill_1 FILLER_62_929 ();
 sg13g2_decap_4 FILLER_62_935 ();
 sg13g2_fill_1 FILLER_62_952 ();
 sg13g2_fill_1 FILLER_62_961 ();
 sg13g2_fill_2 FILLER_62_966 ();
 sg13g2_fill_1 FILLER_62_973 ();
 sg13g2_fill_1 FILLER_62_984 ();
 sg13g2_fill_1 FILLER_62_990 ();
 sg13g2_fill_1 FILLER_62_1017 ();
 sg13g2_fill_2 FILLER_62_1022 ();
 sg13g2_fill_1 FILLER_62_1050 ();
 sg13g2_fill_2 FILLER_62_1061 ();
 sg13g2_decap_4 FILLER_62_1073 ();
 sg13g2_fill_1 FILLER_62_1117 ();
 sg13g2_fill_1 FILLER_62_1146 ();
 sg13g2_decap_8 FILLER_62_1183 ();
 sg13g2_decap_8 FILLER_62_1190 ();
 sg13g2_decap_8 FILLER_62_1197 ();
 sg13g2_decap_8 FILLER_62_1208 ();
 sg13g2_decap_8 FILLER_62_1215 ();
 sg13g2_fill_2 FILLER_62_1222 ();
 sg13g2_fill_2 FILLER_62_1234 ();
 sg13g2_fill_1 FILLER_62_1236 ();
 sg13g2_fill_2 FILLER_62_1273 ();
 sg13g2_fill_1 FILLER_62_1275 ();
 sg13g2_decap_8 FILLER_62_1312 ();
 sg13g2_decap_8 FILLER_62_1319 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_71 ();
 sg13g2_decap_8 FILLER_63_78 ();
 sg13g2_decap_8 FILLER_63_85 ();
 sg13g2_decap_8 FILLER_63_92 ();
 sg13g2_decap_8 FILLER_63_99 ();
 sg13g2_decap_8 FILLER_63_106 ();
 sg13g2_decap_4 FILLER_63_113 ();
 sg13g2_decap_4 FILLER_63_161 ();
 sg13g2_fill_1 FILLER_63_165 ();
 sg13g2_fill_2 FILLER_63_171 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_decap_8 FILLER_63_184 ();
 sg13g2_decap_8 FILLER_63_191 ();
 sg13g2_decap_8 FILLER_63_198 ();
 sg13g2_decap_8 FILLER_63_205 ();
 sg13g2_decap_8 FILLER_63_212 ();
 sg13g2_fill_1 FILLER_63_219 ();
 sg13g2_fill_2 FILLER_63_254 ();
 sg13g2_decap_8 FILLER_63_286 ();
 sg13g2_decap_8 FILLER_63_293 ();
 sg13g2_decap_8 FILLER_63_300 ();
 sg13g2_fill_2 FILLER_63_307 ();
 sg13g2_fill_1 FILLER_63_309 ();
 sg13g2_fill_2 FILLER_63_346 ();
 sg13g2_fill_1 FILLER_63_348 ();
 sg13g2_decap_4 FILLER_63_370 ();
 sg13g2_fill_2 FILLER_63_374 ();
 sg13g2_fill_2 FILLER_63_380 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_decap_4 FILLER_63_397 ();
 sg13g2_decap_8 FILLER_63_409 ();
 sg13g2_decap_8 FILLER_63_416 ();
 sg13g2_decap_8 FILLER_63_423 ();
 sg13g2_decap_4 FILLER_63_430 ();
 sg13g2_fill_2 FILLER_63_468 ();
 sg13g2_decap_4 FILLER_63_491 ();
 sg13g2_fill_2 FILLER_63_500 ();
 sg13g2_decap_4 FILLER_63_523 ();
 sg13g2_fill_2 FILLER_63_574 ();
 sg13g2_decap_8 FILLER_63_590 ();
 sg13g2_decap_8 FILLER_63_597 ();
 sg13g2_decap_8 FILLER_63_604 ();
 sg13g2_decap_8 FILLER_63_611 ();
 sg13g2_fill_2 FILLER_63_618 ();
 sg13g2_fill_1 FILLER_63_620 ();
 sg13g2_fill_2 FILLER_63_630 ();
 sg13g2_decap_4 FILLER_63_706 ();
 sg13g2_decap_4 FILLER_63_719 ();
 sg13g2_fill_2 FILLER_63_727 ();
 sg13g2_fill_1 FILLER_63_729 ();
 sg13g2_fill_2 FILLER_63_756 ();
 sg13g2_decap_8 FILLER_63_762 ();
 sg13g2_decap_8 FILLER_63_769 ();
 sg13g2_decap_8 FILLER_63_776 ();
 sg13g2_decap_4 FILLER_63_783 ();
 sg13g2_fill_1 FILLER_63_787 ();
 sg13g2_decap_4 FILLER_63_792 ();
 sg13g2_fill_1 FILLER_63_796 ();
 sg13g2_fill_2 FILLER_63_807 ();
 sg13g2_decap_8 FILLER_63_829 ();
 sg13g2_fill_2 FILLER_63_836 ();
 sg13g2_fill_1 FILLER_63_838 ();
 sg13g2_fill_1 FILLER_63_848 ();
 sg13g2_decap_8 FILLER_63_853 ();
 sg13g2_fill_1 FILLER_63_860 ();
 sg13g2_fill_2 FILLER_63_865 ();
 sg13g2_fill_1 FILLER_63_913 ();
 sg13g2_fill_2 FILLER_63_974 ();
 sg13g2_fill_1 FILLER_63_981 ();
 sg13g2_fill_2 FILLER_63_993 ();
 sg13g2_fill_1 FILLER_63_995 ();
 sg13g2_decap_8 FILLER_63_1005 ();
 sg13g2_decap_8 FILLER_63_1012 ();
 sg13g2_decap_8 FILLER_63_1019 ();
 sg13g2_decap_4 FILLER_63_1026 ();
 sg13g2_fill_1 FILLER_63_1030 ();
 sg13g2_fill_2 FILLER_63_1057 ();
 sg13g2_fill_1 FILLER_63_1059 ();
 sg13g2_decap_8 FILLER_63_1110 ();
 sg13g2_decap_8 FILLER_63_1117 ();
 sg13g2_fill_1 FILLER_63_1124 ();
 sg13g2_decap_8 FILLER_63_1129 ();
 sg13g2_decap_8 FILLER_63_1136 ();
 sg13g2_fill_1 FILLER_63_1143 ();
 sg13g2_decap_8 FILLER_63_1189 ();
 sg13g2_decap_8 FILLER_63_1196 ();
 sg13g2_decap_4 FILLER_63_1203 ();
 sg13g2_decap_8 FILLER_63_1233 ();
 sg13g2_fill_2 FILLER_63_1240 ();
 sg13g2_fill_2 FILLER_63_1306 ();
 sg13g2_decap_8 FILLER_63_1312 ();
 sg13g2_decap_8 FILLER_63_1319 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_fill_2 FILLER_64_75 ();
 sg13g2_fill_1 FILLER_64_77 ();
 sg13g2_decap_4 FILLER_64_99 ();
 sg13g2_decap_4 FILLER_64_113 ();
 sg13g2_fill_2 FILLER_64_117 ();
 sg13g2_fill_2 FILLER_64_146 ();
 sg13g2_decap_8 FILLER_64_194 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_fill_1 FILLER_64_217 ();
 sg13g2_decap_8 FILLER_64_222 ();
 sg13g2_fill_2 FILLER_64_229 ();
 sg13g2_fill_1 FILLER_64_231 ();
 sg13g2_fill_2 FILLER_64_236 ();
 sg13g2_fill_1 FILLER_64_238 ();
 sg13g2_fill_2 FILLER_64_274 ();
 sg13g2_decap_4 FILLER_64_302 ();
 sg13g2_fill_1 FILLER_64_306 ();
 sg13g2_fill_1 FILLER_64_314 ();
 sg13g2_fill_2 FILLER_64_320 ();
 sg13g2_fill_1 FILLER_64_322 ();
 sg13g2_decap_4 FILLER_64_363 ();
 sg13g2_fill_2 FILLER_64_367 ();
 sg13g2_decap_4 FILLER_64_395 ();
 sg13g2_fill_2 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_4 FILLER_64_417 ();
 sg13g2_fill_1 FILLER_64_421 ();
 sg13g2_decap_4 FILLER_64_427 ();
 sg13g2_fill_2 FILLER_64_431 ();
 sg13g2_fill_1 FILLER_64_442 ();
 sg13g2_fill_1 FILLER_64_512 ();
 sg13g2_decap_8 FILLER_64_527 ();
 sg13g2_decap_4 FILLER_64_565 ();
 sg13g2_fill_2 FILLER_64_569 ();
 sg13g2_decap_8 FILLER_64_592 ();
 sg13g2_decap_8 FILLER_64_599 ();
 sg13g2_decap_8 FILLER_64_606 ();
 sg13g2_decap_8 FILLER_64_613 ();
 sg13g2_decap_4 FILLER_64_620 ();
 sg13g2_fill_1 FILLER_64_624 ();
 sg13g2_fill_1 FILLER_64_628 ();
 sg13g2_fill_2 FILLER_64_633 ();
 sg13g2_fill_1 FILLER_64_656 ();
 sg13g2_fill_2 FILLER_64_681 ();
 sg13g2_fill_1 FILLER_64_687 ();
 sg13g2_decap_8 FILLER_64_696 ();
 sg13g2_decap_8 FILLER_64_703 ();
 sg13g2_decap_8 FILLER_64_710 ();
 sg13g2_decap_4 FILLER_64_717 ();
 sg13g2_fill_2 FILLER_64_721 ();
 sg13g2_fill_2 FILLER_64_749 ();
 sg13g2_fill_2 FILLER_64_763 ();
 sg13g2_fill_1 FILLER_64_765 ();
 sg13g2_decap_8 FILLER_64_814 ();
 sg13g2_decap_8 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_4 FILLER_64_845 ();
 sg13g2_fill_1 FILLER_64_849 ();
 sg13g2_fill_1 FILLER_64_876 ();
 sg13g2_decap_4 FILLER_64_887 ();
 sg13g2_fill_2 FILLER_64_891 ();
 sg13g2_fill_2 FILLER_64_902 ();
 sg13g2_fill_1 FILLER_64_911 ();
 sg13g2_fill_2 FILLER_64_920 ();
 sg13g2_fill_1 FILLER_64_922 ();
 sg13g2_fill_1 FILLER_64_933 ();
 sg13g2_fill_2 FILLER_64_939 ();
 sg13g2_fill_1 FILLER_64_946 ();
 sg13g2_decap_4 FILLER_64_955 ();
 sg13g2_fill_1 FILLER_64_959 ();
 sg13g2_fill_1 FILLER_64_970 ();
 sg13g2_decap_8 FILLER_64_1006 ();
 sg13g2_decap_8 FILLER_64_1013 ();
 sg13g2_decap_8 FILLER_64_1020 ();
 sg13g2_decap_8 FILLER_64_1027 ();
 sg13g2_fill_2 FILLER_64_1034 ();
 sg13g2_fill_1 FILLER_64_1036 ();
 sg13g2_fill_1 FILLER_64_1041 ();
 sg13g2_fill_1 FILLER_64_1046 ();
 sg13g2_decap_4 FILLER_64_1077 ();
 sg13g2_fill_1 FILLER_64_1081 ();
 sg13g2_fill_1 FILLER_64_1092 ();
 sg13g2_decap_4 FILLER_64_1119 ();
 sg13g2_fill_1 FILLER_64_1127 ();
 sg13g2_decap_8 FILLER_64_1138 ();
 sg13g2_decap_8 FILLER_64_1145 ();
 sg13g2_decap_8 FILLER_64_1152 ();
 sg13g2_fill_2 FILLER_64_1159 ();
 sg13g2_fill_2 FILLER_64_1205 ();
 sg13g2_fill_2 FILLER_64_1237 ();
 sg13g2_fill_2 FILLER_64_1275 ();
 sg13g2_fill_1 FILLER_64_1277 ();
 sg13g2_decap_8 FILLER_64_1290 ();
 sg13g2_fill_2 FILLER_64_1297 ();
 sg13g2_fill_1 FILLER_64_1299 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_fill_2 FILLER_65_54 ();
 sg13g2_fill_1 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_83 ();
 sg13g2_fill_1 FILLER_65_85 ();
 sg13g2_decap_8 FILLER_65_107 ();
 sg13g2_decap_8 FILLER_65_114 ();
 sg13g2_decap_8 FILLER_65_121 ();
 sg13g2_decap_4 FILLER_65_128 ();
 sg13g2_fill_1 FILLER_65_132 ();
 sg13g2_fill_2 FILLER_65_141 ();
 sg13g2_fill_2 FILLER_65_168 ();
 sg13g2_fill_2 FILLER_65_199 ();
 sg13g2_fill_2 FILLER_65_205 ();
 sg13g2_fill_1 FILLER_65_207 ();
 sg13g2_fill_1 FILLER_65_213 ();
 sg13g2_decap_8 FILLER_65_228 ();
 sg13g2_decap_4 FILLER_65_235 ();
 sg13g2_fill_1 FILLER_65_239 ();
 sg13g2_decap_8 FILLER_65_258 ();
 sg13g2_decap_8 FILLER_65_265 ();
 sg13g2_fill_2 FILLER_65_272 ();
 sg13g2_fill_2 FILLER_65_295 ();
 sg13g2_fill_1 FILLER_65_297 ();
 sg13g2_fill_1 FILLER_65_310 ();
 sg13g2_fill_1 FILLER_65_323 ();
 sg13g2_fill_1 FILLER_65_334 ();
 sg13g2_fill_1 FILLER_65_361 ();
 sg13g2_decap_4 FILLER_65_377 ();
 sg13g2_fill_2 FILLER_65_381 ();
 sg13g2_fill_2 FILLER_65_387 ();
 sg13g2_fill_1 FILLER_65_389 ();
 sg13g2_decap_4 FILLER_65_394 ();
 sg13g2_fill_1 FILLER_65_480 ();
 sg13g2_fill_1 FILLER_65_485 ();
 sg13g2_fill_2 FILLER_65_494 ();
 sg13g2_fill_2 FILLER_65_512 ();
 sg13g2_fill_1 FILLER_65_514 ();
 sg13g2_decap_4 FILLER_65_554 ();
 sg13g2_fill_1 FILLER_65_558 ();
 sg13g2_decap_4 FILLER_65_564 ();
 sg13g2_fill_2 FILLER_65_568 ();
 sg13g2_decap_8 FILLER_65_606 ();
 sg13g2_decap_8 FILLER_65_613 ();
 sg13g2_decap_8 FILLER_65_620 ();
 sg13g2_fill_2 FILLER_65_627 ();
 sg13g2_fill_1 FILLER_65_629 ();
 sg13g2_fill_1 FILLER_65_634 ();
 sg13g2_decap_8 FILLER_65_651 ();
 sg13g2_decap_8 FILLER_65_658 ();
 sg13g2_decap_4 FILLER_65_665 ();
 sg13g2_decap_4 FILLER_65_674 ();
 sg13g2_fill_1 FILLER_65_682 ();
 sg13g2_fill_2 FILLER_65_713 ();
 sg13g2_fill_1 FILLER_65_755 ();
 sg13g2_fill_2 FILLER_65_790 ();
 sg13g2_decap_4 FILLER_65_830 ();
 sg13g2_fill_2 FILLER_65_838 ();
 sg13g2_decap_8 FILLER_65_850 ();
 sg13g2_fill_1 FILLER_65_857 ();
 sg13g2_decap_4 FILLER_65_862 ();
 sg13g2_fill_1 FILLER_65_866 ();
 sg13g2_fill_1 FILLER_65_871 ();
 sg13g2_decap_4 FILLER_65_876 ();
 sg13g2_fill_1 FILLER_65_880 ();
 sg13g2_fill_2 FILLER_65_901 ();
 sg13g2_fill_1 FILLER_65_903 ();
 sg13g2_fill_1 FILLER_65_908 ();
 sg13g2_fill_1 FILLER_65_914 ();
 sg13g2_fill_1 FILLER_65_919 ();
 sg13g2_fill_1 FILLER_65_925 ();
 sg13g2_fill_1 FILLER_65_942 ();
 sg13g2_fill_1 FILLER_65_948 ();
 sg13g2_fill_1 FILLER_65_962 ();
 sg13g2_fill_2 FILLER_65_1007 ();
 sg13g2_decap_4 FILLER_65_1039 ();
 sg13g2_fill_2 FILLER_65_1043 ();
 sg13g2_decap_8 FILLER_65_1055 ();
 sg13g2_fill_2 FILLER_65_1062 ();
 sg13g2_fill_2 FILLER_65_1094 ();
 sg13g2_fill_1 FILLER_65_1100 ();
 sg13g2_fill_1 FILLER_65_1127 ();
 sg13g2_fill_1 FILLER_65_1138 ();
 sg13g2_decap_4 FILLER_65_1165 ();
 sg13g2_decap_4 FILLER_65_1209 ();
 sg13g2_decap_4 FILLER_65_1221 ();
 sg13g2_fill_2 FILLER_65_1225 ();
 sg13g2_decap_8 FILLER_65_1237 ();
 sg13g2_fill_2 FILLER_65_1244 ();
 sg13g2_fill_1 FILLER_65_1246 ();
 sg13g2_decap_8 FILLER_65_1283 ();
 sg13g2_decap_8 FILLER_65_1290 ();
 sg13g2_decap_8 FILLER_65_1297 ();
 sg13g2_decap_8 FILLER_65_1304 ();
 sg13g2_decap_8 FILLER_65_1311 ();
 sg13g2_decap_8 FILLER_65_1318 ();
 sg13g2_fill_1 FILLER_65_1325 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_4 FILLER_66_21 ();
 sg13g2_fill_1 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_46 ();
 sg13g2_fill_2 FILLER_66_73 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_4 FILLER_66_112 ();
 sg13g2_fill_2 FILLER_66_116 ();
 sg13g2_fill_1 FILLER_66_143 ();
 sg13g2_decap_8 FILLER_66_190 ();
 sg13g2_decap_4 FILLER_66_197 ();
 sg13g2_fill_1 FILLER_66_201 ();
 sg13g2_fill_2 FILLER_66_214 ();
 sg13g2_fill_1 FILLER_66_216 ();
 sg13g2_fill_2 FILLER_66_243 ();
 sg13g2_decap_8 FILLER_66_255 ();
 sg13g2_decap_4 FILLER_66_262 ();
 sg13g2_decap_8 FILLER_66_295 ();
 sg13g2_decap_8 FILLER_66_302 ();
 sg13g2_fill_2 FILLER_66_309 ();
 sg13g2_fill_1 FILLER_66_311 ();
 sg13g2_fill_2 FILLER_66_316 ();
 sg13g2_fill_1 FILLER_66_318 ();
 sg13g2_fill_1 FILLER_66_333 ();
 sg13g2_fill_1 FILLER_66_360 ();
 sg13g2_fill_1 FILLER_66_369 ();
 sg13g2_fill_2 FILLER_66_374 ();
 sg13g2_fill_2 FILLER_66_384 ();
 sg13g2_fill_1 FILLER_66_386 ();
 sg13g2_fill_2 FILLER_66_427 ();
 sg13g2_decap_4 FILLER_66_463 ();
 sg13g2_fill_2 FILLER_66_467 ();
 sg13g2_decap_4 FILLER_66_473 ();
 sg13g2_fill_1 FILLER_66_512 ();
 sg13g2_decap_4 FILLER_66_534 ();
 sg13g2_fill_1 FILLER_66_538 ();
 sg13g2_decap_4 FILLER_66_543 ();
 sg13g2_fill_2 FILLER_66_583 ();
 sg13g2_fill_1 FILLER_66_585 ();
 sg13g2_fill_1 FILLER_66_590 ();
 sg13g2_decap_4 FILLER_66_599 ();
 sg13g2_decap_8 FILLER_66_637 ();
 sg13g2_decap_8 FILLER_66_644 ();
 sg13g2_decap_8 FILLER_66_651 ();
 sg13g2_decap_8 FILLER_66_658 ();
 sg13g2_decap_8 FILLER_66_665 ();
 sg13g2_decap_8 FILLER_66_672 ();
 sg13g2_decap_8 FILLER_66_679 ();
 sg13g2_fill_1 FILLER_66_686 ();
 sg13g2_fill_1 FILLER_66_739 ();
 sg13g2_fill_2 FILLER_66_745 ();
 sg13g2_fill_1 FILLER_66_747 ();
 sg13g2_fill_1 FILLER_66_753 ();
 sg13g2_fill_1 FILLER_66_758 ();
 sg13g2_fill_2 FILLER_66_773 ();
 sg13g2_fill_1 FILLER_66_775 ();
 sg13g2_fill_2 FILLER_66_781 ();
 sg13g2_decap_4 FILLER_66_787 ();
 sg13g2_fill_2 FILLER_66_791 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_fill_2 FILLER_66_857 ();
 sg13g2_fill_2 FILLER_66_863 ();
 sg13g2_fill_1 FILLER_66_865 ();
 sg13g2_decap_8 FILLER_66_896 ();
 sg13g2_decap_8 FILLER_66_903 ();
 sg13g2_decap_4 FILLER_66_910 ();
 sg13g2_fill_2 FILLER_66_918 ();
 sg13g2_fill_1 FILLER_66_929 ();
 sg13g2_fill_1 FILLER_66_934 ();
 sg13g2_fill_2 FILLER_66_969 ();
 sg13g2_fill_1 FILLER_66_986 ();
 sg13g2_fill_1 FILLER_66_992 ();
 sg13g2_fill_2 FILLER_66_996 ();
 sg13g2_fill_2 FILLER_66_1002 ();
 sg13g2_decap_8 FILLER_66_1046 ();
 sg13g2_decap_8 FILLER_66_1053 ();
 sg13g2_decap_4 FILLER_66_1060 ();
 sg13g2_fill_1 FILLER_66_1064 ();
 sg13g2_fill_2 FILLER_66_1069 ();
 sg13g2_fill_1 FILLER_66_1071 ();
 sg13g2_decap_4 FILLER_66_1082 ();
 sg13g2_fill_1 FILLER_66_1086 ();
 sg13g2_decap_4 FILLER_66_1113 ();
 sg13g2_fill_1 FILLER_66_1117 ();
 sg13g2_decap_8 FILLER_66_1156 ();
 sg13g2_decap_4 FILLER_66_1173 ();
 sg13g2_fill_1 FILLER_66_1177 ();
 sg13g2_decap_8 FILLER_66_1182 ();
 sg13g2_decap_8 FILLER_66_1193 ();
 sg13g2_decap_8 FILLER_66_1200 ();
 sg13g2_fill_1 FILLER_66_1207 ();
 sg13g2_decap_4 FILLER_66_1244 ();
 sg13g2_fill_2 FILLER_66_1248 ();
 sg13g2_decap_8 FILLER_66_1276 ();
 sg13g2_decap_8 FILLER_66_1283 ();
 sg13g2_decap_8 FILLER_66_1290 ();
 sg13g2_decap_8 FILLER_66_1297 ();
 sg13g2_decap_8 FILLER_66_1304 ();
 sg13g2_decap_8 FILLER_66_1311 ();
 sg13g2_decap_8 FILLER_66_1318 ();
 sg13g2_fill_1 FILLER_66_1325 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_4 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_25 ();
 sg13g2_fill_1 FILLER_67_67 ();
 sg13g2_fill_2 FILLER_67_115 ();
 sg13g2_fill_1 FILLER_67_117 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_fill_2 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_183 ();
 sg13g2_decap_8 FILLER_67_190 ();
 sg13g2_decap_8 FILLER_67_197 ();
 sg13g2_decap_4 FILLER_67_204 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_decap_4 FILLER_67_329 ();
 sg13g2_fill_1 FILLER_67_337 ();
 sg13g2_fill_1 FILLER_67_342 ();
 sg13g2_fill_1 FILLER_67_347 ();
 sg13g2_fill_1 FILLER_67_353 ();
 sg13g2_fill_1 FILLER_67_359 ();
 sg13g2_fill_1 FILLER_67_364 ();
 sg13g2_fill_1 FILLER_67_375 ();
 sg13g2_fill_2 FILLER_67_402 ();
 sg13g2_decap_4 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_67_433 ();
 sg13g2_decap_4 FILLER_67_456 ();
 sg13g2_decap_4 FILLER_67_496 ();
 sg13g2_decap_4 FILLER_67_531 ();
 sg13g2_fill_1 FILLER_67_535 ();
 sg13g2_fill_2 FILLER_67_572 ();
 sg13g2_fill_1 FILLER_67_574 ();
 sg13g2_decap_4 FILLER_67_587 ();
 sg13g2_decap_4 FILLER_67_607 ();
 sg13g2_fill_1 FILLER_67_611 ();
 sg13g2_fill_2 FILLER_67_616 ();
 sg13g2_fill_1 FILLER_67_652 ();
 sg13g2_decap_8 FILLER_67_657 ();
 sg13g2_decap_8 FILLER_67_664 ();
 sg13g2_decap_8 FILLER_67_671 ();
 sg13g2_decap_8 FILLER_67_678 ();
 sg13g2_decap_8 FILLER_67_685 ();
 sg13g2_fill_2 FILLER_67_696 ();
 sg13g2_fill_2 FILLER_67_702 ();
 sg13g2_fill_1 FILLER_67_704 ();
 sg13g2_decap_4 FILLER_67_708 ();
 sg13g2_fill_1 FILLER_67_712 ();
 sg13g2_decap_8 FILLER_67_723 ();
 sg13g2_fill_2 FILLER_67_743 ();
 sg13g2_decap_4 FILLER_67_750 ();
 sg13g2_fill_2 FILLER_67_754 ();
 sg13g2_fill_1 FILLER_67_835 ();
 sg13g2_decap_8 FILLER_67_867 ();
 sg13g2_decap_8 FILLER_67_874 ();
 sg13g2_decap_8 FILLER_67_881 ();
 sg13g2_decap_8 FILLER_67_888 ();
 sg13g2_decap_8 FILLER_67_921 ();
 sg13g2_decap_8 FILLER_67_928 ();
 sg13g2_decap_4 FILLER_67_943 ();
 sg13g2_fill_2 FILLER_67_957 ();
 sg13g2_fill_1 FILLER_67_959 ();
 sg13g2_decap_4 FILLER_67_965 ();
 sg13g2_fill_1 FILLER_67_969 ();
 sg13g2_decap_8 FILLER_67_974 ();
 sg13g2_decap_8 FILLER_67_981 ();
 sg13g2_decap_8 FILLER_67_988 ();
 sg13g2_decap_4 FILLER_67_995 ();
 sg13g2_fill_1 FILLER_67_999 ();
 sg13g2_decap_4 FILLER_67_1037 ();
 sg13g2_fill_1 FILLER_67_1041 ();
 sg13g2_fill_2 FILLER_67_1050 ();
 sg13g2_fill_2 FILLER_67_1056 ();
 sg13g2_decap_8 FILLER_67_1084 ();
 sg13g2_fill_2 FILLER_67_1091 ();
 sg13g2_fill_1 FILLER_67_1093 ();
 sg13g2_decap_4 FILLER_67_1098 ();
 sg13g2_fill_1 FILLER_67_1102 ();
 sg13g2_fill_1 FILLER_67_1113 ();
 sg13g2_fill_2 FILLER_67_1168 ();
 sg13g2_decap_8 FILLER_67_1196 ();
 sg13g2_decap_4 FILLER_67_1203 ();
 sg13g2_fill_2 FILLER_67_1207 ();
 sg13g2_decap_8 FILLER_67_1245 ();
 sg13g2_fill_1 FILLER_67_1252 ();
 sg13g2_decap_8 FILLER_67_1283 ();
 sg13g2_decap_8 FILLER_67_1290 ();
 sg13g2_decap_8 FILLER_67_1297 ();
 sg13g2_decap_8 FILLER_67_1304 ();
 sg13g2_decap_8 FILLER_67_1311 ();
 sg13g2_decap_8 FILLER_67_1318 ();
 sg13g2_fill_1 FILLER_67_1325 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_4 FILLER_68_35 ();
 sg13g2_fill_2 FILLER_68_55 ();
 sg13g2_fill_1 FILLER_68_57 ();
 sg13g2_decap_8 FILLER_68_72 ();
 sg13g2_decap_8 FILLER_68_79 ();
 sg13g2_decap_8 FILLER_68_86 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_4 FILLER_68_112 ();
 sg13g2_decap_4 FILLER_68_120 ();
 sg13g2_fill_2 FILLER_68_128 ();
 sg13g2_fill_1 FILLER_68_130 ();
 sg13g2_fill_2 FILLER_68_139 ();
 sg13g2_fill_1 FILLER_68_141 ();
 sg13g2_fill_2 FILLER_68_168 ();
 sg13g2_fill_1 FILLER_68_170 ();
 sg13g2_decap_8 FILLER_68_207 ();
 sg13g2_fill_1 FILLER_68_214 ();
 sg13g2_decap_8 FILLER_68_296 ();
 sg13g2_decap_8 FILLER_68_303 ();
 sg13g2_fill_2 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_316 ();
 sg13g2_fill_1 FILLER_68_318 ();
 sg13g2_decap_8 FILLER_68_324 ();
 sg13g2_decap_8 FILLER_68_331 ();
 sg13g2_decap_4 FILLER_68_338 ();
 sg13g2_decap_8 FILLER_68_350 ();
 sg13g2_fill_1 FILLER_68_357 ();
 sg13g2_decap_8 FILLER_68_366 ();
 sg13g2_decap_4 FILLER_68_373 ();
 sg13g2_fill_2 FILLER_68_377 ();
 sg13g2_decap_8 FILLER_68_423 ();
 sg13g2_decap_4 FILLER_68_430 ();
 sg13g2_decap_8 FILLER_68_455 ();
 sg13g2_decap_8 FILLER_68_462 ();
 sg13g2_fill_2 FILLER_68_469 ();
 sg13g2_decap_8 FILLER_68_501 ();
 sg13g2_decap_4 FILLER_68_508 ();
 sg13g2_decap_4 FILLER_68_533 ();
 sg13g2_fill_1 FILLER_68_537 ();
 sg13g2_fill_1 FILLER_68_572 ();
 sg13g2_fill_2 FILLER_68_595 ();
 sg13g2_fill_1 FILLER_68_605 ();
 sg13g2_fill_2 FILLER_68_619 ();
 sg13g2_fill_2 FILLER_68_624 ();
 sg13g2_decap_4 FILLER_68_632 ();
 sg13g2_fill_1 FILLER_68_640 ();
 sg13g2_decap_8 FILLER_68_672 ();
 sg13g2_decap_4 FILLER_68_679 ();
 sg13g2_fill_1 FILLER_68_683 ();
 sg13g2_fill_1 FILLER_68_717 ();
 sg13g2_fill_2 FILLER_68_728 ();
 sg13g2_fill_2 FILLER_68_733 ();
 sg13g2_fill_1 FILLER_68_735 ();
 sg13g2_decap_4 FILLER_68_739 ();
 sg13g2_fill_1 FILLER_68_743 ();
 sg13g2_fill_1 FILLER_68_749 ();
 sg13g2_fill_2 FILLER_68_755 ();
 sg13g2_fill_1 FILLER_68_770 ();
 sg13g2_decap_8 FILLER_68_781 ();
 sg13g2_decap_8 FILLER_68_788 ();
 sg13g2_fill_1 FILLER_68_795 ();
 sg13g2_decap_8 FILLER_68_800 ();
 sg13g2_fill_2 FILLER_68_807 ();
 sg13g2_decap_8 FILLER_68_831 ();
 sg13g2_fill_2 FILLER_68_838 ();
 sg13g2_fill_1 FILLER_68_840 ();
 sg13g2_fill_2 FILLER_68_847 ();
 sg13g2_decap_8 FILLER_68_853 ();
 sg13g2_decap_8 FILLER_68_860 ();
 sg13g2_decap_8 FILLER_68_867 ();
 sg13g2_fill_2 FILLER_68_874 ();
 sg13g2_fill_1 FILLER_68_876 ();
 sg13g2_decap_4 FILLER_68_890 ();
 sg13g2_fill_1 FILLER_68_894 ();
 sg13g2_fill_2 FILLER_68_899 ();
 sg13g2_fill_1 FILLER_68_901 ();
 sg13g2_decap_8 FILLER_68_906 ();
 sg13g2_decap_8 FILLER_68_913 ();
 sg13g2_decap_4 FILLER_68_920 ();
 sg13g2_fill_1 FILLER_68_924 ();
 sg13g2_fill_2 FILLER_68_943 ();
 sg13g2_fill_1 FILLER_68_945 ();
 sg13g2_decap_4 FILLER_68_950 ();
 sg13g2_decap_8 FILLER_68_962 ();
 sg13g2_decap_8 FILLER_68_969 ();
 sg13g2_fill_1 FILLER_68_976 ();
 sg13g2_decap_8 FILLER_68_989 ();
 sg13g2_fill_2 FILLER_68_996 ();
 sg13g2_fill_2 FILLER_68_1038 ();
 sg13g2_fill_2 FILLER_68_1070 ();
 sg13g2_fill_1 FILLER_68_1082 ();
 sg13g2_fill_1 FILLER_68_1093 ();
 sg13g2_fill_2 FILLER_68_1120 ();
 sg13g2_fill_2 FILLER_68_1130 ();
 sg13g2_decap_4 FILLER_68_1136 ();
 sg13g2_decap_4 FILLER_68_1166 ();
 sg13g2_fill_2 FILLER_68_1180 ();
 sg13g2_fill_1 FILLER_68_1182 ();
 sg13g2_decap_8 FILLER_68_1187 ();
 sg13g2_decap_8 FILLER_68_1194 ();
 sg13g2_decap_8 FILLER_68_1201 ();
 sg13g2_decap_8 FILLER_68_1208 ();
 sg13g2_fill_1 FILLER_68_1215 ();
 sg13g2_decap_8 FILLER_68_1220 ();
 sg13g2_decap_8 FILLER_68_1227 ();
 sg13g2_decap_4 FILLER_68_1234 ();
 sg13g2_fill_1 FILLER_68_1238 ();
 sg13g2_decap_4 FILLER_68_1259 ();
 sg13g2_decap_8 FILLER_68_1267 ();
 sg13g2_decap_8 FILLER_68_1274 ();
 sg13g2_decap_8 FILLER_68_1281 ();
 sg13g2_decap_8 FILLER_68_1288 ();
 sg13g2_decap_8 FILLER_68_1295 ();
 sg13g2_decap_8 FILLER_68_1302 ();
 sg13g2_decap_8 FILLER_68_1309 ();
 sg13g2_decap_8 FILLER_68_1316 ();
 sg13g2_fill_2 FILLER_68_1323 ();
 sg13g2_fill_1 FILLER_68_1325 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_fill_2 FILLER_69_28 ();
 sg13g2_fill_1 FILLER_69_30 ();
 sg13g2_decap_4 FILLER_69_35 ();
 sg13g2_fill_1 FILLER_69_60 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_4 FILLER_69_112 ();
 sg13g2_fill_1 FILLER_69_156 ();
 sg13g2_decap_8 FILLER_69_208 ();
 sg13g2_decap_8 FILLER_69_215 ();
 sg13g2_decap_4 FILLER_69_222 ();
 sg13g2_decap_4 FILLER_69_235 ();
 sg13g2_fill_2 FILLER_69_243 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_8 FILLER_69_294 ();
 sg13g2_fill_2 FILLER_69_301 ();
 sg13g2_fill_1 FILLER_69_303 ();
 sg13g2_decap_8 FILLER_69_308 ();
 sg13g2_decap_8 FILLER_69_315 ();
 sg13g2_fill_1 FILLER_69_322 ();
 sg13g2_decap_4 FILLER_69_344 ();
 sg13g2_fill_1 FILLER_69_348 ();
 sg13g2_fill_2 FILLER_69_353 ();
 sg13g2_fill_1 FILLER_69_355 ();
 sg13g2_fill_2 FILLER_69_386 ();
 sg13g2_fill_2 FILLER_69_401 ();
 sg13g2_fill_1 FILLER_69_403 ();
 sg13g2_fill_2 FILLER_69_414 ();
 sg13g2_fill_1 FILLER_69_416 ();
 sg13g2_fill_2 FILLER_69_443 ();
 sg13g2_decap_4 FILLER_69_453 ();
 sg13g2_fill_1 FILLER_69_457 ();
 sg13g2_decap_8 FILLER_69_463 ();
 sg13g2_decap_8 FILLER_69_470 ();
 sg13g2_decap_4 FILLER_69_477 ();
 sg13g2_decap_8 FILLER_69_537 ();
 sg13g2_fill_2 FILLER_69_544 ();
 sg13g2_fill_1 FILLER_69_546 ();
 sg13g2_fill_2 FILLER_69_551 ();
 sg13g2_fill_1 FILLER_69_585 ();
 sg13g2_decap_4 FILLER_69_599 ();
 sg13g2_fill_1 FILLER_69_603 ();
 sg13g2_fill_1 FILLER_69_638 ();
 sg13g2_fill_2 FILLER_69_643 ();
 sg13g2_fill_1 FILLER_69_649 ();
 sg13g2_decap_4 FILLER_69_676 ();
 sg13g2_fill_2 FILLER_69_680 ();
 sg13g2_fill_1 FILLER_69_712 ();
 sg13g2_decap_8 FILLER_69_726 ();
 sg13g2_fill_2 FILLER_69_733 ();
 sg13g2_fill_1 FILLER_69_735 ();
 sg13g2_decap_8 FILLER_69_762 ();
 sg13g2_fill_2 FILLER_69_769 ();
 sg13g2_decap_8 FILLER_69_778 ();
 sg13g2_decap_8 FILLER_69_785 ();
 sg13g2_decap_8 FILLER_69_792 ();
 sg13g2_decap_8 FILLER_69_799 ();
 sg13g2_decap_8 FILLER_69_806 ();
 sg13g2_decap_8 FILLER_69_813 ();
 sg13g2_decap_8 FILLER_69_820 ();
 sg13g2_decap_8 FILLER_69_827 ();
 sg13g2_decap_8 FILLER_69_834 ();
 sg13g2_decap_8 FILLER_69_841 ();
 sg13g2_fill_1 FILLER_69_848 ();
 sg13g2_decap_8 FILLER_69_882 ();
 sg13g2_fill_2 FILLER_69_889 ();
 sg13g2_fill_1 FILLER_69_891 ();
 sg13g2_fill_2 FILLER_69_920 ();
 sg13g2_decap_4 FILLER_69_926 ();
 sg13g2_decap_4 FILLER_69_935 ();
 sg13g2_fill_1 FILLER_69_969 ();
 sg13g2_decap_4 FILLER_69_1005 ();
 sg13g2_decap_4 FILLER_69_1022 ();
 sg13g2_decap_4 FILLER_69_1034 ();
 sg13g2_fill_1 FILLER_69_1038 ();
 sg13g2_decap_4 FILLER_69_1043 ();
 sg13g2_decap_4 FILLER_69_1051 ();
 sg13g2_fill_2 FILLER_69_1081 ();
 sg13g2_fill_1 FILLER_69_1083 ();
 sg13g2_decap_8 FILLER_69_1114 ();
 sg13g2_decap_8 FILLER_69_1121 ();
 sg13g2_decap_8 FILLER_69_1128 ();
 sg13g2_decap_4 FILLER_69_1135 ();
 sg13g2_fill_1 FILLER_69_1139 ();
 sg13g2_decap_8 FILLER_69_1154 ();
 sg13g2_decap_4 FILLER_69_1161 ();
 sg13g2_fill_2 FILLER_69_1165 ();
 sg13g2_decap_8 FILLER_69_1197 ();
 sg13g2_decap_8 FILLER_69_1204 ();
 sg13g2_decap_8 FILLER_69_1211 ();
 sg13g2_decap_8 FILLER_69_1218 ();
 sg13g2_decap_8 FILLER_69_1225 ();
 sg13g2_decap_8 FILLER_69_1232 ();
 sg13g2_fill_2 FILLER_69_1239 ();
 sg13g2_decap_8 FILLER_69_1267 ();
 sg13g2_decap_8 FILLER_69_1274 ();
 sg13g2_decap_8 FILLER_69_1281 ();
 sg13g2_decap_8 FILLER_69_1288 ();
 sg13g2_decap_8 FILLER_69_1295 ();
 sg13g2_decap_8 FILLER_69_1302 ();
 sg13g2_decap_8 FILLER_69_1309 ();
 sg13g2_decap_8 FILLER_69_1316 ();
 sg13g2_fill_2 FILLER_69_1323 ();
 sg13g2_fill_1 FILLER_69_1325 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_4 FILLER_70_14 ();
 sg13g2_fill_1 FILLER_70_18 ();
 sg13g2_fill_1 FILLER_70_23 ();
 sg13g2_fill_2 FILLER_70_127 ();
 sg13g2_fill_2 FILLER_70_148 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_166 ();
 sg13g2_fill_1 FILLER_70_168 ();
 sg13g2_fill_1 FILLER_70_173 ();
 sg13g2_fill_2 FILLER_70_195 ();
 sg13g2_fill_1 FILLER_70_197 ();
 sg13g2_decap_8 FILLER_70_202 ();
 sg13g2_decap_4 FILLER_70_209 ();
 sg13g2_fill_1 FILLER_70_213 ();
 sg13g2_decap_8 FILLER_70_244 ();
 sg13g2_decap_8 FILLER_70_251 ();
 sg13g2_decap_8 FILLER_70_258 ();
 sg13g2_decap_8 FILLER_70_265 ();
 sg13g2_fill_1 FILLER_70_272 ();
 sg13g2_fill_2 FILLER_70_277 ();
 sg13g2_decap_8 FILLER_70_324 ();
 sg13g2_decap_8 FILLER_70_331 ();
 sg13g2_fill_2 FILLER_70_359 ();
 sg13g2_decap_8 FILLER_70_391 ();
 sg13g2_decap_8 FILLER_70_398 ();
 sg13g2_fill_1 FILLER_70_405 ();
 sg13g2_decap_4 FILLER_70_410 ();
 sg13g2_fill_2 FILLER_70_425 ();
 sg13g2_fill_1 FILLER_70_427 ();
 sg13g2_decap_8 FILLER_70_470 ();
 sg13g2_decap_8 FILLER_70_477 ();
 sg13g2_decap_4 FILLER_70_484 ();
 sg13g2_fill_2 FILLER_70_488 ();
 sg13g2_decap_8 FILLER_70_516 ();
 sg13g2_decap_8 FILLER_70_523 ();
 sg13g2_decap_8 FILLER_70_530 ();
 sg13g2_decap_8 FILLER_70_537 ();
 sg13g2_decap_8 FILLER_70_544 ();
 sg13g2_fill_1 FILLER_70_551 ();
 sg13g2_fill_2 FILLER_70_578 ();
 sg13g2_fill_1 FILLER_70_584 ();
 sg13g2_fill_1 FILLER_70_593 ();
 sg13g2_fill_1 FILLER_70_598 ();
 sg13g2_fill_1 FILLER_70_632 ();
 sg13g2_decap_4 FILLER_70_637 ();
 sg13g2_fill_2 FILLER_70_641 ();
 sg13g2_fill_2 FILLER_70_651 ();
 sg13g2_fill_2 FILLER_70_657 ();
 sg13g2_fill_1 FILLER_70_663 ();
 sg13g2_decap_4 FILLER_70_668 ();
 sg13g2_decap_8 FILLER_70_677 ();
 sg13g2_fill_2 FILLER_70_684 ();
 sg13g2_fill_1 FILLER_70_690 ();
 sg13g2_fill_1 FILLER_70_717 ();
 sg13g2_fill_1 FILLER_70_724 ();
 sg13g2_fill_1 FILLER_70_728 ();
 sg13g2_fill_1 FILLER_70_734 ();
 sg13g2_decap_4 FILLER_70_739 ();
 sg13g2_fill_1 FILLER_70_743 ();
 sg13g2_fill_2 FILLER_70_758 ();
 sg13g2_fill_1 FILLER_70_760 ();
 sg13g2_decap_4 FILLER_70_764 ();
 sg13g2_fill_1 FILLER_70_811 ();
 sg13g2_decap_8 FILLER_70_816 ();
 sg13g2_fill_2 FILLER_70_823 ();
 sg13g2_fill_2 FILLER_70_834 ();
 sg13g2_fill_2 FILLER_70_896 ();
 sg13g2_decap_4 FILLER_70_950 ();
 sg13g2_decap_8 FILLER_70_958 ();
 sg13g2_decap_8 FILLER_70_965 ();
 sg13g2_decap_8 FILLER_70_972 ();
 sg13g2_decap_4 FILLER_70_979 ();
 sg13g2_fill_1 FILLER_70_983 ();
 sg13g2_fill_1 FILLER_70_989 ();
 sg13g2_decap_8 FILLER_70_999 ();
 sg13g2_fill_2 FILLER_70_1023 ();
 sg13g2_decap_8 FILLER_70_1033 ();
 sg13g2_decap_8 FILLER_70_1040 ();
 sg13g2_decap_8 FILLER_70_1047 ();
 sg13g2_fill_1 FILLER_70_1054 ();
 sg13g2_decap_8 FILLER_70_1058 ();
 sg13g2_decap_8 FILLER_70_1065 ();
 sg13g2_decap_8 FILLER_70_1072 ();
 sg13g2_fill_2 FILLER_70_1079 ();
 sg13g2_fill_1 FILLER_70_1081 ();
 sg13g2_fill_1 FILLER_70_1100 ();
 sg13g2_fill_2 FILLER_70_1105 ();
 sg13g2_fill_2 FILLER_70_1117 ();
 sg13g2_fill_2 FILLER_70_1123 ();
 sg13g2_decap_8 FILLER_70_1161 ();
 sg13g2_decap_4 FILLER_70_1168 ();
 sg13g2_fill_1 FILLER_70_1172 ();
 sg13g2_decap_8 FILLER_70_1217 ();
 sg13g2_decap_8 FILLER_70_1224 ();
 sg13g2_decap_8 FILLER_70_1231 ();
 sg13g2_decap_8 FILLER_70_1238 ();
 sg13g2_decap_8 FILLER_70_1249 ();
 sg13g2_decap_8 FILLER_70_1256 ();
 sg13g2_decap_8 FILLER_70_1263 ();
 sg13g2_decap_8 FILLER_70_1270 ();
 sg13g2_decap_8 FILLER_70_1277 ();
 sg13g2_decap_8 FILLER_70_1284 ();
 sg13g2_decap_8 FILLER_70_1291 ();
 sg13g2_decap_8 FILLER_70_1298 ();
 sg13g2_decap_8 FILLER_70_1305 ();
 sg13g2_decap_8 FILLER_70_1312 ();
 sg13g2_decap_8 FILLER_70_1319 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_fill_2 FILLER_71_14 ();
 sg13g2_fill_1 FILLER_71_16 ();
 sg13g2_fill_2 FILLER_71_93 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_4 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_decap_8 FILLER_71_142 ();
 sg13g2_decap_8 FILLER_71_195 ();
 sg13g2_decap_8 FILLER_71_202 ();
 sg13g2_fill_2 FILLER_71_209 ();
 sg13g2_fill_1 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_240 ();
 sg13g2_decap_8 FILLER_71_268 ();
 sg13g2_decap_8 FILLER_71_275 ();
 sg13g2_fill_1 FILLER_71_339 ();
 sg13g2_fill_2 FILLER_71_344 ();
 sg13g2_fill_1 FILLER_71_346 ();
 sg13g2_fill_2 FILLER_71_367 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_385 ();
 sg13g2_fill_1 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_397 ();
 sg13g2_fill_2 FILLER_71_440 ();
 sg13g2_decap_4 FILLER_71_468 ();
 sg13g2_fill_1 FILLER_71_472 ();
 sg13g2_decap_4 FILLER_71_494 ();
 sg13g2_fill_1 FILLER_71_498 ();
 sg13g2_decap_8 FILLER_71_503 ();
 sg13g2_decap_8 FILLER_71_510 ();
 sg13g2_decap_4 FILLER_71_517 ();
 sg13g2_fill_2 FILLER_71_521 ();
 sg13g2_decap_8 FILLER_71_549 ();
 sg13g2_decap_4 FILLER_71_556 ();
 sg13g2_decap_8 FILLER_71_564 ();
 sg13g2_decap_4 FILLER_71_571 ();
 sg13g2_fill_1 FILLER_71_575 ();
 sg13g2_fill_1 FILLER_71_583 ();
 sg13g2_decap_4 FILLER_71_590 ();
 sg13g2_decap_8 FILLER_71_636 ();
 sg13g2_fill_2 FILLER_71_643 ();
 sg13g2_decap_8 FILLER_71_662 ();
 sg13g2_fill_2 FILLER_71_669 ();
 sg13g2_fill_1 FILLER_71_697 ();
 sg13g2_fill_1 FILLER_71_702 ();
 sg13g2_fill_1 FILLER_71_707 ();
 sg13g2_fill_1 FILLER_71_712 ();
 sg13g2_fill_2 FILLER_71_723 ();
 sg13g2_decap_8 FILLER_71_765 ();
 sg13g2_fill_2 FILLER_71_772 ();
 sg13g2_fill_1 FILLER_71_774 ();
 sg13g2_fill_1 FILLER_71_779 ();
 sg13g2_fill_1 FILLER_71_791 ();
 sg13g2_fill_1 FILLER_71_796 ();
 sg13g2_fill_1 FILLER_71_828 ();
 sg13g2_fill_2 FILLER_71_855 ();
 sg13g2_fill_1 FILLER_71_857 ();
 sg13g2_fill_2 FILLER_71_884 ();
 sg13g2_decap_4 FILLER_71_890 ();
 sg13g2_fill_2 FILLER_71_894 ();
 sg13g2_fill_2 FILLER_71_901 ();
 sg13g2_fill_1 FILLER_71_903 ();
 sg13g2_decap_4 FILLER_71_941 ();
 sg13g2_decap_4 FILLER_71_948 ();
 sg13g2_fill_2 FILLER_71_952 ();
 sg13g2_decap_8 FILLER_71_958 ();
 sg13g2_decap_8 FILLER_71_965 ();
 sg13g2_fill_2 FILLER_71_989 ();
 sg13g2_fill_1 FILLER_71_999 ();
 sg13g2_fill_1 FILLER_71_1005 ();
 sg13g2_fill_1 FILLER_71_1014 ();
 sg13g2_fill_2 FILLER_71_1019 ();
 sg13g2_fill_1 FILLER_71_1021 ();
 sg13g2_decap_4 FILLER_71_1048 ();
 sg13g2_fill_1 FILLER_71_1052 ();
 sg13g2_decap_8 FILLER_71_1083 ();
 sg13g2_decap_8 FILLER_71_1090 ();
 sg13g2_decap_8 FILLER_71_1097 ();
 sg13g2_decap_8 FILLER_71_1104 ();
 sg13g2_decap_8 FILLER_71_1111 ();
 sg13g2_decap_4 FILLER_71_1118 ();
 sg13g2_fill_1 FILLER_71_1122 ();
 sg13g2_decap_4 FILLER_71_1163 ();
 sg13g2_fill_1 FILLER_71_1167 ();
 sg13g2_decap_8 FILLER_71_1178 ();
 sg13g2_decap_4 FILLER_71_1185 ();
 sg13g2_fill_1 FILLER_71_1189 ();
 sg13g2_decap_8 FILLER_71_1194 ();
 sg13g2_decap_8 FILLER_71_1201 ();
 sg13g2_decap_8 FILLER_71_1208 ();
 sg13g2_decap_8 FILLER_71_1215 ();
 sg13g2_decap_8 FILLER_71_1222 ();
 sg13g2_decap_8 FILLER_71_1229 ();
 sg13g2_decap_8 FILLER_71_1236 ();
 sg13g2_decap_8 FILLER_71_1243 ();
 sg13g2_decap_8 FILLER_71_1250 ();
 sg13g2_decap_8 FILLER_71_1257 ();
 sg13g2_decap_8 FILLER_71_1264 ();
 sg13g2_decap_8 FILLER_71_1271 ();
 sg13g2_decap_8 FILLER_71_1278 ();
 sg13g2_decap_8 FILLER_71_1285 ();
 sg13g2_decap_8 FILLER_71_1292 ();
 sg13g2_decap_8 FILLER_71_1299 ();
 sg13g2_decap_8 FILLER_71_1306 ();
 sg13g2_decap_8 FILLER_71_1313 ();
 sg13g2_decap_4 FILLER_71_1320 ();
 sg13g2_fill_2 FILLER_71_1324 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_fill_2 FILLER_72_21 ();
 sg13g2_fill_1 FILLER_72_23 ();
 sg13g2_fill_2 FILLER_72_28 ();
 sg13g2_fill_1 FILLER_72_30 ();
 sg13g2_fill_1 FILLER_72_41 ();
 sg13g2_decap_8 FILLER_72_46 ();
 sg13g2_decap_8 FILLER_72_53 ();
 sg13g2_fill_1 FILLER_72_60 ();
 sg13g2_decap_4 FILLER_72_74 ();
 sg13g2_fill_1 FILLER_72_78 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_fill_2 FILLER_72_119 ();
 sg13g2_fill_1 FILLER_72_157 ();
 sg13g2_decap_4 FILLER_72_168 ();
 sg13g2_fill_2 FILLER_72_172 ();
 sg13g2_fill_2 FILLER_72_195 ();
 sg13g2_fill_1 FILLER_72_197 ();
 sg13g2_decap_8 FILLER_72_208 ();
 sg13g2_fill_2 FILLER_72_215 ();
 sg13g2_fill_1 FILLER_72_217 ();
 sg13g2_decap_4 FILLER_72_222 ();
 sg13g2_fill_2 FILLER_72_226 ();
 sg13g2_decap_8 FILLER_72_285 ();
 sg13g2_decap_4 FILLER_72_292 ();
 sg13g2_fill_2 FILLER_72_296 ();
 sg13g2_decap_4 FILLER_72_302 ();
 sg13g2_fill_1 FILLER_72_373 ();
 sg13g2_fill_2 FILLER_72_405 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_fill_2 FILLER_72_434 ();
 sg13g2_decap_8 FILLER_72_503 ();
 sg13g2_decap_8 FILLER_72_510 ();
 sg13g2_fill_2 FILLER_72_517 ();
 sg13g2_decap_4 FILLER_72_522 ();
 sg13g2_fill_1 FILLER_72_526 ();
 sg13g2_decap_8 FILLER_72_531 ();
 sg13g2_fill_2 FILLER_72_538 ();
 sg13g2_fill_1 FILLER_72_540 ();
 sg13g2_decap_8 FILLER_72_546 ();
 sg13g2_fill_1 FILLER_72_553 ();
 sg13g2_decap_8 FILLER_72_558 ();
 sg13g2_decap_4 FILLER_72_565 ();
 sg13g2_fill_1 FILLER_72_569 ();
 sg13g2_decap_8 FILLER_72_574 ();
 sg13g2_decap_8 FILLER_72_581 ();
 sg13g2_decap_8 FILLER_72_588 ();
 sg13g2_decap_4 FILLER_72_595 ();
 sg13g2_fill_2 FILLER_72_599 ();
 sg13g2_fill_2 FILLER_72_609 ();
 sg13g2_fill_1 FILLER_72_615 ();
 sg13g2_decap_8 FILLER_72_630 ();
 sg13g2_decap_8 FILLER_72_637 ();
 sg13g2_decap_8 FILLER_72_644 ();
 sg13g2_fill_1 FILLER_72_651 ();
 sg13g2_decap_8 FILLER_72_656 ();
 sg13g2_decap_8 FILLER_72_663 ();
 sg13g2_decap_4 FILLER_72_670 ();
 sg13g2_fill_1 FILLER_72_674 ();
 sg13g2_decap_8 FILLER_72_683 ();
 sg13g2_decap_8 FILLER_72_690 ();
 sg13g2_decap_4 FILLER_72_697 ();
 sg13g2_fill_1 FILLER_72_701 ();
 sg13g2_fill_1 FILLER_72_708 ();
 sg13g2_fill_1 FILLER_72_730 ();
 sg13g2_fill_1 FILLER_72_741 ();
 sg13g2_fill_2 FILLER_72_747 ();
 sg13g2_fill_2 FILLER_72_754 ();
 sg13g2_decap_4 FILLER_72_760 ();
 sg13g2_fill_2 FILLER_72_764 ();
 sg13g2_fill_1 FILLER_72_784 ();
 sg13g2_fill_1 FILLER_72_795 ();
 sg13g2_fill_2 FILLER_72_801 ();
 sg13g2_fill_1 FILLER_72_827 ();
 sg13g2_fill_1 FILLER_72_833 ();
 sg13g2_fill_1 FILLER_72_839 ();
 sg13g2_fill_2 FILLER_72_845 ();
 sg13g2_fill_1 FILLER_72_847 ();
 sg13g2_fill_2 FILLER_72_852 ();
 sg13g2_fill_1 FILLER_72_854 ();
 sg13g2_decap_4 FILLER_72_863 ();
 sg13g2_decap_8 FILLER_72_887 ();
 sg13g2_fill_2 FILLER_72_894 ();
 sg13g2_decap_4 FILLER_72_905 ();
 sg13g2_fill_2 FILLER_72_918 ();
 sg13g2_fill_1 FILLER_72_920 ();
 sg13g2_fill_1 FILLER_72_925 ();
 sg13g2_fill_1 FILLER_72_963 ();
 sg13g2_fill_2 FILLER_72_1007 ();
 sg13g2_fill_1 FILLER_72_1013 ();
 sg13g2_decap_8 FILLER_72_1087 ();
 sg13g2_decap_8 FILLER_72_1094 ();
 sg13g2_decap_8 FILLER_72_1101 ();
 sg13g2_decap_8 FILLER_72_1108 ();
 sg13g2_decap_8 FILLER_72_1115 ();
 sg13g2_decap_8 FILLER_72_1122 ();
 sg13g2_fill_1 FILLER_72_1129 ();
 sg13g2_fill_2 FILLER_72_1156 ();
 sg13g2_fill_1 FILLER_72_1158 ();
 sg13g2_decap_8 FILLER_72_1189 ();
 sg13g2_decap_8 FILLER_72_1196 ();
 sg13g2_decap_8 FILLER_72_1203 ();
 sg13g2_decap_8 FILLER_72_1210 ();
 sg13g2_decap_8 FILLER_72_1217 ();
 sg13g2_decap_8 FILLER_72_1224 ();
 sg13g2_decap_8 FILLER_72_1231 ();
 sg13g2_decap_8 FILLER_72_1238 ();
 sg13g2_decap_8 FILLER_72_1245 ();
 sg13g2_decap_8 FILLER_72_1252 ();
 sg13g2_decap_8 FILLER_72_1259 ();
 sg13g2_decap_8 FILLER_72_1266 ();
 sg13g2_decap_8 FILLER_72_1273 ();
 sg13g2_decap_8 FILLER_72_1280 ();
 sg13g2_decap_8 FILLER_72_1287 ();
 sg13g2_decap_8 FILLER_72_1294 ();
 sg13g2_decap_8 FILLER_72_1301 ();
 sg13g2_decap_8 FILLER_72_1308 ();
 sg13g2_decap_8 FILLER_72_1315 ();
 sg13g2_decap_4 FILLER_72_1322 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_fill_1 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_40 ();
 sg13g2_decap_8 FILLER_73_47 ();
 sg13g2_decap_8 FILLER_73_54 ();
 sg13g2_decap_8 FILLER_73_61 ();
 sg13g2_decap_8 FILLER_73_68 ();
 sg13g2_decap_8 FILLER_73_75 ();
 sg13g2_fill_1 FILLER_73_82 ();
 sg13g2_decap_8 FILLER_73_87 ();
 sg13g2_fill_2 FILLER_73_94 ();
 sg13g2_fill_1 FILLER_73_96 ();
 sg13g2_decap_4 FILLER_73_118 ();
 sg13g2_fill_2 FILLER_73_122 ();
 sg13g2_fill_2 FILLER_73_134 ();
 sg13g2_decap_8 FILLER_73_209 ();
 sg13g2_decap_4 FILLER_73_216 ();
 sg13g2_fill_1 FILLER_73_220 ();
 sg13g2_decap_8 FILLER_73_225 ();
 sg13g2_fill_2 FILLER_73_232 ();
 sg13g2_fill_1 FILLER_73_234 ();
 sg13g2_fill_1 FILLER_73_277 ();
 sg13g2_decap_4 FILLER_73_299 ();
 sg13g2_fill_2 FILLER_73_303 ();
 sg13g2_fill_2 FILLER_73_326 ();
 sg13g2_fill_1 FILLER_73_342 ();
 sg13g2_decap_8 FILLER_73_369 ();
 sg13g2_fill_2 FILLER_73_397 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_fill_1 FILLER_73_435 ();
 sg13g2_fill_1 FILLER_73_440 ();
 sg13g2_fill_1 FILLER_73_477 ();
 sg13g2_decap_8 FILLER_73_499 ();
 sg13g2_decap_8 FILLER_73_506 ();
 sg13g2_decap_4 FILLER_73_513 ();
 sg13g2_fill_1 FILLER_73_517 ();
 sg13g2_fill_1 FILLER_73_524 ();
 sg13g2_fill_1 FILLER_73_539 ();
 sg13g2_fill_1 FILLER_73_545 ();
 sg13g2_fill_1 FILLER_73_584 ();
 sg13g2_fill_1 FILLER_73_605 ();
 sg13g2_decap_8 FILLER_73_610 ();
 sg13g2_decap_4 FILLER_73_617 ();
 sg13g2_fill_1 FILLER_73_628 ();
 sg13g2_decap_4 FILLER_73_634 ();
 sg13g2_fill_2 FILLER_73_664 ();
 sg13g2_fill_1 FILLER_73_700 ();
 sg13g2_fill_2 FILLER_73_725 ();
 sg13g2_decap_8 FILLER_73_750 ();
 sg13g2_decap_8 FILLER_73_761 ();
 sg13g2_decap_8 FILLER_73_768 ();
 sg13g2_decap_8 FILLER_73_775 ();
 sg13g2_fill_1 FILLER_73_782 ();
 sg13g2_fill_1 FILLER_73_786 ();
 sg13g2_fill_2 FILLER_73_792 ();
 sg13g2_fill_2 FILLER_73_802 ();
 sg13g2_fill_1 FILLER_73_809 ();
 sg13g2_fill_1 FILLER_73_814 ();
 sg13g2_fill_1 FILLER_73_820 ();
 sg13g2_fill_1 FILLER_73_825 ();
 sg13g2_decap_4 FILLER_73_834 ();
 sg13g2_fill_2 FILLER_73_838 ();
 sg13g2_decap_8 FILLER_73_845 ();
 sg13g2_decap_8 FILLER_73_888 ();
 sg13g2_decap_8 FILLER_73_895 ();
 sg13g2_decap_8 FILLER_73_906 ();
 sg13g2_fill_1 FILLER_73_913 ();
 sg13g2_decap_4 FILLER_73_918 ();
 sg13g2_decap_4 FILLER_73_927 ();
 sg13g2_fill_1 FILLER_73_931 ();
 sg13g2_fill_1 FILLER_73_936 ();
 sg13g2_fill_2 FILLER_73_987 ();
 sg13g2_fill_2 FILLER_73_1028 ();
 sg13g2_fill_2 FILLER_73_1034 ();
 sg13g2_decap_8 FILLER_73_1091 ();
 sg13g2_decap_8 FILLER_73_1098 ();
 sg13g2_decap_8 FILLER_73_1105 ();
 sg13g2_decap_8 FILLER_73_1112 ();
 sg13g2_decap_8 FILLER_73_1119 ();
 sg13g2_decap_8 FILLER_73_1126 ();
 sg13g2_fill_2 FILLER_73_1137 ();
 sg13g2_fill_2 FILLER_73_1149 ();
 sg13g2_fill_1 FILLER_73_1151 ();
 sg13g2_fill_2 FILLER_73_1162 ();
 sg13g2_fill_1 FILLER_73_1164 ();
 sg13g2_fill_2 FILLER_73_1169 ();
 sg13g2_decap_8 FILLER_73_1197 ();
 sg13g2_decap_8 FILLER_73_1204 ();
 sg13g2_decap_8 FILLER_73_1211 ();
 sg13g2_decap_8 FILLER_73_1218 ();
 sg13g2_decap_8 FILLER_73_1225 ();
 sg13g2_decap_8 FILLER_73_1232 ();
 sg13g2_decap_8 FILLER_73_1239 ();
 sg13g2_decap_8 FILLER_73_1246 ();
 sg13g2_decap_8 FILLER_73_1253 ();
 sg13g2_decap_8 FILLER_73_1260 ();
 sg13g2_decap_8 FILLER_73_1267 ();
 sg13g2_decap_8 FILLER_73_1274 ();
 sg13g2_decap_8 FILLER_73_1281 ();
 sg13g2_decap_8 FILLER_73_1288 ();
 sg13g2_decap_8 FILLER_73_1295 ();
 sg13g2_decap_8 FILLER_73_1302 ();
 sg13g2_decap_8 FILLER_73_1309 ();
 sg13g2_decap_8 FILLER_73_1316 ();
 sg13g2_fill_2 FILLER_73_1323 ();
 sg13g2_fill_1 FILLER_73_1325 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_4 FILLER_74_14 ();
 sg13g2_fill_1 FILLER_74_18 ();
 sg13g2_decap_8 FILLER_74_55 ();
 sg13g2_decap_8 FILLER_74_62 ();
 sg13g2_decap_8 FILLER_74_69 ();
 sg13g2_fill_2 FILLER_74_76 ();
 sg13g2_fill_2 FILLER_74_99 ();
 sg13g2_fill_2 FILLER_74_122 ();
 sg13g2_fill_1 FILLER_74_124 ();
 sg13g2_decap_8 FILLER_74_150 ();
 sg13g2_fill_1 FILLER_74_157 ();
 sg13g2_fill_2 FILLER_74_170 ();
 sg13g2_fill_1 FILLER_74_172 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_decap_8 FILLER_74_201 ();
 sg13g2_decap_8 FILLER_74_208 ();
 sg13g2_decap_4 FILLER_74_215 ();
 sg13g2_fill_2 FILLER_74_219 ();
 sg13g2_fill_1 FILLER_74_278 ();
 sg13g2_decap_8 FILLER_74_283 ();
 sg13g2_decap_8 FILLER_74_290 ();
 sg13g2_decap_4 FILLER_74_297 ();
 sg13g2_decap_8 FILLER_74_326 ();
 sg13g2_decap_8 FILLER_74_333 ();
 sg13g2_decap_4 FILLER_74_340 ();
 sg13g2_fill_1 FILLER_74_344 ();
 sg13g2_fill_1 FILLER_74_353 ();
 sg13g2_decap_8 FILLER_74_358 ();
 sg13g2_decap_4 FILLER_74_365 ();
 sg13g2_fill_2 FILLER_74_369 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_decap_4 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_410 ();
 sg13g2_fill_1 FILLER_74_420 ();
 sg13g2_fill_1 FILLER_74_461 ();
 sg13g2_decap_4 FILLER_74_466 ();
 sg13g2_fill_1 FILLER_74_470 ();
 sg13g2_decap_8 FILLER_74_492 ();
 sg13g2_decap_8 FILLER_74_499 ();
 sg13g2_decap_4 FILLER_74_506 ();
 sg13g2_fill_1 FILLER_74_510 ();
 sg13g2_decap_4 FILLER_74_519 ();
 sg13g2_decap_8 FILLER_74_543 ();
 sg13g2_fill_2 FILLER_74_595 ();
 sg13g2_decap_8 FILLER_74_609 ();
 sg13g2_decap_8 FILLER_74_616 ();
 sg13g2_decap_8 FILLER_74_623 ();
 sg13g2_decap_8 FILLER_74_630 ();
 sg13g2_fill_1 FILLER_74_637 ();
 sg13g2_fill_1 FILLER_74_659 ();
 sg13g2_decap_8 FILLER_74_664 ();
 sg13g2_fill_2 FILLER_74_671 ();
 sg13g2_fill_1 FILLER_74_673 ();
 sg13g2_fill_1 FILLER_74_711 ();
 sg13g2_fill_1 FILLER_74_733 ();
 sg13g2_decap_8 FILLER_74_738 ();
 sg13g2_decap_8 FILLER_74_745 ();
 sg13g2_decap_8 FILLER_74_752 ();
 sg13g2_decap_8 FILLER_74_759 ();
 sg13g2_fill_2 FILLER_74_766 ();
 sg13g2_fill_2 FILLER_74_800 ();
 sg13g2_fill_1 FILLER_74_802 ();
 sg13g2_fill_1 FILLER_74_813 ();
 sg13g2_decap_8 FILLER_74_849 ();
 sg13g2_decap_4 FILLER_74_856 ();
 sg13g2_fill_1 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_74_887 ();
 sg13g2_fill_2 FILLER_74_894 ();
 sg13g2_fill_1 FILLER_74_906 ();
 sg13g2_fill_1 FILLER_74_913 ();
 sg13g2_fill_1 FILLER_74_922 ();
 sg13g2_fill_1 FILLER_74_929 ();
 sg13g2_fill_2 FILLER_74_934 ();
 sg13g2_fill_2 FILLER_74_964 ();
 sg13g2_fill_2 FILLER_74_1004 ();
 sg13g2_fill_1 FILLER_74_1006 ();
 sg13g2_decap_8 FILLER_74_1015 ();
 sg13g2_decap_8 FILLER_74_1022 ();
 sg13g2_decap_8 FILLER_74_1029 ();
 sg13g2_decap_8 FILLER_74_1036 ();
 sg13g2_decap_8 FILLER_74_1043 ();
 sg13g2_decap_4 FILLER_74_1050 ();
 sg13g2_decap_8 FILLER_74_1058 ();
 sg13g2_fill_2 FILLER_74_1078 ();
 sg13g2_decap_8 FILLER_74_1084 ();
 sg13g2_decap_8 FILLER_74_1091 ();
 sg13g2_decap_8 FILLER_74_1098 ();
 sg13g2_decap_8 FILLER_74_1105 ();
 sg13g2_decap_8 FILLER_74_1112 ();
 sg13g2_decap_8 FILLER_74_1119 ();
 sg13g2_decap_8 FILLER_74_1126 ();
 sg13g2_decap_8 FILLER_74_1133 ();
 sg13g2_decap_8 FILLER_74_1140 ();
 sg13g2_decap_8 FILLER_74_1147 ();
 sg13g2_decap_8 FILLER_74_1154 ();
 sg13g2_decap_8 FILLER_74_1161 ();
 sg13g2_decap_8 FILLER_74_1168 ();
 sg13g2_decap_8 FILLER_74_1175 ();
 sg13g2_decap_8 FILLER_74_1182 ();
 sg13g2_decap_8 FILLER_74_1189 ();
 sg13g2_decap_8 FILLER_74_1196 ();
 sg13g2_decap_8 FILLER_74_1203 ();
 sg13g2_decap_8 FILLER_74_1210 ();
 sg13g2_decap_8 FILLER_74_1217 ();
 sg13g2_decap_8 FILLER_74_1224 ();
 sg13g2_decap_8 FILLER_74_1231 ();
 sg13g2_decap_8 FILLER_74_1238 ();
 sg13g2_decap_8 FILLER_74_1245 ();
 sg13g2_decap_8 FILLER_74_1252 ();
 sg13g2_decap_8 FILLER_74_1259 ();
 sg13g2_decap_8 FILLER_74_1266 ();
 sg13g2_decap_8 FILLER_74_1273 ();
 sg13g2_decap_8 FILLER_74_1280 ();
 sg13g2_decap_8 FILLER_74_1287 ();
 sg13g2_decap_8 FILLER_74_1294 ();
 sg13g2_decap_8 FILLER_74_1301 ();
 sg13g2_decap_8 FILLER_74_1308 ();
 sg13g2_decap_8 FILLER_74_1315 ();
 sg13g2_decap_4 FILLER_74_1322 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_26 ();
 sg13g2_fill_2 FILLER_75_33 ();
 sg13g2_fill_1 FILLER_75_61 ();
 sg13g2_fill_2 FILLER_75_88 ();
 sg13g2_fill_1 FILLER_75_90 ();
 sg13g2_decap_4 FILLER_75_95 ();
 sg13g2_fill_1 FILLER_75_99 ();
 sg13g2_decap_8 FILLER_75_121 ();
 sg13g2_decap_8 FILLER_75_128 ();
 sg13g2_fill_2 FILLER_75_135 ();
 sg13g2_decap_8 FILLER_75_181 ();
 sg13g2_decap_8 FILLER_75_188 ();
 sg13g2_decap_4 FILLER_75_195 ();
 sg13g2_fill_1 FILLER_75_199 ();
 sg13g2_fill_1 FILLER_75_230 ();
 sg13g2_decap_4 FILLER_75_265 ();
 sg13g2_fill_1 FILLER_75_269 ();
 sg13g2_fill_2 FILLER_75_274 ();
 sg13g2_decap_8 FILLER_75_290 ();
 sg13g2_decap_4 FILLER_75_297 ();
 sg13g2_fill_1 FILLER_75_301 ();
 sg13g2_fill_2 FILLER_75_323 ();
 sg13g2_decap_8 FILLER_75_335 ();
 sg13g2_decap_4 FILLER_75_346 ();
 sg13g2_decap_8 FILLER_75_360 ();
 sg13g2_decap_8 FILLER_75_367 ();
 sg13g2_fill_2 FILLER_75_374 ();
 sg13g2_decap_8 FILLER_75_397 ();
 sg13g2_decap_8 FILLER_75_404 ();
 sg13g2_decap_8 FILLER_75_411 ();
 sg13g2_decap_8 FILLER_75_418 ();
 sg13g2_decap_8 FILLER_75_425 ();
 sg13g2_decap_8 FILLER_75_432 ();
 sg13g2_decap_4 FILLER_75_443 ();
 sg13g2_fill_1 FILLER_75_447 ();
 sg13g2_decap_8 FILLER_75_458 ();
 sg13g2_decap_8 FILLER_75_465 ();
 sg13g2_decap_8 FILLER_75_472 ();
 sg13g2_decap_8 FILLER_75_479 ();
 sg13g2_decap_4 FILLER_75_486 ();
 sg13g2_fill_1 FILLER_75_516 ();
 sg13g2_fill_2 FILLER_75_540 ();
 sg13g2_fill_1 FILLER_75_542 ();
 sg13g2_fill_1 FILLER_75_552 ();
 sg13g2_fill_1 FILLER_75_565 ();
 sg13g2_decap_8 FILLER_75_591 ();
 sg13g2_decap_8 FILLER_75_598 ();
 sg13g2_fill_2 FILLER_75_605 ();
 sg13g2_decap_4 FILLER_75_641 ();
 sg13g2_fill_1 FILLER_75_667 ();
 sg13g2_decap_8 FILLER_75_672 ();
 sg13g2_fill_2 FILLER_75_679 ();
 sg13g2_fill_1 FILLER_75_681 ();
 sg13g2_decap_8 FILLER_75_686 ();
 sg13g2_decap_8 FILLER_75_693 ();
 sg13g2_decap_8 FILLER_75_700 ();
 sg13g2_fill_1 FILLER_75_707 ();
 sg13g2_fill_1 FILLER_75_728 ();
 sg13g2_fill_1 FILLER_75_739 ();
 sg13g2_fill_2 FILLER_75_744 ();
 sg13g2_decap_8 FILLER_75_755 ();
 sg13g2_decap_4 FILLER_75_762 ();
 sg13g2_fill_2 FILLER_75_766 ();
 sg13g2_fill_1 FILLER_75_773 ();
 sg13g2_fill_2 FILLER_75_778 ();
 sg13g2_fill_1 FILLER_75_785 ();
 sg13g2_fill_1 FILLER_75_791 ();
 sg13g2_fill_2 FILLER_75_796 ();
 sg13g2_fill_1 FILLER_75_848 ();
 sg13g2_fill_1 FILLER_75_853 ();
 sg13g2_fill_1 FILLER_75_858 ();
 sg13g2_fill_1 FILLER_75_885 ();
 sg13g2_decap_8 FILLER_75_912 ();
 sg13g2_fill_2 FILLER_75_919 ();
 sg13g2_fill_1 FILLER_75_921 ();
 sg13g2_decap_8 FILLER_75_958 ();
 sg13g2_decap_8 FILLER_75_965 ();
 sg13g2_decap_8 FILLER_75_972 ();
 sg13g2_fill_1 FILLER_75_979 ();
 sg13g2_decap_8 FILLER_75_996 ();
 sg13g2_decap_8 FILLER_75_1008 ();
 sg13g2_decap_8 FILLER_75_1015 ();
 sg13g2_decap_8 FILLER_75_1022 ();
 sg13g2_decap_8 FILLER_75_1029 ();
 sg13g2_decap_4 FILLER_75_1036 ();
 sg13g2_fill_1 FILLER_75_1046 ();
 sg13g2_fill_2 FILLER_75_1051 ();
 sg13g2_fill_1 FILLER_75_1062 ();
 sg13g2_decap_8 FILLER_75_1068 ();
 sg13g2_decap_8 FILLER_75_1075 ();
 sg13g2_decap_8 FILLER_75_1082 ();
 sg13g2_decap_8 FILLER_75_1089 ();
 sg13g2_decap_8 FILLER_75_1096 ();
 sg13g2_decap_8 FILLER_75_1103 ();
 sg13g2_decap_8 FILLER_75_1110 ();
 sg13g2_decap_8 FILLER_75_1117 ();
 sg13g2_decap_8 FILLER_75_1124 ();
 sg13g2_decap_8 FILLER_75_1131 ();
 sg13g2_decap_8 FILLER_75_1138 ();
 sg13g2_decap_8 FILLER_75_1145 ();
 sg13g2_decap_8 FILLER_75_1152 ();
 sg13g2_decap_8 FILLER_75_1159 ();
 sg13g2_decap_8 FILLER_75_1166 ();
 sg13g2_decap_8 FILLER_75_1173 ();
 sg13g2_decap_8 FILLER_75_1180 ();
 sg13g2_decap_8 FILLER_75_1187 ();
 sg13g2_decap_8 FILLER_75_1194 ();
 sg13g2_decap_8 FILLER_75_1201 ();
 sg13g2_decap_8 FILLER_75_1208 ();
 sg13g2_decap_8 FILLER_75_1215 ();
 sg13g2_decap_8 FILLER_75_1222 ();
 sg13g2_decap_8 FILLER_75_1229 ();
 sg13g2_decap_8 FILLER_75_1236 ();
 sg13g2_decap_8 FILLER_75_1243 ();
 sg13g2_decap_8 FILLER_75_1250 ();
 sg13g2_decap_8 FILLER_75_1257 ();
 sg13g2_decap_8 FILLER_75_1264 ();
 sg13g2_decap_8 FILLER_75_1271 ();
 sg13g2_decap_8 FILLER_75_1278 ();
 sg13g2_decap_8 FILLER_75_1285 ();
 sg13g2_decap_8 FILLER_75_1292 ();
 sg13g2_decap_8 FILLER_75_1299 ();
 sg13g2_decap_8 FILLER_75_1306 ();
 sg13g2_decap_8 FILLER_75_1313 ();
 sg13g2_decap_4 FILLER_75_1320 ();
 sg13g2_fill_2 FILLER_75_1324 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_fill_2 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_30 ();
 sg13g2_decap_4 FILLER_76_49 ();
 sg13g2_fill_1 FILLER_76_53 ();
 sg13g2_fill_1 FILLER_76_94 ();
 sg13g2_decap_8 FILLER_76_116 ();
 sg13g2_decap_8 FILLER_76_123 ();
 sg13g2_decap_8 FILLER_76_130 ();
 sg13g2_fill_1 FILLER_76_137 ();
 sg13g2_decap_8 FILLER_76_142 ();
 sg13g2_fill_2 FILLER_76_149 ();
 sg13g2_decap_4 FILLER_76_155 ();
 sg13g2_fill_2 FILLER_76_163 ();
 sg13g2_fill_1 FILLER_76_165 ();
 sg13g2_decap_4 FILLER_76_170 ();
 sg13g2_decap_4 FILLER_76_203 ();
 sg13g2_fill_2 FILLER_76_207 ();
 sg13g2_decap_8 FILLER_76_248 ();
 sg13g2_decap_8 FILLER_76_255 ();
 sg13g2_decap_4 FILLER_76_262 ();
 sg13g2_fill_2 FILLER_76_278 ();
 sg13g2_decap_8 FILLER_76_335 ();
 sg13g2_decap_8 FILLER_76_342 ();
 sg13g2_decap_4 FILLER_76_349 ();
 sg13g2_fill_1 FILLER_76_353 ();
 sg13g2_fill_1 FILLER_76_358 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_fill_1 FILLER_76_409 ();
 sg13g2_fill_2 FILLER_76_418 ();
 sg13g2_decap_4 FILLER_76_424 ();
 sg13g2_fill_1 FILLER_76_428 ();
 sg13g2_decap_4 FILLER_76_436 ();
 sg13g2_decap_8 FILLER_76_487 ();
 sg13g2_fill_1 FILLER_76_494 ();
 sg13g2_decap_8 FILLER_76_499 ();
 sg13g2_fill_1 FILLER_76_519 ();
 sg13g2_fill_2 FILLER_76_525 ();
 sg13g2_fill_2 FILLER_76_532 ();
 sg13g2_decap_4 FILLER_76_548 ();
 sg13g2_fill_1 FILLER_76_552 ();
 sg13g2_fill_1 FILLER_76_561 ();
 sg13g2_fill_2 FILLER_76_566 ();
 sg13g2_fill_1 FILLER_76_572 ();
 sg13g2_fill_2 FILLER_76_577 ();
 sg13g2_decap_4 FILLER_76_583 ();
 sg13g2_fill_1 FILLER_76_587 ();
 sg13g2_fill_1 FILLER_76_592 ();
 sg13g2_fill_1 FILLER_76_619 ();
 sg13g2_fill_1 FILLER_76_650 ();
 sg13g2_fill_1 FILLER_76_664 ();
 sg13g2_decap_8 FILLER_76_671 ();
 sg13g2_decap_8 FILLER_76_678 ();
 sg13g2_decap_8 FILLER_76_685 ();
 sg13g2_decap_8 FILLER_76_692 ();
 sg13g2_decap_4 FILLER_76_699 ();
 sg13g2_fill_2 FILLER_76_703 ();
 sg13g2_fill_1 FILLER_76_728 ();
 sg13g2_fill_1 FILLER_76_733 ();
 sg13g2_fill_1 FILLER_76_764 ();
 sg13g2_fill_1 FILLER_76_786 ();
 sg13g2_decap_8 FILLER_76_805 ();
 sg13g2_fill_2 FILLER_76_812 ();
 sg13g2_fill_1 FILLER_76_814 ();
 sg13g2_decap_8 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_834 ();
 sg13g2_decap_8 FILLER_76_841 ();
 sg13g2_decap_4 FILLER_76_848 ();
 sg13g2_fill_2 FILLER_76_852 ();
 sg13g2_decap_8 FILLER_76_871 ();
 sg13g2_decap_4 FILLER_76_878 ();
 sg13g2_fill_2 FILLER_76_882 ();
 sg13g2_decap_4 FILLER_76_888 ();
 sg13g2_decap_4 FILLER_76_896 ();
 sg13g2_fill_2 FILLER_76_900 ();
 sg13g2_fill_1 FILLER_76_906 ();
 sg13g2_fill_2 FILLER_76_917 ();
 sg13g2_decap_8 FILLER_76_927 ();
 sg13g2_decap_8 FILLER_76_938 ();
 sg13g2_fill_1 FILLER_76_945 ();
 sg13g2_decap_8 FILLER_76_950 ();
 sg13g2_decap_8 FILLER_76_957 ();
 sg13g2_decap_8 FILLER_76_964 ();
 sg13g2_decap_4 FILLER_76_971 ();
 sg13g2_decap_8 FILLER_76_985 ();
 sg13g2_decap_4 FILLER_76_992 ();
 sg13g2_fill_2 FILLER_76_996 ();
 sg13g2_fill_1 FILLER_76_1001 ();
 sg13g2_fill_1 FILLER_76_1007 ();
 sg13g2_fill_1 FILLER_76_1034 ();
 sg13g2_fill_2 FILLER_76_1065 ();
 sg13g2_decap_8 FILLER_76_1093 ();
 sg13g2_decap_8 FILLER_76_1100 ();
 sg13g2_decap_8 FILLER_76_1107 ();
 sg13g2_decap_8 FILLER_76_1114 ();
 sg13g2_decap_8 FILLER_76_1121 ();
 sg13g2_decap_8 FILLER_76_1128 ();
 sg13g2_decap_8 FILLER_76_1135 ();
 sg13g2_decap_8 FILLER_76_1142 ();
 sg13g2_decap_8 FILLER_76_1149 ();
 sg13g2_decap_8 FILLER_76_1156 ();
 sg13g2_decap_8 FILLER_76_1163 ();
 sg13g2_decap_8 FILLER_76_1170 ();
 sg13g2_decap_8 FILLER_76_1177 ();
 sg13g2_decap_8 FILLER_76_1184 ();
 sg13g2_decap_8 FILLER_76_1191 ();
 sg13g2_decap_8 FILLER_76_1198 ();
 sg13g2_decap_8 FILLER_76_1205 ();
 sg13g2_decap_8 FILLER_76_1212 ();
 sg13g2_decap_8 FILLER_76_1219 ();
 sg13g2_decap_8 FILLER_76_1226 ();
 sg13g2_decap_8 FILLER_76_1233 ();
 sg13g2_decap_8 FILLER_76_1240 ();
 sg13g2_decap_8 FILLER_76_1247 ();
 sg13g2_decap_8 FILLER_76_1254 ();
 sg13g2_decap_8 FILLER_76_1261 ();
 sg13g2_decap_8 FILLER_76_1268 ();
 sg13g2_decap_8 FILLER_76_1275 ();
 sg13g2_decap_8 FILLER_76_1282 ();
 sg13g2_decap_8 FILLER_76_1289 ();
 sg13g2_decap_8 FILLER_76_1296 ();
 sg13g2_decap_8 FILLER_76_1303 ();
 sg13g2_decap_8 FILLER_76_1310 ();
 sg13g2_decap_8 FILLER_76_1317 ();
 sg13g2_fill_2 FILLER_76_1324 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_4 FILLER_77_49 ();
 sg13g2_fill_1 FILLER_77_53 ();
 sg13g2_fill_1 FILLER_77_68 ();
 sg13g2_decap_8 FILLER_77_121 ();
 sg13g2_decap_8 FILLER_77_128 ();
 sg13g2_decap_4 FILLER_77_135 ();
 sg13g2_fill_2 FILLER_77_139 ();
 sg13g2_fill_1 FILLER_77_197 ();
 sg13g2_decap_8 FILLER_77_204 ();
 sg13g2_fill_2 FILLER_77_211 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_fill_1 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_249 ();
 sg13g2_decap_8 FILLER_77_256 ();
 sg13g2_fill_2 FILLER_77_263 ();
 sg13g2_fill_1 FILLER_77_265 ();
 sg13g2_fill_2 FILLER_77_312 ();
 sg13g2_fill_1 FILLER_77_314 ();
 sg13g2_fill_1 FILLER_77_375 ();
 sg13g2_fill_2 FILLER_77_384 ();
 sg13g2_fill_1 FILLER_77_386 ();
 sg13g2_fill_1 FILLER_77_396 ();
 sg13g2_decap_4 FILLER_77_453 ();
 sg13g2_fill_1 FILLER_77_457 ();
 sg13g2_decap_8 FILLER_77_466 ();
 sg13g2_decap_8 FILLER_77_473 ();
 sg13g2_decap_8 FILLER_77_480 ();
 sg13g2_decap_8 FILLER_77_487 ();
 sg13g2_decap_8 FILLER_77_494 ();
 sg13g2_fill_2 FILLER_77_501 ();
 sg13g2_fill_1 FILLER_77_503 ();
 sg13g2_decap_4 FILLER_77_509 ();
 sg13g2_fill_2 FILLER_77_513 ();
 sg13g2_fill_1 FILLER_77_529 ();
 sg13g2_decap_4 FILLER_77_558 ();
 sg13g2_fill_2 FILLER_77_587 ();
 sg13g2_fill_1 FILLER_77_619 ();
 sg13g2_decap_8 FILLER_77_625 ();
 sg13g2_fill_1 FILLER_77_632 ();
 sg13g2_fill_1 FILLER_77_637 ();
 sg13g2_decap_8 FILLER_77_642 ();
 sg13g2_decap_8 FILLER_77_669 ();
 sg13g2_decap_8 FILLER_77_676 ();
 sg13g2_decap_8 FILLER_77_683 ();
 sg13g2_decap_8 FILLER_77_690 ();
 sg13g2_decap_4 FILLER_77_697 ();
 sg13g2_fill_2 FILLER_77_701 ();
 sg13g2_fill_1 FILLER_77_723 ();
 sg13g2_fill_1 FILLER_77_729 ();
 sg13g2_fill_1 FILLER_77_756 ();
 sg13g2_fill_1 FILLER_77_762 ();
 sg13g2_fill_1 FILLER_77_777 ();
 sg13g2_fill_1 FILLER_77_801 ();
 sg13g2_decap_8 FILLER_77_827 ();
 sg13g2_fill_2 FILLER_77_834 ();
 sg13g2_decap_8 FILLER_77_885 ();
 sg13g2_fill_1 FILLER_77_892 ();
 sg13g2_fill_1 FILLER_77_909 ();
 sg13g2_fill_1 FILLER_77_918 ();
 sg13g2_fill_2 FILLER_77_923 ();
 sg13g2_fill_1 FILLER_77_929 ();
 sg13g2_decap_4 FILLER_77_942 ();
 sg13g2_fill_2 FILLER_77_946 ();
 sg13g2_decap_4 FILLER_77_952 ();
 sg13g2_fill_2 FILLER_77_956 ();
 sg13g2_fill_1 FILLER_77_962 ();
 sg13g2_fill_1 FILLER_77_1012 ();
 sg13g2_fill_1 FILLER_77_1026 ();
 sg13g2_fill_2 FILLER_77_1066 ();
 sg13g2_decap_8 FILLER_77_1081 ();
 sg13g2_decap_8 FILLER_77_1088 ();
 sg13g2_decap_8 FILLER_77_1095 ();
 sg13g2_decap_8 FILLER_77_1102 ();
 sg13g2_decap_8 FILLER_77_1109 ();
 sg13g2_decap_8 FILLER_77_1116 ();
 sg13g2_decap_8 FILLER_77_1123 ();
 sg13g2_decap_8 FILLER_77_1130 ();
 sg13g2_decap_8 FILLER_77_1137 ();
 sg13g2_decap_8 FILLER_77_1144 ();
 sg13g2_decap_8 FILLER_77_1151 ();
 sg13g2_decap_8 FILLER_77_1158 ();
 sg13g2_decap_8 FILLER_77_1165 ();
 sg13g2_decap_8 FILLER_77_1172 ();
 sg13g2_decap_8 FILLER_77_1179 ();
 sg13g2_decap_8 FILLER_77_1186 ();
 sg13g2_decap_8 FILLER_77_1193 ();
 sg13g2_decap_8 FILLER_77_1200 ();
 sg13g2_decap_8 FILLER_77_1207 ();
 sg13g2_decap_8 FILLER_77_1214 ();
 sg13g2_decap_8 FILLER_77_1221 ();
 sg13g2_decap_8 FILLER_77_1228 ();
 sg13g2_decap_8 FILLER_77_1235 ();
 sg13g2_decap_8 FILLER_77_1242 ();
 sg13g2_decap_8 FILLER_77_1249 ();
 sg13g2_decap_8 FILLER_77_1256 ();
 sg13g2_decap_8 FILLER_77_1263 ();
 sg13g2_decap_8 FILLER_77_1270 ();
 sg13g2_decap_8 FILLER_77_1277 ();
 sg13g2_decap_8 FILLER_77_1284 ();
 sg13g2_decap_8 FILLER_77_1291 ();
 sg13g2_decap_8 FILLER_77_1298 ();
 sg13g2_decap_8 FILLER_77_1305 ();
 sg13g2_decap_8 FILLER_77_1312 ();
 sg13g2_decap_8 FILLER_77_1319 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_fill_2 FILLER_78_70 ();
 sg13g2_fill_1 FILLER_78_72 ();
 sg13g2_fill_1 FILLER_78_77 ();
 sg13g2_decap_4 FILLER_78_119 ();
 sg13g2_fill_1 FILLER_78_123 ();
 sg13g2_fill_2 FILLER_78_128 ();
 sg13g2_fill_1 FILLER_78_130 ();
 sg13g2_fill_2 FILLER_78_135 ();
 sg13g2_fill_1 FILLER_78_137 ();
 sg13g2_decap_8 FILLER_78_263 ();
 sg13g2_decap_8 FILLER_78_270 ();
 sg13g2_decap_4 FILLER_78_354 ();
 sg13g2_fill_1 FILLER_78_368 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_decap_4 FILLER_78_402 ();
 sg13g2_fill_1 FILLER_78_456 ();
 sg13g2_decap_8 FILLER_78_487 ();
 sg13g2_fill_2 FILLER_78_494 ();
 sg13g2_decap_8 FILLER_78_500 ();
 sg13g2_fill_2 FILLER_78_507 ();
 sg13g2_fill_1 FILLER_78_509 ();
 sg13g2_fill_2 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_551 ();
 sg13g2_decap_4 FILLER_78_558 ();
 sg13g2_fill_2 FILLER_78_568 ();
 sg13g2_fill_1 FILLER_78_596 ();
 sg13g2_decap_8 FILLER_78_626 ();
 sg13g2_fill_2 FILLER_78_633 ();
 sg13g2_decap_8 FILLER_78_661 ();
 sg13g2_decap_8 FILLER_78_668 ();
 sg13g2_decap_8 FILLER_78_675 ();
 sg13g2_decap_8 FILLER_78_682 ();
 sg13g2_decap_4 FILLER_78_689 ();
 sg13g2_fill_1 FILLER_78_727 ();
 sg13g2_fill_2 FILLER_78_737 ();
 sg13g2_decap_8 FILLER_78_743 ();
 sg13g2_fill_2 FILLER_78_750 ();
 sg13g2_fill_1 FILLER_78_756 ();
 sg13g2_fill_2 FILLER_78_782 ();
 sg13g2_fill_2 FILLER_78_793 ();
 sg13g2_fill_1 FILLER_78_800 ();
 sg13g2_fill_1 FILLER_78_806 ();
 sg13g2_fill_2 FILLER_78_845 ();
 sg13g2_decap_4 FILLER_78_885 ();
 sg13g2_fill_1 FILLER_78_889 ();
 sg13g2_fill_1 FILLER_78_921 ();
 sg13g2_fill_2 FILLER_78_986 ();
 sg13g2_fill_1 FILLER_78_1027 ();
 sg13g2_decap_8 FILLER_78_1066 ();
 sg13g2_decap_8 FILLER_78_1073 ();
 sg13g2_decap_8 FILLER_78_1080 ();
 sg13g2_decap_8 FILLER_78_1087 ();
 sg13g2_decap_8 FILLER_78_1094 ();
 sg13g2_decap_8 FILLER_78_1101 ();
 sg13g2_decap_8 FILLER_78_1108 ();
 sg13g2_decap_8 FILLER_78_1115 ();
 sg13g2_decap_8 FILLER_78_1122 ();
 sg13g2_decap_8 FILLER_78_1129 ();
 sg13g2_decap_8 FILLER_78_1136 ();
 sg13g2_decap_8 FILLER_78_1143 ();
 sg13g2_decap_8 FILLER_78_1150 ();
 sg13g2_decap_8 FILLER_78_1157 ();
 sg13g2_decap_8 FILLER_78_1164 ();
 sg13g2_decap_8 FILLER_78_1171 ();
 sg13g2_decap_8 FILLER_78_1178 ();
 sg13g2_decap_8 FILLER_78_1185 ();
 sg13g2_decap_8 FILLER_78_1192 ();
 sg13g2_decap_8 FILLER_78_1199 ();
 sg13g2_decap_8 FILLER_78_1206 ();
 sg13g2_decap_8 FILLER_78_1213 ();
 sg13g2_decap_8 FILLER_78_1220 ();
 sg13g2_decap_8 FILLER_78_1227 ();
 sg13g2_decap_8 FILLER_78_1234 ();
 sg13g2_decap_8 FILLER_78_1241 ();
 sg13g2_decap_8 FILLER_78_1248 ();
 sg13g2_decap_8 FILLER_78_1255 ();
 sg13g2_decap_8 FILLER_78_1262 ();
 sg13g2_decap_8 FILLER_78_1269 ();
 sg13g2_decap_8 FILLER_78_1276 ();
 sg13g2_decap_8 FILLER_78_1283 ();
 sg13g2_decap_8 FILLER_78_1290 ();
 sg13g2_decap_8 FILLER_78_1297 ();
 sg13g2_decap_8 FILLER_78_1304 ();
 sg13g2_decap_8 FILLER_78_1311 ();
 sg13g2_decap_8 FILLER_78_1318 ();
 sg13g2_fill_1 FILLER_78_1325 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_4 FILLER_79_84 ();
 sg13g2_fill_2 FILLER_79_92 ();
 sg13g2_fill_1 FILLER_79_94 ();
 sg13g2_fill_2 FILLER_79_99 ();
 sg13g2_fill_1 FILLER_79_167 ();
 sg13g2_fill_1 FILLER_79_178 ();
 sg13g2_fill_1 FILLER_79_183 ();
 sg13g2_fill_2 FILLER_79_188 ();
 sg13g2_fill_2 FILLER_79_211 ();
 sg13g2_fill_1 FILLER_79_223 ();
 sg13g2_fill_1 FILLER_79_228 ();
 sg13g2_decap_4 FILLER_79_272 ();
 sg13g2_fill_2 FILLER_79_276 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_fill_1 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_341 ();
 sg13g2_decap_4 FILLER_79_348 ();
 sg13g2_fill_1 FILLER_79_362 ();
 sg13g2_fill_2 FILLER_79_397 ();
 sg13g2_fill_1 FILLER_79_399 ();
 sg13g2_fill_2 FILLER_79_440 ();
 sg13g2_decap_4 FILLER_79_446 ();
 sg13g2_decap_8 FILLER_79_460 ();
 sg13g2_fill_2 FILLER_79_467 ();
 sg13g2_decap_8 FILLER_79_473 ();
 sg13g2_decap_8 FILLER_79_480 ();
 sg13g2_fill_2 FILLER_79_487 ();
 sg13g2_fill_1 FILLER_79_489 ();
 sg13g2_decap_4 FILLER_79_516 ();
 sg13g2_fill_1 FILLER_79_520 ();
 sg13g2_decap_8 FILLER_79_530 ();
 sg13g2_fill_2 FILLER_79_537 ();
 sg13g2_decap_8 FILLER_79_599 ();
 sg13g2_decap_8 FILLER_79_606 ();
 sg13g2_decap_8 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_654 ();
 sg13g2_decap_8 FILLER_79_661 ();
 sg13g2_decap_8 FILLER_79_668 ();
 sg13g2_decap_8 FILLER_79_675 ();
 sg13g2_decap_8 FILLER_79_682 ();
 sg13g2_decap_8 FILLER_79_689 ();
 sg13g2_decap_4 FILLER_79_696 ();
 sg13g2_fill_1 FILLER_79_700 ();
 sg13g2_fill_2 FILLER_79_705 ();
 sg13g2_fill_1 FILLER_79_707 ();
 sg13g2_fill_2 FILLER_79_734 ();
 sg13g2_fill_1 FILLER_79_736 ();
 sg13g2_fill_1 FILLER_79_794 ();
 sg13g2_fill_2 FILLER_79_859 ();
 sg13g2_fill_2 FILLER_79_874 ();
 sg13g2_fill_1 FILLER_79_876 ();
 sg13g2_decap_8 FILLER_79_882 ();
 sg13g2_decap_8 FILLER_79_919 ();
 sg13g2_decap_8 FILLER_79_926 ();
 sg13g2_decap_4 FILLER_79_933 ();
 sg13g2_fill_1 FILLER_79_1040 ();
 sg13g2_decap_8 FILLER_79_1067 ();
 sg13g2_decap_8 FILLER_79_1074 ();
 sg13g2_decap_8 FILLER_79_1081 ();
 sg13g2_decap_8 FILLER_79_1088 ();
 sg13g2_decap_8 FILLER_79_1095 ();
 sg13g2_decap_8 FILLER_79_1102 ();
 sg13g2_decap_8 FILLER_79_1109 ();
 sg13g2_decap_8 FILLER_79_1116 ();
 sg13g2_decap_8 FILLER_79_1123 ();
 sg13g2_decap_8 FILLER_79_1130 ();
 sg13g2_decap_8 FILLER_79_1137 ();
 sg13g2_decap_8 FILLER_79_1144 ();
 sg13g2_decap_8 FILLER_79_1151 ();
 sg13g2_decap_8 FILLER_79_1158 ();
 sg13g2_decap_8 FILLER_79_1165 ();
 sg13g2_decap_8 FILLER_79_1172 ();
 sg13g2_decap_8 FILLER_79_1179 ();
 sg13g2_decap_8 FILLER_79_1186 ();
 sg13g2_decap_8 FILLER_79_1193 ();
 sg13g2_decap_8 FILLER_79_1200 ();
 sg13g2_decap_8 FILLER_79_1207 ();
 sg13g2_decap_8 FILLER_79_1214 ();
 sg13g2_decap_8 FILLER_79_1221 ();
 sg13g2_decap_8 FILLER_79_1228 ();
 sg13g2_decap_8 FILLER_79_1235 ();
 sg13g2_decap_8 FILLER_79_1242 ();
 sg13g2_decap_8 FILLER_79_1249 ();
 sg13g2_decap_8 FILLER_79_1256 ();
 sg13g2_decap_8 FILLER_79_1263 ();
 sg13g2_decap_8 FILLER_79_1270 ();
 sg13g2_decap_8 FILLER_79_1277 ();
 sg13g2_decap_8 FILLER_79_1284 ();
 sg13g2_decap_8 FILLER_79_1291 ();
 sg13g2_decap_8 FILLER_79_1298 ();
 sg13g2_decap_8 FILLER_79_1305 ();
 sg13g2_decap_8 FILLER_79_1312 ();
 sg13g2_decap_8 FILLER_79_1319 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_fill_2 FILLER_80_80 ();
 sg13g2_fill_1 FILLER_80_82 ();
 sg13g2_fill_1 FILLER_80_91 ();
 sg13g2_fill_2 FILLER_80_96 ();
 sg13g2_fill_2 FILLER_80_102 ();
 sg13g2_fill_2 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_118 ();
 sg13g2_fill_2 FILLER_80_122 ();
 sg13g2_decap_8 FILLER_80_132 ();
 sg13g2_fill_1 FILLER_80_155 ();
 sg13g2_fill_1 FILLER_80_164 ();
 sg13g2_fill_2 FILLER_80_173 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_decap_4 FILLER_80_184 ();
 sg13g2_fill_2 FILLER_80_188 ();
 sg13g2_fill_1 FILLER_80_241 ();
 sg13g2_fill_1 FILLER_80_246 ();
 sg13g2_fill_1 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_260 ();
 sg13g2_decap_8 FILLER_80_267 ();
 sg13g2_decap_8 FILLER_80_274 ();
 sg13g2_decap_8 FILLER_80_281 ();
 sg13g2_fill_1 FILLER_80_288 ();
 sg13g2_decap_8 FILLER_80_293 ();
 sg13g2_decap_8 FILLER_80_304 ();
 sg13g2_decap_8 FILLER_80_311 ();
 sg13g2_decap_8 FILLER_80_318 ();
 sg13g2_decap_8 FILLER_80_325 ();
 sg13g2_decap_8 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_339 ();
 sg13g2_decap_8 FILLER_80_346 ();
 sg13g2_decap_4 FILLER_80_353 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_decap_4 FILLER_80_398 ();
 sg13g2_fill_2 FILLER_80_402 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_fill_1 FILLER_80_415 ();
 sg13g2_decap_8 FILLER_80_424 ();
 sg13g2_decap_8 FILLER_80_431 ();
 sg13g2_decap_8 FILLER_80_438 ();
 sg13g2_decap_8 FILLER_80_445 ();
 sg13g2_decap_8 FILLER_80_452 ();
 sg13g2_decap_8 FILLER_80_459 ();
 sg13g2_decap_8 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_473 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_fill_1 FILLER_80_529 ();
 sg13g2_fill_2 FILLER_80_534 ();
 sg13g2_decap_8 FILLER_80_562 ();
 sg13g2_decap_8 FILLER_80_569 ();
 sg13g2_decap_4 FILLER_80_576 ();
 sg13g2_decap_8 FILLER_80_584 ();
 sg13g2_decap_8 FILLER_80_591 ();
 sg13g2_decap_8 FILLER_80_598 ();
 sg13g2_fill_1 FILLER_80_605 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_4 FILLER_80_711 ();
 sg13g2_fill_2 FILLER_80_715 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_fill_2 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_748 ();
 sg13g2_decap_8 FILLER_80_755 ();
 sg13g2_decap_8 FILLER_80_762 ();
 sg13g2_fill_1 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_774 ();
 sg13g2_decap_4 FILLER_80_784 ();
 sg13g2_fill_1 FILLER_80_788 ();
 sg13g2_decap_8 FILLER_80_792 ();
 sg13g2_decap_4 FILLER_80_799 ();
 sg13g2_fill_2 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_4 FILLER_80_830 ();
 sg13g2_fill_2 FILLER_80_834 ();
 sg13g2_fill_2 FILLER_80_840 ();
 sg13g2_fill_1 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_856 ();
 sg13g2_decap_8 FILLER_80_863 ();
 sg13g2_decap_8 FILLER_80_870 ();
 sg13g2_decap_8 FILLER_80_877 ();
 sg13g2_decap_8 FILLER_80_884 ();
 sg13g2_decap_8 FILLER_80_891 ();
 sg13g2_decap_8 FILLER_80_906 ();
 sg13g2_decap_8 FILLER_80_913 ();
 sg13g2_decap_8 FILLER_80_920 ();
 sg13g2_decap_8 FILLER_80_927 ();
 sg13g2_decap_8 FILLER_80_934 ();
 sg13g2_decap_8 FILLER_80_941 ();
 sg13g2_fill_1 FILLER_80_948 ();
 sg13g2_fill_2 FILLER_80_953 ();
 sg13g2_decap_8 FILLER_80_959 ();
 sg13g2_decap_8 FILLER_80_966 ();
 sg13g2_decap_8 FILLER_80_981 ();
 sg13g2_decap_8 FILLER_80_988 ();
 sg13g2_decap_4 FILLER_80_995 ();
 sg13g2_decap_8 FILLER_80_1003 ();
 sg13g2_decap_8 FILLER_80_1014 ();
 sg13g2_decap_8 FILLER_80_1021 ();
 sg13g2_decap_8 FILLER_80_1028 ();
 sg13g2_fill_2 FILLER_80_1035 ();
 sg13g2_fill_1 FILLER_80_1049 ();
 sg13g2_decap_8 FILLER_80_1054 ();
 sg13g2_decap_8 FILLER_80_1061 ();
 sg13g2_decap_8 FILLER_80_1068 ();
 sg13g2_decap_8 FILLER_80_1075 ();
 sg13g2_decap_8 FILLER_80_1082 ();
 sg13g2_decap_8 FILLER_80_1089 ();
 sg13g2_decap_8 FILLER_80_1096 ();
 sg13g2_decap_8 FILLER_80_1103 ();
 sg13g2_decap_8 FILLER_80_1110 ();
 sg13g2_decap_8 FILLER_80_1117 ();
 sg13g2_decap_8 FILLER_80_1124 ();
 sg13g2_decap_8 FILLER_80_1131 ();
 sg13g2_decap_8 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_decap_8 FILLER_80_1152 ();
 sg13g2_decap_8 FILLER_80_1159 ();
 sg13g2_decap_8 FILLER_80_1166 ();
 sg13g2_decap_8 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_decap_8 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1201 ();
 sg13g2_decap_8 FILLER_80_1208 ();
 sg13g2_decap_8 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1222 ();
 sg13g2_decap_8 FILLER_80_1229 ();
 sg13g2_decap_8 FILLER_80_1236 ();
 sg13g2_decap_8 FILLER_80_1243 ();
 sg13g2_decap_8 FILLER_80_1250 ();
 sg13g2_decap_8 FILLER_80_1257 ();
 sg13g2_decap_8 FILLER_80_1264 ();
 sg13g2_decap_8 FILLER_80_1271 ();
 sg13g2_decap_8 FILLER_80_1278 ();
 sg13g2_decap_8 FILLER_80_1285 ();
 sg13g2_decap_8 FILLER_80_1292 ();
 sg13g2_decap_8 FILLER_80_1299 ();
 sg13g2_decap_8 FILLER_80_1306 ();
 sg13g2_decap_8 FILLER_80_1313 ();
 sg13g2_decap_4 FILLER_80_1320 ();
 sg13g2_fill_2 FILLER_80_1324 ();
endmodule
