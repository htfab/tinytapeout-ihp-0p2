module tt_um_NicklausThompson_SkyKing (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire BNC_trig;
 wire \BNC_x[0] ;
 wire \BNC_x[1] ;
 wire \BNC_x[2] ;
 wire \BNC_x[3] ;
 wire \BNC_x[4] ;
 wire \BNC_x[5] ;
 wire \BNC_x[6] ;
 wire \BNC_x[7] ;
 wire \BNC_y[0] ;
 wire \BNC_y[1] ;
 wire \BNC_y[2] ;
 wire \BNC_y[3] ;
 wire \BNC_y[4] ;
 wire \BNC_y[5] ;
 wire \BNC_y[6] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire clknet_0_clk;
 wire \bnc_image_generator.counter[0] ;
 wire \bnc_image_generator.counter[1] ;
 wire \bnc_image_generator.counter[2] ;
 wire \bnc_image_generator.counter[4] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \vga_image_generator.character_hold[0] ;
 wire \vga_image_generator.character_hold[10] ;
 wire \vga_image_generator.character_hold[11] ;
 wire \vga_image_generator.character_hold[12] ;
 wire \vga_image_generator.character_hold[13] ;
 wire \vga_image_generator.character_hold[14] ;
 wire \vga_image_generator.character_hold[15] ;
 wire \vga_image_generator.character_hold[16] ;
 wire \vga_image_generator.character_hold[17] ;
 wire \vga_image_generator.character_hold[1] ;
 wire \vga_image_generator.character_hold[2] ;
 wire \vga_image_generator.character_hold[3] ;
 wire \vga_image_generator.character_hold[4] ;
 wire \vga_image_generator.character_hold[5] ;
 wire \vga_image_generator.character_hold[6] ;
 wire \vga_image_generator.character_hold[7] ;
 wire \vga_image_generator.character_hold[8] ;
 wire \vga_image_generator.character_hold[9] ;
 wire \vga_image_generator.counter[0] ;
 wire \vga_image_generator.counter[10] ;
 wire \vga_image_generator.counter[11] ;
 wire \vga_image_generator.counter[12] ;
 wire \vga_image_generator.counter[13] ;
 wire \vga_image_generator.counter[14] ;
 wire \vga_image_generator.counter[15] ;
 wire \vga_image_generator.counter[16] ;
 wire \vga_image_generator.counter[17] ;
 wire \vga_image_generator.counter[18] ;
 wire \vga_image_generator.counter[19] ;
 wire \vga_image_generator.counter[1] ;
 wire \vga_image_generator.counter[20] ;
 wire \vga_image_generator.counter[21] ;
 wire \vga_image_generator.counter[22] ;
 wire \vga_image_generator.counter[23] ;
 wire \vga_image_generator.counter[24] ;
 wire \vga_image_generator.counter[25] ;
 wire \vga_image_generator.counter[26] ;
 wire \vga_image_generator.counter[27] ;
 wire \vga_image_generator.counter[2] ;
 wire \vga_image_generator.counter[3] ;
 wire \vga_image_generator.counter[4] ;
 wire \vga_image_generator.counter[5] ;
 wire \vga_image_generator.counter[6] ;
 wire \vga_image_generator.counter[7] ;
 wire \vga_image_generator.counter[8] ;
 wire \vga_image_generator.counter[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net163;

 sg13g2_buf_1 _0919_ (.A(\hvsync_gen.vpos[4] ),
    .X(_0154_));
 sg13g2_buf_2 _0920_ (.A(\hvsync_gen.vpos[5] ),
    .X(_0155_));
 sg13g2_nor2b_2 _0921_ (.A(net63),
    .B_N(_0155_),
    .Y(_0156_));
 sg13g2_buf_1 _0922_ (.A(\hvsync_gen.vpos[0] ),
    .X(_0157_));
 sg13g2_buf_1 _0923_ (.A(\hvsync_gen.vpos[2] ),
    .X(_0158_));
 sg13g2_buf_1 _0924_ (.A(\hvsync_gen.vpos[3] ),
    .X(_0159_));
 sg13g2_nor2b_1 _0925_ (.A(_0158_),
    .B_N(net60),
    .Y(_0160_));
 sg13g2_nand2b_1 _0926_ (.Y(_0161_),
    .B(_0160_),
    .A_N(_0157_));
 sg13g2_o21ai_1 _0927_ (.B1(_0161_),
    .Y(_0162_),
    .A1(_0021_),
    .A2(_0020_));
 sg13g2_buf_2 _0928_ (.A(\hvsync_gen.vpos[8] ),
    .X(_0163_));
 sg13g2_inv_1 _0929_ (.Y(_0164_),
    .A(_0163_));
 sg13g2_buf_2 _0930_ (.A(\hvsync_gen.vpos[9] ),
    .X(_0165_));
 sg13g2_buf_1 _0931_ (.A(\hvsync_gen.vpos[7] ),
    .X(_0166_));
 sg13g2_buf_1 _0932_ (.A(\hvsync_gen.vpos[6] ),
    .X(_0167_));
 sg13g2_nand2_2 _0933_ (.Y(_0168_),
    .A(net59),
    .B(net58));
 sg13g2_nor3_1 _0934_ (.A(_0164_),
    .B(_0165_),
    .C(_0168_),
    .Y(_0169_));
 sg13g2_buf_1 _0935_ (.A(_0158_),
    .X(_0170_));
 sg13g2_inv_1 _0936_ (.Y(_0171_),
    .A(_0170_));
 sg13g2_nor2_1 _0937_ (.A(_0171_),
    .B(_0020_),
    .Y(_0172_));
 sg13g2_buf_1 _0938_ (.A(\hvsync_gen.vpos[1] ),
    .X(_0173_));
 sg13g2_nand2b_2 _0939_ (.Y(_0174_),
    .B(_0155_),
    .A_N(\hvsync_gen.vpos[4] ));
 sg13g2_nor3_1 _0940_ (.A(net57),
    .B(net47),
    .C(_0174_),
    .Y(_0175_));
 sg13g2_buf_1 _0941_ (.A(\hvsync_gen.vpos[3] ),
    .X(_0176_));
 sg13g2_o21ai_1 _0942_ (.B1(_0176_),
    .Y(_0177_),
    .A1(_0172_),
    .A2(_0175_));
 sg13g2_and4_1 _0943_ (.A(_0156_),
    .B(_0162_),
    .C(_0169_),
    .D(_0177_),
    .X(_0016_));
 sg13g2_buf_1 _0944_ (.A(_0022_),
    .X(_0178_));
 sg13g2_inv_1 _0945_ (.Y(_0179_),
    .A(_0178_));
 sg13g2_buf_2 _0946_ (.A(\hvsync_gen.hpos[8] ),
    .X(_0180_));
 sg13g2_inv_2 _0947_ (.Y(_0181_),
    .A(_0180_));
 sg13g2_buf_2 _0948_ (.A(\hvsync_gen.hpos[5] ),
    .X(_0182_));
 sg13g2_buf_1 _0949_ (.A(_0182_),
    .X(_0183_));
 sg13g2_buf_1 _0950_ (.A(\hvsync_gen.hpos[4] ),
    .X(_0184_));
 sg13g2_buf_1 _0951_ (.A(\hvsync_gen.hpos[6] ),
    .X(_0185_));
 sg13g2_nand3_1 _0952_ (.B(net55),
    .C(net54),
    .A(net46),
    .Y(_0186_));
 sg13g2_nand2_1 _0953_ (.Y(_0187_),
    .A(_0181_),
    .B(_0186_));
 sg13g2_buf_1 _0954_ (.A(net54),
    .X(_0188_));
 sg13g2_or2_1 _0955_ (.X(_0189_),
    .B(net55),
    .A(_0182_));
 sg13g2_buf_2 _0956_ (.A(_0189_),
    .X(_0190_));
 sg13g2_buf_1 _0957_ (.A(\hvsync_gen.hpos[7] ),
    .X(_0191_));
 sg13g2_buf_1 _0958_ (.A(_0191_),
    .X(_0192_));
 sg13g2_o21ai_1 _0959_ (.B1(net44),
    .Y(_0193_),
    .A1(net45),
    .A2(_0190_));
 sg13g2_buf_1 _0960_ (.A(\hvsync_gen.hpos[9] ),
    .X(_0194_));
 sg13g2_inv_1 _0961_ (.Y(_0195_),
    .A(_0194_));
 sg13g2_a221oi_1 _0962_ (.B2(_0181_),
    .C1(_0195_),
    .B1(_0193_),
    .A1(_0179_),
    .Y(_0015_),
    .A2(_0187_));
 sg13g2_buf_1 _0963_ (.A(BNC_trig),
    .X(_0196_));
 sg13g2_buf_1 _0964_ (.A(_0196_),
    .X(_0197_));
 sg13g2_buf_1 _0965_ (.A(net43),
    .X(_0198_));
 sg13g2_buf_1 _0966_ (.A(\bnc_image_generator.counter[0] ),
    .X(_0199_));
 sg13g2_buf_1 _0967_ (.A(net53),
    .X(_0200_));
 sg13g2_buf_1 _0968_ (.A(\bnc_image_generator.counter[2] ),
    .X(_0201_));
 sg13g2_inv_2 _0969_ (.Y(_0202_),
    .A(_0201_));
 sg13g2_buf_1 _0970_ (.A(\bnc_image_generator.counter[4] ),
    .X(_0203_));
 sg13g2_buf_1 _0971_ (.A(_0203_),
    .X(_0204_));
 sg13g2_nand2_2 _0972_ (.Y(_0205_),
    .A(_0202_),
    .B(net41));
 sg13g2_buf_1 _0973_ (.A(_0201_),
    .X(_0206_));
 sg13g2_nand2b_1 _0974_ (.Y(_0207_),
    .B(net40),
    .A_N(_0203_));
 sg13g2_nand3_1 _0975_ (.B(_0205_),
    .C(_0207_),
    .A(net42),
    .Y(_0208_));
 sg13g2_o21ai_1 _0976_ (.B1(_0208_),
    .Y(_0209_),
    .A1(net42),
    .A2(_0205_));
 sg13g2_buf_1 _0977_ (.A(\bnc_image_generator.counter[1] ),
    .X(_0210_));
 sg13g2_buf_1 _0978_ (.A(net52),
    .X(_0211_));
 sg13g2_buf_1 _0979_ (.A(_0196_),
    .X(_0212_));
 sg13g2_nand2b_1 _0980_ (.Y(_0213_),
    .B(_0201_),
    .A_N(net53));
 sg13g2_nand2_2 _0981_ (.Y(_0214_),
    .A(net53),
    .B(_0202_));
 sg13g2_a22oi_1 _0982_ (.Y(_0215_),
    .B1(_0213_),
    .B2(_0214_),
    .A2(net41),
    .A1(net38));
 sg13g2_inv_2 _0983_ (.Y(_0216_),
    .A(net52));
 sg13g2_or2_1 _0984_ (.X(_0217_),
    .B(_0213_),
    .A(_0216_));
 sg13g2_inv_1 _0985_ (.Y(_0218_),
    .A(_0196_));
 sg13g2_nand2b_1 _0986_ (.Y(_0219_),
    .B(net37),
    .A_N(_0217_));
 sg13g2_o21ai_1 _0987_ (.B1(_0219_),
    .Y(_0220_),
    .A1(net39),
    .A2(_0215_));
 sg13g2_a21oi_1 _0988_ (.A1(net24),
    .A2(_0209_),
    .Y(_0000_),
    .B1(_0220_));
 sg13g2_a21oi_1 _0989_ (.A1(_0205_),
    .A2(_0207_),
    .Y(_0221_),
    .B1(_0216_));
 sg13g2_nand2_1 _0990_ (.Y(_0222_),
    .A(net40),
    .B(net41));
 sg13g2_nor2_1 _0991_ (.A(net39),
    .B(_0222_),
    .Y(_0223_));
 sg13g2_nor2_1 _0992_ (.A(_0221_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_nor2_1 _0993_ (.A(_0202_),
    .B(_0203_),
    .Y(_0225_));
 sg13g2_a22oi_1 _0994_ (.Y(_0226_),
    .B1(_0225_),
    .B2(net39),
    .A2(net41),
    .A1(net43));
 sg13g2_nor2_1 _0995_ (.A(net42),
    .B(_0226_),
    .Y(_0227_));
 sg13g2_buf_1 _0996_ (.A(net40),
    .X(_0228_));
 sg13g2_nand2_2 _0997_ (.Y(_0229_),
    .A(_0216_),
    .B(net53));
 sg13g2_nor3_1 _0998_ (.A(net23),
    .B(net41),
    .C(_0229_),
    .Y(_0230_));
 sg13g2_nor2_1 _0999_ (.A(net52),
    .B(_0203_),
    .Y(_0231_));
 sg13g2_nand2_1 _1000_ (.Y(_0232_),
    .A(_0213_),
    .B(_0231_));
 sg13g2_a21oi_1 _1001_ (.A1(_0214_),
    .A2(_0232_),
    .Y(_0233_),
    .B1(net38));
 sg13g2_nor3_1 _1002_ (.A(_0227_),
    .B(_0230_),
    .C(_0233_),
    .Y(_0234_));
 sg13g2_o21ai_1 _1003_ (.B1(_0234_),
    .Y(_0001_),
    .A1(net37),
    .A2(_0224_));
 sg13g2_buf_1 _1004_ (.A(_0204_),
    .X(_0235_));
 sg13g2_and2_1 _1005_ (.A(\bnc_image_generator.counter[1] ),
    .B(_0199_),
    .X(_0236_));
 sg13g2_buf_1 _1006_ (.A(_0236_),
    .X(_0237_));
 sg13g2_xnor2_1 _1007_ (.Y(_0238_),
    .A(net40),
    .B(_0237_));
 sg13g2_nand2b_2 _1008_ (.Y(_0239_),
    .B(net52),
    .A_N(net53));
 sg13g2_a21oi_1 _1009_ (.A1(_0229_),
    .A2(_0239_),
    .Y(_0240_),
    .B1(_0018_));
 sg13g2_nor2_1 _1010_ (.A(net38),
    .B(_0240_),
    .Y(_0241_));
 sg13g2_a21oi_1 _1011_ (.A1(net24),
    .A2(_0238_),
    .Y(_0242_),
    .B1(_0241_));
 sg13g2_buf_1 _1012_ (.A(net41),
    .X(_0243_));
 sg13g2_nand2_1 _1013_ (.Y(_0244_),
    .A(_0210_),
    .B(net42));
 sg13g2_nor2_1 _1014_ (.A(net40),
    .B(_0244_),
    .Y(_0245_));
 sg13g2_a21oi_1 _1015_ (.A1(_0217_),
    .A2(_0229_),
    .Y(_0246_),
    .B1(net38));
 sg13g2_and3_1 _1016_ (.X(_0247_),
    .A(net43),
    .B(net23),
    .C(_0019_));
 sg13g2_nor4_1 _1017_ (.A(net21),
    .B(_0245_),
    .C(_0246_),
    .D(_0247_),
    .Y(_0248_));
 sg13g2_a21oi_1 _1018_ (.A1(net22),
    .A2(_0242_),
    .Y(_0002_),
    .B1(_0248_));
 sg13g2_inv_1 _1019_ (.Y(_0249_),
    .A(_0030_));
 sg13g2_nor2_1 _1020_ (.A(\bnc_image_generator.counter[1] ),
    .B(net53),
    .Y(_0250_));
 sg13g2_nor2_1 _1021_ (.A(_0201_),
    .B(_0250_),
    .Y(_0251_));
 sg13g2_nor2_1 _1022_ (.A(_0196_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_a221oi_1 _1023_ (.B2(net38),
    .C1(_0252_),
    .B1(_0245_),
    .A1(_0228_),
    .Y(_0253_),
    .A2(_0249_));
 sg13g2_o21ai_1 _1024_ (.B1(_0200_),
    .Y(_0254_),
    .A1(net52),
    .A2(net40));
 sg13g2_nor2_1 _1025_ (.A(_0199_),
    .B(_0201_),
    .Y(_0255_));
 sg13g2_a221oi_1 _1026_ (.B2(net39),
    .C1(net21),
    .B1(_0255_),
    .A1(_0212_),
    .Y(_0256_),
    .A2(_0254_));
 sg13g2_a21o_1 _1027_ (.A2(_0253_),
    .A1(net22),
    .B1(_0256_),
    .X(_0003_));
 sg13g2_nor2_1 _1028_ (.A(net37),
    .B(net21),
    .Y(_0257_));
 sg13g2_nor3_1 _1029_ (.A(net38),
    .B(net42),
    .C(_0205_),
    .Y(_0258_));
 sg13g2_o21ai_1 _1030_ (.B1(_0211_),
    .Y(_0259_),
    .A1(_0257_),
    .A2(_0258_));
 sg13g2_nor2_1 _1031_ (.A(net52),
    .B(_0214_),
    .Y(_0260_));
 sg13g2_a21o_1 _1032_ (.A2(_0019_),
    .A1(net23),
    .B1(_0260_),
    .X(_0261_));
 sg13g2_nand3_1 _1033_ (.B(net21),
    .C(_0261_),
    .A(net24),
    .Y(_0262_));
 sg13g2_a21oi_1 _1034_ (.A1(_0197_),
    .A2(_0255_),
    .Y(_0263_),
    .B1(_0252_));
 sg13g2_or2_1 _1035_ (.X(_0264_),
    .B(_0263_),
    .A(net21));
 sg13g2_nand3_1 _1036_ (.B(_0262_),
    .C(_0264_),
    .A(_0259_),
    .Y(_0004_));
 sg13g2_inv_1 _1037_ (.Y(_0265_),
    .A(_0255_));
 sg13g2_nand2_1 _1038_ (.Y(_0266_),
    .A(net42),
    .B(_0206_));
 sg13g2_o21ai_1 _1039_ (.B1(_0266_),
    .Y(_0267_),
    .A1(_0216_),
    .A2(_0265_));
 sg13g2_nor3_1 _1040_ (.A(net43),
    .B(_0211_),
    .C(_0214_),
    .Y(_0268_));
 sg13g2_a21oi_1 _1041_ (.A1(net24),
    .A2(_0267_),
    .Y(_0269_),
    .B1(_0268_));
 sg13g2_xor2_1 _1042_ (.B(_0269_),
    .A(net22),
    .X(_0005_));
 sg13g2_nor2b_1 _1043_ (.A(_0196_),
    .B_N(_0203_),
    .Y(_0270_));
 sg13g2_a21o_1 _1044_ (.A2(_0237_),
    .A1(net41),
    .B1(_0231_),
    .X(_0271_));
 sg13g2_a22oi_1 _1045_ (.Y(_0272_),
    .B1(_0271_),
    .B2(net24),
    .A2(_0270_),
    .A1(_0250_));
 sg13g2_a22oi_1 _1046_ (.Y(_0273_),
    .B1(_0265_),
    .B2(net37),
    .A2(_0214_),
    .A1(net39));
 sg13g2_nand4_1 _1047_ (.B(_0206_),
    .C(_0204_),
    .A(_0197_),
    .Y(_0274_),
    .D(_0019_));
 sg13g2_o21ai_1 _1048_ (.B1(_0274_),
    .Y(_0275_),
    .A1(net21),
    .A2(_0273_));
 sg13g2_inv_1 _1049_ (.Y(_0276_),
    .A(_0275_));
 sg13g2_o21ai_1 _1050_ (.B1(_0276_),
    .Y(_0006_),
    .A1(net23),
    .A2(_0272_));
 sg13g2_nand3_1 _1051_ (.B(net39),
    .C(net23),
    .A(net38),
    .Y(_0277_));
 sg13g2_nand2_1 _1052_ (.Y(_0278_),
    .A(net52),
    .B(net40));
 sg13g2_o21ai_1 _1053_ (.B1(net21),
    .Y(_0279_),
    .A1(_0017_),
    .A2(_0278_));
 sg13g2_o21ai_1 _1054_ (.B1(_0279_),
    .Y(_0280_),
    .A1(net22),
    .A2(_0277_));
 sg13g2_inv_1 _1055_ (.Y(_0007_),
    .A(_0280_));
 sg13g2_nor2b_2 _1056_ (.A(net53),
    .B_N(_0203_),
    .Y(_0281_));
 sg13g2_nor2_1 _1057_ (.A(net23),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_a22oi_1 _1058_ (.Y(_0283_),
    .B1(_0282_),
    .B2(net24),
    .A2(_0270_),
    .A1(_0265_));
 sg13g2_nand2b_1 _1059_ (.Y(_0284_),
    .B(net43),
    .A_N(net42));
 sg13g2_o21ai_1 _1060_ (.B1(_0205_),
    .Y(_0285_),
    .A1(_0207_),
    .A2(_0284_));
 sg13g2_a21oi_1 _1061_ (.A1(_0019_),
    .A2(_0225_),
    .Y(_0286_),
    .B1(_0260_));
 sg13g2_nor2_1 _1062_ (.A(net38),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_a21oi_1 _1063_ (.A1(_0216_),
    .A2(_0285_),
    .Y(_0288_),
    .B1(_0287_));
 sg13g2_o21ai_1 _1064_ (.B1(_0288_),
    .Y(_0008_),
    .A1(_0216_),
    .A2(_0283_));
 sg13g2_xnor2_1 _1065_ (.Y(_0289_),
    .A(net40),
    .B(_0281_));
 sg13g2_nor2b_1 _1066_ (.A(_0203_),
    .B_N(net53),
    .Y(_0290_));
 sg13g2_nor3_1 _1067_ (.A(net52),
    .B(_0281_),
    .C(_0290_),
    .Y(_0291_));
 sg13g2_a21oi_1 _1068_ (.A1(net39),
    .A2(_0289_),
    .Y(_0292_),
    .B1(_0291_));
 sg13g2_a21oi_1 _1069_ (.A1(_0018_),
    .A2(_0281_),
    .Y(_0293_),
    .B1(_0225_));
 sg13g2_mux2_1 _1070_ (.A0(_0292_),
    .A1(_0293_),
    .S(net37),
    .X(_0294_));
 sg13g2_o21ai_1 _1071_ (.B1(_0294_),
    .Y(_0009_),
    .A1(net22),
    .A2(_0244_));
 sg13g2_o21ai_1 _1072_ (.B1(_0207_),
    .Y(_0295_),
    .A1(_0205_),
    .A2(_0239_));
 sg13g2_a21oi_1 _1073_ (.A1(_0237_),
    .A2(_0270_),
    .Y(_0296_),
    .B1(_0231_));
 sg13g2_nor2_1 _1074_ (.A(_0030_),
    .B(_0222_),
    .Y(_0297_));
 sg13g2_nor2_1 _1075_ (.A(net42),
    .B(net41),
    .Y(_0298_));
 sg13g2_o21ai_1 _1076_ (.B1(net37),
    .Y(_0299_),
    .A1(_0297_),
    .A2(_0298_));
 sg13g2_o21ai_1 _1077_ (.B1(_0299_),
    .Y(_0300_),
    .A1(net23),
    .A2(_0296_));
 sg13g2_a21oi_1 _1078_ (.A1(net24),
    .A2(_0295_),
    .Y(_0010_),
    .B1(_0300_));
 sg13g2_inv_1 _1079_ (.Y(_0301_),
    .A(_0251_));
 sg13g2_a221oi_1 _1080_ (.B2(_0212_),
    .C1(_0268_),
    .B1(_0301_),
    .A1(net23),
    .Y(_0302_),
    .A2(_0019_));
 sg13g2_o21ai_1 _1081_ (.B1(_0239_),
    .Y(_0303_),
    .A1(net37),
    .A2(_0229_));
 sg13g2_nand2_1 _1082_ (.Y(_0304_),
    .A(_0216_),
    .B(_0265_));
 sg13g2_a221oi_1 _1083_ (.B2(net37),
    .C1(_0243_),
    .B1(_0304_),
    .A1(_0202_),
    .Y(_0305_),
    .A2(_0303_));
 sg13g2_a21oi_1 _1084_ (.A1(_0235_),
    .A2(_0302_),
    .Y(_0011_),
    .B1(_0305_));
 sg13g2_a21oi_1 _1085_ (.A1(_0198_),
    .A2(_0229_),
    .Y(_0306_),
    .B1(_0267_));
 sg13g2_nor2_1 _1086_ (.A(net43),
    .B(_0202_),
    .Y(_0307_));
 sg13g2_nand2_1 _1087_ (.Y(_0308_),
    .A(_0218_),
    .B(_0239_));
 sg13g2_nand2_1 _1088_ (.Y(_0309_),
    .A(_0229_),
    .B(_0308_));
 sg13g2_a221oi_1 _1089_ (.B2(_0202_),
    .C1(_0243_),
    .B1(_0309_),
    .A1(_0030_),
    .Y(_0310_),
    .A2(_0307_));
 sg13g2_a21oi_1 _1090_ (.A1(_0235_),
    .A2(_0306_),
    .Y(_0012_),
    .B1(_0310_));
 sg13g2_o21ai_1 _1091_ (.B1(_0196_),
    .Y(_0311_),
    .A1(_0210_),
    .A2(_0200_));
 sg13g2_o21ai_1 _1092_ (.B1(_0311_),
    .Y(_0312_),
    .A1(net39),
    .A2(_0202_));
 sg13g2_or2_1 _1093_ (.X(_0313_),
    .B(_0312_),
    .A(_0245_));
 sg13g2_nand2b_1 _1094_ (.Y(_0314_),
    .B(_0307_),
    .A_N(_0019_));
 sg13g2_nor2_1 _1095_ (.A(net43),
    .B(_0237_),
    .Y(_0315_));
 sg13g2_o21ai_1 _1096_ (.B1(_0202_),
    .Y(_0316_),
    .A1(_0250_),
    .A2(_0315_));
 sg13g2_nand3_1 _1097_ (.B(_0314_),
    .C(_0316_),
    .A(net22),
    .Y(_0317_));
 sg13g2_o21ai_1 _1098_ (.B1(_0317_),
    .Y(_0013_),
    .A1(net22),
    .A2(_0313_));
 sg13g2_a21oi_1 _1099_ (.A1(_0017_),
    .A2(_0278_),
    .Y(_0318_),
    .B1(net22));
 sg13g2_a21oi_1 _1100_ (.A1(_0270_),
    .A2(_0278_),
    .Y(_0014_),
    .B1(_0318_));
 sg13g2_nor2_1 _1101_ (.A(net57),
    .B(net62),
    .Y(_0319_));
 sg13g2_nor2_1 _1102_ (.A(_0155_),
    .B(net63),
    .Y(_0320_));
 sg13g2_nand3_1 _1103_ (.B(_0165_),
    .C(_0320_),
    .A(_0164_),
    .Y(_0321_));
 sg13g2_nand2_1 _1104_ (.Y(_0322_),
    .A(net47),
    .B(net60));
 sg13g2_nor4_1 _1105_ (.A(net59),
    .B(net58),
    .C(_0321_),
    .D(_0322_),
    .Y(_0323_));
 sg13g2_inv_1 _1106_ (.Y(_0324_),
    .A(net1));
 sg13g2_a21o_1 _1107_ (.A2(_0323_),
    .A1(_0319_),
    .B1(_0324_),
    .X(_0325_));
 sg13g2_buf_1 _1108_ (.A(_0325_),
    .X(_0326_));
 sg13g2_buf_1 _1109_ (.A(_0180_),
    .X(_0327_));
 sg13g2_buf_1 _1110_ (.A(_0194_),
    .X(_0328_));
 sg13g2_buf_1 _1111_ (.A(\hvsync_gen.hpos[1] ),
    .X(_0329_));
 sg13g2_buf_2 _1112_ (.A(\hvsync_gen.hpos[0] ),
    .X(_0330_));
 sg13g2_and2_1 _1113_ (.A(net51),
    .B(_0330_),
    .X(_0331_));
 sg13g2_buf_1 _1114_ (.A(_0331_),
    .X(_0332_));
 sg13g2_buf_1 _1115_ (.A(\hvsync_gen.hpos[2] ),
    .X(_0333_));
 sg13g2_buf_1 _1116_ (.A(\hvsync_gen.hpos[3] ),
    .X(_0334_));
 sg13g2_and2_1 _1117_ (.A(net50),
    .B(net49),
    .X(_0335_));
 sg13g2_buf_1 _1118_ (.A(_0335_),
    .X(_0336_));
 sg13g2_nand2_1 _1119_ (.Y(_0337_),
    .A(_0332_),
    .B(_0336_));
 sg13g2_nand2b_1 _1120_ (.Y(_0338_),
    .B(net55),
    .A_N(_0182_));
 sg13g2_nor2_1 _1121_ (.A(_0337_),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_nor2_1 _1122_ (.A(net54),
    .B(_0192_),
    .Y(_0340_));
 sg13g2_nand4_1 _1123_ (.B(net35),
    .C(_0339_),
    .A(net36),
    .Y(_0341_),
    .D(_0340_));
 sg13g2_inv_1 _1124_ (.Y(_0342_),
    .A(_0341_));
 sg13g2_nand2_1 _1125_ (.Y(_0343_),
    .A(_0029_),
    .B(_0342_));
 sg13g2_nand3_1 _1126_ (.B(_0157_),
    .C(_0341_),
    .A(net1),
    .Y(_0344_));
 sg13g2_o21ai_1 _1127_ (.B1(_0344_),
    .Y(_0047_),
    .A1(_0326_),
    .A2(_0343_));
 sg13g2_nand2_1 _1128_ (.Y(_0345_),
    .A(net62),
    .B(_0342_));
 sg13g2_xnor2_1 _1129_ (.Y(_0346_),
    .A(net57),
    .B(_0345_));
 sg13g2_and2_1 _1130_ (.A(net1),
    .B(_0346_),
    .X(_0048_));
 sg13g2_nand3_1 _1131_ (.B(net62),
    .C(_0171_),
    .A(net57),
    .Y(_0347_));
 sg13g2_or2_1 _1132_ (.X(_0348_),
    .B(_0326_),
    .A(_0341_));
 sg13g2_buf_2 _1133_ (.A(_0348_),
    .X(_0349_));
 sg13g2_buf_1 _1134_ (.A(_0324_),
    .X(_0350_));
 sg13g2_nor2_2 _1135_ (.A(_0350_),
    .B(_0342_),
    .Y(_0351_));
 sg13g2_a21oi_1 _1136_ (.A1(_0173_),
    .A2(net62),
    .Y(_0352_),
    .B1(net19));
 sg13g2_o21ai_1 _1137_ (.B1(_0170_),
    .Y(_0353_),
    .A1(_0351_),
    .A2(_0352_));
 sg13g2_o21ai_1 _1138_ (.B1(_0353_),
    .Y(_0049_),
    .A1(_0347_),
    .A2(_0349_));
 sg13g2_nand3_1 _1139_ (.B(\hvsync_gen.vpos[0] ),
    .C(net61),
    .A(\hvsync_gen.vpos[1] ),
    .Y(_0354_));
 sg13g2_buf_1 _1140_ (.A(_0354_),
    .X(_0355_));
 sg13g2_or2_1 _1141_ (.X(_0356_),
    .B(_0355_),
    .A(net56));
 sg13g2_nor2b_1 _1142_ (.A(net19),
    .B_N(_0355_),
    .Y(_0357_));
 sg13g2_o21ai_1 _1143_ (.B1(_0176_),
    .Y(_0358_),
    .A1(_0351_),
    .A2(_0357_));
 sg13g2_o21ai_1 _1144_ (.B1(_0358_),
    .Y(_0050_),
    .A1(_0349_),
    .A2(_0356_));
 sg13g2_buf_1 _1145_ (.A(_0154_),
    .X(_0359_));
 sg13g2_inv_1 _1146_ (.Y(_0360_),
    .A(net34));
 sg13g2_and4_1 _1147_ (.A(_0173_),
    .B(net62),
    .C(net61),
    .D(net60),
    .X(_0361_));
 sg13g2_buf_1 _1148_ (.A(_0361_),
    .X(_0362_));
 sg13g2_nand2_1 _1149_ (.Y(_0363_),
    .A(_0360_),
    .B(_0362_));
 sg13g2_nand2_2 _1150_ (.Y(_0364_),
    .A(net1),
    .B(_0341_));
 sg13g2_o21ai_1 _1151_ (.B1(_0364_),
    .Y(_0365_),
    .A1(net19),
    .A2(_0362_));
 sg13g2_nand2_1 _1152_ (.Y(_0366_),
    .A(_0359_),
    .B(_0365_));
 sg13g2_o21ai_1 _1153_ (.B1(_0366_),
    .Y(_0051_),
    .A1(_0349_),
    .A2(_0363_));
 sg13g2_buf_1 _1154_ (.A(_0155_),
    .X(_0367_));
 sg13g2_inv_1 _1155_ (.Y(_0368_),
    .A(net33));
 sg13g2_nand3_1 _1156_ (.B(net34),
    .C(_0362_),
    .A(_0368_),
    .Y(_0369_));
 sg13g2_a21oi_1 _1157_ (.A1(net34),
    .A2(_0362_),
    .Y(_0370_),
    .B1(net19));
 sg13g2_o21ai_1 _1158_ (.B1(_0367_),
    .Y(_0371_),
    .A1(_0351_),
    .A2(_0370_));
 sg13g2_o21ai_1 _1159_ (.B1(_0371_),
    .Y(_0052_),
    .A1(_0349_),
    .A2(_0369_));
 sg13g2_and3_1 _1160_ (.X(_0372_),
    .A(_0367_),
    .B(_0359_),
    .C(_0362_));
 sg13g2_buf_2 _1161_ (.A(_0372_),
    .X(_0373_));
 sg13g2_nand2b_1 _1162_ (.Y(_0374_),
    .B(_0373_),
    .A_N(_0349_));
 sg13g2_o21ai_1 _1163_ (.B1(_0364_),
    .Y(_0375_),
    .A1(net19),
    .A2(_0373_));
 sg13g2_nand2_1 _1164_ (.Y(_0376_),
    .A(net58),
    .B(_0375_));
 sg13g2_o21ai_1 _1165_ (.B1(_0376_),
    .Y(_0053_),
    .A1(net58),
    .A2(_0374_));
 sg13g2_nand3b_1 _1166_ (.B(_0167_),
    .C(_0373_),
    .Y(_0377_),
    .A_N(net59));
 sg13g2_a21oi_1 _1167_ (.A1(_0167_),
    .A2(_0373_),
    .Y(_0378_),
    .B1(net19));
 sg13g2_o21ai_1 _1168_ (.B1(net59),
    .Y(_0379_),
    .A1(_0351_),
    .A2(_0378_));
 sg13g2_o21ai_1 _1169_ (.B1(_0379_),
    .Y(_0054_),
    .A1(_0349_),
    .A2(_0377_));
 sg13g2_nand2b_1 _1170_ (.Y(_0380_),
    .B(_0373_),
    .A_N(_0168_));
 sg13g2_nor3_1 _1171_ (.A(_0163_),
    .B(_0349_),
    .C(_0380_),
    .Y(_0381_));
 sg13g2_nand2b_1 _1172_ (.Y(_0382_),
    .B(_0380_),
    .A_N(net19));
 sg13g2_a21oi_1 _1173_ (.A1(_0364_),
    .A2(_0382_),
    .Y(_0383_),
    .B1(_0164_));
 sg13g2_or2_1 _1174_ (.X(_0055_),
    .B(_0383_),
    .A(_0381_));
 sg13g2_nand2_1 _1175_ (.Y(_0384_),
    .A(_0169_),
    .B(_0373_));
 sg13g2_nor2_1 _1176_ (.A(_0164_),
    .B(_0168_),
    .Y(_0385_));
 sg13g2_a21oi_1 _1177_ (.A1(_0385_),
    .A2(_0373_),
    .Y(_0386_),
    .B1(net19));
 sg13g2_o21ai_1 _1178_ (.B1(_0165_),
    .Y(_0387_),
    .A1(_0351_),
    .A2(_0386_));
 sg13g2_o21ai_1 _1179_ (.B1(_0387_),
    .Y(_0056_),
    .A1(_0349_),
    .A2(_0384_));
 sg13g2_and2_1 _1180_ (.A(_0028_),
    .B(_0351_),
    .X(_0037_));
 sg13g2_nand2b_1 _1181_ (.Y(_0388_),
    .B(_0330_),
    .A_N(net51));
 sg13g2_nand2b_1 _1182_ (.Y(_0389_),
    .B(net51),
    .A_N(_0330_));
 sg13g2_a21oi_1 _1183_ (.A1(_0388_),
    .A2(_0389_),
    .Y(_0038_),
    .B1(net48));
 sg13g2_buf_1 _1184_ (.A(net48),
    .X(_0390_));
 sg13g2_buf_1 _1185_ (.A(net50),
    .X(_0391_));
 sg13g2_xnor2_1 _1186_ (.Y(_0392_),
    .A(net31),
    .B(_0332_));
 sg13g2_nor2_1 _1187_ (.A(net32),
    .B(_0392_),
    .Y(_0039_));
 sg13g2_inv_2 _1188_ (.Y(_0393_),
    .A(net49));
 sg13g2_nand3_1 _1189_ (.B(_0330_),
    .C(net50),
    .A(net51),
    .Y(_0394_));
 sg13g2_xnor2_1 _1190_ (.Y(_0395_),
    .A(_0393_),
    .B(_0394_));
 sg13g2_nor2_1 _1191_ (.A(net32),
    .B(_0395_),
    .Y(_0040_));
 sg13g2_inv_1 _1192_ (.Y(_0396_),
    .A(net55));
 sg13g2_xnor2_1 _1193_ (.Y(_0397_),
    .A(_0396_),
    .B(_0337_));
 sg13g2_nor2_1 _1194_ (.A(net32),
    .B(_0397_),
    .Y(_0041_));
 sg13g2_nand2_1 _1195_ (.Y(_0398_),
    .A(net51),
    .B(_0330_));
 sg13g2_buf_1 _1196_ (.A(net49),
    .X(_0399_));
 sg13g2_buf_1 _1197_ (.A(net55),
    .X(_0400_));
 sg13g2_nand3_1 _1198_ (.B(net30),
    .C(net29),
    .A(net50),
    .Y(_0401_));
 sg13g2_nor2_2 _1199_ (.A(_0398_),
    .B(_0401_),
    .Y(_0402_));
 sg13g2_xnor2_1 _1200_ (.Y(_0403_),
    .A(net46),
    .B(_0402_));
 sg13g2_nor2_1 _1201_ (.A(_0364_),
    .B(_0403_),
    .Y(_0042_));
 sg13g2_nand2_1 _1202_ (.Y(_0404_),
    .A(net46),
    .B(_0402_));
 sg13g2_xor2_1 _1203_ (.B(_0404_),
    .A(net45),
    .X(_0405_));
 sg13g2_nor2_1 _1204_ (.A(_0364_),
    .B(_0405_),
    .Y(_0043_));
 sg13g2_and2_1 _1205_ (.A(_0182_),
    .B(net54),
    .X(_0406_));
 sg13g2_buf_1 _1206_ (.A(_0406_),
    .X(_0407_));
 sg13g2_nand2_1 _1207_ (.Y(_0408_),
    .A(_0402_),
    .B(_0407_));
 sg13g2_xor2_1 _1208_ (.B(_0408_),
    .A(net44),
    .X(_0409_));
 sg13g2_nor2_1 _1209_ (.A(_0364_),
    .B(_0409_),
    .Y(_0044_));
 sg13g2_nand3_1 _1210_ (.B(_0402_),
    .C(_0407_),
    .A(net44),
    .Y(_0410_));
 sg13g2_xnor2_1 _1211_ (.Y(_0411_),
    .A(_0181_),
    .B(_0410_));
 sg13g2_nor2_1 _1212_ (.A(_0364_),
    .B(_0411_),
    .Y(_0045_));
 sg13g2_or2_1 _1213_ (.X(_0412_),
    .B(_0410_),
    .A(_0181_));
 sg13g2_xnor2_1 _1214_ (.Y(_0413_),
    .A(_0195_),
    .B(_0412_));
 sg13g2_nor2_1 _1215_ (.A(_0364_),
    .B(_0413_),
    .Y(_0046_));
 sg13g2_nor2_1 _1216_ (.A(net32),
    .B(_0249_),
    .Y(_0032_));
 sg13g2_a21oi_1 _1217_ (.A1(_0229_),
    .A2(_0239_),
    .Y(_0033_),
    .B1(net48));
 sg13g2_nor2_1 _1218_ (.A(net32),
    .B(_0238_),
    .Y(_0034_));
 sg13g2_nor2_1 _1219_ (.A(_0030_),
    .B(_0278_),
    .Y(_0414_));
 sg13g2_xnor2_1 _1220_ (.Y(_0415_),
    .A(_0198_),
    .B(_0414_));
 sg13g2_nor2_1 _1221_ (.A(net32),
    .B(_0415_),
    .Y(_0035_));
 sg13g2_nand3_1 _1222_ (.B(_0228_),
    .C(_0237_),
    .A(net43),
    .Y(_0416_));
 sg13g2_xor2_1 _1223_ (.B(_0416_),
    .A(net21),
    .X(_0417_));
 sg13g2_nor2_1 _1224_ (.A(net32),
    .B(_0417_),
    .Y(_0036_));
 sg13g2_inv_2 _1225_ (.Y(_0418_),
    .A(\vga_image_generator.counter[24] ));
 sg13g2_buf_2 _1226_ (.A(\vga_image_generator.counter[25] ),
    .X(_0419_));
 sg13g2_nand2_1 _1227_ (.Y(_0420_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_nand2b_1 _1228_ (.Y(_0421_),
    .B(\vga_image_generator.counter[26] ),
    .A_N(\vga_image_generator.counter[27] ));
 sg13g2_nor2_1 _1229_ (.A(_0420_),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_buf_2 _1230_ (.A(\vga_image_generator.counter[21] ),
    .X(_0423_));
 sg13g2_buf_2 _1231_ (.A(\vga_image_generator.counter[20] ),
    .X(_0424_));
 sg13g2_buf_2 _1232_ (.A(\vga_image_generator.counter[22] ),
    .X(_0425_));
 sg13g2_nor4_2 _1233_ (.A(_0423_),
    .B(_0424_),
    .C(\vga_image_generator.counter[23] ),
    .Y(_0426_),
    .D(_0425_));
 sg13g2_a21oi_1 _1234_ (.A1(_0422_),
    .A2(_0426_),
    .Y(_0427_),
    .B1(\vga_image_generator.character_hold[0] ));
 sg13g2_nor2_1 _1235_ (.A(_0390_),
    .B(_0427_),
    .Y(_0057_));
 sg13g2_nand2b_1 _1236_ (.Y(_0428_),
    .B(\vga_image_generator.counter[27] ),
    .A_N(\vga_image_generator.counter[26] ));
 sg13g2_nor3_2 _1237_ (.A(\vga_image_generator.counter[24] ),
    .B(_0419_),
    .C(_0428_),
    .Y(_0429_));
 sg13g2_inv_1 _1238_ (.Y(_0430_),
    .A(\vga_image_generator.counter[23] ));
 sg13g2_nor4_2 _1239_ (.A(_0423_),
    .B(_0424_),
    .C(_0430_),
    .Y(_0431_),
    .D(_0425_));
 sg13g2_a21oi_1 _1240_ (.A1(_0429_),
    .A2(_0431_),
    .Y(_0432_),
    .B1(\vga_image_generator.character_hold[10] ));
 sg13g2_nor2_1 _1241_ (.A(net32),
    .B(_0432_),
    .Y(_0058_));
 sg13g2_nand2_1 _1242_ (.Y(_0433_),
    .A(\vga_image_generator.counter[23] ),
    .B(_0425_));
 sg13g2_nor3_2 _1243_ (.A(_0423_),
    .B(_0424_),
    .C(_0433_),
    .Y(_0434_));
 sg13g2_a21oi_1 _1244_ (.A1(_0429_),
    .A2(_0434_),
    .Y(_0435_),
    .B1(\vga_image_generator.character_hold[11] ));
 sg13g2_nor2_1 _1245_ (.A(_0390_),
    .B(_0435_),
    .Y(_0059_));
 sg13g2_buf_1 _1246_ (.A(net48),
    .X(_0436_));
 sg13g2_nor3_2 _1247_ (.A(_0418_),
    .B(_0419_),
    .C(_0428_),
    .Y(_0437_));
 sg13g2_a21oi_1 _1248_ (.A1(_0426_),
    .A2(_0437_),
    .Y(_0438_),
    .B1(\vga_image_generator.character_hold[12] ));
 sg13g2_nor2_1 _1249_ (.A(net28),
    .B(_0438_),
    .Y(_0060_));
 sg13g2_inv_1 _1250_ (.Y(_0439_),
    .A(_0425_));
 sg13g2_nor4_2 _1251_ (.A(_0423_),
    .B(_0424_),
    .C(\vga_image_generator.counter[23] ),
    .Y(_0440_),
    .D(_0439_));
 sg13g2_a21oi_1 _1252_ (.A1(_0437_),
    .A2(_0440_),
    .Y(_0441_),
    .B1(\vga_image_generator.character_hold[13] ));
 sg13g2_nor2_1 _1253_ (.A(net28),
    .B(_0441_),
    .Y(_0061_));
 sg13g2_a21oi_1 _1254_ (.A1(_0431_),
    .A2(_0437_),
    .Y(_0442_),
    .B1(\vga_image_generator.character_hold[14] ));
 sg13g2_nor2_1 _1255_ (.A(net28),
    .B(_0442_),
    .Y(_0062_));
 sg13g2_a21oi_1 _1256_ (.A1(_0434_),
    .A2(_0437_),
    .Y(_0443_),
    .B1(\vga_image_generator.character_hold[15] ));
 sg13g2_nor2_1 _1257_ (.A(_0436_),
    .B(_0443_),
    .Y(_0063_));
 sg13g2_nor2_1 _1258_ (.A(_0420_),
    .B(_0428_),
    .Y(_0444_));
 sg13g2_a21oi_1 _1259_ (.A1(_0426_),
    .A2(_0444_),
    .Y(_0445_),
    .B1(\vga_image_generator.character_hold[16] ));
 sg13g2_nor2_1 _1260_ (.A(net28),
    .B(_0445_),
    .Y(_0064_));
 sg13g2_a21oi_1 _1261_ (.A1(_0440_),
    .A2(_0444_),
    .Y(_0446_),
    .B1(\vga_image_generator.character_hold[17] ));
 sg13g2_nor2_1 _1262_ (.A(net28),
    .B(_0446_),
    .Y(_0065_));
 sg13g2_a21oi_1 _1263_ (.A1(_0422_),
    .A2(_0440_),
    .Y(_0447_),
    .B1(\vga_image_generator.character_hold[1] ));
 sg13g2_nor2_1 _1264_ (.A(net28),
    .B(_0447_),
    .Y(_0066_));
 sg13g2_a21oi_1 _1265_ (.A1(_0422_),
    .A2(_0431_),
    .Y(_0448_),
    .B1(\vga_image_generator.character_hold[2] ));
 sg13g2_nor2_1 _1266_ (.A(net28),
    .B(_0448_),
    .Y(_0067_));
 sg13g2_a21oi_1 _1267_ (.A1(_0422_),
    .A2(_0434_),
    .Y(_0449_),
    .B1(\vga_image_generator.character_hold[3] ));
 sg13g2_nor2_1 _1268_ (.A(net28),
    .B(_0449_),
    .Y(_0068_));
 sg13g2_inv_1 _1269_ (.Y(_0450_),
    .A(_0419_));
 sg13g2_nor3_2 _1270_ (.A(_0418_),
    .B(_0450_),
    .C(_0421_),
    .Y(_0451_));
 sg13g2_a21oi_1 _1271_ (.A1(_0426_),
    .A2(_0451_),
    .Y(_0452_),
    .B1(\vga_image_generator.character_hold[4] ));
 sg13g2_nor2_1 _1272_ (.A(_0436_),
    .B(_0452_),
    .Y(_0069_));
 sg13g2_buf_1 _1273_ (.A(net48),
    .X(_0453_));
 sg13g2_a21oi_1 _1274_ (.A1(_0440_),
    .A2(_0451_),
    .Y(_0454_),
    .B1(\vga_image_generator.character_hold[5] ));
 sg13g2_nor2_1 _1275_ (.A(net27),
    .B(_0454_),
    .Y(_0070_));
 sg13g2_a21oi_1 _1276_ (.A1(_0431_),
    .A2(_0451_),
    .Y(_0455_),
    .B1(\vga_image_generator.character_hold[6] ));
 sg13g2_nor2_1 _1277_ (.A(net27),
    .B(_0455_),
    .Y(_0071_));
 sg13g2_a21oi_1 _1278_ (.A1(_0434_),
    .A2(_0451_),
    .Y(_0456_),
    .B1(\vga_image_generator.character_hold[7] ));
 sg13g2_nor2_1 _1279_ (.A(net27),
    .B(_0456_),
    .Y(_0072_));
 sg13g2_a21oi_1 _1280_ (.A1(_0426_),
    .A2(_0429_),
    .Y(_0457_),
    .B1(\vga_image_generator.character_hold[8] ));
 sg13g2_nor2_1 _1281_ (.A(_0453_),
    .B(_0457_),
    .Y(_0073_));
 sg13g2_a21oi_1 _1282_ (.A1(_0429_),
    .A2(_0440_),
    .Y(_0458_),
    .B1(\vga_image_generator.character_hold[9] ));
 sg13g2_nor2_1 _1283_ (.A(_0453_),
    .B(_0458_),
    .Y(_0074_));
 sg13g2_and2_1 _1284_ (.A(net1),
    .B(_0031_),
    .X(_0075_));
 sg13g2_inv_1 _1285_ (.Y(_0459_),
    .A(\vga_image_generator.counter[7] ));
 sg13g2_and4_1 _1286_ (.A(\vga_image_generator.counter[1] ),
    .B(\vga_image_generator.counter[0] ),
    .C(\vga_image_generator.counter[2] ),
    .D(\vga_image_generator.counter[3] ),
    .X(_0460_));
 sg13g2_buf_1 _1287_ (.A(_0460_),
    .X(_0461_));
 sg13g2_nand4_1 _1288_ (.B(\vga_image_generator.counter[5] ),
    .C(\vga_image_generator.counter[6] ),
    .A(\vga_image_generator.counter[4] ),
    .Y(_0462_),
    .D(_0461_));
 sg13g2_nor2_1 _1289_ (.A(_0459_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_and2_1 _1290_ (.A(\vga_image_generator.counter[8] ),
    .B(_0463_),
    .X(_0464_));
 sg13g2_buf_1 _1291_ (.A(_0464_),
    .X(_0465_));
 sg13g2_nand2_1 _1292_ (.Y(_0466_),
    .A(\vga_image_generator.counter[9] ),
    .B(_0465_));
 sg13g2_xor2_1 _1293_ (.B(_0466_),
    .A(\vga_image_generator.counter[10] ),
    .X(_0467_));
 sg13g2_nor2_1 _1294_ (.A(net27),
    .B(_0467_),
    .Y(_0076_));
 sg13g2_nand3_1 _1295_ (.B(\vga_image_generator.counter[10] ),
    .C(_0465_),
    .A(\vga_image_generator.counter[9] ),
    .Y(_0468_));
 sg13g2_xor2_1 _1296_ (.B(_0468_),
    .A(\vga_image_generator.counter[11] ),
    .X(_0469_));
 sg13g2_nor2_1 _1297_ (.A(net27),
    .B(_0469_),
    .Y(_0077_));
 sg13g2_inv_1 _1298_ (.Y(_0470_),
    .A(\vga_image_generator.counter[12] ));
 sg13g2_nand4_1 _1299_ (.B(\vga_image_generator.counter[10] ),
    .C(\vga_image_generator.counter[11] ),
    .A(\vga_image_generator.counter[9] ),
    .Y(_0471_),
    .D(_0465_));
 sg13g2_xnor2_1 _1300_ (.Y(_0472_),
    .A(_0470_),
    .B(_0471_));
 sg13g2_nor2_1 _1301_ (.A(net27),
    .B(_0472_),
    .Y(_0078_));
 sg13g2_nand4_1 _1302_ (.B(\vga_image_generator.counter[9] ),
    .C(\vga_image_generator.counter[10] ),
    .A(\vga_image_generator.counter[8] ),
    .Y(_0473_),
    .D(\vga_image_generator.counter[11] ));
 sg13g2_nor4_2 _1303_ (.A(_0459_),
    .B(_0470_),
    .C(_0462_),
    .Y(_0474_),
    .D(_0473_));
 sg13g2_xnor2_1 _1304_ (.Y(_0475_),
    .A(\vga_image_generator.counter[13] ),
    .B(_0474_));
 sg13g2_nor2_1 _1305_ (.A(net27),
    .B(_0475_),
    .Y(_0079_));
 sg13g2_nand2_1 _1306_ (.Y(_0476_),
    .A(\vga_image_generator.counter[13] ),
    .B(_0474_));
 sg13g2_xor2_1 _1307_ (.B(_0476_),
    .A(\vga_image_generator.counter[14] ),
    .X(_0477_));
 sg13g2_nor2_1 _1308_ (.A(net27),
    .B(_0477_),
    .Y(_0080_));
 sg13g2_buf_1 _1309_ (.A(net48),
    .X(_0478_));
 sg13g2_and3_1 _1310_ (.X(_0479_),
    .A(\vga_image_generator.counter[13] ),
    .B(\vga_image_generator.counter[14] ),
    .C(_0474_));
 sg13g2_xnor2_1 _1311_ (.Y(_0480_),
    .A(\vga_image_generator.counter[15] ),
    .B(_0479_));
 sg13g2_nor2_1 _1312_ (.A(net26),
    .B(_0480_),
    .Y(_0081_));
 sg13g2_and2_1 _1313_ (.A(\vga_image_generator.counter[15] ),
    .B(_0479_),
    .X(_0481_));
 sg13g2_buf_8 _1314_ (.A(_0481_),
    .X(_0482_));
 sg13g2_xnor2_1 _1315_ (.Y(_0483_),
    .A(\vga_image_generator.counter[16] ),
    .B(_0482_));
 sg13g2_nor2_1 _1316_ (.A(net26),
    .B(_0483_),
    .Y(_0082_));
 sg13g2_nand2_1 _1317_ (.Y(_0484_),
    .A(\vga_image_generator.counter[16] ),
    .B(_0482_));
 sg13g2_xor2_1 _1318_ (.B(_0484_),
    .A(\vga_image_generator.counter[17] ),
    .X(_0485_));
 sg13g2_nor2_1 _1319_ (.A(net26),
    .B(_0485_),
    .Y(_0083_));
 sg13g2_nand3_1 _1320_ (.B(\vga_image_generator.counter[17] ),
    .C(_0482_),
    .A(\vga_image_generator.counter[16] ),
    .Y(_0486_));
 sg13g2_xor2_1 _1321_ (.B(_0486_),
    .A(\vga_image_generator.counter[18] ),
    .X(_0487_));
 sg13g2_nor2_1 _1322_ (.A(net26),
    .B(_0487_),
    .Y(_0084_));
 sg13g2_nand4_1 _1323_ (.B(\vga_image_generator.counter[17] ),
    .C(\vga_image_generator.counter[18] ),
    .A(\vga_image_generator.counter[16] ),
    .Y(_0488_),
    .D(_0482_));
 sg13g2_xor2_1 _1324_ (.B(_0488_),
    .A(\vga_image_generator.counter[19] ),
    .X(_0489_));
 sg13g2_nor2_1 _1325_ (.A(net26),
    .B(_0489_),
    .Y(_0085_));
 sg13g2_xnor2_1 _1326_ (.Y(_0490_),
    .A(\vga_image_generator.counter[1] ),
    .B(\vga_image_generator.counter[0] ));
 sg13g2_nor2_1 _1327_ (.A(net26),
    .B(_0490_),
    .Y(_0086_));
 sg13g2_nand2_1 _1328_ (.Y(_0491_),
    .A(\vga_image_generator.counter[15] ),
    .B(_0479_));
 sg13g2_nand4_1 _1329_ (.B(\vga_image_generator.counter[17] ),
    .C(\vga_image_generator.counter[18] ),
    .A(\vga_image_generator.counter[16] ),
    .Y(_0492_),
    .D(\vga_image_generator.counter[19] ));
 sg13g2_nor2_1 _1330_ (.A(_0491_),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_xnor2_1 _1331_ (.Y(_0494_),
    .A(_0424_),
    .B(_0493_));
 sg13g2_nor2_1 _1332_ (.A(_0478_),
    .B(_0494_),
    .Y(_0087_));
 sg13g2_nand4_1 _1333_ (.B(\vga_image_generator.counter[13] ),
    .C(\vga_image_generator.counter[14] ),
    .A(_0424_),
    .Y(_0495_),
    .D(\vga_image_generator.counter[15] ));
 sg13g2_nor2_1 _1334_ (.A(_0492_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_and2_1 _1335_ (.A(_0474_),
    .B(_0496_),
    .X(_0497_));
 sg13g2_buf_2 _1336_ (.A(_0497_),
    .X(_0498_));
 sg13g2_xnor2_1 _1337_ (.Y(_0499_),
    .A(_0423_),
    .B(_0498_));
 sg13g2_nor2_1 _1338_ (.A(net26),
    .B(_0499_),
    .Y(_0088_));
 sg13g2_nand2_1 _1339_ (.Y(_0500_),
    .A(_0423_),
    .B(_0498_));
 sg13g2_xnor2_1 _1340_ (.Y(_0501_),
    .A(_0439_),
    .B(_0500_));
 sg13g2_nor2_1 _1341_ (.A(_0478_),
    .B(_0501_),
    .Y(_0089_));
 sg13g2_nand3_1 _1342_ (.B(_0425_),
    .C(_0498_),
    .A(_0423_),
    .Y(_0502_));
 sg13g2_xnor2_1 _1343_ (.Y(_0503_),
    .A(_0430_),
    .B(_0502_));
 sg13g2_nor2_1 _1344_ (.A(net26),
    .B(_0503_),
    .Y(_0090_));
 sg13g2_buf_1 _1345_ (.A(_0350_),
    .X(_0504_));
 sg13g2_or2_1 _1346_ (.X(_0505_),
    .B(_0500_),
    .A(_0433_));
 sg13g2_xnor2_1 _1347_ (.Y(_0506_),
    .A(_0418_),
    .B(_0505_));
 sg13g2_nor2_1 _1348_ (.A(net25),
    .B(_0506_),
    .Y(_0091_));
 sg13g2_o21ai_1 _1349_ (.B1(_0419_),
    .Y(_0507_),
    .A1(_0418_),
    .A2(_0505_));
 sg13g2_inv_1 _1350_ (.Y(_0508_),
    .A(_0423_));
 sg13g2_nor3_1 _1351_ (.A(_0508_),
    .B(_0418_),
    .C(_0433_),
    .Y(_0509_));
 sg13g2_nand3_1 _1352_ (.B(_0498_),
    .C(_0509_),
    .A(_0450_),
    .Y(_0510_));
 sg13g2_a21oi_1 _1353_ (.A1(_0507_),
    .A2(_0510_),
    .Y(_0092_),
    .B1(net48));
 sg13g2_and3_1 _1354_ (.X(_0511_),
    .A(_0419_),
    .B(_0498_),
    .C(_0509_));
 sg13g2_xnor2_1 _1355_ (.Y(_0512_),
    .A(\vga_image_generator.counter[26] ),
    .B(_0511_));
 sg13g2_nor2_1 _1356_ (.A(net25),
    .B(_0512_),
    .Y(_0093_));
 sg13g2_nand2_1 _1357_ (.Y(_0513_),
    .A(\vga_image_generator.counter[26] ),
    .B(_0511_));
 sg13g2_xor2_1 _1358_ (.B(_0513_),
    .A(\vga_image_generator.counter[27] ),
    .X(_0514_));
 sg13g2_nor2_1 _1359_ (.A(_0504_),
    .B(_0514_),
    .Y(_0094_));
 sg13g2_nand2_1 _1360_ (.Y(_0515_),
    .A(\vga_image_generator.counter[1] ),
    .B(\vga_image_generator.counter[0] ));
 sg13g2_xor2_1 _1361_ (.B(_0515_),
    .A(\vga_image_generator.counter[2] ),
    .X(_0516_));
 sg13g2_nor2_1 _1362_ (.A(net25),
    .B(_0516_),
    .Y(_0095_));
 sg13g2_nand3_1 _1363_ (.B(\vga_image_generator.counter[0] ),
    .C(\vga_image_generator.counter[2] ),
    .A(\vga_image_generator.counter[1] ),
    .Y(_0517_));
 sg13g2_xor2_1 _1364_ (.B(_0517_),
    .A(\vga_image_generator.counter[3] ),
    .X(_0518_));
 sg13g2_nor2_1 _1365_ (.A(_0504_),
    .B(_0518_),
    .Y(_0096_));
 sg13g2_xnor2_1 _1366_ (.Y(_0519_),
    .A(\vga_image_generator.counter[4] ),
    .B(_0461_));
 sg13g2_nor2_1 _1367_ (.A(net25),
    .B(_0519_),
    .Y(_0097_));
 sg13g2_nand2_1 _1368_ (.Y(_0520_),
    .A(\vga_image_generator.counter[4] ),
    .B(_0461_));
 sg13g2_xor2_1 _1369_ (.B(_0520_),
    .A(\vga_image_generator.counter[5] ),
    .X(_0521_));
 sg13g2_nor2_1 _1370_ (.A(net25),
    .B(_0521_),
    .Y(_0098_));
 sg13g2_nand3_1 _1371_ (.B(\vga_image_generator.counter[5] ),
    .C(_0461_),
    .A(\vga_image_generator.counter[4] ),
    .Y(_0522_));
 sg13g2_xor2_1 _1372_ (.B(_0522_),
    .A(\vga_image_generator.counter[6] ),
    .X(_0523_));
 sg13g2_nor2_1 _1373_ (.A(net25),
    .B(_0523_),
    .Y(_0099_));
 sg13g2_xnor2_1 _1374_ (.Y(_0524_),
    .A(_0459_),
    .B(_0462_));
 sg13g2_nor2_1 _1375_ (.A(net25),
    .B(_0524_),
    .Y(_0100_));
 sg13g2_xnor2_1 _1376_ (.Y(_0525_),
    .A(\vga_image_generator.counter[8] ),
    .B(_0463_));
 sg13g2_nor2_1 _1377_ (.A(net25),
    .B(_0525_),
    .Y(_0101_));
 sg13g2_xnor2_1 _1378_ (.Y(_0526_),
    .A(\vga_image_generator.counter[9] ),
    .B(_0465_));
 sg13g2_nor2_1 _1379_ (.A(net48),
    .B(_0526_),
    .Y(_0102_));
 sg13g2_buf_1 _1380_ (.A(ui_in[1]),
    .X(_0527_));
 sg13g2_buf_2 _1381_ (.A(net66),
    .X(_0528_));
 sg13g2_and2_1 _1382_ (.A(net163),
    .B(\BNC_x[0] ),
    .X(net3));
 sg13g2_and2_1 _1383_ (.A(net163),
    .B(\BNC_x[2] ),
    .X(net4));
 sg13g2_and2_1 _1384_ (.A(net163),
    .B(\BNC_x[4] ),
    .X(net5));
 sg13g2_and2_1 _1385_ (.A(_0528_),
    .B(\BNC_x[6] ),
    .X(net6));
 sg13g2_and2_1 _1386_ (.A(net163),
    .B(\BNC_x[1] ),
    .X(net7));
 sg13g2_and2_1 _1387_ (.A(net163),
    .B(\BNC_x[3] ),
    .X(net8));
 sg13g2_and2_1 _1388_ (.A(net163),
    .B(\BNC_x[5] ),
    .X(net9));
 sg13g2_and2_1 _1389_ (.A(net163),
    .B(\BNC_x[7] ),
    .X(net10));
 sg13g2_buf_1 _1390_ (.A(net2),
    .X(_0529_));
 sg13g2_inv_1 _1391_ (.Y(_0530_),
    .A(net65));
 sg13g2_nor2_1 _1392_ (.A(_0218_),
    .B(net66),
    .Y(_0531_));
 sg13g2_a21oi_1 _1393_ (.A1(\BNC_y[0] ),
    .A2(_0527_),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_nor4_2 _1394_ (.A(net59),
    .B(net58),
    .C(_0164_),
    .Y(_0533_),
    .D(_0165_));
 sg13g2_inv_1 _1395_ (.Y(_0534_),
    .A(_0533_));
 sg13g2_o21ai_1 _1396_ (.B1(_0156_),
    .Y(_0535_),
    .A1(_0319_),
    .A2(_0322_));
 sg13g2_nor2b_1 _1397_ (.A(_0020_),
    .B_N(_0535_),
    .Y(_0536_));
 sg13g2_nand2_1 _1398_ (.Y(_0537_),
    .A(_0155_),
    .B(net63));
 sg13g2_nor2_2 _1399_ (.A(net61),
    .B(net60),
    .Y(_0538_));
 sg13g2_inv_1 _1400_ (.Y(_0539_),
    .A(net58));
 sg13g2_o21ai_1 _1401_ (.B1(_0539_),
    .Y(_0540_),
    .A1(_0537_),
    .A2(_0538_));
 sg13g2_nor2_2 _1402_ (.A(_0163_),
    .B(_0165_),
    .Y(_0541_));
 sg13g2_nand3_1 _1403_ (.B(_0540_),
    .C(_0541_),
    .A(net59),
    .Y(_0542_));
 sg13g2_o21ai_1 _1404_ (.B1(_0542_),
    .Y(_0543_),
    .A1(_0534_),
    .A2(_0536_));
 sg13g2_and2_1 _1405_ (.A(_0182_),
    .B(net55),
    .X(_0544_));
 sg13g2_buf_2 _1406_ (.A(_0544_),
    .X(_0545_));
 sg13g2_or2_1 _1407_ (.X(_0546_),
    .B(_0191_),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_buf_1 _1408_ (.A(_0546_),
    .X(_0547_));
 sg13g2_a21oi_2 _1409_ (.B1(net35),
    .Y(_0548_),
    .A2(_0547_),
    .A1(net36));
 sg13g2_nand2_1 _1410_ (.Y(_0549_),
    .A(_0545_),
    .B(_0548_));
 sg13g2_nand2b_1 _1411_ (.Y(_0550_),
    .B(_0180_),
    .A_N(_0194_));
 sg13g2_nor2_1 _1412_ (.A(_0547_),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_nand2b_1 _1413_ (.Y(_0552_),
    .B(net31),
    .A_N(net30));
 sg13g2_nor2_1 _1414_ (.A(_0389_),
    .B(_0552_),
    .Y(_0553_));
 sg13g2_nand2_2 _1415_ (.Y(_0554_),
    .A(_0181_),
    .B(_0195_));
 sg13g2_nand2_1 _1416_ (.Y(_0555_),
    .A(_0393_),
    .B(_0394_));
 sg13g2_a22oi_1 _1417_ (.Y(_0556_),
    .B1(_0554_),
    .B2(_0555_),
    .A2(_0553_),
    .A1(_0551_));
 sg13g2_nand2b_2 _1418_ (.Y(_0557_),
    .B(\hvsync_gen.hpos[6] ),
    .A_N(_0191_));
 sg13g2_nor2_2 _1419_ (.A(_0550_),
    .B(_0557_),
    .Y(_0558_));
 sg13g2_nor4_1 _1420_ (.A(net31),
    .B(_0393_),
    .C(_0190_),
    .D(_0332_),
    .Y(_0559_));
 sg13g2_nand2b_2 _1421_ (.Y(_0560_),
    .B(_0180_),
    .A_N(_0191_));
 sg13g2_nand2b_1 _1422_ (.Y(_0561_),
    .B(net54),
    .A_N(net49));
 sg13g2_nor4_1 _1423_ (.A(net35),
    .B(_0190_),
    .C(_0560_),
    .D(_0561_),
    .Y(_0562_));
 sg13g2_a21oi_1 _1424_ (.A1(_0558_),
    .A2(_0559_),
    .Y(_0563_),
    .B1(_0562_));
 sg13g2_o21ai_1 _1425_ (.B1(_0563_),
    .Y(_0564_),
    .A1(_0549_),
    .A2(_0556_));
 sg13g2_nor2_1 _1426_ (.A(net31),
    .B(_0398_),
    .Y(_0565_));
 sg13g2_a22oi_1 _1427_ (.Y(_0566_),
    .B1(_0554_),
    .B2(net31),
    .A2(_0551_),
    .A1(_0565_));
 sg13g2_nand3_1 _1428_ (.B(_0545_),
    .C(_0548_),
    .A(net30),
    .Y(_0567_));
 sg13g2_nand2b_1 _1429_ (.Y(_0568_),
    .B(net31),
    .A_N(_0024_));
 sg13g2_nor3_1 _1430_ (.A(_0190_),
    .B(_0388_),
    .C(_0552_),
    .Y(_0569_));
 sg13g2_a22oi_1 _1431_ (.Y(_0570_),
    .B1(_0569_),
    .B2(_0558_),
    .A2(_0568_),
    .A1(_0562_));
 sg13g2_o21ai_1 _1432_ (.B1(_0570_),
    .Y(_0571_),
    .A1(_0566_),
    .A2(_0567_));
 sg13g2_or2_1 _1433_ (.X(_0572_),
    .B(_0165_),
    .A(_0163_));
 sg13g2_buf_1 _1434_ (.A(_0572_),
    .X(_0573_));
 sg13g2_nor2b_1 _1435_ (.A(net60),
    .B_N(net63),
    .Y(_0574_));
 sg13g2_o21ai_1 _1436_ (.B1(net61),
    .Y(_0575_),
    .A1(\hvsync_gen.vpos[1] ),
    .A2(net62));
 sg13g2_and2_1 _1437_ (.A(_0574_),
    .B(_0575_),
    .X(_0576_));
 sg13g2_a21oi_1 _1438_ (.A1(_0360_),
    .A2(_0362_),
    .Y(_0577_),
    .B1(_0576_));
 sg13g2_nand3b_1 _1439_ (.B(_0166_),
    .C(_0155_),
    .Y(_0578_),
    .A_N(net58));
 sg13g2_nor3_1 _1440_ (.A(_0573_),
    .B(_0577_),
    .C(_0578_),
    .Y(_0579_));
 sg13g2_a22oi_1 _1441_ (.Y(_0580_),
    .B1(_0571_),
    .B2(_0579_),
    .A2(_0564_),
    .A1(_0543_));
 sg13g2_or2_1 _1442_ (.X(_0581_),
    .B(_0550_),
    .A(_0547_));
 sg13g2_buf_1 _1443_ (.A(_0581_),
    .X(_0582_));
 sg13g2_nor2_1 _1444_ (.A(_0182_),
    .B(net54),
    .Y(_0583_));
 sg13g2_nor2_1 _1445_ (.A(_0191_),
    .B(_0194_),
    .Y(_0584_));
 sg13g2_nor2_1 _1446_ (.A(_0180_),
    .B(_0194_),
    .Y(_0585_));
 sg13g2_a21oi_2 _1447_ (.B1(_0585_),
    .Y(_0586_),
    .A2(_0584_),
    .A1(_0583_));
 sg13g2_o21ai_1 _1448_ (.B1(_0586_),
    .Y(_0587_),
    .A1(net29),
    .A2(_0582_));
 sg13g2_nor2_1 _1449_ (.A(net51),
    .B(_0330_),
    .Y(_0588_));
 sg13g2_nor2b_2 _1450_ (.A(net55),
    .B_N(_0182_),
    .Y(_0589_));
 sg13g2_nand4_1 _1451_ (.B(_0551_),
    .C(_0588_),
    .A(_0336_),
    .Y(_0590_),
    .D(_0589_));
 sg13g2_or2_1 _1452_ (.X(_0591_),
    .B(_0330_),
    .A(_0329_));
 sg13g2_buf_1 _1453_ (.A(_0591_),
    .X(_0592_));
 sg13g2_nand3_1 _1454_ (.B(_0586_),
    .C(_0592_),
    .A(_0336_),
    .Y(_0593_));
 sg13g2_nand3_1 _1455_ (.B(_0590_),
    .C(_0593_),
    .A(_0587_),
    .Y(_0594_));
 sg13g2_nor2_1 _1456_ (.A(_0020_),
    .B(_0541_),
    .Y(_0595_));
 sg13g2_nor2_1 _1457_ (.A(net56),
    .B(_0355_),
    .Y(_0596_));
 sg13g2_o21ai_1 _1458_ (.B1(_0360_),
    .Y(_0597_),
    .A1(_0021_),
    .A2(_0596_));
 sg13g2_nand2_1 _1459_ (.Y(_0598_),
    .A(net33),
    .B(_0533_));
 sg13g2_a21oi_1 _1460_ (.A1(_0595_),
    .A2(_0597_),
    .Y(_0599_),
    .B1(_0598_));
 sg13g2_nand2b_1 _1461_ (.Y(_0600_),
    .B(net54),
    .A_N(net46));
 sg13g2_nor3_1 _1462_ (.A(net35),
    .B(_0560_),
    .C(_0600_),
    .Y(_0601_));
 sg13g2_and2_1 _1463_ (.A(net50),
    .B(net55),
    .X(_0602_));
 sg13g2_and2_1 _1464_ (.A(net49),
    .B(_0184_),
    .X(_0603_));
 sg13g2_a21oi_1 _1465_ (.A1(_0592_),
    .A2(_0602_),
    .Y(_0604_),
    .B1(_0603_));
 sg13g2_a21oi_1 _1466_ (.A1(_0601_),
    .A2(_0604_),
    .Y(_0605_),
    .B1(_0548_));
 sg13g2_nor2_1 _1467_ (.A(net60),
    .B(net63),
    .Y(_0606_));
 sg13g2_nor2b_1 _1468_ (.A(net57),
    .B_N(net62),
    .Y(_0607_));
 sg13g2_a22oi_1 _1469_ (.Y(_0608_),
    .B1(_0606_),
    .B2(_0607_),
    .A2(_0573_),
    .A1(net57));
 sg13g2_or2_1 _1470_ (.X(_0609_),
    .B(_0606_),
    .A(_0541_));
 sg13g2_o21ai_1 _1471_ (.B1(_0609_),
    .Y(_0610_),
    .A1(_0171_),
    .A2(_0608_));
 sg13g2_nor2b_1 _1472_ (.A(_0605_),
    .B_N(_0610_),
    .Y(_0611_));
 sg13g2_nand3_1 _1473_ (.B(_0599_),
    .C(_0611_),
    .A(_0594_),
    .Y(_0612_));
 sg13g2_nand2_1 _1474_ (.Y(_0613_),
    .A(net33),
    .B(_0385_));
 sg13g2_nor2_1 _1475_ (.A(net44),
    .B(net36),
    .Y(_0614_));
 sg13g2_nor2_1 _1476_ (.A(_0195_),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_nor3_1 _1477_ (.A(_0165_),
    .B(net2),
    .C(_0615_),
    .Y(_0616_));
 sg13g2_nor4_1 _1478_ (.A(\hvsync_gen.vpos[1] ),
    .B(net61),
    .C(net60),
    .D(_0155_),
    .Y(_0617_));
 sg13g2_nor4_1 _1479_ (.A(_0168_),
    .B(_0320_),
    .C(_0573_),
    .D(_0617_),
    .Y(_0618_));
 sg13g2_nand2b_1 _1480_ (.Y(_0619_),
    .B(_0388_),
    .A_N(_0024_));
 sg13g2_nand2b_1 _1481_ (.Y(_0620_),
    .B(net46),
    .A_N(net29));
 sg13g2_or2_1 _1482_ (.X(_0621_),
    .B(_0334_),
    .A(net50));
 sg13g2_nor2_1 _1483_ (.A(_0620_),
    .B(_0621_),
    .Y(_0622_));
 sg13g2_nand4_1 _1484_ (.B(_0618_),
    .C(_0619_),
    .A(_0558_),
    .Y(_0623_),
    .D(_0622_));
 sg13g2_nand3_1 _1485_ (.B(_0616_),
    .C(_0623_),
    .A(_0613_),
    .Y(_0624_));
 sg13g2_nand4_1 _1486_ (.B(_0407_),
    .C(_0592_),
    .A(_0391_),
    .Y(_0625_),
    .D(_0603_));
 sg13g2_nor2_2 _1487_ (.A(_0183_),
    .B(net29),
    .Y(_0626_));
 sg13g2_nor2_2 _1488_ (.A(net50),
    .B(net49),
    .Y(_0627_));
 sg13g2_nand3b_1 _1489_ (.B(_0626_),
    .C(_0627_),
    .Y(_0628_),
    .A_N(_0188_));
 sg13g2_nand2b_1 _1490_ (.Y(_0629_),
    .B(net33),
    .A_N(net35));
 sg13g2_nor4_1 _1491_ (.A(_0168_),
    .B(_0573_),
    .C(_0560_),
    .D(_0629_),
    .Y(_0630_));
 sg13g2_nand3_1 _1492_ (.B(_0628_),
    .C(_0630_),
    .A(_0625_),
    .Y(_0631_));
 sg13g2_a21o_1 _1493_ (.A2(net47),
    .A1(net57),
    .B1(net56),
    .X(_0632_));
 sg13g2_nor3_1 _1494_ (.A(net57),
    .B(net62),
    .C(net47),
    .Y(_0633_));
 sg13g2_a22oi_1 _1495_ (.Y(_0634_),
    .B1(_0633_),
    .B2(_0574_),
    .A2(_0632_),
    .A1(_0360_));
 sg13g2_a21o_1 _1496_ (.A2(_0627_),
    .A1(_0398_),
    .B1(_0186_),
    .X(_0635_));
 sg13g2_nand3_1 _1497_ (.B(_0333_),
    .C(net30),
    .A(net51),
    .Y(_0636_));
 sg13g2_nand3b_1 _1498_ (.B(_0626_),
    .C(_0636_),
    .Y(_0637_),
    .A_N(net45));
 sg13g2_nand4_1 _1499_ (.B(_0630_),
    .C(_0635_),
    .A(_0576_),
    .Y(_0638_),
    .D(_0637_));
 sg13g2_o21ai_1 _1500_ (.B1(_0638_),
    .Y(_0639_),
    .A1(_0631_),
    .A2(_0634_));
 sg13g2_nor2b_1 _1501_ (.A(_0021_),
    .B_N(_0575_),
    .Y(_0640_));
 sg13g2_a21oi_1 _1502_ (.A1(_0021_),
    .A2(_0355_),
    .Y(_0641_),
    .B1(net56));
 sg13g2_a21oi_1 _1503_ (.A1(_0595_),
    .A2(_0640_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_nand2_1 _1504_ (.Y(_0643_),
    .A(_0393_),
    .B(_0589_));
 sg13g2_nor4_1 _1505_ (.A(net51),
    .B(_0391_),
    .C(_0582_),
    .D(_0643_),
    .Y(_0644_));
 sg13g2_o21ai_1 _1506_ (.B1(_0355_),
    .Y(_0645_),
    .A1(_0020_),
    .A2(_0541_));
 sg13g2_nand4_1 _1507_ (.B(_0533_),
    .C(_0586_),
    .A(_0156_),
    .Y(_0646_),
    .D(_0645_));
 sg13g2_nor2_1 _1508_ (.A(_0332_),
    .B(_0401_),
    .Y(_0647_));
 sg13g2_a21o_1 _1509_ (.A2(net54),
    .A1(net46),
    .B1(net44),
    .X(_0648_));
 sg13g2_a21oi_1 _1510_ (.A1(net36),
    .A2(_0648_),
    .Y(_0649_),
    .B1(net35));
 sg13g2_and3_1 _1511_ (.X(_0650_),
    .A(_0333_),
    .B(net30),
    .C(_0184_));
 sg13g2_nand3_1 _1512_ (.B(_0650_),
    .C(_0547_),
    .A(net36),
    .Y(_0651_));
 sg13g2_a22oi_1 _1513_ (.Y(_0652_),
    .B1(_0649_),
    .B2(_0651_),
    .A2(_0647_),
    .A1(_0601_));
 sg13g2_nor4_1 _1514_ (.A(_0642_),
    .B(_0644_),
    .C(_0646_),
    .D(_0652_),
    .Y(_0653_));
 sg13g2_nor3_1 _1515_ (.A(_0624_),
    .B(_0639_),
    .C(_0653_),
    .Y(_0654_));
 sg13g2_nand3_1 _1516_ (.B(_0612_),
    .C(_0654_),
    .A(_0580_),
    .Y(_0655_));
 sg13g2_a21oi_1 _1517_ (.A1(_0336_),
    .A2(_0592_),
    .Y(_0656_),
    .B1(net29));
 sg13g2_nor2b_1 _1518_ (.A(_0182_),
    .B_N(\hvsync_gen.hpos[4] ),
    .Y(_0657_));
 sg13g2_buf_1 _1519_ (.A(_0657_),
    .X(_0658_));
 sg13g2_nor2b_1 _1520_ (.A(net50),
    .B_N(\hvsync_gen.hpos[3] ),
    .Y(_0659_));
 sg13g2_buf_2 _1521_ (.A(_0659_),
    .X(_0660_));
 sg13g2_nand2_1 _1522_ (.Y(_0661_),
    .A(net20),
    .B(_0660_));
 sg13g2_nor3_1 _1523_ (.A(_0586_),
    .B(_0592_),
    .C(_0661_),
    .Y(_0662_));
 sg13g2_a21oi_1 _1524_ (.A1(_0586_),
    .A2(_0656_),
    .Y(_0663_),
    .B1(_0662_));
 sg13g2_or4_1 _1525_ (.A(_0396_),
    .B(_0025_),
    .C(_0585_),
    .D(_0586_),
    .X(_0664_));
 sg13g2_o21ai_1 _1526_ (.B1(_0664_),
    .Y(_0665_),
    .A1(_0582_),
    .A2(_0663_));
 sg13g2_nor2b_1 _1527_ (.A(net49),
    .B_N(\hvsync_gen.hpos[2] ),
    .Y(_0666_));
 sg13g2_buf_2 _1528_ (.A(_0666_),
    .X(_0667_));
 sg13g2_nand3_1 _1529_ (.B(_0667_),
    .C(_0588_),
    .A(net20),
    .Y(_0668_));
 sg13g2_nand2b_1 _1530_ (.Y(_0669_),
    .B(_0668_),
    .A_N(_0605_));
 sg13g2_a21oi_1 _1531_ (.A1(_0660_),
    .A2(_0588_),
    .Y(_0670_),
    .B1(_0025_));
 sg13g2_nor2b_1 _1532_ (.A(_0548_),
    .B_N(net46),
    .Y(_0671_));
 sg13g2_o21ai_1 _1533_ (.B1(_0671_),
    .Y(_0672_),
    .A1(net29),
    .A2(_0670_));
 sg13g2_and3_1 _1534_ (.X(_0673_),
    .A(_0558_),
    .B(_0669_),
    .C(_0672_));
 sg13g2_nand2_1 _1535_ (.Y(_0674_),
    .A(_0368_),
    .B(net34));
 sg13g2_a21oi_1 _1536_ (.A1(net56),
    .A2(net34),
    .Y(_0675_),
    .B1(net33));
 sg13g2_o21ai_1 _1537_ (.B1(_0541_),
    .Y(_0676_),
    .A1(_0168_),
    .A2(_0675_));
 sg13g2_nand2_1 _1538_ (.Y(_0677_),
    .A(net56),
    .B(_0633_));
 sg13g2_nand2_1 _1539_ (.Y(_0678_),
    .A(_0676_),
    .B(_0677_));
 sg13g2_o21ai_1 _1540_ (.B1(_0678_),
    .Y(_0679_),
    .A1(_0596_),
    .A2(_0676_));
 sg13g2_nor4_1 _1541_ (.A(_0168_),
    .B(_0674_),
    .C(_0573_),
    .D(_0679_),
    .Y(_0680_));
 sg13g2_o21ai_1 _1542_ (.B1(_0680_),
    .Y(_0681_),
    .A1(_0665_),
    .A2(_0673_));
 sg13g2_nand4_1 _1543_ (.B(net20),
    .C(_0558_),
    .A(_0332_),
    .Y(_0682_),
    .D(_0660_));
 sg13g2_o21ai_1 _1544_ (.B1(_0682_),
    .Y(_0683_),
    .A1(_0401_),
    .A2(_0548_));
 sg13g2_nor2_1 _1545_ (.A(net30),
    .B(_0620_),
    .Y(_0684_));
 sg13g2_nand2b_1 _1546_ (.Y(_0685_),
    .B(_0388_),
    .A_N(_0568_));
 sg13g2_a21oi_1 _1547_ (.A1(_0684_),
    .A2(_0685_),
    .Y(_0686_),
    .B1(_0023_));
 sg13g2_o21ai_1 _1548_ (.B1(_0554_),
    .Y(_0687_),
    .A1(_0582_),
    .A2(_0686_));
 sg13g2_a21o_1 _1549_ (.A2(_0551_),
    .A1(_0339_),
    .B1(_0586_),
    .X(_0688_));
 sg13g2_a22oi_1 _1550_ (.Y(_0689_),
    .B1(_0687_),
    .B2(_0688_),
    .A2(_0683_),
    .A1(_0649_));
 sg13g2_nand2b_1 _1551_ (.Y(_0690_),
    .B(_0618_),
    .A_N(_0689_));
 sg13g2_nand3b_1 _1552_ (.B(_0681_),
    .C(_0690_),
    .Y(_0691_),
    .A_N(_0655_));
 sg13g2_buf_1 _1553_ (.A(_0691_),
    .X(_0692_));
 sg13g2_o21ai_1 _1554_ (.B1(_0692_),
    .Y(net11),
    .A1(_0530_),
    .A2(_0532_));
 sg13g2_mux2_1 _1555_ (.A0(\BNC_y[5] ),
    .A1(\BNC_y[2] ),
    .S(_0527_),
    .X(_0693_));
 sg13g2_nand2_1 _1556_ (.Y(_0694_),
    .A(net65),
    .B(_0693_));
 sg13g2_inv_1 _1557_ (.Y(_0695_),
    .A(_0027_));
 sg13g2_nor2b_2 _1558_ (.A(_0185_),
    .B_N(_0191_),
    .Y(_0696_));
 sg13g2_nand4_1 _1559_ (.B(\vga_image_generator.character_hold[16] ),
    .C(_0545_),
    .A(_0695_),
    .Y(_0697_),
    .D(_0696_));
 sg13g2_or2_1 _1560_ (.X(_0698_),
    .B(_0660_),
    .A(_0667_));
 sg13g2_buf_1 _1561_ (.A(_0698_),
    .X(_0699_));
 sg13g2_nand2b_1 _1562_ (.Y(_0700_),
    .B(\hvsync_gen.vpos[7] ),
    .A_N(\hvsync_gen.vpos[6] ));
 sg13g2_buf_2 _1563_ (.A(_0700_),
    .X(_0701_));
 sg13g2_nand2b_1 _1564_ (.Y(_0702_),
    .B(_0155_),
    .A_N(\hvsync_gen.vpos[3] ));
 sg13g2_nand2b_1 _1565_ (.Y(_0703_),
    .B(_0163_),
    .A_N(_0154_));
 sg13g2_nor3_2 _1566_ (.A(_0701_),
    .B(_0702_),
    .C(_0703_),
    .Y(_0704_));
 sg13g2_buf_2 _1567_ (.A(_0026_),
    .X(_0705_));
 sg13g2_or2_1 _1568_ (.X(_0706_),
    .B(\hvsync_gen.vpos[3] ),
    .A(net61));
 sg13g2_buf_1 _1569_ (.A(_0706_),
    .X(_0707_));
 sg13g2_or4_1 _1570_ (.A(_0705_),
    .B(_0537_),
    .C(_0707_),
    .D(_0701_),
    .X(_0708_));
 sg13g2_nor2b_1 _1571_ (.A(net58),
    .B_N(_0166_),
    .Y(_0709_));
 sg13g2_nor2b_1 _1572_ (.A(\hvsync_gen.vpos[4] ),
    .B_N(_0163_),
    .Y(_0710_));
 sg13g2_nand4_1 _1573_ (.B(net33),
    .C(_0709_),
    .A(net56),
    .Y(_0711_),
    .D(_0710_));
 sg13g2_nand3_1 _1574_ (.B(_0711_),
    .C(_0699_),
    .A(_0708_),
    .Y(_0712_));
 sg13g2_o21ai_1 _1575_ (.B1(_0712_),
    .Y(_0713_),
    .A1(_0699_),
    .A2(_0704_));
 sg13g2_or2_1 _1576_ (.X(_0714_),
    .B(_0713_),
    .A(_0697_));
 sg13g2_nand2_1 _1577_ (.Y(_0715_),
    .A(_0399_),
    .B(net20));
 sg13g2_nor3_2 _1578_ (.A(_0705_),
    .B(_0174_),
    .C(_0701_),
    .Y(_0716_));
 sg13g2_nand2_1 _1579_ (.Y(_0717_),
    .A(_0160_),
    .B(_0716_));
 sg13g2_nand2_1 _1580_ (.Y(_0718_),
    .A(_0667_),
    .B(_0589_));
 sg13g2_nand2b_1 _1581_ (.Y(_0719_),
    .B(_0704_),
    .A_N(_0718_));
 sg13g2_nand2b_1 _1582_ (.Y(_0720_),
    .B(_0181_),
    .A_N(_0557_));
 sg13g2_or2_1 _1583_ (.X(_0721_),
    .B(_0720_),
    .A(_0179_));
 sg13g2_buf_1 _1584_ (.A(_0721_),
    .X(_0722_));
 sg13g2_a221oi_1 _1585_ (.B2(_0719_),
    .C1(_0722_),
    .B1(_0717_),
    .A1(_0643_),
    .Y(_0723_),
    .A2(_0715_));
 sg13g2_nor3_1 _1586_ (.A(_0554_),
    .B(_0557_),
    .C(_0661_),
    .Y(_0724_));
 sg13g2_a22oi_1 _1587_ (.Y(_0725_),
    .B1(_0589_),
    .B2(_0627_),
    .A2(net20),
    .A1(_0336_));
 sg13g2_a21oi_1 _1588_ (.A1(_0708_),
    .A2(_0711_),
    .Y(_0726_),
    .B1(_0725_));
 sg13g2_nor2_1 _1589_ (.A(_0179_),
    .B(_0720_),
    .Y(_0727_));
 sg13g2_buf_1 _1590_ (.A(ui_in[3]),
    .X(_0728_));
 sg13g2_inv_1 _1591_ (.Y(_0729_),
    .A(net64));
 sg13g2_a221oi_1 _1592_ (.B2(_0727_),
    .C1(_0729_),
    .B1(_0726_),
    .A1(_0704_),
    .Y(_0730_),
    .A2(_0724_));
 sg13g2_nand2b_1 _1593_ (.Y(_0731_),
    .B(_0730_),
    .A_N(_0723_));
 sg13g2_inv_1 _1594_ (.Y(_0732_),
    .A(_0705_));
 sg13g2_nand2b_1 _1595_ (.Y(_0733_),
    .B(_0732_),
    .A_N(_0578_));
 sg13g2_nor2_1 _1596_ (.A(_0707_),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_o21ai_1 _1597_ (.B1(_0643_),
    .Y(_0735_),
    .A1(_0715_),
    .A2(_0708_));
 sg13g2_nand3_1 _1598_ (.B(_0156_),
    .C(_0709_),
    .A(_0732_),
    .Y(_0736_));
 sg13g2_a21oi_1 _1599_ (.A1(_0661_),
    .A2(_0718_),
    .Y(_0737_),
    .B1(_0736_));
 sg13g2_a21oi_1 _1600_ (.A1(_0734_),
    .A2(_0735_),
    .Y(_0738_),
    .B1(_0737_));
 sg13g2_nor4_2 _1601_ (.A(net35),
    .B(_0705_),
    .C(_0174_),
    .Y(_0739_),
    .D(_0701_));
 sg13g2_nand3_1 _1602_ (.B(_0603_),
    .C(_0614_),
    .A(_0538_),
    .Y(_0740_));
 sg13g2_nor2_1 _1603_ (.A(_0600_),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_a21oi_1 _1604_ (.A1(_0739_),
    .A2(_0741_),
    .Y(_0742_),
    .B1(net64));
 sg13g2_o21ai_1 _1605_ (.B1(_0742_),
    .Y(_0743_),
    .A1(_0722_),
    .A2(_0738_));
 sg13g2_nand3_1 _1606_ (.B(_0731_),
    .C(_0743_),
    .A(\vga_image_generator.character_hold[3] ),
    .Y(_0744_));
 sg13g2_o21ai_1 _1607_ (.B1(_0661_),
    .Y(_0745_),
    .A1(_0728_),
    .A2(_0718_));
 sg13g2_nor3_1 _1608_ (.A(net35),
    .B(_0707_),
    .C(_0643_),
    .Y(_0746_));
 sg13g2_a21o_1 _1609_ (.A2(_0745_),
    .A1(_0178_),
    .B1(_0746_),
    .X(_0747_));
 sg13g2_nor2_1 _1610_ (.A(_0327_),
    .B(_0547_),
    .Y(_0748_));
 sg13g2_nand4_1 _1611_ (.B(_0747_),
    .C(_0716_),
    .A(\vga_image_generator.character_hold[1] ),
    .Y(_0749_),
    .D(_0748_));
 sg13g2_and2_1 _1612_ (.A(_0181_),
    .B(_0696_),
    .X(_0750_));
 sg13g2_nor4_1 _1613_ (.A(_0701_),
    .B(_0621_),
    .C(_0702_),
    .D(_0703_),
    .Y(_0751_));
 sg13g2_and4_1 _1614_ (.A(_0159_),
    .B(net33),
    .C(_0709_),
    .D(_0710_),
    .X(_0752_));
 sg13g2_and2_1 _1615_ (.A(_0159_),
    .B(net63),
    .X(_0753_));
 sg13g2_nor2_1 _1616_ (.A(net47),
    .B(_0753_),
    .Y(_0754_));
 sg13g2_nor2_2 _1617_ (.A(_0705_),
    .B(_0578_),
    .Y(_0755_));
 sg13g2_a22oi_1 _1618_ (.Y(_0756_),
    .B1(_0754_),
    .B2(_0755_),
    .A2(_0752_),
    .A1(_0650_));
 sg13g2_nand2b_1 _1619_ (.Y(_0757_),
    .B(_0756_),
    .A_N(_0751_));
 sg13g2_nand4_1 _1620_ (.B(_0545_),
    .C(_0750_),
    .A(\vga_image_generator.character_hold[6] ),
    .Y(_0758_),
    .D(_0757_));
 sg13g2_nor2b_1 _1621_ (.A(net64),
    .B_N(_0178_),
    .Y(_0759_));
 sg13g2_nand2b_1 _1622_ (.Y(_0760_),
    .B(net44),
    .A_N(_0180_));
 sg13g2_or4_1 _1623_ (.A(_0399_),
    .B(net45),
    .C(_0338_),
    .D(_0760_),
    .X(_0761_));
 sg13g2_nand4_1 _1624_ (.B(_0667_),
    .C(_0752_),
    .A(net20),
    .Y(_0762_),
    .D(_0750_));
 sg13g2_o21ai_1 _1625_ (.B1(_0762_),
    .Y(_0763_),
    .A1(_0717_),
    .A2(_0761_));
 sg13g2_nand3_1 _1626_ (.B(_0759_),
    .C(_0763_),
    .A(\vga_image_generator.character_hold[5] ),
    .Y(_0764_));
 sg13g2_and3_1 _1627_ (.X(_0765_),
    .A(_0695_),
    .B(\vga_image_generator.character_hold[15] ),
    .C(_0696_));
 sg13g2_nor2b_1 _1628_ (.A(_0180_),
    .B_N(net44),
    .Y(_0766_));
 sg13g2_and4_1 _1629_ (.A(\vga_image_generator.character_hold[5] ),
    .B(_0583_),
    .C(_0716_),
    .D(_0766_),
    .X(_0767_));
 sg13g2_nand2b_1 _1630_ (.Y(_0768_),
    .B(_0328_),
    .A_N(net64));
 sg13g2_nand3_1 _1631_ (.B(_0660_),
    .C(_0768_),
    .A(_0396_),
    .Y(_0769_));
 sg13g2_nand3_1 _1632_ (.B(net64),
    .C(_0667_),
    .A(net29),
    .Y(_0770_));
 sg13g2_nand2_1 _1633_ (.Y(_0771_),
    .A(_0769_),
    .B(_0770_));
 sg13g2_inv_1 _1634_ (.Y(_0772_),
    .A(\vga_image_generator.character_hold[11] ));
 sg13g2_nand2_1 _1635_ (.Y(_0773_),
    .A(_0538_),
    .B(_0755_));
 sg13g2_nor2b_1 _1636_ (.A(_0188_),
    .B_N(_0183_),
    .Y(_0774_));
 sg13g2_nor2_1 _1637_ (.A(_0190_),
    .B(_0561_),
    .Y(_0775_));
 sg13g2_a21oi_1 _1638_ (.A1(_0603_),
    .A2(_0774_),
    .Y(_0776_),
    .B1(_0775_));
 sg13g2_nor4_1 _1639_ (.A(_0772_),
    .B(_0560_),
    .C(_0773_),
    .D(_0776_),
    .Y(_0777_));
 sg13g2_a221oi_1 _1640_ (.B2(_0771_),
    .C1(_0777_),
    .B1(_0767_),
    .A1(_0765_),
    .Y(_0778_),
    .A2(_0737_));
 sg13g2_and4_1 _1641_ (.A(_0749_),
    .B(_0758_),
    .C(_0764_),
    .D(_0778_),
    .X(_0779_));
 sg13g2_nand2_1 _1642_ (.Y(_0780_),
    .A(_0327_),
    .B(_0696_));
 sg13g2_nand3_1 _1643_ (.B(_0160_),
    .C(_0545_),
    .A(\vga_image_generator.character_hold[16] ),
    .Y(_0781_));
 sg13g2_and3_1 _1644_ (.X(_0782_),
    .A(\vga_image_generator.character_hold[4] ),
    .B(_0407_),
    .C(_0614_));
 sg13g2_nand3_1 _1645_ (.B(_0650_),
    .C(_0782_),
    .A(_0178_),
    .Y(_0783_));
 sg13g2_o21ai_1 _1646_ (.B1(_0783_),
    .Y(_0784_),
    .A1(_0780_),
    .A2(_0781_));
 sg13g2_nand4_1 _1647_ (.B(\vga_image_generator.character_hold[14] ),
    .C(_0626_),
    .A(_0695_),
    .Y(_0785_),
    .D(_0696_));
 sg13g2_nor3_1 _1648_ (.A(_0753_),
    .B(_0733_),
    .C(_0785_),
    .Y(_0786_));
 sg13g2_o21ai_1 _1649_ (.B1(net47),
    .Y(_0787_),
    .A1(net34),
    .A2(_0699_));
 sg13g2_a21oi_1 _1650_ (.A1(_0360_),
    .A2(_0627_),
    .Y(_0788_),
    .B1(_0754_));
 sg13g2_nand4_1 _1651_ (.B(\vga_image_generator.character_hold[10] ),
    .C(_0658_),
    .A(_0695_),
    .Y(_0789_),
    .D(_0340_));
 sg13g2_nor3_1 _1652_ (.A(_0733_),
    .B(_0788_),
    .C(_0789_),
    .Y(_0790_));
 sg13g2_nand2_1 _1653_ (.Y(_0791_),
    .A(net34),
    .B(_0707_));
 sg13g2_nand2_1 _1654_ (.Y(_0792_),
    .A(\vga_image_generator.character_hold[13] ),
    .B(_0407_));
 sg13g2_nor3_1 _1655_ (.A(_0192_),
    .B(_0027_),
    .C(_0792_),
    .Y(_0793_));
 sg13g2_nand2_1 _1656_ (.Y(_0794_),
    .A(net30),
    .B(_0396_));
 sg13g2_nand3_1 _1657_ (.B(_0393_),
    .C(net29),
    .A(net31),
    .Y(_0795_));
 sg13g2_o21ai_1 _1658_ (.B1(_0795_),
    .Y(_0796_),
    .A1(net31),
    .A2(_0794_));
 sg13g2_nand4_1 _1659_ (.B(_0791_),
    .C(_0793_),
    .A(_0755_),
    .Y(_0797_),
    .D(_0796_));
 sg13g2_nand2_1 _1660_ (.Y(_0798_),
    .A(\vga_image_generator.character_hold[9] ),
    .B(_0766_));
 sg13g2_nand4_1 _1661_ (.B(\vga_image_generator.character_hold[11] ),
    .C(_0545_),
    .A(_0695_),
    .Y(_0799_),
    .D(_0340_));
 sg13g2_o21ai_1 _1662_ (.B1(_0799_),
    .Y(_0800_),
    .A1(_0186_),
    .A2(_0798_));
 sg13g2_nand3_1 _1663_ (.B(_0716_),
    .C(_0800_),
    .A(_0660_),
    .Y(_0801_));
 sg13g2_nand3b_1 _1664_ (.B(_0797_),
    .C(_0801_),
    .Y(_0802_),
    .A_N(_0790_));
 sg13g2_a221oi_1 _1665_ (.B2(_0787_),
    .C1(_0802_),
    .B1(_0786_),
    .A1(_0716_),
    .Y(_0803_),
    .A2(_0784_));
 sg13g2_and4_1 _1666_ (.A(_0714_),
    .B(_0744_),
    .C(_0779_),
    .D(_0803_),
    .X(_0804_));
 sg13g2_buf_2 _1667_ (.A(_0804_),
    .X(_0805_));
 sg13g2_and2_1 _1668_ (.A(_0626_),
    .B(_0660_),
    .X(_0806_));
 sg13g2_nand4_1 _1669_ (.B(_0806_),
    .C(_0755_),
    .A(net45),
    .Y(_0807_),
    .D(_0791_));
 sg13g2_and3_1 _1670_ (.X(_0808_),
    .A(net45),
    .B(net20),
    .C(_0667_));
 sg13g2_nor4_1 _1671_ (.A(net61),
    .B(_0705_),
    .C(_0174_),
    .D(_0701_),
    .Y(_0809_));
 sg13g2_xnor2_1 _1672_ (.Y(_0810_),
    .A(net49),
    .B(_0400_));
 sg13g2_nor2_1 _1673_ (.A(_0600_),
    .B(_0810_),
    .Y(_0811_));
 sg13g2_a22oi_1 _1674_ (.Y(_0812_),
    .B1(_0809_),
    .B2(_0811_),
    .A2(_0808_),
    .A1(_0704_));
 sg13g2_nand2_1 _1675_ (.Y(_0813_),
    .A(\vga_image_generator.character_hold[7] ),
    .B(_0766_));
 sg13g2_a21oi_1 _1676_ (.A1(_0807_),
    .A2(_0812_),
    .Y(_0814_),
    .B1(_0813_));
 sg13g2_mux2_1 _1677_ (.A0(net20),
    .A1(_0589_),
    .S(_0393_),
    .X(_0815_));
 sg13g2_nand3b_1 _1678_ (.B(net64),
    .C(net56),
    .Y(_0816_),
    .A_N(net63));
 sg13g2_nand2b_1 _1679_ (.Y(_0817_),
    .B(_0816_),
    .A_N(_0574_));
 sg13g2_nor4_1 _1680_ (.A(net47),
    .B(net36),
    .C(_0179_),
    .D(_0547_),
    .Y(_0818_));
 sg13g2_and4_1 _1681_ (.A(_0755_),
    .B(_0815_),
    .C(_0817_),
    .D(_0818_),
    .X(_0819_));
 sg13g2_or2_1 _1682_ (.X(_0820_),
    .B(_0185_),
    .A(net46));
 sg13g2_nor4_1 _1683_ (.A(_0179_),
    .B(_0820_),
    .C(_0736_),
    .D(_0740_),
    .Y(_0821_));
 sg13g2_o21ai_1 _1684_ (.B1(\vga_image_generator.character_hold[1] ),
    .Y(_0822_),
    .A1(_0819_),
    .A2(_0821_));
 sg13g2_nor2b_1 _1685_ (.A(_0814_),
    .B_N(_0822_),
    .Y(_0823_));
 sg13g2_xnor2_1 _1686_ (.Y(_0824_),
    .A(net60),
    .B(_0334_));
 sg13g2_and4_1 _1687_ (.A(net47),
    .B(_0400_),
    .C(_0759_),
    .D(_0824_),
    .X(_0825_));
 sg13g2_nor2_1 _1688_ (.A(_0667_),
    .B(_0660_),
    .Y(_0826_));
 sg13g2_inv_1 _1689_ (.Y(_0827_),
    .A(\vga_image_generator.character_hold[12] ));
 sg13g2_nor4_1 _1690_ (.A(_0027_),
    .B(_0827_),
    .C(_0338_),
    .D(_0557_),
    .Y(_0828_));
 sg13g2_a22oi_1 _1691_ (.Y(_0829_),
    .B1(_0826_),
    .B2(_0828_),
    .A2(_0825_),
    .A1(_0782_));
 sg13g2_nor2_1 _1692_ (.A(_0736_),
    .B(_0829_),
    .Y(_0830_));
 sg13g2_a21oi_1 _1693_ (.A1(_0538_),
    .A2(_0739_),
    .Y(_0831_),
    .B1(_0178_));
 sg13g2_or2_1 _1694_ (.X(_0832_),
    .B(net63),
    .A(net61));
 sg13g2_a221oi_1 _1695_ (.B2(_0707_),
    .C1(_0368_),
    .B1(_0832_),
    .A1(_0328_),
    .Y(_0833_),
    .A2(_0606_));
 sg13g2_nor2_1 _1696_ (.A(_0705_),
    .B(_0701_),
    .Y(_0834_));
 sg13g2_a221oi_1 _1697_ (.B2(_0834_),
    .C1(_0751_),
    .B1(_0833_),
    .A1(_0336_),
    .Y(_0835_),
    .A2(_0752_));
 sg13g2_nand3_1 _1698_ (.B(_0626_),
    .C(_0748_),
    .A(\vga_image_generator.character_hold[0] ),
    .Y(_0836_));
 sg13g2_nor3_1 _1699_ (.A(_0831_),
    .B(_0835_),
    .C(_0836_),
    .Y(_0837_));
 sg13g2_nor4_1 _1700_ (.A(_0560_),
    .B(_0810_),
    .C(_0711_),
    .D(_0792_),
    .Y(_0838_));
 sg13g2_nand4_1 _1701_ (.B(net44),
    .C(net36),
    .A(_0425_),
    .Y(_0839_),
    .D(\vga_image_generator.character_hold[17] ));
 sg13g2_nor4_2 _1702_ (.A(_0705_),
    .B(_0537_),
    .C(_0707_),
    .Y(_0840_),
    .D(_0701_));
 sg13g2_nand2_1 _1703_ (.Y(_0841_),
    .A(_0840_),
    .B(_0811_));
 sg13g2_mux2_1 _1704_ (.A0(_0759_),
    .A1(_0768_),
    .S(net34),
    .X(_0842_));
 sg13g2_nand2_1 _1705_ (.Y(_0843_),
    .A(net33),
    .B(\vga_image_generator.character_hold[5] ));
 sg13g2_nor4_1 _1706_ (.A(_0820_),
    .B(_0760_),
    .C(_0810_),
    .D(_0843_),
    .Y(_0844_));
 sg13g2_nand4_1 _1707_ (.B(_0834_),
    .C(_0842_),
    .A(_0538_),
    .Y(_0103_),
    .D(_0844_));
 sg13g2_o21ai_1 _1708_ (.B1(_0103_),
    .Y(_0104_),
    .A1(_0839_),
    .A2(_0841_));
 sg13g2_nor4_1 _1709_ (.A(_0830_),
    .B(_0837_),
    .C(_0838_),
    .D(_0104_),
    .Y(_0105_));
 sg13g2_nor4_1 _1710_ (.A(net30),
    .B(net45),
    .C(_0190_),
    .D(_0560_),
    .Y(_0106_));
 sg13g2_nor3_1 _1711_ (.A(_0393_),
    .B(_0186_),
    .C(_0760_),
    .Y(_0107_));
 sg13g2_o21ai_1 _1712_ (.B1(\vga_image_generator.character_hold[9] ),
    .Y(_0108_),
    .A1(_0106_),
    .A2(_0107_));
 sg13g2_and3_1 _1713_ (.X(_0109_),
    .A(net36),
    .B(\vga_image_generator.character_hold[15] ),
    .C(_0696_));
 sg13g2_a21oi_1 _1714_ (.A1(_0815_),
    .A2(_0109_),
    .Y(_0110_),
    .B1(_0828_));
 sg13g2_a21oi_1 _1715_ (.A1(_0108_),
    .A2(_0110_),
    .Y(_0111_),
    .B1(_0773_));
 sg13g2_nand2_1 _1716_ (.Y(_0112_),
    .A(\vga_image_generator.character_hold[4] ),
    .B(_0545_));
 sg13g2_nor4_1 _1717_ (.A(_0729_),
    .B(_0773_),
    .C(_0722_),
    .D(_0112_),
    .Y(_0113_));
 sg13g2_nor4_1 _1718_ (.A(net64),
    .B(_0717_),
    .C(_0722_),
    .D(_0112_),
    .Y(_0114_));
 sg13g2_a22oi_1 _1719_ (.Y(_0115_),
    .B1(_0739_),
    .B2(_0627_),
    .A2(_0759_),
    .A1(_0840_));
 sg13g2_nor4_1 _1720_ (.A(_0699_),
    .B(_0720_),
    .C(_0112_),
    .D(_0115_),
    .Y(_0116_));
 sg13g2_nor4_1 _1721_ (.A(_0111_),
    .B(_0113_),
    .C(_0114_),
    .D(_0116_),
    .Y(_0117_));
 sg13g2_a21oi_1 _1722_ (.A1(_0156_),
    .A2(_0627_),
    .Y(_0118_),
    .B1(_0833_));
 sg13g2_nand4_1 _1723_ (.B(_0545_),
    .C(_0834_),
    .A(_0728_),
    .Y(_0119_),
    .D(_0748_));
 sg13g2_nor3_1 _1724_ (.A(_0831_),
    .B(_0118_),
    .C(_0119_),
    .Y(_0120_));
 sg13g2_or2_1 _1725_ (.X(_0121_),
    .B(_0809_),
    .A(_0826_));
 sg13g2_and4_1 _1726_ (.A(net45),
    .B(_0755_),
    .C(_0791_),
    .D(_0121_),
    .X(_0122_));
 sg13g2_and3_1 _1727_ (.X(_0123_),
    .A(\vga_image_generator.character_hold[8] ),
    .B(_0589_),
    .C(_0766_));
 sg13g2_nand3_1 _1728_ (.B(_0627_),
    .C(_0716_),
    .A(_0585_),
    .Y(_0124_));
 sg13g2_nand3_1 _1729_ (.B(_0027_),
    .C(_0840_),
    .A(_0178_),
    .Y(_0125_));
 sg13g2_nor3_1 _1730_ (.A(net64),
    .B(_0190_),
    .C(_0557_),
    .Y(_0126_));
 sg13g2_nand2_1 _1731_ (.Y(_0127_),
    .A(\vga_image_generator.character_hold[2] ),
    .B(_0126_));
 sg13g2_a21oi_1 _1732_ (.A1(_0124_),
    .A2(_0125_),
    .Y(_0128_),
    .B1(_0127_));
 sg13g2_a221oi_1 _1733_ (.B2(_0123_),
    .C1(_0128_),
    .B1(_0122_),
    .A1(\vga_image_generator.character_hold[2] ),
    .Y(_0129_),
    .A2(_0120_));
 sg13g2_nand4_1 _1734_ (.B(_0105_),
    .C(_0117_),
    .A(_0823_),
    .Y(_0130_),
    .D(_0129_));
 sg13g2_buf_1 _1735_ (.A(_0130_),
    .X(_0131_));
 sg13g2_nand2_1 _1736_ (.Y(_0132_),
    .A(_0163_),
    .B(_0694_));
 sg13g2_nor2_1 _1737_ (.A(_0131_),
    .B(_0132_),
    .Y(_0133_));
 sg13g2_a22oi_1 _1738_ (.Y(net12),
    .B1(_0805_),
    .B2(_0133_),
    .A2(_0694_),
    .A1(_0692_));
 sg13g2_mux2_1 _1739_ (.A0(\BNC_x[7] ),
    .A1(\BNC_y[4] ),
    .S(net66),
    .X(_0134_));
 sg13g2_nand2_1 _1740_ (.Y(_0135_),
    .A(net65),
    .B(_0134_));
 sg13g2_nor2b_1 _1741_ (.A(_0131_),
    .B_N(_0135_),
    .Y(_0136_));
 sg13g2_a22oi_1 _1742_ (.Y(net13),
    .B1(_0136_),
    .B2(_0805_),
    .A2(_0135_),
    .A1(_0692_));
 sg13g2_nor2b_1 _1743_ (.A(net66),
    .B_N(\BNC_x[5] ),
    .Y(_0137_));
 sg13g2_a21oi_1 _1744_ (.A1(_0528_),
    .A2(\BNC_y[6] ),
    .Y(_0138_),
    .B1(_0137_));
 sg13g2_nor2_1 _1745_ (.A(_0529_),
    .B(\hvsync_gen.vsync ),
    .Y(_0139_));
 sg13g2_a21oi_1 _1746_ (.A1(_0529_),
    .A2(_0138_),
    .Y(net14),
    .B1(_0139_));
 sg13g2_mux2_1 _1747_ (.A0(\BNC_y[6] ),
    .A1(\BNC_y[1] ),
    .S(net66),
    .X(_0140_));
 sg13g2_nand2_1 _1748_ (.Y(_0141_),
    .A(net65),
    .B(_0140_));
 sg13g2_nand3_1 _1749_ (.B(_0163_),
    .C(_0141_),
    .A(net59),
    .Y(_0142_));
 sg13g2_nor2_1 _1750_ (.A(_0131_),
    .B(_0142_),
    .Y(_0143_));
 sg13g2_a22oi_1 _1751_ (.Y(net15),
    .B1(_0143_),
    .B2(_0805_),
    .A2(_0141_),
    .A1(_0692_));
 sg13g2_mux2_1 _1752_ (.A0(\BNC_y[4] ),
    .A1(\BNC_y[3] ),
    .S(net66),
    .X(_0144_));
 sg13g2_nand2_1 _1753_ (.Y(_0145_),
    .A(net65),
    .B(_0144_));
 sg13g2_nand2_1 _1754_ (.Y(_0146_),
    .A(net59),
    .B(_0145_));
 sg13g2_nor2_1 _1755_ (.A(_0131_),
    .B(_0146_),
    .Y(_0147_));
 sg13g2_a22oi_1 _1756_ (.Y(net16),
    .B1(_0147_),
    .B2(_0805_),
    .A2(_0145_),
    .A1(_0655_));
 sg13g2_mux2_1 _1757_ (.A0(\BNC_x[6] ),
    .A1(\BNC_y[5] ),
    .S(net66),
    .X(_0148_));
 sg13g2_nand2_1 _1758_ (.Y(_0149_),
    .A(net65),
    .B(_0148_));
 sg13g2_nor2b_1 _1759_ (.A(_0131_),
    .B_N(_0149_),
    .Y(_0150_));
 sg13g2_a22oi_1 _1760_ (.Y(net17),
    .B1(_0150_),
    .B2(_0805_),
    .A2(_0149_),
    .A1(_0692_));
 sg13g2_nor2b_1 _1761_ (.A(net66),
    .B_N(\BNC_x[4] ),
    .Y(_0151_));
 sg13g2_a21oi_1 _1762_ (.A1(net24),
    .A2(net163),
    .Y(_0152_),
    .B1(_0151_));
 sg13g2_nor2_1 _1763_ (.A(net65),
    .B(hsync),
    .Y(_0153_));
 sg13g2_a21oi_1 _1764_ (.A1(net65),
    .A2(_0152_),
    .Y(net18),
    .B1(_0153_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _1766_ (.A(net67),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1767_ (.A(net68),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1768_ (.A(net69),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1769_ (.A(net70),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1770_ (.A(net71),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1771_ (.A(net72),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1772_ (.A(net73),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1773_ (.A(net74),
    .X(uio_oe[7]));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[0]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net75),
    .D(_0000_),
    .Q_N(_0903_),
    .Q(\BNC_x[0] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[1]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net76),
    .D(_0001_),
    .Q_N(_0904_),
    .Q(\BNC_x[1] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[2]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net77),
    .D(_0002_),
    .Q_N(_0905_),
    .Q(\BNC_x[2] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[3]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net78),
    .D(_0003_),
    .Q_N(_0906_),
    .Q(\BNC_x[3] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[4]$_DFF_P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net79),
    .D(_0004_),
    .Q_N(_0907_),
    .Q(\BNC_x[4] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[5]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net80),
    .D(_0005_),
    .Q_N(_0908_),
    .Q(\BNC_x[5] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[6]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net81),
    .D(_0006_),
    .Q_N(_0909_),
    .Q(\BNC_x[6] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[7]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net82),
    .D(_0007_),
    .Q_N(_0910_),
    .Q(\BNC_x[7] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[0]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net83),
    .D(_0008_),
    .Q_N(_0911_),
    .Q(\BNC_y[0] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[1]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net84),
    .D(_0009_),
    .Q_N(_0912_),
    .Q(\BNC_y[1] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[2]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net85),
    .D(_0010_),
    .Q_N(_0913_),
    .Q(\BNC_y[2] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[3]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net86),
    .D(_0011_),
    .Q_N(_0914_),
    .Q(\BNC_y[3] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[4]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net87),
    .D(_0012_),
    .Q_N(_0915_),
    .Q(\BNC_y[4] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[5]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net88),
    .D(_0013_),
    .Q_N(_0916_),
    .Q(\BNC_y[5] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[6]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net89),
    .D(_0014_),
    .Q_N(_0902_),
    .Q(\BNC_y[6] ));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[0]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net90),
    .D(_0032_),
    .Q_N(_0030_),
    .Q(\bnc_image_generator.counter[0] ));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[1]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net91),
    .D(_0033_),
    .Q_N(_0019_),
    .Q(\bnc_image_generator.counter[1] ));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[2]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net92),
    .D(_0034_),
    .Q_N(_0018_),
    .Q(\bnc_image_generator.counter[2] ));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[3]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net93),
    .D(_0035_),
    .Q_N(_0017_),
    .Q(BNC_trig));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[4]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net94),
    .D(_0036_),
    .Q_N(_0901_),
    .Q(\bnc_image_generator.counter[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net95),
    .D(_0037_),
    .Q_N(_0028_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net96),
    .D(_0038_),
    .Q_N(_0024_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net97),
    .D(_0039_),
    .Q_N(_0900_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net98),
    .D(_0040_),
    .Q_N(_0025_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net99),
    .D(_0041_),
    .Q_N(_0899_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net100),
    .D(_0042_),
    .Q_N(_0023_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net101),
    .D(_0043_),
    .Q_N(_0898_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net102),
    .D(_0044_),
    .Q_N(_0897_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(_0045_),
    .Q_N(_0027_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net104),
    .D(_0046_),
    .Q_N(_0022_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hsync$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net105),
    .D(_0015_),
    .Q_N(_0896_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net106),
    .D(_0047_),
    .Q_N(_0029_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net107),
    .D(_0048_),
    .Q_N(_0895_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net108),
    .D(_0049_),
    .Q_N(_0894_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net109),
    .D(_0050_),
    .Q_N(_0021_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net110),
    .D(_0051_),
    .Q_N(_0893_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net111),
    .D(_0052_),
    .Q_N(_0020_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net112),
    .D(_0053_),
    .Q_N(_0892_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net113),
    .D(_0054_),
    .Q_N(_0891_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net114),
    .D(_0055_),
    .Q_N(_0026_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net115),
    .D(_0056_),
    .Q_N(_0917_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.vsync$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net116),
    .D(_0016_),
    .Q_N(_0890_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[0]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net117),
    .D(_0057_),
    .Q_N(_0889_),
    .Q(\vga_image_generator.character_hold[0] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[10]$_SDFFE_PN0N_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net118),
    .D(_0058_),
    .Q_N(_0888_),
    .Q(\vga_image_generator.character_hold[10] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[11]$_SDFFE_PN0N_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net119),
    .D(_0059_),
    .Q_N(_0887_),
    .Q(\vga_image_generator.character_hold[11] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[12]$_SDFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net120),
    .D(_0060_),
    .Q_N(_0886_),
    .Q(\vga_image_generator.character_hold[12] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[13]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net121),
    .D(_0061_),
    .Q_N(_0885_),
    .Q(\vga_image_generator.character_hold[13] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[14]$_SDFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net122),
    .D(_0062_),
    .Q_N(_0884_),
    .Q(\vga_image_generator.character_hold[14] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[15]$_SDFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net123),
    .D(_0063_),
    .Q_N(_0883_),
    .Q(\vga_image_generator.character_hold[15] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[16]$_SDFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net124),
    .D(_0064_),
    .Q_N(_0882_),
    .Q(\vga_image_generator.character_hold[16] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[17]$_SDFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net125),
    .D(_0065_),
    .Q_N(_0881_),
    .Q(\vga_image_generator.character_hold[17] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[1]$_SDFFE_PN0N_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net126),
    .D(_0066_),
    .Q_N(_0880_),
    .Q(\vga_image_generator.character_hold[1] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[2]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net127),
    .D(_0067_),
    .Q_N(_0879_),
    .Q(\vga_image_generator.character_hold[2] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[3]$_SDFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net128),
    .D(_0068_),
    .Q_N(_0878_),
    .Q(\vga_image_generator.character_hold[3] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[4]$_SDFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net129),
    .D(_0069_),
    .Q_N(_0877_),
    .Q(\vga_image_generator.character_hold[4] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[5]$_SDFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net130),
    .D(_0070_),
    .Q_N(_0876_),
    .Q(\vga_image_generator.character_hold[5] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[6]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net131),
    .D(_0071_),
    .Q_N(_0875_),
    .Q(\vga_image_generator.character_hold[6] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[7]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net132),
    .D(_0072_),
    .Q_N(_0874_),
    .Q(\vga_image_generator.character_hold[7] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[8]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net133),
    .D(_0073_),
    .Q_N(_0873_),
    .Q(\vga_image_generator.character_hold[8] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[9]$_SDFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net134),
    .D(_0074_),
    .Q_N(_0872_),
    .Q(\vga_image_generator.character_hold[9] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[0]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net135),
    .D(_0075_),
    .Q_N(_0031_),
    .Q(\vga_image_generator.counter[0] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[10]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net136),
    .D(_0076_),
    .Q_N(_0871_),
    .Q(\vga_image_generator.counter[10] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[11]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net137),
    .D(_0077_),
    .Q_N(_0870_),
    .Q(\vga_image_generator.counter[11] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[12]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net138),
    .D(_0078_),
    .Q_N(_0869_),
    .Q(\vga_image_generator.counter[12] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[13]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net139),
    .D(_0079_),
    .Q_N(_0868_),
    .Q(\vga_image_generator.counter[13] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[14]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net140),
    .D(_0080_),
    .Q_N(_0867_),
    .Q(\vga_image_generator.counter[14] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[15]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net141),
    .D(_0081_),
    .Q_N(_0866_),
    .Q(\vga_image_generator.counter[15] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[16]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net142),
    .D(_0082_),
    .Q_N(_0865_),
    .Q(\vga_image_generator.counter[16] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[17]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net143),
    .D(_0083_),
    .Q_N(_0864_),
    .Q(\vga_image_generator.counter[17] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[18]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net144),
    .D(_0084_),
    .Q_N(_0863_),
    .Q(\vga_image_generator.counter[18] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[19]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net145),
    .D(_0085_),
    .Q_N(_0862_),
    .Q(\vga_image_generator.counter[19] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[1]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net146),
    .D(_0086_),
    .Q_N(_0861_),
    .Q(\vga_image_generator.counter[1] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[20]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net147),
    .D(_0087_),
    .Q_N(_0860_),
    .Q(\vga_image_generator.counter[20] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[21]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net148),
    .D(_0088_),
    .Q_N(_0859_),
    .Q(\vga_image_generator.counter[21] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[22]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net149),
    .D(_0089_),
    .Q_N(_0858_),
    .Q(\vga_image_generator.counter[22] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[23]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net150),
    .D(_0090_),
    .Q_N(_0857_),
    .Q(\vga_image_generator.counter[23] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[24]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net151),
    .D(_0091_),
    .Q_N(_0856_),
    .Q(\vga_image_generator.counter[24] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[25]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net152),
    .D(_0092_),
    .Q_N(_0855_),
    .Q(\vga_image_generator.counter[25] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[26]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net153),
    .D(_0093_),
    .Q_N(_0854_),
    .Q(\vga_image_generator.counter[26] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[27]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net154),
    .D(_0094_),
    .Q_N(_0853_),
    .Q(\vga_image_generator.counter[27] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[2]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net155),
    .D(_0095_),
    .Q_N(_0852_),
    .Q(\vga_image_generator.counter[2] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[3]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net156),
    .D(_0096_),
    .Q_N(_0851_),
    .Q(\vga_image_generator.counter[3] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[4]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net157),
    .D(_0097_),
    .Q_N(_0850_),
    .Q(\vga_image_generator.counter[4] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[5]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net158),
    .D(_0098_),
    .Q_N(_0849_),
    .Q(\vga_image_generator.counter[5] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[6]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net159),
    .D(_0099_),
    .Q_N(_0848_),
    .Q(\vga_image_generator.counter[6] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[7]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net160),
    .D(_0100_),
    .Q_N(_0847_),
    .Q(\vga_image_generator.counter[7] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[8]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net161),
    .D(_0101_),
    .Q_N(_0846_),
    .Q(\vga_image_generator.counter[8] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[9]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net162),
    .D(_0102_),
    .Q_N(_0845_),
    .Q(\vga_image_generator.counter[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout19 (.A(_0326_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0658_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0243_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0235_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0228_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0198_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0504_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0478_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0453_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0436_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0400_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0399_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0391_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0390_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0367_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0359_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0328_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0327_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0218_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0212_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0211_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0206_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0204_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0200_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0197_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0192_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0188_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0183_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0170_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0350_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0334_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0333_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0329_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0210_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0199_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0185_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0184_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0176_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0173_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0167_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0166_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0159_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0158_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0157_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0154_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0728_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0529_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0527_),
    .X(net66));
 sg13g2_tiehi _1766__67 (.L_HI(net67));
 sg13g2_tiehi _1767__68 (.L_HI(net68));
 sg13g2_tiehi _1768__69 (.L_HI(net69));
 sg13g2_tiehi _1769__70 (.L_HI(net70));
 sg13g2_tiehi _1770__71 (.L_HI(net71));
 sg13g2_tiehi _1771__72 (.L_HI(net72));
 sg13g2_tiehi _1772__73 (.L_HI(net73));
 sg13g2_tiehi _1773__74 (.L_HI(net74));
 sg13g2_tiehi \bnc_image_generator.BNC_x[0]$_DFF_P__75  (.L_HI(net75));
 sg13g2_tiehi \bnc_image_generator.BNC_x[1]$_DFF_P__76  (.L_HI(net76));
 sg13g2_tiehi \bnc_image_generator.BNC_x[2]$_DFF_P__77  (.L_HI(net77));
 sg13g2_tiehi \bnc_image_generator.BNC_x[3]$_DFF_P__78  (.L_HI(net78));
 sg13g2_tiehi \bnc_image_generator.BNC_x[4]$_DFF_P__79  (.L_HI(net79));
 sg13g2_tiehi \bnc_image_generator.BNC_x[5]$_DFF_P__80  (.L_HI(net80));
 sg13g2_tiehi \bnc_image_generator.BNC_x[6]$_DFF_P__81  (.L_HI(net81));
 sg13g2_tiehi \bnc_image_generator.BNC_x[7]$_DFF_P__82  (.L_HI(net82));
 sg13g2_tiehi \bnc_image_generator.BNC_y[0]$_DFF_P__83  (.L_HI(net83));
 sg13g2_tiehi \bnc_image_generator.BNC_y[1]$_DFF_P__84  (.L_HI(net84));
 sg13g2_tiehi \bnc_image_generator.BNC_y[2]$_DFF_P__85  (.L_HI(net85));
 sg13g2_tiehi \bnc_image_generator.BNC_y[3]$_DFF_P__86  (.L_HI(net86));
 sg13g2_tiehi \bnc_image_generator.BNC_y[4]$_DFF_P__87  (.L_HI(net87));
 sg13g2_tiehi \bnc_image_generator.BNC_y[5]$_DFF_P__88  (.L_HI(net88));
 sg13g2_tiehi \bnc_image_generator.BNC_y[6]$_DFF_P__89  (.L_HI(net89));
 sg13g2_tiehi \bnc_image_generator.counter[0]$_SDFF_PN0__90  (.L_HI(net90));
 sg13g2_tiehi \bnc_image_generator.counter[1]$_SDFF_PN0__91  (.L_HI(net91));
 sg13g2_tiehi \bnc_image_generator.counter[2]$_SDFF_PN0__92  (.L_HI(net92));
 sg13g2_tiehi \bnc_image_generator.counter[3]$_SDFF_PN0__93  (.L_HI(net93));
 sg13g2_tiehi \bnc_image_generator.counter[4]$_SDFF_PN0__94  (.L_HI(net94));
 sg13g2_tiehi \hvsync_gen.hpos[0]$_SDFF_PP0__95  (.L_HI(net95));
 sg13g2_tiehi \hvsync_gen.hpos[1]$_SDFF_PP0__96  (.L_HI(net96));
 sg13g2_tiehi \hvsync_gen.hpos[2]$_SDFF_PP0__97  (.L_HI(net97));
 sg13g2_tiehi \hvsync_gen.hpos[3]$_SDFF_PP0__98  (.L_HI(net98));
 sg13g2_tiehi \hvsync_gen.hpos[4]$_SDFF_PP0__99  (.L_HI(net99));
 sg13g2_tiehi \hvsync_gen.hpos[5]$_SDFF_PP0__100  (.L_HI(net100));
 sg13g2_tiehi \hvsync_gen.hpos[6]$_SDFF_PP0__101  (.L_HI(net101));
 sg13g2_tiehi \hvsync_gen.hpos[7]$_SDFF_PP0__102  (.L_HI(net102));
 sg13g2_tiehi \hvsync_gen.hpos[8]$_SDFF_PP0__103  (.L_HI(net103));
 sg13g2_tiehi \hvsync_gen.hpos[9]$_SDFF_PP0__104  (.L_HI(net104));
 sg13g2_tiehi \hvsync_gen.hsync$_DFF_P__105  (.L_HI(net105));
 sg13g2_tiehi \hvsync_gen.vpos[0]$_SDFFCE_PP0P__106  (.L_HI(net106));
 sg13g2_tiehi \hvsync_gen.vpos[1]$_SDFFCE_PP0P__107  (.L_HI(net107));
 sg13g2_tiehi \hvsync_gen.vpos[2]$_SDFFCE_PP0P__108  (.L_HI(net108));
 sg13g2_tiehi \hvsync_gen.vpos[3]$_SDFFCE_PP0P__109  (.L_HI(net109));
 sg13g2_tiehi \hvsync_gen.vpos[4]$_SDFFCE_PP0P__110  (.L_HI(net110));
 sg13g2_tiehi \hvsync_gen.vpos[5]$_SDFFCE_PP0P__111  (.L_HI(net111));
 sg13g2_tiehi \hvsync_gen.vpos[6]$_SDFFCE_PP0P__112  (.L_HI(net112));
 sg13g2_tiehi \hvsync_gen.vpos[7]$_SDFFCE_PP0P__113  (.L_HI(net113));
 sg13g2_tiehi \hvsync_gen.vpos[8]$_SDFFCE_PP0P__114  (.L_HI(net114));
 sg13g2_tiehi \hvsync_gen.vpos[9]$_SDFFCE_PP0P__115  (.L_HI(net115));
 sg13g2_tiehi \hvsync_gen.vsync$_DFF_P__116  (.L_HI(net116));
 sg13g2_tiehi \vga_image_generator.character_hold[0]$_SDFFE_PN0N__117  (.L_HI(net117));
 sg13g2_tiehi \vga_image_generator.character_hold[10]$_SDFFE_PN0N__118  (.L_HI(net118));
 sg13g2_tiehi \vga_image_generator.character_hold[11]$_SDFFE_PN0N__119  (.L_HI(net119));
 sg13g2_tiehi \vga_image_generator.character_hold[12]$_SDFFE_PN0N__120  (.L_HI(net120));
 sg13g2_tiehi \vga_image_generator.character_hold[13]$_SDFFE_PN0N__121  (.L_HI(net121));
 sg13g2_tiehi \vga_image_generator.character_hold[14]$_SDFFE_PN0N__122  (.L_HI(net122));
 sg13g2_tiehi \vga_image_generator.character_hold[15]$_SDFFE_PN0N__123  (.L_HI(net123));
 sg13g2_tiehi \vga_image_generator.character_hold[16]$_SDFFE_PN0N__124  (.L_HI(net124));
 sg13g2_tiehi \vga_image_generator.character_hold[17]$_SDFFE_PN0N__125  (.L_HI(net125));
 sg13g2_tiehi \vga_image_generator.character_hold[1]$_SDFFE_PN0N__126  (.L_HI(net126));
 sg13g2_tiehi \vga_image_generator.character_hold[2]$_SDFFE_PN0N__127  (.L_HI(net127));
 sg13g2_tiehi \vga_image_generator.character_hold[3]$_SDFFE_PN0N__128  (.L_HI(net128));
 sg13g2_tiehi \vga_image_generator.character_hold[4]$_SDFFE_PN0N__129  (.L_HI(net129));
 sg13g2_tiehi \vga_image_generator.character_hold[5]$_SDFFE_PN0N__130  (.L_HI(net130));
 sg13g2_tiehi \vga_image_generator.character_hold[6]$_SDFFE_PN0N__131  (.L_HI(net131));
 sg13g2_tiehi \vga_image_generator.character_hold[7]$_SDFFE_PN0N__132  (.L_HI(net132));
 sg13g2_tiehi \vga_image_generator.character_hold[8]$_SDFFE_PN0N__133  (.L_HI(net133));
 sg13g2_tiehi \vga_image_generator.character_hold[9]$_SDFFE_PN0N__134  (.L_HI(net134));
 sg13g2_tiehi \vga_image_generator.counter[0]$_SDFF_PN0__135  (.L_HI(net135));
 sg13g2_tiehi \vga_image_generator.counter[10]$_SDFF_PN0__136  (.L_HI(net136));
 sg13g2_tiehi \vga_image_generator.counter[11]$_SDFF_PN0__137  (.L_HI(net137));
 sg13g2_tiehi \vga_image_generator.counter[12]$_SDFF_PN0__138  (.L_HI(net138));
 sg13g2_tiehi \vga_image_generator.counter[13]$_SDFF_PN0__139  (.L_HI(net139));
 sg13g2_tiehi \vga_image_generator.counter[14]$_SDFF_PN0__140  (.L_HI(net140));
 sg13g2_tiehi \vga_image_generator.counter[15]$_SDFF_PN0__141  (.L_HI(net141));
 sg13g2_tiehi \vga_image_generator.counter[16]$_SDFF_PN0__142  (.L_HI(net142));
 sg13g2_tiehi \vga_image_generator.counter[17]$_SDFF_PN0__143  (.L_HI(net143));
 sg13g2_tiehi \vga_image_generator.counter[18]$_SDFF_PN0__144  (.L_HI(net144));
 sg13g2_tiehi \vga_image_generator.counter[19]$_SDFF_PN0__145  (.L_HI(net145));
 sg13g2_tiehi \vga_image_generator.counter[1]$_SDFF_PN0__146  (.L_HI(net146));
 sg13g2_tiehi \vga_image_generator.counter[20]$_SDFF_PN0__147  (.L_HI(net147));
 sg13g2_tiehi \vga_image_generator.counter[21]$_SDFF_PN0__148  (.L_HI(net148));
 sg13g2_tiehi \vga_image_generator.counter[22]$_SDFF_PN0__149  (.L_HI(net149));
 sg13g2_tiehi \vga_image_generator.counter[23]$_SDFF_PN0__150  (.L_HI(net150));
 sg13g2_tiehi \vga_image_generator.counter[24]$_SDFF_PN0__151  (.L_HI(net151));
 sg13g2_tiehi \vga_image_generator.counter[25]$_SDFF_PN0__152  (.L_HI(net152));
 sg13g2_tiehi \vga_image_generator.counter[26]$_SDFF_PN0__153  (.L_HI(net153));
 sg13g2_tiehi \vga_image_generator.counter[27]$_SDFF_PN0__154  (.L_HI(net154));
 sg13g2_tiehi \vga_image_generator.counter[2]$_SDFF_PN0__155  (.L_HI(net155));
 sg13g2_tiehi \vga_image_generator.counter[3]$_SDFF_PN0__156  (.L_HI(net156));
 sg13g2_tiehi \vga_image_generator.counter[4]$_SDFF_PN0__157  (.L_HI(net157));
 sg13g2_tiehi \vga_image_generator.counter[5]$_SDFF_PN0__158  (.L_HI(net158));
 sg13g2_tiehi \vga_image_generator.counter[6]$_SDFF_PN0__159  (.L_HI(net159));
 sg13g2_tiehi \vga_image_generator.counter[7]$_SDFF_PN0__160  (.L_HI(net160));
 sg13g2_tiehi \vga_image_generator.counter[8]$_SDFF_PN0__161  (.L_HI(net161));
 sg13g2_tiehi \vga_image_generator.counter[9]$_SDFF_PN0__162  (.L_HI(net162));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_15_0_clk));
 sg13g2_buf_1 fanout1 (.A(_0528_),
    .X(net163));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_4 FILLER_3_217 ();
 sg13g2_fill_2 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_227 ();
 sg13g2_decap_8 FILLER_3_234 ();
 sg13g2_fill_2 FILLER_3_241 ();
 sg13g2_fill_1 FILLER_3_243 ();
 sg13g2_fill_1 FILLER_3_248 ();
 sg13g2_decap_8 FILLER_3_257 ();
 sg13g2_decap_8 FILLER_3_264 ();
 sg13g2_decap_8 FILLER_3_271 ();
 sg13g2_decap_8 FILLER_3_278 ();
 sg13g2_decap_8 FILLER_3_285 ();
 sg13g2_decap_8 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_299 ();
 sg13g2_decap_8 FILLER_3_306 ();
 sg13g2_decap_8 FILLER_3_313 ();
 sg13g2_decap_8 FILLER_3_320 ();
 sg13g2_decap_8 FILLER_3_327 ();
 sg13g2_decap_8 FILLER_3_334 ();
 sg13g2_decap_8 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_8 FILLER_3_404 ();
 sg13g2_decap_8 FILLER_3_411 ();
 sg13g2_decap_8 FILLER_3_418 ();
 sg13g2_decap_4 FILLER_3_425 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_fill_2 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_170 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_fill_2 FILLER_4_210 ();
 sg13g2_fill_2 FILLER_4_250 ();
 sg13g2_fill_1 FILLER_4_252 ();
 sg13g2_fill_2 FILLER_4_287 ();
 sg13g2_fill_1 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_316 ();
 sg13g2_fill_2 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_decap_8 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_4_414 ();
 sg13g2_decap_8 FILLER_4_421 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_fill_2 FILLER_5_161 ();
 sg13g2_fill_1 FILLER_5_163 ();
 sg13g2_decap_4 FILLER_5_190 ();
 sg13g2_fill_2 FILLER_5_194 ();
 sg13g2_decap_4 FILLER_5_208 ();
 sg13g2_fill_1 FILLER_5_212 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_fill_1 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_254 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_decap_8 FILLER_5_268 ();
 sg13g2_decap_8 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_282 ();
 sg13g2_fill_1 FILLER_5_289 ();
 sg13g2_decap_4 FILLER_5_294 ();
 sg13g2_fill_1 FILLER_5_302 ();
 sg13g2_fill_2 FILLER_5_311 ();
 sg13g2_fill_1 FILLER_5_321 ();
 sg13g2_fill_2 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_decap_8 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_5_414 ();
 sg13g2_decap_8 FILLER_5_421 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_4 FILLER_6_126 ();
 sg13g2_fill_1 FILLER_6_130 ();
 sg13g2_fill_1 FILLER_6_157 ();
 sg13g2_fill_1 FILLER_6_170 ();
 sg13g2_fill_1 FILLER_6_179 ();
 sg13g2_fill_1 FILLER_6_196 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_fill_1 FILLER_6_234 ();
 sg13g2_decap_4 FILLER_6_269 ();
 sg13g2_fill_1 FILLER_6_303 ();
 sg13g2_fill_1 FILLER_6_312 ();
 sg13g2_fill_2 FILLER_6_318 ();
 sg13g2_decap_8 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_6_331 ();
 sg13g2_decap_4 FILLER_6_338 ();
 sg13g2_fill_1 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_decap_8 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_4 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_141 ();
 sg13g2_decap_8 FILLER_7_148 ();
 sg13g2_fill_1 FILLER_7_155 ();
 sg13g2_fill_2 FILLER_7_177 ();
 sg13g2_fill_1 FILLER_7_179 ();
 sg13g2_decap_8 FILLER_7_188 ();
 sg13g2_decap_8 FILLER_7_195 ();
 sg13g2_fill_2 FILLER_7_202 ();
 sg13g2_fill_1 FILLER_7_204 ();
 sg13g2_decap_4 FILLER_7_217 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_fill_2 FILLER_7_230 ();
 sg13g2_decap_4 FILLER_7_236 ();
 sg13g2_fill_2 FILLER_7_244 ();
 sg13g2_fill_1 FILLER_7_249 ();
 sg13g2_decap_8 FILLER_7_254 ();
 sg13g2_decap_8 FILLER_7_261 ();
 sg13g2_decap_8 FILLER_7_268 ();
 sg13g2_decap_8 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_282 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_4 FILLER_7_294 ();
 sg13g2_fill_2 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_fill_1 FILLER_7_318 ();
 sg13g2_decap_4 FILLER_7_349 ();
 sg13g2_fill_1 FILLER_7_353 ();
 sg13g2_decap_4 FILLER_7_358 ();
 sg13g2_fill_1 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_8 FILLER_7_403 ();
 sg13g2_decap_8 FILLER_7_410 ();
 sg13g2_decap_8 FILLER_7_417 ();
 sg13g2_decap_4 FILLER_7_424 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_4 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_169 ();
 sg13g2_decap_4 FILLER_8_176 ();
 sg13g2_fill_1 FILLER_8_180 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_fill_1 FILLER_8_221 ();
 sg13g2_fill_2 FILLER_8_252 ();
 sg13g2_fill_1 FILLER_8_254 ();
 sg13g2_fill_2 FILLER_8_281 ();
 sg13g2_fill_1 FILLER_8_283 ();
 sg13g2_fill_2 FILLER_8_319 ();
 sg13g2_decap_4 FILLER_8_345 ();
 sg13g2_fill_2 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_8 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_8_412 ();
 sg13g2_decap_8 FILLER_8_419 ();
 sg13g2_decap_4 FILLER_8_426 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_150 ();
 sg13g2_decap_4 FILLER_9_157 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_197 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_4 FILLER_9_215 ();
 sg13g2_fill_1 FILLER_9_219 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_4 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_235 ();
 sg13g2_decap_4 FILLER_9_241 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_4 FILLER_9_273 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_decap_4 FILLER_9_291 ();
 sg13g2_fill_1 FILLER_9_295 ();
 sg13g2_fill_2 FILLER_9_308 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_fill_2 FILLER_9_315 ();
 sg13g2_fill_1 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_4 FILLER_9_424 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_152 ();
 sg13g2_decap_8 FILLER_10_159 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_decap_8 FILLER_10_177 ();
 sg13g2_decap_4 FILLER_10_184 ();
 sg13g2_fill_2 FILLER_10_188 ();
 sg13g2_fill_2 FILLER_10_202 ();
 sg13g2_fill_1 FILLER_10_204 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_fill_1 FILLER_10_274 ();
 sg13g2_decap_4 FILLER_10_292 ();
 sg13g2_fill_2 FILLER_10_296 ();
 sg13g2_fill_1 FILLER_10_308 ();
 sg13g2_fill_2 FILLER_10_313 ();
 sg13g2_fill_1 FILLER_10_318 ();
 sg13g2_decap_4 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_341 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_fill_2 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_10_409 ();
 sg13g2_decap_8 FILLER_10_416 ();
 sg13g2_decap_8 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_4 FILLER_11_119 ();
 sg13g2_fill_1 FILLER_11_123 ();
 sg13g2_decap_4 FILLER_11_150 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_fill_1 FILLER_11_215 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_fill_2 FILLER_11_242 ();
 sg13g2_fill_1 FILLER_11_244 ();
 sg13g2_decap_4 FILLER_11_254 ();
 sg13g2_decap_4 FILLER_11_268 ();
 sg13g2_decap_4 FILLER_11_275 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_decap_4 FILLER_11_292 ();
 sg13g2_fill_2 FILLER_11_296 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_fill_1 FILLER_11_342 ();
 sg13g2_fill_2 FILLER_11_348 ();
 sg13g2_fill_1 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_fill_2 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_4 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_fill_1 FILLER_12_142 ();
 sg13g2_decap_8 FILLER_12_155 ();
 sg13g2_fill_1 FILLER_12_162 ();
 sg13g2_fill_2 FILLER_12_167 ();
 sg13g2_fill_2 FILLER_12_182 ();
 sg13g2_fill_1 FILLER_12_184 ();
 sg13g2_fill_2 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_205 ();
 sg13g2_decap_8 FILLER_12_212 ();
 sg13g2_decap_4 FILLER_12_219 ();
 sg13g2_fill_1 FILLER_12_223 ();
 sg13g2_decap_8 FILLER_12_229 ();
 sg13g2_decap_4 FILLER_12_236 ();
 sg13g2_fill_1 FILLER_12_240 ();
 sg13g2_decap_4 FILLER_12_249 ();
 sg13g2_fill_2 FILLER_12_285 ();
 sg13g2_fill_1 FILLER_12_287 ();
 sg13g2_decap_4 FILLER_12_292 ();
 sg13g2_fill_2 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_fill_2 FILLER_12_338 ();
 sg13g2_fill_1 FILLER_12_349 ();
 sg13g2_fill_1 FILLER_12_380 ();
 sg13g2_fill_1 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_fill_1 FILLER_12_403 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_135 ();
 sg13g2_fill_2 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_fill_2 FILLER_13_151 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_fill_2 FILLER_13_166 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_173 ();
 sg13g2_decap_8 FILLER_13_180 ();
 sg13g2_decap_8 FILLER_13_187 ();
 sg13g2_fill_2 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_204 ();
 sg13g2_fill_1 FILLER_13_231 ();
 sg13g2_decap_4 FILLER_13_258 ();
 sg13g2_fill_1 FILLER_13_262 ();
 sg13g2_fill_2 FILLER_13_267 ();
 sg13g2_fill_1 FILLER_13_269 ();
 sg13g2_decap_4 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_4 FILLER_13_338 ();
 sg13g2_fill_1 FILLER_13_342 ();
 sg13g2_decap_4 FILLER_13_381 ();
 sg13g2_fill_1 FILLER_13_385 ();
 sg13g2_decap_4 FILLER_13_425 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_fill_2 FILLER_14_145 ();
 sg13g2_fill_1 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_188 ();
 sg13g2_decap_8 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_202 ();
 sg13g2_decap_4 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_239 ();
 sg13g2_decap_4 FILLER_14_246 ();
 sg13g2_fill_2 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_291 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_330 ();
 sg13g2_decap_8 FILLER_14_337 ();
 sg13g2_fill_1 FILLER_14_344 ();
 sg13g2_fill_2 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_fill_2 FILLER_14_364 ();
 sg13g2_fill_2 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_fill_2 FILLER_14_384 ();
 sg13g2_fill_1 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_153 ();
 sg13g2_decap_8 FILLER_15_160 ();
 sg13g2_decap_8 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_174 ();
 sg13g2_decap_8 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_188 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_decap_8 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_208 ();
 sg13g2_decap_8 FILLER_15_215 ();
 sg13g2_decap_8 FILLER_15_222 ();
 sg13g2_decap_8 FILLER_15_233 ();
 sg13g2_decap_4 FILLER_15_240 ();
 sg13g2_decap_4 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_fill_1 FILLER_15_339 ();
 sg13g2_fill_1 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_15_355 ();
 sg13g2_fill_2 FILLER_15_383 ();
 sg13g2_decap_4 FILLER_15_399 ();
 sg13g2_decap_4 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_fill_1 FILLER_16_261 ();
 sg13g2_decap_4 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_decap_4 FILLER_16_296 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_333 ();
 sg13g2_fill_2 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_fill_1 FILLER_16_383 ();
 sg13g2_decap_4 FILLER_16_388 ();
 sg13g2_fill_2 FILLER_16_392 ();
 sg13g2_decap_4 FILLER_16_398 ();
 sg13g2_fill_2 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_fill_2 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_157 ();
 sg13g2_decap_8 FILLER_17_164 ();
 sg13g2_decap_8 FILLER_17_171 ();
 sg13g2_decap_8 FILLER_17_178 ();
 sg13g2_decap_8 FILLER_17_185 ();
 sg13g2_decap_4 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_196 ();
 sg13g2_decap_4 FILLER_17_201 ();
 sg13g2_fill_2 FILLER_17_205 ();
 sg13g2_decap_8 FILLER_17_215 ();
 sg13g2_fill_1 FILLER_17_222 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_4 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_307 ();
 sg13g2_decap_4 FILLER_17_320 ();
 sg13g2_decap_4 FILLER_17_354 ();
 sg13g2_fill_2 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_4 FILLER_17_382 ();
 sg13g2_fill_1 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_4 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_176 ();
 sg13g2_decap_8 FILLER_18_183 ();
 sg13g2_decap_4 FILLER_18_221 ();
 sg13g2_fill_1 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_fill_2 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_decap_4 FILLER_18_258 ();
 sg13g2_fill_1 FILLER_18_271 ();
 sg13g2_fill_2 FILLER_18_280 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_fill_2 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_4 FILLER_18_341 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_361 ();
 sg13g2_fill_1 FILLER_18_363 ();
 sg13g2_decap_4 FILLER_18_390 ();
 sg13g2_fill_2 FILLER_18_394 ();
 sg13g2_decap_4 FILLER_18_426 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_4 FILLER_19_161 ();
 sg13g2_decap_4 FILLER_19_191 ();
 sg13g2_fill_2 FILLER_19_195 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_219 ();
 sg13g2_decap_8 FILLER_19_225 ();
 sg13g2_decap_8 FILLER_19_232 ();
 sg13g2_fill_2 FILLER_19_239 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_decap_4 FILLER_19_268 ();
 sg13g2_fill_2 FILLER_19_298 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_309 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_decap_4 FILLER_19_332 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_fill_1 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_19_409 ();
 sg13g2_decap_8 FILLER_19_416 ();
 sg13g2_decap_8 FILLER_19_423 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_fill_2 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_181 ();
 sg13g2_decap_8 FILLER_20_187 ();
 sg13g2_decap_4 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_212 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_232 ();
 sg13g2_decap_4 FILLER_20_242 ();
 sg13g2_decap_4 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_259 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_287 ();
 sg13g2_decap_4 FILLER_20_299 ();
 sg13g2_fill_1 FILLER_20_303 ();
 sg13g2_fill_2 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_fill_2 FILLER_20_349 ();
 sg13g2_fill_2 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_fill_2 FILLER_20_383 ();
 sg13g2_fill_1 FILLER_20_385 ();
 sg13g2_fill_2 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_403 ();
 sg13g2_decap_8 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_4 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_decap_8 FILLER_21_164 ();
 sg13g2_fill_2 FILLER_21_171 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_199 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_decap_4 FILLER_21_214 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_247 ();
 sg13g2_decap_4 FILLER_21_256 ();
 sg13g2_fill_2 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_2 FILLER_21_308 ();
 sg13g2_fill_2 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_322 ();
 sg13g2_decap_4 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_4 FILLER_21_386 ();
 sg13g2_fill_1 FILLER_21_390 ();
 sg13g2_fill_2 FILLER_21_400 ();
 sg13g2_fill_1 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_21_415 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_fill_2 FILLER_22_183 ();
 sg13g2_fill_2 FILLER_22_199 ();
 sg13g2_fill_1 FILLER_22_201 ();
 sg13g2_fill_2 FILLER_22_226 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_239 ();
 sg13g2_decap_4 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_257 ();
 sg13g2_fill_2 FILLER_22_277 ();
 sg13g2_fill_1 FILLER_22_279 ();
 sg13g2_decap_8 FILLER_22_285 ();
 sg13g2_decap_8 FILLER_22_292 ();
 sg13g2_decap_4 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_324 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_4 FILLER_22_354 ();
 sg13g2_fill_2 FILLER_22_358 ();
 sg13g2_fill_1 FILLER_22_370 ();
 sg13g2_fill_1 FILLER_22_379 ();
 sg13g2_decap_4 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_4 FILLER_22_424 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_fill_2 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_fill_2 FILLER_23_191 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_fill_2 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_205 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_255 ();
 sg13g2_fill_2 FILLER_23_278 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_312 ();
 sg13g2_fill_2 FILLER_23_319 ();
 sg13g2_fill_1 FILLER_23_321 ();
 sg13g2_decap_4 FILLER_23_333 ();
 sg13g2_fill_1 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_4 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_fill_2 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_fill_2 FILLER_23_391 ();
 sg13g2_decap_4 FILLER_23_426 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_decap_8 FILLER_24_176 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_226 ();
 sg13g2_decap_4 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_243 ();
 sg13g2_decap_4 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_302 ();
 sg13g2_fill_2 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_24_378 ();
 sg13g2_fill_1 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_4 FILLER_24_425 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_4 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_78 ();
 sg13g2_decap_8 FILLER_25_85 ();
 sg13g2_decap_8 FILLER_25_92 ();
 sg13g2_decap_8 FILLER_25_99 ();
 sg13g2_decap_8 FILLER_25_106 ();
 sg13g2_decap_8 FILLER_25_113 ();
 sg13g2_decap_8 FILLER_25_120 ();
 sg13g2_decap_8 FILLER_25_127 ();
 sg13g2_decap_8 FILLER_25_134 ();
 sg13g2_decap_4 FILLER_25_141 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_152 ();
 sg13g2_fill_2 FILLER_25_157 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_fill_2 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_decap_4 FILLER_25_240 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_decap_4 FILLER_25_280 ();
 sg13g2_decap_4 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_320 ();
 sg13g2_decap_4 FILLER_25_332 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_fill_1 FILLER_25_376 ();
 sg13g2_fill_2 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_25_386 ();
 sg13g2_fill_2 FILLER_25_392 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_fill_2 FILLER_25_403 ();
 sg13g2_fill_1 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_25_416 ();
 sg13g2_decap_8 FILLER_25_423 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_decap_4 FILLER_26_94 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_4 FILLER_26_109 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_131 ();
 sg13g2_decap_8 FILLER_26_138 ();
 sg13g2_decap_8 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_254 ();
 sg13g2_decap_4 FILLER_26_261 ();
 sg13g2_fill_1 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_fill_2 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_decap_4 FILLER_26_370 ();
 sg13g2_fill_2 FILLER_26_379 ();
 sg13g2_fill_2 FILLER_26_386 ();
 sg13g2_fill_2 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_decap_4 FILLER_27_68 ();
 sg13g2_decap_8 FILLER_27_76 ();
 sg13g2_decap_4 FILLER_27_83 ();
 sg13g2_fill_1 FILLER_27_87 ();
 sg13g2_fill_2 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_decap_8 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_195 ();
 sg13g2_fill_1 FILLER_27_201 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_218 ();
 sg13g2_fill_2 FILLER_27_225 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_244 ();
 sg13g2_decap_8 FILLER_27_257 ();
 sg13g2_decap_8 FILLER_27_276 ();
 sg13g2_decap_4 FILLER_27_283 ();
 sg13g2_decap_4 FILLER_27_292 ();
 sg13g2_fill_1 FILLER_27_296 ();
 sg13g2_decap_4 FILLER_27_305 ();
 sg13g2_decap_4 FILLER_27_312 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_350 ();
 sg13g2_fill_1 FILLER_27_371 ();
 sg13g2_decap_4 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_36 ();
 sg13g2_decap_8 FILLER_28_43 ();
 sg13g2_fill_1 FILLER_28_50 ();
 sg13g2_fill_2 FILLER_28_64 ();
 sg13g2_decap_8 FILLER_28_82 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_121 ();
 sg13g2_decap_8 FILLER_28_127 ();
 sg13g2_fill_2 FILLER_28_134 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_decap_8 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_decap_8 FILLER_28_254 ();
 sg13g2_decap_8 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_decap_8 FILLER_28_276 ();
 sg13g2_decap_4 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_293 ();
 sg13g2_decap_4 FILLER_28_300 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_376 ();
 sg13g2_fill_1 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_34 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_fill_2 FILLER_29_52 ();
 sg13g2_fill_1 FILLER_29_54 ();
 sg13g2_fill_2 FILLER_29_64 ();
 sg13g2_fill_1 FILLER_29_75 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_fill_2 FILLER_29_149 ();
 sg13g2_fill_1 FILLER_29_151 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_176 ();
 sg13g2_decap_4 FILLER_29_183 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_224 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_fill_1 FILLER_29_234 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_decap_4 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_decap_4 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_312 ();
 sg13g2_fill_2 FILLER_29_319 ();
 sg13g2_fill_1 FILLER_29_325 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_4 FILLER_29_338 ();
 sg13g2_decap_4 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_396 ();
 sg13g2_fill_1 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_425 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_57 ();
 sg13g2_fill_1 FILLER_30_59 ();
 sg13g2_fill_2 FILLER_30_64 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_1 FILLER_30_81 ();
 sg13g2_fill_2 FILLER_30_100 ();
 sg13g2_fill_1 FILLER_30_102 ();
 sg13g2_fill_2 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_127 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_decap_4 FILLER_30_138 ();
 sg13g2_decap_4 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_151 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_decap_4 FILLER_30_228 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_298 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_314 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_fill_1 FILLER_30_330 ();
 sg13g2_fill_2 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_340 ();
 sg13g2_fill_2 FILLER_30_352 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_fill_2 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_379 ();
 sg13g2_fill_1 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_4 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_30_410 ();
 sg13g2_decap_8 FILLER_30_417 ();
 sg13g2_decap_4 FILLER_30_424 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_23 ();
 sg13g2_fill_2 FILLER_31_33 ();
 sg13g2_fill_1 FILLER_31_54 ();
 sg13g2_fill_2 FILLER_31_60 ();
 sg13g2_fill_1 FILLER_31_79 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_121 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_decap_4 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_decap_4 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_decap_4 FILLER_31_188 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_decap_4 FILLER_31_197 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_decap_8 FILLER_31_206 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_fill_2 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_277 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_301 ();
 sg13g2_decap_4 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_decap_4 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_331 ();
 sg13g2_decap_4 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_341 ();
 sg13g2_decap_4 FILLER_31_352 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_fill_1 FILLER_31_381 ();
 sg13g2_fill_2 FILLER_31_428 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_21 ();
 sg13g2_fill_1 FILLER_32_23 ();
 sg13g2_fill_1 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_decap_8 FILLER_32_148 ();
 sg13g2_decap_4 FILLER_32_155 ();
 sg13g2_fill_1 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_decap_4 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_335 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_fill_2 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_4 FILLER_32_382 ();
 sg13g2_fill_1 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_fill_2 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_fill_1 FILLER_33_31 ();
 sg13g2_fill_2 FILLER_33_52 ();
 sg13g2_decap_4 FILLER_33_64 ();
 sg13g2_decap_4 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_decap_4 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_130 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_decap_4 FILLER_33_200 ();
 sg13g2_fill_2 FILLER_33_204 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_decap_8 FILLER_33_241 ();
 sg13g2_decap_8 FILLER_33_248 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_decap_4 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_345 ();
 sg13g2_decap_8 FILLER_33_351 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_decap_4 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_42 ();
 sg13g2_fill_2 FILLER_34_48 ();
 sg13g2_fill_2 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_1 FILLER_34_80 ();
 sg13g2_decap_4 FILLER_34_86 ();
 sg13g2_fill_2 FILLER_34_90 ();
 sg13g2_fill_1 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_decap_4 FILLER_34_130 ();
 sg13g2_fill_2 FILLER_34_134 ();
 sg13g2_decap_8 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_decap_8 FILLER_34_157 ();
 sg13g2_decap_8 FILLER_34_164 ();
 sg13g2_decap_8 FILLER_34_171 ();
 sg13g2_decap_4 FILLER_34_178 ();
 sg13g2_decap_8 FILLER_34_208 ();
 sg13g2_decap_8 FILLER_34_215 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_251 ();
 sg13g2_decap_4 FILLER_34_258 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_fill_1 FILLER_34_280 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_319 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_fill_2 FILLER_34_352 ();
 sg13g2_decap_4 FILLER_34_365 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_382 ();
 sg13g2_fill_2 FILLER_34_387 ();
 sg13g2_fill_1 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_414 ();
 sg13g2_decap_8 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_38 ();
 sg13g2_decap_4 FILLER_35_45 ();
 sg13g2_decap_8 FILLER_35_54 ();
 sg13g2_fill_2 FILLER_35_61 ();
 sg13g2_fill_1 FILLER_35_63 ();
 sg13g2_decap_4 FILLER_35_83 ();
 sg13g2_fill_1 FILLER_35_87 ();
 sg13g2_decap_4 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_104 ();
 sg13g2_decap_4 FILLER_35_111 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_decap_8 FILLER_35_128 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_decap_8 FILLER_35_141 ();
 sg13g2_decap_4 FILLER_35_148 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_186 ();
 sg13g2_decap_4 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_decap_8 FILLER_35_216 ();
 sg13g2_fill_1 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_decap_4 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_260 ();
 sg13g2_decap_8 FILLER_35_267 ();
 sg13g2_decap_8 FILLER_35_274 ();
 sg13g2_decap_8 FILLER_35_281 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_fill_1 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_339 ();
 sg13g2_decap_4 FILLER_35_346 ();
 sg13g2_decap_8 FILLER_35_355 ();
 sg13g2_decap_4 FILLER_35_362 ();
 sg13g2_fill_2 FILLER_35_366 ();
 sg13g2_decap_4 FILLER_35_382 ();
 sg13g2_fill_1 FILLER_35_395 ();
 sg13g2_fill_2 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_48 ();
 sg13g2_decap_8 FILLER_36_54 ();
 sg13g2_decap_8 FILLER_36_61 ();
 sg13g2_decap_8 FILLER_36_68 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_decap_8 FILLER_36_90 ();
 sg13g2_decap_8 FILLER_36_97 ();
 sg13g2_decap_8 FILLER_36_108 ();
 sg13g2_decap_8 FILLER_36_115 ();
 sg13g2_decap_8 FILLER_36_122 ();
 sg13g2_fill_1 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_165 ();
 sg13g2_decap_8 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_197 ();
 sg13g2_decap_4 FILLER_36_219 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_fill_2 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_fill_2 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_253 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_fill_1 FILLER_36_384 ();
 sg13g2_decap_4 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_394 ();
 sg13g2_fill_1 FILLER_36_403 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_decap_4 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_149 ();
 sg13g2_fill_1 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_decap_4 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_193 ();
 sg13g2_decap_4 FILLER_37_199 ();
 sg13g2_fill_2 FILLER_37_212 ();
 sg13g2_fill_1 FILLER_37_218 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_229 ();
 sg13g2_fill_1 FILLER_37_236 ();
 sg13g2_decap_4 FILLER_37_270 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_decap_8 FILLER_37_284 ();
 sg13g2_decap_8 FILLER_37_291 ();
 sg13g2_decap_4 FILLER_37_364 ();
 sg13g2_fill_2 FILLER_37_368 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_419 ();
 sg13g2_decap_4 FILLER_37_426 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_fill_1 FILLER_38_158 ();
 sg13g2_fill_1 FILLER_38_164 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_fill_2 FILLER_38_231 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_326 ();
 sg13g2_fill_2 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_377 ();
 sg13g2_decap_4 FILLER_38_384 ();
 sg13g2_fill_2 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_421 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
