module tt_um_silice (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire _4601_;
 wire _4602_;
 wire _4603_;
 wire _4604_;
 wire _4605_;
 wire _4606_;
 wire _4607_;
 wire _4608_;
 wire _4609_;
 wire _4610_;
 wire _4611_;
 wire _4612_;
 wire _4613_;
 wire _4614_;
 wire _4615_;
 wire _4616_;
 wire _4617_;
 wire _4618_;
 wire _4619_;
 wire _4620_;
 wire _4621_;
 wire _4622_;
 wire _4623_;
 wire _4624_;
 wire _4625_;
 wire _4626_;
 wire _4627_;
 wire _4628_;
 wire _4629_;
 wire _4630_;
 wire _4631_;
 wire _4632_;
 wire _4633_;
 wire _4634_;
 wire clknet_leaf_0_clk;
 wire net92;
 wire \main._w_demo_audio1 ;
 wire \main._w_demo_video_hs ;
 wire \main._w_demo_video_vs ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[1] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[2] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[3] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[4] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[6] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[7] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[0] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[10] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[7] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[8] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[9] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[0] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[10] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[1] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[2] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[3] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[4] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[5] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[6] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[7] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[8] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[9] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[1] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[2] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[3] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[4] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[5] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[6] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[7] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[0] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[10] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[7] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[8] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[9] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[1] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[2] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[3] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[4] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[5] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[6] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[7] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[0] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[10] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[7] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[8] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[9] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[0] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[1] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[2] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[3] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[4] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[5] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_h[0] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_h[1] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_h[2] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_l[0] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_l[1] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[9] ;
 wire \main.demo._d_prev_b[0] ;
 wire \main.demo._d_prev_b[1] ;
 wire \main.demo._d_prev_b[2] ;
 wire \main.demo._d_prev_b[3] ;
 wire \main.demo._d_prev_b[4] ;
 wire \main.demo._d_prev_b[5] ;
 wire \main.demo._d_prev_b[6] ;
 wire \main.demo._d_prev_b[7] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[0] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[10] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[1] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[2] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[3] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[4] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[5] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[6] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[7] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[8] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[9] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[0] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[10] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[1] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[2] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[3] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[4] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[5] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[6] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[7] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[8] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[9] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[1] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[2] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[3] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[4] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[6] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[7] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[0] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[10] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[1] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[2] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[3] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[4] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[5] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[6] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[7] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[8] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[9] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[0] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[10] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[1] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[2] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[3] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[4] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[5] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[6] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[7] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[8] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[9] ;
 wire \main.demo._q_effect[0] ;
 wire \main.demo._q_effect[1] ;
 wire \main.demo._q_frame[0] ;
 wire \main.demo._q_frame[10] ;
 wire \main.demo._q_frame[11] ;
 wire \main.demo._q_frame[12] ;
 wire \main.demo._q_frame[13] ;
 wire \main.demo._q_frame[14] ;
 wire \main.demo._q_frame[1] ;
 wire \main.demo._q_frame[2] ;
 wire \main.demo._q_frame[3] ;
 wire \main.demo._q_frame[4] ;
 wire \main.demo._q_frame[5] ;
 wire \main.demo._q_frame[6] ;
 wire \main.demo._q_frame[7] ;
 wire \main.demo._q_frame[8] ;
 wire \main.demo._q_frame[9] ;
 wire \main.demo._q_go ;
 wire \main.demo._q_prev_b[6] ;
 wire \main.demo._q_prev_b[7] ;
 wire \main.demo._q_prev_vs ;
 wire \main.demo._q_rot_en ;
 wire \main.demo._q_speed[0] ;
 wire \main.demo._q_speed[10] ;
 wire \main.demo._q_speed[11] ;
 wire \main.demo._q_speed[12] ;
 wire \main.demo._q_speed[13] ;
 wire \main.demo._q_speed[14] ;
 wire \main.demo._q_speed[15] ;
 wire \main.demo._q_speed[1] ;
 wire \main.demo._q_speed[2] ;
 wire \main.demo._q_speed[3] ;
 wire \main.demo._q_speed[4] ;
 wire \main.demo._q_speed[5] ;
 wire \main.demo._q_speed[6] ;
 wire \main.demo._q_speed[7] ;
 wire \main.demo._q_speed[8] ;
 wire \main.demo._q_speed[9] ;
 wire \main.demo._q_th[0] ;
 wire \main.demo._q_th[1] ;
 wire \main.demo._q_th[2] ;
 wire \main.demo._q_th[3] ;
 wire \main.demo._q_th[4] ;
 wire \main.demo._q_th[5] ;
 wire \main.demo._q_th[6] ;
 wire \main.demo._q_th[7] ;
 wire \main.demo._q_th[8] ;
 wire \main.demo._t___block_68_frag[0] ;
 wire \main.demo._t___block_68_frag[1] ;
 wire \main.demo._t___block_68_frag[2] ;
 wire \main.demo._t___block_68_frag[3] ;
 wire \main.demo._t___block_68_frag[4] ;
 wire \main.demo._t___block_68_frag[5] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_a[6] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_a[7] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[0] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[10] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[1] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[2] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[3] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[4] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[5] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[6] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[7] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[8] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[9] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[0] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[10] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[1] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[2] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[3] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[4] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[5] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[6] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[7] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[8] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[9] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_h[0] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_h[1] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_h[2] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_l[0] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_l[1] ;
 wire \main.demo._t___stage___block_3_x[0] ;
 wire \main.demo._t___stage___block_3_x[1] ;
 wire \main.demo._t___stage___block_3_x[2] ;
 wire \main.demo._t___stage___block_3_y[0] ;
 wire \main.demo._t___stage___block_3_y[1] ;
 wire \main.demo._t___stage___block_3_y[2] ;
 wire \main.demo._w_vga_active ;
 wire \main.demo._w_vga_vga_x[10] ;
 wire \main.demo._w_vga_vga_x[3] ;
 wire \main.demo._w_vga_vga_x[4] ;
 wire \main.demo._w_vga_vga_x[5] ;
 wire \main.demo._w_vga_vga_x[6] ;
 wire \main.demo._w_vga_vga_x[7] ;
 wire \main.demo._w_vga_vga_x[8] ;
 wire \main.demo._w_vga_vga_x[9] ;
 wire \main.demo._w_vga_vga_y[10] ;
 wire \main.demo._w_vga_vga_y[3] ;
 wire \main.demo._w_vga_vga_y[4] ;
 wire \main.demo._w_vga_vga_y[5] ;
 wire \main.demo._w_vga_vga_y[6] ;
 wire \main.demo._w_vga_vga_y[7] ;
 wire \main.demo._w_vga_vga_y[8] ;
 wire \main.demo.vga._d_active ;
 wire \main.demo.vga._d_vblank ;
 wire \main.demo.vga._q_active_h ;
 wire \main.demo.vga._q_active_v ;
 wire \main.demo.vga._q_xcount[0] ;
 wire \main.demo.vga._q_xcount[10] ;
 wire \main.demo.vga._q_xcount[1] ;
 wire \main.demo.vga._q_xcount[2] ;
 wire \main.demo.vga._q_xcount[3] ;
 wire \main.demo.vga._q_xcount[4] ;
 wire \main.demo.vga._q_xcount[5] ;
 wire \main.demo.vga._q_xcount[6] ;
 wire \main.demo.vga._q_xcount[7] ;
 wire \main.demo.vga._q_xcount[8] ;
 wire \main.demo.vga._q_xcount[9] ;
 wire \main.demo.vga._q_ycount[0] ;
 wire \main.demo.vga._q_ycount[1] ;
 wire \main.demo.vga._q_ycount[2] ;
 wire \main.demo.vga._q_ycount[3] ;
 wire \main.demo.vga._q_ycount[4] ;
 wire \main.demo.vga._q_ycount[5] ;
 wire \main.demo.vga._q_ycount[6] ;
 wire \main.demo.vga._q_ycount[7] ;
 wire \main.demo.vga._q_ycount[8] ;
 wire \main.demo.zic._q_clock_count[0] ;
 wire \main.demo.zic._q_clock_count[1] ;
 wire \main.demo.zic._q_clock_count[2] ;
 wire \main.demo.zic._q_clock_count[3] ;
 wire \main.demo.zic._q_clock_count[4] ;
 wire \main.demo.zic._q_clock_count[5] ;
 wire \main.demo.zic._q_clock_count[6] ;
 wire \main.demo.zic._q_clock_count[7] ;
 wire \main.demo.zic._q_clock_count[8] ;
 wire \main.demo.zic._q_drum_inc[0] ;
 wire \main.demo.zic._q_drum_inc[1] ;
 wire \main.demo.zic._q_drum_inc[2] ;
 wire \main.demo.zic._q_drum_inc[3] ;
 wire \main.demo.zic._q_idx[0] ;
 wire \main.demo.zic._q_idx[1] ;
 wire \main.demo.zic._q_idx[2] ;
 wire \main.demo.zic._q_idx[3] ;
 wire \main.demo.zic._q_idx[4] ;
 wire \main.demo.zic._q_idx[5] ;
 wire \main.demo.zic._q_idx[6] ;
 wire \main.demo.zic._q_qpos[0] ;
 wire \main.demo.zic._q_qpos[10] ;
 wire \main.demo.zic._q_qpos[11] ;
 wire \main.demo.zic._q_qpos[12] ;
 wire \main.demo.zic._q_qpos[1] ;
 wire \main.demo.zic._q_qpos[2] ;
 wire \main.demo.zic._q_qpos[3] ;
 wire \main.demo.zic._q_qpos[4] ;
 wire \main.demo.zic._q_qpos[5] ;
 wire \main.demo.zic._q_qpos[6] ;
 wire \main.demo.zic._q_qpos[7] ;
 wire \main.demo.zic._q_qpos[8] ;
 wire \main.demo.zic._q_qpos[9] ;
 wire \main.demo.zic._q_rythm_count[0] ;
 wire \main.demo.zic._q_rythm_count[10] ;
 wire \main.demo.zic._q_rythm_count[11] ;
 wire \main.demo.zic._q_rythm_count[12] ;
 wire \main.demo.zic._q_rythm_count[1] ;
 wire \main.demo.zic._q_rythm_count[2] ;
 wire \main.demo.zic._q_rythm_count[3] ;
 wire \main.demo.zic._q_rythm_count[4] ;
 wire \main.demo.zic._q_rythm_count[5] ;
 wire \main.demo.zic._q_rythm_count[6] ;
 wire \main.demo.zic._q_rythm_count[7] ;
 wire \main.demo.zic._q_rythm_count[8] ;
 wire \main.demo.zic._q_rythm_count[9] ;
 wire \main.demo.zic._q_squ_env[0] ;
 wire \main.demo.zic._q_squ_env[1] ;
 wire \main.demo.zic._q_squ_env[2] ;
 wire \main.demo.zic._q_squ_env[3] ;
 wire \main.demo.zic._q_squ_env[4] ;
 wire \main.demo.zic._q_squ_env[5] ;
 wire \main.demo.zic._q_tpos[0] ;
 wire \main.demo.zic._q_tpos[10] ;
 wire \main.demo.zic._q_tpos[11] ;
 wire \main.demo.zic._q_tpos[1] ;
 wire \main.demo.zic._q_tpos[2] ;
 wire \main.demo.zic._q_tpos[3] ;
 wire \main.demo.zic._q_tpos[4] ;
 wire \main.demo.zic._q_tpos[5] ;
 wire \main.demo.zic._q_tpos[6] ;
 wire \main.demo.zic._q_tpos[7] ;
 wire \main.demo.zic._q_tpos[8] ;
 wire \main.demo.zic._q_tpos[9] ;
 wire rst_n_q;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_inv_1 _4637_ (.Y(_4031_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[10] ));
 sg13g2_inv_1 _4638_ (.Y(_4032_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ));
 sg13g2_nor2_1 _4639_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ),
    .B(_4032_),
    .Y(_4033_));
 sg13g2_nand2_1 _4640_ (.Y(_4034_),
    .A(_4032_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ));
 sg13g2_inv_1 _4641_ (.Y(_4035_),
    .A(_4034_));
 sg13g2_nor2_1 _4642_ (.A(_4033_),
    .B(_4035_),
    .Y(_4036_));
 sg13g2_inv_1 _4643_ (.Y(_4037_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ));
 sg13g2_inv_1 _4644_ (.Y(_4038_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ));
 sg13g2_inv_1 _4645_ (.Y(_4039_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ));
 sg13g2_inv_1 _4646_ (.Y(_4040_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ));
 sg13g2_inv_1 _4647_ (.Y(_4041_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ));
 sg13g2_inv_1 _4648_ (.Y(_4042_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ));
 sg13g2_inv_1 _4649_ (.Y(_4043_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ));
 sg13g2_inv_1 _4650_ (.Y(_4044_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_inv_1 _4651_ (.Y(_4045_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ));
 sg13g2_inv_1 _4652_ (.Y(_4046_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ));
 sg13g2_inv_1 _4653_ (.Y(_4047_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ));
 sg13g2_inv_1 _4654_ (.Y(_4048_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ));
 sg13g2_inv_1 _4655_ (.Y(_4049_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ));
 sg13g2_inv_1 _4656_ (.Y(_4050_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ));
 sg13g2_nand2_1 _4657_ (.Y(_4051_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ));
 sg13g2_inv_1 _4658_ (.Y(_4052_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ));
 sg13g2_nor2_1 _4659_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ),
    .B(_4052_),
    .Y(_4053_));
 sg13g2_inv_1 _4660_ (.Y(_4054_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ));
 sg13g2_nor2_1 _4661_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ),
    .B(_4054_),
    .Y(_4055_));
 sg13g2_nor2_2 _4662_ (.A(_4053_),
    .B(_4055_),
    .Y(_4056_));
 sg13g2_nand2_1 _4663_ (.Y(_4057_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ));
 sg13g2_o21ai_1 _4664_ (.B1(_4057_),
    .Y(_4058_),
    .A1(_4051_),
    .A2(_4056_));
 sg13g2_nor2_1 _4665_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ),
    .B(_4049_),
    .Y(_4059_));
 sg13g2_nor2_1 _4666_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ),
    .B(_4050_),
    .Y(_4060_));
 sg13g2_nor2_1 _4667_ (.A(_4059_),
    .B(_4060_),
    .Y(_4061_));
 sg13g2_inv_1 _4668_ (.Y(_4062_),
    .A(_4061_));
 sg13g2_nand2_1 _4669_ (.Y(_4063_),
    .A(_4058_),
    .B(_4062_));
 sg13g2_o21ai_1 _4670_ (.B1(_4063_),
    .Y(_4064_),
    .A1(_4049_),
    .A2(_4050_));
 sg13g2_nor2_2 _4671_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ),
    .B(_4048_),
    .Y(_4065_));
 sg13g2_nor2_2 _4672_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ),
    .B(_4047_),
    .Y(_4066_));
 sg13g2_nor2_2 _4673_ (.A(_4065_),
    .B(_4066_),
    .Y(_4067_));
 sg13g2_inv_1 _4674_ (.Y(_4068_),
    .A(_4067_));
 sg13g2_nand2_1 _4675_ (.Y(_4069_),
    .A(_4064_),
    .B(_4068_));
 sg13g2_o21ai_1 _4676_ (.B1(_4069_),
    .Y(_4070_),
    .A1(_4047_),
    .A2(_4048_));
 sg13g2_nor2_1 _4677_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ),
    .B(_4046_),
    .Y(_4071_));
 sg13g2_nor2_1 _4678_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ),
    .B(_4045_),
    .Y(_4072_));
 sg13g2_nor2_2 _4679_ (.A(_4071_),
    .B(_4072_),
    .Y(_4073_));
 sg13g2_inv_1 _4680_ (.Y(_4074_),
    .A(_4073_));
 sg13g2_nand2_1 _4681_ (.Y(_4075_),
    .A(_4070_),
    .B(_4074_));
 sg13g2_o21ai_1 _4682_ (.B1(_4075_),
    .Y(_4076_),
    .A1(_4045_),
    .A2(_4046_));
 sg13g2_nor2_1 _4683_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ),
    .B(_4044_),
    .Y(_4077_));
 sg13g2_nor2_1 _4684_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ),
    .B(_4043_),
    .Y(_4078_));
 sg13g2_nor2_1 _4685_ (.A(_4077_),
    .B(_4078_),
    .Y(_4079_));
 sg13g2_buf_2 _4686_ (.A(_4079_),
    .X(_4080_));
 sg13g2_inv_1 _4687_ (.Y(_4081_),
    .A(_4080_));
 sg13g2_nand2_1 _4688_ (.Y(_4082_),
    .A(_4076_),
    .B(_4081_));
 sg13g2_o21ai_1 _4689_ (.B1(_4082_),
    .Y(_4083_),
    .A1(_4043_),
    .A2(_4044_));
 sg13g2_nor2_1 _4690_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ),
    .B(_4042_),
    .Y(_4084_));
 sg13g2_nor2_1 _4691_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ),
    .B(_4041_),
    .Y(_4085_));
 sg13g2_nor2_2 _4692_ (.A(_4084_),
    .B(_4085_),
    .Y(_4086_));
 sg13g2_inv_1 _4693_ (.Y(_4087_),
    .A(_4086_));
 sg13g2_nand2_1 _4694_ (.Y(_4088_),
    .A(_4083_),
    .B(_4087_));
 sg13g2_o21ai_1 _4695_ (.B1(_4088_),
    .Y(_4089_),
    .A1(_4041_),
    .A2(_4042_));
 sg13g2_nor2_1 _4696_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ),
    .B(_4040_),
    .Y(_4090_));
 sg13g2_nor2_1 _4697_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ),
    .B(_4039_),
    .Y(_4091_));
 sg13g2_nor2_2 _4698_ (.A(_4090_),
    .B(_4091_),
    .Y(_4092_));
 sg13g2_inv_2 _4699_ (.Y(_4093_),
    .A(_4092_));
 sg13g2_nand2_1 _4700_ (.Y(_4094_),
    .A(_4089_),
    .B(_4093_));
 sg13g2_o21ai_1 _4701_ (.B1(_4094_),
    .Y(_4095_),
    .A1(_4039_),
    .A2(_4040_));
 sg13g2_nor2_1 _4702_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ),
    .B(_4038_),
    .Y(_4096_));
 sg13g2_nor2_1 _4703_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ),
    .B(_4037_),
    .Y(_4097_));
 sg13g2_nor2_1 _4704_ (.A(_4096_),
    .B(_4097_),
    .Y(_4098_));
 sg13g2_buf_2 _4705_ (.A(_4098_),
    .X(_4099_));
 sg13g2_inv_1 _4706_ (.Y(_4100_),
    .A(_4099_));
 sg13g2_nand2_1 _4707_ (.Y(_4101_),
    .A(_4095_),
    .B(_4100_));
 sg13g2_o21ai_1 _4708_ (.B1(_4101_),
    .Y(_4102_),
    .A1(_4037_),
    .A2(_4038_));
 sg13g2_nor2b_1 _4709_ (.A(_4036_),
    .B_N(_4102_),
    .Y(_4103_));
 sg13g2_a21oi_1 _4710_ (.A1(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ),
    .A2(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ),
    .Y(_4104_),
    .B1(_4103_));
 sg13g2_inv_1 _4711_ (.Y(_4105_),
    .A(_4036_));
 sg13g2_nor2_1 _4712_ (.A(_4100_),
    .B(_4105_),
    .Y(_4106_));
 sg13g2_a21oi_1 _4713_ (.A1(_4092_),
    .A2(_4084_),
    .Y(_4107_),
    .B1(_4090_));
 sg13g2_inv_1 _4714_ (.Y(_4108_),
    .A(_4107_));
 sg13g2_inv_1 _4715_ (.Y(_4109_),
    .A(_4066_));
 sg13g2_inv_1 _4716_ (.Y(_4110_),
    .A(_4059_));
 sg13g2_a21oi_1 _4717_ (.A1(_4109_),
    .A2(_4110_),
    .Y(_4111_),
    .B1(_4065_));
 sg13g2_inv_1 _4718_ (.Y(_4112_),
    .A(_4111_));
 sg13g2_nor2_1 _4719_ (.A(_4081_),
    .B(_4074_),
    .Y(_4113_));
 sg13g2_inv_1 _4720_ (.Y(_4114_),
    .A(_4113_));
 sg13g2_a21oi_1 _4721_ (.A1(_4080_),
    .A2(_4071_),
    .Y(_4115_),
    .B1(_4077_));
 sg13g2_o21ai_1 _4722_ (.B1(_4115_),
    .Y(_4116_),
    .A1(_4112_),
    .A2(_4114_));
 sg13g2_nor2_1 _4723_ (.A(_4093_),
    .B(_4087_),
    .Y(_4117_));
 sg13g2_and2_1 _4724_ (.A(_4106_),
    .B(_4117_),
    .X(_4118_));
 sg13g2_buf_1 _4725_ (.A(_4118_),
    .X(_4119_));
 sg13g2_a21o_1 _4726_ (.A2(_4034_),
    .A1(_4096_),
    .B1(_4033_),
    .X(_4120_));
 sg13g2_a221oi_1 _4727_ (.B2(_4119_),
    .C1(_4120_),
    .B1(_4116_),
    .A1(_4106_),
    .Y(_4121_),
    .A2(_4108_));
 sg13g2_nor2_1 _4728_ (.A(_4068_),
    .B(_4062_),
    .Y(_4122_));
 sg13g2_inv_1 _4729_ (.Y(_4123_),
    .A(_4122_));
 sg13g2_nor2_1 _4730_ (.A(_4114_),
    .B(_4123_),
    .Y(_4124_));
 sg13g2_inv_1 _4731_ (.Y(_4125_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ));
 sg13g2_nor2_1 _4732_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ),
    .B(_4125_),
    .Y(_4126_));
 sg13g2_inv_1 _4733_ (.Y(_4127_),
    .A(_4126_));
 sg13g2_nand2_1 _4734_ (.Y(_4128_),
    .A(_4056_),
    .B(_4127_));
 sg13g2_inv_1 _4735_ (.Y(_4129_),
    .A(_4053_));
 sg13g2_nand2_2 _4736_ (.Y(_4130_),
    .A(_4128_),
    .B(_4129_));
 sg13g2_nand3_1 _4737_ (.B(_4124_),
    .C(_4130_),
    .A(_4119_),
    .Y(_4131_));
 sg13g2_buf_1 _4738_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[10] ),
    .X(_4132_));
 sg13g2_a21o_1 _4739_ (.A2(_4131_),
    .A1(_4121_),
    .B1(net77),
    .X(_4133_));
 sg13g2_o21ai_1 _4740_ (.B1(_4133_),
    .Y(_4134_),
    .A1(_4031_),
    .A2(_4104_));
 sg13g2_nand2b_1 _4741_ (.Y(_4135_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ),
    .A_N(_4134_));
 sg13g2_nand2b_1 _4742_ (.Y(_4136_),
    .B(_4134_),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ));
 sg13g2_nand2_1 _4743_ (.Y(_4137_),
    .A(_4135_),
    .B(_4136_));
 sg13g2_buf_2 _4744_ (.A(_4137_),
    .X(_4138_));
 sg13g2_buf_1 _4745_ (.A(_4138_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ));
 sg13g2_buf_2 _4746_ (.A(\main.demo._q_rot_en ),
    .X(_4139_));
 sg13g2_buf_1 _4747_ (.A(\main.demo._q_frame[6] ),
    .X(_4140_));
 sg13g2_buf_1 _4748_ (.A(\main.demo._w_vga_vga_y[8] ),
    .X(_4141_));
 sg13g2_a21oi_1 _4749_ (.A1(_4139_),
    .A2(_4140_),
    .Y(_4142_),
    .B1(_4141_));
 sg13g2_nand2_1 _4750_ (.Y(_4143_),
    .A(_4139_),
    .B(_4140_));
 sg13g2_xnor2_1 _4751_ (.Y(_4144_),
    .A(\main.demo._w_vga_vga_y[10] ),
    .B(_4143_));
 sg13g2_nor2_1 _4752_ (.A(_4142_),
    .B(_4144_),
    .Y(_4145_));
 sg13g2_buf_2 _4753_ (.A(\main.demo._q_frame[4] ),
    .X(_4146_));
 sg13g2_inv_1 _4754_ (.Y(_4147_),
    .A(_4140_));
 sg13g2_buf_1 _4755_ (.A(\main.demo._q_frame[5] ),
    .X(_4148_));
 sg13g2_inv_1 _4756_ (.Y(_4149_),
    .A(_4148_));
 sg13g2_nand2_1 _4757_ (.Y(_4150_),
    .A(_4147_),
    .B(_4149_));
 sg13g2_nand2_1 _4758_ (.Y(_4151_),
    .A(_4140_),
    .B(_4148_));
 sg13g2_nand2_1 _4759_ (.Y(_4152_),
    .A(_4150_),
    .B(_4151_));
 sg13g2_inv_1 _4760_ (.Y(_4153_),
    .A(_4152_));
 sg13g2_buf_1 _4761_ (.A(_4153_),
    .X(_4154_));
 sg13g2_inv_2 _4762_ (.Y(_4155_),
    .A(_4139_));
 sg13g2_a21oi_1 _4763_ (.A1(net42),
    .A2(_4146_),
    .Y(_4156_),
    .B1(_4155_));
 sg13g2_o21ai_1 _4764_ (.B1(_4156_),
    .Y(_4157_),
    .A1(_4146_),
    .A2(net42));
 sg13g2_xnor2_1 _4765_ (.Y(_4158_),
    .A(_0008_),
    .B(_4157_));
 sg13g2_buf_1 _4766_ (.A(\main.demo._q_frame[3] ),
    .X(_4159_));
 sg13g2_a21oi_1 _4767_ (.A1(net42),
    .A2(_4159_),
    .Y(_4160_),
    .B1(_4155_));
 sg13g2_o21ai_1 _4768_ (.B1(_4160_),
    .Y(_4161_),
    .A1(_4159_),
    .A2(net42));
 sg13g2_nor2_1 _4769_ (.A(_0009_),
    .B(_4161_),
    .Y(_4162_));
 sg13g2_inv_1 _4770_ (.Y(_4163_),
    .A(_4162_));
 sg13g2_buf_2 _4771_ (.A(\main.demo._q_frame[0] ),
    .X(_4164_));
 sg13g2_nor2b_1 _4772_ (.A(_4152_),
    .B_N(_4164_),
    .Y(_4165_));
 sg13g2_nor2_1 _4773_ (.A(_4164_),
    .B(_4153_),
    .Y(_4166_));
 sg13g2_nor3_1 _4774_ (.A(_4155_),
    .B(_4165_),
    .C(_4166_),
    .Y(_4167_));
 sg13g2_nor2b_1 _4775_ (.A(_0011_),
    .B_N(_4167_),
    .Y(_4168_));
 sg13g2_inv_1 _4776_ (.Y(_4169_),
    .A(_4168_));
 sg13g2_buf_1 _4777_ (.A(\main.demo._w_vga_vga_y[4] ),
    .X(_4170_));
 sg13g2_buf_1 _4778_ (.A(\main.demo._q_frame[1] ),
    .X(_4171_));
 sg13g2_a21oi_1 _4779_ (.A1(net42),
    .A2(_4171_),
    .Y(_4172_),
    .B1(_4155_));
 sg13g2_o21ai_1 _4780_ (.B1(_4172_),
    .Y(_4173_),
    .A1(_4171_),
    .A2(net42));
 sg13g2_xnor2_1 _4781_ (.Y(_4174_),
    .A(_4170_),
    .B(_4173_));
 sg13g2_nor2_1 _4782_ (.A(_4169_),
    .B(_4174_),
    .Y(_4175_));
 sg13g2_inv_1 _4783_ (.Y(_4176_),
    .A(_4175_));
 sg13g2_inv_1 _4784_ (.Y(_4177_),
    .A(_4170_));
 sg13g2_nand2_1 _4785_ (.Y(_4178_),
    .A(_4173_),
    .B(_4177_));
 sg13g2_buf_1 _4786_ (.A(\main.demo._q_frame[2] ),
    .X(_4179_));
 sg13g2_a21oi_1 _4787_ (.A1(net42),
    .A2(_4179_),
    .Y(_4180_),
    .B1(_4155_));
 sg13g2_o21ai_1 _4788_ (.B1(_4180_),
    .Y(_4181_),
    .A1(_4179_),
    .A2(net42));
 sg13g2_xnor2_1 _4789_ (.Y(_4182_),
    .A(_0010_),
    .B(_4181_));
 sg13g2_xor2_1 _4790_ (.B(_4182_),
    .A(_4178_),
    .X(_4183_));
 sg13g2_nand2b_1 _4791_ (.Y(_4184_),
    .B(_4178_),
    .A_N(_4182_));
 sg13g2_o21ai_1 _4792_ (.B1(_4184_),
    .Y(_4185_),
    .A1(_4176_),
    .A2(_4183_));
 sg13g2_xnor2_1 _4793_ (.Y(_4186_),
    .A(_0009_),
    .B(_4161_));
 sg13g2_nor2_1 _4794_ (.A(_0010_),
    .B(_4181_),
    .Y(_4187_));
 sg13g2_inv_1 _4795_ (.Y(_4188_),
    .A(_4187_));
 sg13g2_nand2_1 _4796_ (.Y(_4189_),
    .A(_4186_),
    .B(_4188_));
 sg13g2_nor2_1 _4797_ (.A(_4188_),
    .B(_4186_),
    .Y(_4190_));
 sg13g2_a21o_1 _4798_ (.A2(_4189_),
    .A1(_4185_),
    .B1(_4190_),
    .X(_4191_));
 sg13g2_xnor2_1 _4799_ (.Y(_4192_),
    .A(_4162_),
    .B(_4158_));
 sg13g2_nand2_1 _4800_ (.Y(_4193_),
    .A(_4191_),
    .B(_4192_));
 sg13g2_o21ai_1 _4801_ (.B1(_4193_),
    .Y(_4194_),
    .A1(_4158_),
    .A2(_4163_));
 sg13g2_xnor2_1 _4802_ (.Y(_4195_),
    .A(_4141_),
    .B(_4143_));
 sg13g2_nor2_1 _4803_ (.A(_0008_),
    .B(_4157_),
    .Y(_4196_));
 sg13g2_xnor2_1 _4804_ (.Y(_4197_),
    .A(_4195_),
    .B(_4196_));
 sg13g2_nor3_1 _4805_ (.A(_0008_),
    .B(_4195_),
    .C(_4157_),
    .Y(_4198_));
 sg13g2_a21oi_1 _4806_ (.A1(_4194_),
    .A2(_4197_),
    .Y(_4199_),
    .B1(_4198_));
 sg13g2_inv_1 _4807_ (.Y(_4200_),
    .A(_4199_));
 sg13g2_nand2_1 _4808_ (.Y(_4201_),
    .A(_4144_),
    .B(_4142_));
 sg13g2_o21ai_1 _4809_ (.B1(_4201_),
    .Y(_4202_),
    .A1(_4145_),
    .A2(_4200_));
 sg13g2_nor2_1 _4810_ (.A(_0007_),
    .B(_4143_),
    .Y(_4203_));
 sg13g2_nand2b_1 _4811_ (.Y(_4204_),
    .B(_4203_),
    .A_N(_4202_));
 sg13g2_nand2b_1 _4812_ (.Y(_4205_),
    .B(_4202_),
    .A_N(_4203_));
 sg13g2_nand2_1 _4813_ (.Y(_4206_),
    .A(_4204_),
    .B(_4205_));
 sg13g2_inv_1 _4814_ (.Y(_4207_),
    .A(_4206_));
 sg13g2_buf_1 _4815_ (.A(_4207_),
    .X(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ));
 sg13g2_inv_1 _4816_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ),
    .A(_4138_));
 sg13g2_buf_1 _4817_ (.A(\main.demo._q_speed[10] ),
    .X(_4208_));
 sg13g2_inv_1 _4818_ (.Y(_4209_),
    .A(_4208_));
 sg13g2_buf_2 _4819_ (.A(\main.demo._q_speed[9] ),
    .X(_4210_));
 sg13g2_buf_1 _4820_ (.A(\main.demo._q_speed[15] ),
    .X(_4211_));
 sg13g2_xor2_1 _4821_ (.B(_4211_),
    .A(_4210_),
    .X(_4212_));
 sg13g2_inv_1 _4822_ (.Y(_4213_),
    .A(_4212_));
 sg13g2_buf_2 _4823_ (.A(\main.demo._q_speed[8] ),
    .X(_4214_));
 sg13g2_buf_2 _4824_ (.A(\main.demo._q_speed[14] ),
    .X(_4215_));
 sg13g2_nor2_1 _4825_ (.A(_4214_),
    .B(_4215_),
    .Y(_4216_));
 sg13g2_buf_2 _4826_ (.A(\main.demo._q_speed[7] ),
    .X(_4217_));
 sg13g2_buf_1 _4827_ (.A(\main.demo._q_speed[13] ),
    .X(_4218_));
 sg13g2_nor2_1 _4828_ (.A(_4217_),
    .B(_4218_),
    .Y(_4219_));
 sg13g2_buf_1 _4829_ (.A(\main.demo._q_speed[4] ),
    .X(_4220_));
 sg13g2_xor2_1 _4830_ (.B(_4220_),
    .A(_4208_),
    .X(_4221_));
 sg13g2_inv_1 _4831_ (.Y(_4222_),
    .A(_4221_));
 sg13g2_buf_2 _4832_ (.A(\main.demo._q_speed[3] ),
    .X(_4223_));
 sg13g2_xor2_1 _4833_ (.B(_4210_),
    .A(_4223_),
    .X(_4224_));
 sg13g2_inv_1 _4834_ (.Y(_4225_),
    .A(_4224_));
 sg13g2_buf_2 _4835_ (.A(\main.demo._q_speed[2] ),
    .X(_4226_));
 sg13g2_xor2_1 _4836_ (.B(_4214_),
    .A(_4226_),
    .X(_4227_));
 sg13g2_inv_1 _4837_ (.Y(_4228_),
    .A(_4227_));
 sg13g2_buf_2 _4838_ (.A(\main.demo._q_speed[1] ),
    .X(_4229_));
 sg13g2_buf_1 _4839_ (.A(\main.demo._q_speed[0] ),
    .X(_4230_));
 sg13g2_buf_2 _4840_ (.A(\main.demo._q_speed[6] ),
    .X(_4231_));
 sg13g2_nor2_1 _4841_ (.A(_4230_),
    .B(_4231_),
    .Y(_4232_));
 sg13g2_xor2_1 _4842_ (.B(_4229_),
    .A(_4217_),
    .X(_4233_));
 sg13g2_inv_1 _4843_ (.Y(_4234_),
    .A(_4233_));
 sg13g2_nor2_1 _4844_ (.A(_4232_),
    .B(_4234_),
    .Y(_4235_));
 sg13g2_a21oi_1 _4845_ (.A1(_4217_),
    .A2(_4229_),
    .Y(_4236_),
    .B1(_4235_));
 sg13g2_nor2_1 _4846_ (.A(_4228_),
    .B(_4236_),
    .Y(_4237_));
 sg13g2_a21oi_1 _4847_ (.A1(_4226_),
    .A2(_4214_),
    .Y(_4238_),
    .B1(_4237_));
 sg13g2_nor2_1 _4848_ (.A(_4225_),
    .B(_4238_),
    .Y(_4239_));
 sg13g2_a21o_1 _4849_ (.A2(_4210_),
    .A1(_4223_),
    .B1(_4239_),
    .X(_4240_));
 sg13g2_inv_1 _4850_ (.Y(_4241_),
    .A(_4240_));
 sg13g2_nor2_1 _4851_ (.A(_4222_),
    .B(_4241_),
    .Y(_4242_));
 sg13g2_inv_1 _4852_ (.Y(_4243_),
    .A(_4242_));
 sg13g2_nand2_1 _4853_ (.Y(_4244_),
    .A(_4208_),
    .B(_4220_));
 sg13g2_nand2_1 _4854_ (.Y(_4245_),
    .A(_4243_),
    .B(_4244_));
 sg13g2_inv_1 _4855_ (.Y(_4246_),
    .A(_4245_));
 sg13g2_buf_8 _4856_ (.A(\main.demo._q_speed[5] ),
    .X(_4247_));
 sg13g2_nand2_1 _4857_ (.Y(_4248_),
    .A(\main.demo._q_speed[11] ),
    .B(_4247_));
 sg13g2_nor2_1 _4858_ (.A(\main.demo._q_speed[11] ),
    .B(_4247_),
    .Y(_4249_));
 sg13g2_a21oi_1 _4859_ (.A1(_4246_),
    .A2(_4248_),
    .Y(_4250_),
    .B1(_4249_));
 sg13g2_buf_1 _4860_ (.A(\main.demo._q_speed[12] ),
    .X(_4251_));
 sg13g2_nor2_1 _4861_ (.A(_4231_),
    .B(_4251_),
    .Y(_4252_));
 sg13g2_inv_1 _4862_ (.Y(_4253_),
    .A(_4252_));
 sg13g2_nand2_1 _4863_ (.Y(_4254_),
    .A(_4231_),
    .B(_4251_));
 sg13g2_inv_1 _4864_ (.Y(_4255_),
    .A(_4254_));
 sg13g2_a21oi_1 _4865_ (.A1(_4250_),
    .A2(_4253_),
    .Y(_4256_),
    .B1(_4255_));
 sg13g2_nand2_1 _4866_ (.Y(_4257_),
    .A(_4217_),
    .B(_4218_));
 sg13g2_o21ai_1 _4867_ (.B1(_4257_),
    .Y(_4258_),
    .A1(_4219_),
    .A2(_4256_));
 sg13g2_inv_1 _4868_ (.Y(_4259_),
    .A(_4258_));
 sg13g2_nand2_1 _4869_ (.Y(_4260_),
    .A(_4214_),
    .B(_4215_));
 sg13g2_o21ai_1 _4870_ (.B1(_4260_),
    .Y(_4261_),
    .A1(_4216_),
    .A2(_4259_));
 sg13g2_inv_1 _4871_ (.Y(_4262_),
    .A(_4261_));
 sg13g2_nor2_1 _4872_ (.A(_4213_),
    .B(_4262_),
    .Y(_4263_));
 sg13g2_a21o_1 _4873_ (.A2(_4211_),
    .A1(_4210_),
    .B1(_4263_),
    .X(_4264_));
 sg13g2_inv_1 _4874_ (.Y(_4265_),
    .A(_4264_));
 sg13g2_nor2_1 _4875_ (.A(_4209_),
    .B(_4265_),
    .Y(_4266_));
 sg13g2_inv_1 _4876_ (.Y(_4267_),
    .A(_4266_));
 sg13g2_nand2_1 _4877_ (.Y(_4268_),
    .A(_4265_),
    .B(_4209_));
 sg13g2_nor2b_1 _4878_ (.A(\main._w_demo_video_vs ),
    .B_N(\main.demo._q_prev_vs ),
    .Y(_4269_));
 sg13g2_buf_2 _4879_ (.A(_4269_),
    .X(_4270_));
 sg13g2_inv_2 _4880_ (.Y(_4271_),
    .A(_4270_));
 sg13g2_inv_1 _4881_ (.Y(_4272_),
    .A(\main.demo._q_go ));
 sg13g2_buf_1 _4882_ (.A(\main.demo._q_effect[0] ),
    .X(_4273_));
 sg13g2_buf_8 _4883_ (.A(\main.demo._q_effect[1] ),
    .X(_4274_));
 sg13g2_inv_1 _4884_ (.Y(_4275_),
    .A(_4274_));
 sg13g2_nor2_1 _4885_ (.A(_4273_),
    .B(_4275_),
    .Y(_4276_));
 sg13g2_inv_1 _4886_ (.Y(_4277_),
    .A(_4276_));
 sg13g2_nor2_2 _4887_ (.A(_4272_),
    .B(_4277_),
    .Y(_4278_));
 sg13g2_inv_2 _4888_ (.Y(_4279_),
    .A(_4278_));
 sg13g2_nor2_1 _4889_ (.A(_4271_),
    .B(_4279_),
    .Y(_4280_));
 sg13g2_buf_1 _4890_ (.A(_4280_),
    .X(_4281_));
 sg13g2_buf_1 _4891_ (.A(_4281_),
    .X(_4282_));
 sg13g2_nand3_1 _4892_ (.B(_4268_),
    .C(net31),
    .A(_4267_),
    .Y(_4283_));
 sg13g2_nor2_1 _4893_ (.A(_4270_),
    .B(_4279_),
    .Y(_4284_));
 sg13g2_buf_1 _4894_ (.A(_4284_),
    .X(_4285_));
 sg13g2_buf_1 _4895_ (.A(_4285_),
    .X(_4286_));
 sg13g2_buf_1 _4896_ (.A(_4279_),
    .X(_4287_));
 sg13g2_buf_2 _4897_ (.A(\main.demo._q_frame[7] ),
    .X(_4288_));
 sg13g2_nand2_1 _4898_ (.Y(_4289_),
    .A(_4288_),
    .B(_4140_));
 sg13g2_nand2_1 _4899_ (.Y(_4290_),
    .A(_4159_),
    .B(_4179_));
 sg13g2_nand2_1 _4900_ (.Y(_4291_),
    .A(_4171_),
    .B(_4164_));
 sg13g2_nor3_2 _4901_ (.A(_4290_),
    .B(_4291_),
    .C(_4271_),
    .Y(_4292_));
 sg13g2_nand2_2 _4902_ (.Y(_4293_),
    .A(_4292_),
    .B(_4146_));
 sg13g2_nor3_1 _4903_ (.A(_4149_),
    .B(_4289_),
    .C(_4293_),
    .Y(_4294_));
 sg13g2_inv_1 _4904_ (.Y(_4295_),
    .A(_4294_));
 sg13g2_buf_1 _4905_ (.A(\main.demo._q_frame[8] ),
    .X(_4296_));
 sg13g2_nor2b_1 _4906_ (.A(_4295_),
    .B_N(_4296_),
    .Y(_4297_));
 sg13g2_xor2_1 _4907_ (.B(_4297_),
    .A(\main.demo._q_frame[9] ),
    .X(_4298_));
 sg13g2_a22oi_1 _4908_ (.Y(_4299_),
    .B1(net35),
    .B2(_4298_),
    .A2(net30),
    .A1(_4208_));
 sg13g2_nand2_1 _4909_ (.Y(_0098_),
    .A(_4283_),
    .B(_4299_));
 sg13g2_inv_1 _4910_ (.Y(_4300_),
    .A(\main.demo._q_speed[11] ));
 sg13g2_nor2_1 _4911_ (.A(_0019_),
    .B(_4265_),
    .Y(_4301_));
 sg13g2_inv_1 _4912_ (.Y(_4302_),
    .A(_4301_));
 sg13g2_nor2_1 _4913_ (.A(_4300_),
    .B(_4302_),
    .Y(_4303_));
 sg13g2_inv_1 _4914_ (.Y(_4304_),
    .A(_4303_));
 sg13g2_nand2_1 _4915_ (.Y(_4305_),
    .A(_4302_),
    .B(_4300_));
 sg13g2_nand3_1 _4916_ (.B(net31),
    .C(_4305_),
    .A(_4304_),
    .Y(_4306_));
 sg13g2_nand2_1 _4917_ (.Y(_4307_),
    .A(_4297_),
    .B(\main.demo._q_frame[9] ));
 sg13g2_xnor2_1 _4918_ (.Y(_4308_),
    .A(\main.demo._q_frame[10] ),
    .B(_4307_));
 sg13g2_a22oi_1 _4919_ (.Y(_4309_),
    .B1(net35),
    .B2(_4308_),
    .A2(net30),
    .A1(\main.demo._q_speed[11] ));
 sg13g2_nand2_1 _4920_ (.Y(_0099_),
    .A(_4306_),
    .B(_4309_));
 sg13g2_inv_1 _4921_ (.Y(_4310_),
    .A(_4251_));
 sg13g2_nor2_1 _4922_ (.A(_4300_),
    .B(_4267_),
    .Y(_4311_));
 sg13g2_inv_1 _4923_ (.Y(_4312_),
    .A(_4311_));
 sg13g2_nor2_1 _4924_ (.A(_4310_),
    .B(_4312_),
    .Y(_4313_));
 sg13g2_inv_1 _4925_ (.Y(_4314_),
    .A(_4313_));
 sg13g2_nand2_1 _4926_ (.Y(_4315_),
    .A(_4312_),
    .B(_4310_));
 sg13g2_nand3_1 _4927_ (.B(net31),
    .C(_4315_),
    .A(_4314_),
    .Y(_4316_));
 sg13g2_nor2b_1 _4928_ (.A(_4307_),
    .B_N(\main.demo._q_frame[10] ),
    .Y(_4317_));
 sg13g2_xor2_1 _4929_ (.B(_4317_),
    .A(\main.demo._q_frame[11] ),
    .X(_4318_));
 sg13g2_a22oi_1 _4930_ (.Y(_4319_),
    .B1(net35),
    .B2(_4318_),
    .A2(net30),
    .A1(_4251_));
 sg13g2_nand2_1 _4931_ (.Y(_0100_),
    .A(_4316_),
    .B(_4319_));
 sg13g2_inv_1 _4932_ (.Y(_4320_),
    .A(_4218_));
 sg13g2_nor3_1 _4933_ (.A(_4310_),
    .B(_4320_),
    .C(_4304_),
    .Y(_4321_));
 sg13g2_o21ai_1 _4934_ (.B1(_4320_),
    .Y(_4322_),
    .A1(_4310_),
    .A2(_4304_));
 sg13g2_nand2_1 _4935_ (.Y(_4323_),
    .A(_4322_),
    .B(net31));
 sg13g2_nand2_1 _4936_ (.Y(_4324_),
    .A(_4317_),
    .B(\main.demo._q_frame[11] ));
 sg13g2_xnor2_1 _4937_ (.Y(_4325_),
    .A(\main.demo._q_frame[12] ),
    .B(_4324_));
 sg13g2_a22oi_1 _4938_ (.Y(_4326_),
    .B1(_4287_),
    .B2(_4325_),
    .A2(_4285_),
    .A1(_4218_));
 sg13g2_o21ai_1 _4939_ (.B1(_4326_),
    .Y(_0101_),
    .A1(_4321_),
    .A2(_4323_));
 sg13g2_a21oi_1 _4940_ (.A1(_4313_),
    .A2(_4218_),
    .Y(_4327_),
    .B1(_4215_));
 sg13g2_nand3_1 _4941_ (.B(_4218_),
    .C(_4215_),
    .A(_4313_),
    .Y(_4328_));
 sg13g2_nand3b_1 _4942_ (.B(net31),
    .C(_4328_),
    .Y(_4329_),
    .A_N(_4327_));
 sg13g2_nand2_1 _4943_ (.Y(_4330_),
    .A(net30),
    .B(_4215_));
 sg13g2_nor2b_1 _4944_ (.A(_4324_),
    .B_N(\main.demo._q_frame[12] ),
    .Y(_4331_));
 sg13g2_xnor2_1 _4945_ (.Y(_4332_),
    .A(\main.demo._q_frame[13] ),
    .B(_4331_));
 sg13g2_nand2b_1 _4946_ (.Y(_4333_),
    .B(_4279_),
    .A_N(_4332_));
 sg13g2_nand3_1 _4947_ (.B(_4330_),
    .C(_4333_),
    .A(_4329_),
    .Y(_0102_));
 sg13g2_a21oi_1 _4948_ (.A1(_4321_),
    .A2(_4215_),
    .Y(_4334_),
    .B1(_4211_));
 sg13g2_nand3_1 _4949_ (.B(_4215_),
    .C(_4211_),
    .A(_4321_),
    .Y(_4335_));
 sg13g2_nand2_1 _4950_ (.Y(_4336_),
    .A(_4335_),
    .B(_4282_));
 sg13g2_nand2_1 _4951_ (.Y(_4337_),
    .A(_4331_),
    .B(\main.demo._q_frame[13] ));
 sg13g2_xnor2_1 _4952_ (.Y(_4338_),
    .A(\main.demo._q_frame[14] ),
    .B(_4337_));
 sg13g2_a22oi_1 _4953_ (.Y(_4339_),
    .B1(_4287_),
    .B2(_4338_),
    .A2(_4285_),
    .A1(_4211_));
 sg13g2_o21ai_1 _4954_ (.B1(_4339_),
    .Y(_0103_),
    .A1(_4334_),
    .A2(_4336_));
 sg13g2_nand2_1 _4955_ (.Y(_4340_),
    .A(_4234_),
    .B(_4232_));
 sg13g2_nand3b_1 _4956_ (.B(net31),
    .C(_4340_),
    .Y(_4341_),
    .A_N(_4235_));
 sg13g2_nand2_1 _4957_ (.Y(_4342_),
    .A(net30),
    .B(_4229_));
 sg13g2_xnor2_1 _4958_ (.Y(_4343_),
    .A(_4164_),
    .B(_4270_));
 sg13g2_nand2b_1 _4959_ (.Y(_4344_),
    .B(_4279_),
    .A_N(_4343_));
 sg13g2_nand3_1 _4960_ (.B(_4342_),
    .C(_4344_),
    .A(_4341_),
    .Y(_0104_));
 sg13g2_inv_1 _4961_ (.Y(_4345_),
    .A(_4236_));
 sg13g2_o21ai_1 _4962_ (.B1(_4281_),
    .Y(_4346_),
    .A1(_4227_),
    .A2(_4345_));
 sg13g2_nor2_2 _4963_ (.A(_4291_),
    .B(_4271_),
    .Y(_4347_));
 sg13g2_a21oi_1 _4964_ (.A1(_4270_),
    .A2(_4164_),
    .Y(_4348_),
    .B1(_4171_));
 sg13g2_nor2_1 _4965_ (.A(_4347_),
    .B(_4348_),
    .Y(_4349_));
 sg13g2_a22oi_1 _4966_ (.Y(_4350_),
    .B1(net35),
    .B2(_4349_),
    .A2(_4226_),
    .A1(net30));
 sg13g2_o21ai_1 _4967_ (.B1(_4350_),
    .Y(_0105_),
    .A1(_4237_),
    .A2(_4346_));
 sg13g2_nand2_1 _4968_ (.Y(_4351_),
    .A(_4238_),
    .B(_4225_));
 sg13g2_nand2_1 _4969_ (.Y(_4352_),
    .A(_4351_),
    .B(_4281_));
 sg13g2_inv_1 _4970_ (.Y(_4353_),
    .A(_4179_));
 sg13g2_xnor2_1 _4971_ (.Y(_4354_),
    .A(_4353_),
    .B(_4347_));
 sg13g2_a22oi_1 _4972_ (.Y(_4355_),
    .B1(net35),
    .B2(_4354_),
    .A2(_4285_),
    .A1(_4223_));
 sg13g2_o21ai_1 _4973_ (.B1(_4355_),
    .Y(_0106_),
    .A1(_4239_),
    .A2(_4352_));
 sg13g2_nand2_1 _4974_ (.Y(_4356_),
    .A(_4241_),
    .B(_4222_));
 sg13g2_nand3_1 _4975_ (.B(net31),
    .C(_4356_),
    .A(_4243_),
    .Y(_4357_));
 sg13g2_a21oi_1 _4976_ (.A1(_4347_),
    .A2(_4179_),
    .Y(_4358_),
    .B1(_4159_));
 sg13g2_nor2_1 _4977_ (.A(_4292_),
    .B(_4358_),
    .Y(_4359_));
 sg13g2_a22oi_1 _4978_ (.Y(_4360_),
    .B1(net35),
    .B2(_4359_),
    .A2(net30),
    .A1(_4220_));
 sg13g2_nand2_1 _4979_ (.Y(_0107_),
    .A(_4357_),
    .B(_4360_));
 sg13g2_inv_1 _4980_ (.Y(_4361_),
    .A(_4146_));
 sg13g2_xnor2_1 _4981_ (.Y(_4362_),
    .A(_4361_),
    .B(_4292_));
 sg13g2_inv_1 _4982_ (.Y(_4363_),
    .A(_4362_));
 sg13g2_nand2b_1 _4983_ (.Y(_4364_),
    .B(_4248_),
    .A_N(_4249_));
 sg13g2_xnor2_1 _4984_ (.Y(_4365_),
    .A(_4364_),
    .B(_4245_));
 sg13g2_a22oi_1 _4985_ (.Y(_4366_),
    .B1(net31),
    .B2(_4365_),
    .A2(_4285_),
    .A1(_4247_));
 sg13g2_o21ai_1 _4986_ (.B1(_4366_),
    .Y(_0108_),
    .A1(_4278_),
    .A2(_4363_));
 sg13g2_nor2_1 _4987_ (.A(_4252_),
    .B(_4255_),
    .Y(_4367_));
 sg13g2_o21ai_1 _4988_ (.B1(_4281_),
    .Y(_4368_),
    .A1(_4367_),
    .A2(_4250_));
 sg13g2_a21oi_1 _4989_ (.A1(_4250_),
    .A2(_4367_),
    .Y(_4369_),
    .B1(_4368_));
 sg13g2_xnor2_1 _4990_ (.Y(_4370_),
    .A(_4148_),
    .B(_4293_));
 sg13g2_a22oi_1 _4991_ (.Y(_4371_),
    .B1(net35),
    .B2(_4370_),
    .A2(net30),
    .A1(_4231_));
 sg13g2_nand2b_1 _4992_ (.Y(_0109_),
    .B(_4371_),
    .A_N(_4369_));
 sg13g2_nor2b_1 _4993_ (.A(_4219_),
    .B_N(_4257_),
    .Y(_4372_));
 sg13g2_nor2b_1 _4994_ (.A(_4256_),
    .B_N(_4372_),
    .Y(_4373_));
 sg13g2_nand2b_1 _4995_ (.Y(_4374_),
    .B(_4256_),
    .A_N(_4372_));
 sg13g2_nand2_1 _4996_ (.Y(_4375_),
    .A(_4374_),
    .B(_4281_));
 sg13g2_nor2_1 _4997_ (.A(_4149_),
    .B(_4293_),
    .Y(_4376_));
 sg13g2_xnor2_1 _4998_ (.Y(_4377_),
    .A(_4147_),
    .B(_4376_));
 sg13g2_a22oi_1 _4999_ (.Y(_4378_),
    .B1(_4279_),
    .B2(_4377_),
    .A2(_4285_),
    .A1(_4217_));
 sg13g2_o21ai_1 _5000_ (.B1(_4378_),
    .Y(_0110_),
    .A1(_4373_),
    .A2(_4375_));
 sg13g2_nor2b_1 _5001_ (.A(_4216_),
    .B_N(_4260_),
    .Y(_4379_));
 sg13g2_nand2b_1 _5002_ (.Y(_4380_),
    .B(_4259_),
    .A_N(_4379_));
 sg13g2_nand2_1 _5003_ (.Y(_4381_),
    .A(_4258_),
    .B(_4379_));
 sg13g2_nand3_1 _5004_ (.B(_4381_),
    .C(_4282_),
    .A(_4380_),
    .Y(_4382_));
 sg13g2_nand2_1 _5005_ (.Y(_4383_),
    .A(_4286_),
    .B(_4214_));
 sg13g2_inv_1 _5006_ (.Y(_4384_),
    .A(_4288_));
 sg13g2_o21ai_1 _5007_ (.B1(_4384_),
    .Y(_4385_),
    .A1(_4151_),
    .A2(_4293_));
 sg13g2_nand3_1 _5008_ (.B(_4295_),
    .C(_4279_),
    .A(_4385_),
    .Y(_4386_));
 sg13g2_nand3_1 _5009_ (.B(_4383_),
    .C(_4386_),
    .A(_4382_),
    .Y(_0111_));
 sg13g2_nand2_1 _5010_ (.Y(_4387_),
    .A(_4262_),
    .B(_4213_));
 sg13g2_nand2_1 _5011_ (.Y(_4388_),
    .A(_4387_),
    .B(_4281_));
 sg13g2_xnor2_1 _5012_ (.Y(_4389_),
    .A(_4296_),
    .B(_4294_));
 sg13g2_nor2_1 _5013_ (.A(_4278_),
    .B(_4389_),
    .Y(_4390_));
 sg13g2_a21oi_1 _5014_ (.A1(_4210_),
    .A2(_4286_),
    .Y(_4391_),
    .B1(_4390_));
 sg13g2_o21ai_1 _5015_ (.B1(_4391_),
    .Y(_0112_),
    .A1(_4263_),
    .A2(_4388_));
 sg13g2_inv_1 _5016_ (.Y(_4392_),
    .A(\main.demo.zic._q_rythm_count[5] ));
 sg13g2_inv_1 _5017_ (.Y(_4393_),
    .A(\main.demo.zic._q_rythm_count[6] ));
 sg13g2_nand2_1 _5018_ (.Y(_4394_),
    .A(_4392_),
    .B(_4393_));
 sg13g2_inv_1 _5019_ (.Y(_4395_),
    .A(\main.demo.zic._q_rythm_count[1] ));
 sg13g2_inv_1 _5020_ (.Y(_4396_),
    .A(\main.demo.zic._q_rythm_count[0] ));
 sg13g2_inv_1 _5021_ (.Y(_4397_),
    .A(\main.demo.zic._q_rythm_count[3] ));
 sg13g2_inv_1 _5022_ (.Y(_4398_),
    .A(\main.demo.zic._q_rythm_count[2] ));
 sg13g2_nand4_1 _5023_ (.B(_4396_),
    .C(_4397_),
    .A(_4395_),
    .Y(_4399_),
    .D(_4398_));
 sg13g2_nor4_1 _5024_ (.A(\main.demo.zic._q_rythm_count[4] ),
    .B(\main.demo.zic._q_rythm_count[7] ),
    .C(_4394_),
    .D(_4399_),
    .Y(_4400_));
 sg13g2_nor2_1 _5025_ (.A(\main.demo.zic._q_clock_count[1] ),
    .B(\main.demo.zic._q_clock_count[0] ),
    .Y(_4401_));
 sg13g2_buf_1 _5026_ (.A(\main.demo.zic._q_clock_count[3] ),
    .X(_4402_));
 sg13g2_buf_1 _5027_ (.A(\main.demo.zic._q_clock_count[2] ),
    .X(_4403_));
 sg13g2_nor2_1 _5028_ (.A(_4402_),
    .B(_4403_),
    .Y(_4404_));
 sg13g2_inv_1 _5029_ (.Y(_4405_),
    .A(\main.demo.zic._q_clock_count[5] ));
 sg13g2_buf_1 _5030_ (.A(\main.demo.zic._q_clock_count[4] ),
    .X(_4406_));
 sg13g2_inv_1 _5031_ (.Y(_4407_),
    .A(_4406_));
 sg13g2_nand4_1 _5032_ (.B(_4404_),
    .C(_4405_),
    .A(_4401_),
    .Y(_4408_),
    .D(_4407_));
 sg13g2_nor3_1 _5033_ (.A(\main.demo.zic._q_clock_count[7] ),
    .B(\main.demo.zic._q_clock_count[6] ),
    .C(\main.demo.zic._q_clock_count[8] ),
    .Y(_4409_));
 sg13g2_nor2b_1 _5034_ (.A(_4408_),
    .B_N(_4409_),
    .Y(_4410_));
 sg13g2_buf_1 _5035_ (.A(_4410_),
    .X(_4411_));
 sg13g2_nand2_2 _5036_ (.Y(_4412_),
    .A(_4400_),
    .B(net45));
 sg13g2_inv_1 _5037_ (.Y(_4413_),
    .A(_4412_));
 sg13g2_buf_1 _5038_ (.A(\main.demo.zic._q_drum_inc[3] ),
    .X(_4414_));
 sg13g2_buf_1 _5039_ (.A(\main.demo.zic._q_drum_inc[2] ),
    .X(_4415_));
 sg13g2_buf_1 _5040_ (.A(\main.demo.zic._q_drum_inc[1] ),
    .X(_4416_));
 sg13g2_nor2_1 _5041_ (.A(\main.demo.zic._q_drum_inc[0] ),
    .B(_4416_),
    .Y(_4417_));
 sg13g2_inv_1 _5042_ (.Y(_4418_),
    .A(_4417_));
 sg13g2_nor3_1 _5043_ (.A(_4414_),
    .B(_4415_),
    .C(_4418_),
    .Y(_4419_));
 sg13g2_nor2_1 _5044_ (.A(\main.demo.zic._q_rythm_count[9] ),
    .B(\main.demo.zic._q_rythm_count[8] ),
    .Y(_4420_));
 sg13g2_inv_1 _5045_ (.Y(_4421_),
    .A(\main.demo.zic._q_rythm_count[11] ));
 sg13g2_nand4_1 _5046_ (.B(_4421_),
    .C(\main.demo.zic._q_rythm_count[10] ),
    .A(_4420_),
    .Y(_4422_),
    .D(\main.demo.zic._q_rythm_count[12] ));
 sg13g2_buf_1 _5047_ (.A(_4422_),
    .X(_4423_));
 sg13g2_inv_1 _5048_ (.Y(_4424_),
    .A(net62));
 sg13g2_nor2_1 _5049_ (.A(_4419_),
    .B(net52),
    .Y(_4425_));
 sg13g2_inv_1 _5050_ (.Y(_4426_),
    .A(\main.demo.zic._q_drum_inc[0] ));
 sg13g2_nor2_1 _5051_ (.A(_4426_),
    .B(_4424_),
    .Y(_4427_));
 sg13g2_a21oi_1 _5052_ (.A1(_4413_),
    .A2(_4425_),
    .Y(_4428_),
    .B1(_4427_));
 sg13g2_nor2_1 _5053_ (.A(_4426_),
    .B(_4412_),
    .Y(_4429_));
 sg13g2_buf_1 _5054_ (.A(\main.demo.zic._q_idx[4] ),
    .X(_4430_));
 sg13g2_inv_2 _5055_ (.Y(_4431_),
    .A(_4430_));
 sg13g2_buf_2 _5056_ (.A(\main.demo.zic._q_idx[1] ),
    .X(_4432_));
 sg13g2_buf_1 _5057_ (.A(\main.demo.zic._q_idx[0] ),
    .X(_4433_));
 sg13g2_nand2_1 _5058_ (.Y(_4434_),
    .A(_4432_),
    .B(_4433_));
 sg13g2_buf_1 _5059_ (.A(_4434_),
    .X(_4435_));
 sg13g2_buf_2 _5060_ (.A(\main.demo.zic._q_idx[3] ),
    .X(_4436_));
 sg13g2_buf_1 _5061_ (.A(\main.demo.zic._q_idx[2] ),
    .X(_4437_));
 sg13g2_nand2_2 _5062_ (.Y(_4438_),
    .A(_4436_),
    .B(_4437_));
 sg13g2_nor2_2 _5063_ (.A(_4435_),
    .B(_4438_),
    .Y(_4439_));
 sg13g2_nand2_1 _5064_ (.Y(_4440_),
    .A(net52),
    .B(_4439_));
 sg13g2_xnor2_1 _5065_ (.Y(_4441_),
    .A(_4431_),
    .B(_4440_));
 sg13g2_inv_1 _5066_ (.Y(_4442_),
    .A(_4441_));
 sg13g2_buf_2 _5067_ (.A(\main.demo.zic._q_idx[5] ),
    .X(_4443_));
 sg13g2_inv_1 _5068_ (.Y(_0232_),
    .A(_4443_));
 sg13g2_inv_1 _5069_ (.Y(_0233_),
    .A(_4439_));
 sg13g2_nor2_1 _5070_ (.A(_4431_),
    .B(_0233_),
    .Y(_0234_));
 sg13g2_nand2_1 _5071_ (.Y(_0235_),
    .A(net52),
    .B(_0234_));
 sg13g2_xnor2_1 _5072_ (.Y(_0236_),
    .A(_0232_),
    .B(_0235_));
 sg13g2_inv_1 _5073_ (.Y(_0237_),
    .A(_0236_));
 sg13g2_inv_1 _5074_ (.Y(_0238_),
    .A(_4437_));
 sg13g2_inv_1 _5075_ (.Y(_0239_),
    .A(_4435_));
 sg13g2_nand2_1 _5076_ (.Y(_0240_),
    .A(net52),
    .B(_0239_));
 sg13g2_xnor2_1 _5077_ (.Y(_0241_),
    .A(_0238_),
    .B(_0240_));
 sg13g2_inv_1 _5078_ (.Y(_0242_),
    .A(_4436_));
 sg13g2_nand3b_1 _5079_ (.B(_4437_),
    .C(_4432_),
    .Y(_0243_),
    .A_N(_0045_));
 sg13g2_xnor2_1 _5080_ (.Y(_0244_),
    .A(_0242_),
    .B(_0243_));
 sg13g2_inv_1 _5081_ (.Y(_0245_),
    .A(_0244_));
 sg13g2_inv_1 _5082_ (.Y(_0246_),
    .A(\main.demo.zic._q_idx[6] ));
 sg13g2_nor3_1 _5083_ (.A(_4443_),
    .B(_4431_),
    .C(_0246_),
    .Y(_0247_));
 sg13g2_buf_2 _5084_ (.A(_0247_),
    .X(_0248_));
 sg13g2_a21oi_2 _5085_ (.B1(net62),
    .Y(_0249_),
    .A2(_0248_),
    .A1(_4439_));
 sg13g2_a22oi_1 _5086_ (.Y(_0250_),
    .B1(_0245_),
    .B2(_0249_),
    .A2(net62),
    .A1(_4436_));
 sg13g2_buf_1 _5087_ (.A(_0250_),
    .X(_0251_));
 sg13g2_nor2_1 _5088_ (.A(_0241_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_nand2_1 _5089_ (.Y(_0253_),
    .A(_4443_),
    .B(_0044_));
 sg13g2_nor2_2 _5090_ (.A(_4431_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_inv_1 _5091_ (.Y(_0255_),
    .A(_0254_));
 sg13g2_a21o_1 _5092_ (.A2(_4443_),
    .A1(_0234_),
    .B1(_0044_),
    .X(_0256_));
 sg13g2_o21ai_1 _5093_ (.B1(_0256_),
    .Y(_0257_),
    .A1(_0233_),
    .A2(_0255_));
 sg13g2_a22oi_1 _5094_ (.Y(_0258_),
    .B1(_0249_),
    .B2(_0257_),
    .A2(net62),
    .A1(\main.demo.zic._q_idx[6] ));
 sg13g2_buf_1 _5095_ (.A(_0258_),
    .X(_0259_));
 sg13g2_inv_1 _5096_ (.Y(_0260_),
    .A(_0259_));
 sg13g2_nor4_1 _5097_ (.A(_4442_),
    .B(_0237_),
    .C(_0252_),
    .D(_0260_),
    .Y(_0261_));
 sg13g2_nor2_1 _5098_ (.A(_4432_),
    .B(_4433_),
    .Y(_0262_));
 sg13g2_nor2_1 _5099_ (.A(_0262_),
    .B(_0239_),
    .Y(_0263_));
 sg13g2_nor2b_1 _5100_ (.A(net62),
    .B_N(_0263_),
    .Y(_0264_));
 sg13g2_a21oi_2 _5101_ (.B1(_0264_),
    .Y(_0265_),
    .A2(net62),
    .A1(_4432_));
 sg13g2_inv_1 _5102_ (.Y(_0266_),
    .A(_0265_));
 sg13g2_nand2_1 _5103_ (.Y(_0267_),
    .A(_0252_),
    .B(_0266_));
 sg13g2_nor3_1 _5104_ (.A(_0237_),
    .B(_0267_),
    .C(_0260_),
    .Y(_0268_));
 sg13g2_nand3_1 _5105_ (.B(_4441_),
    .C(_0237_),
    .A(_0259_),
    .Y(_0269_));
 sg13g2_nor2_1 _5106_ (.A(_4442_),
    .B(_0237_),
    .Y(_0270_));
 sg13g2_nand2_1 _5107_ (.Y(_0271_),
    .A(_0260_),
    .B(_0270_));
 sg13g2_a21oi_1 _5108_ (.A1(_0269_),
    .A2(_0271_),
    .Y(_0272_),
    .B1(_0265_));
 sg13g2_nor3_1 _5109_ (.A(_0261_),
    .B(_0268_),
    .C(_0272_),
    .Y(_0273_));
 sg13g2_xnor2_1 _5110_ (.Y(_0274_),
    .A(_0241_),
    .B(_0251_));
 sg13g2_nand2_1 _5111_ (.Y(_0275_),
    .A(_4442_),
    .B(_0232_));
 sg13g2_nor2_1 _5112_ (.A(_0275_),
    .B(_0259_),
    .Y(_0276_));
 sg13g2_nand2b_1 _5113_ (.Y(_0277_),
    .B(_0276_),
    .A_N(_0274_));
 sg13g2_nand2_1 _5114_ (.Y(_0278_),
    .A(_0276_),
    .B(_0274_));
 sg13g2_nand3_1 _5115_ (.B(_4443_),
    .C(_4442_),
    .A(_0259_),
    .Y(_0279_));
 sg13g2_nand3_1 _5116_ (.B(_0278_),
    .C(_0279_),
    .A(_0277_),
    .Y(_0280_));
 sg13g2_nand2_1 _5117_ (.Y(_0281_),
    .A(_0280_),
    .B(_0266_));
 sg13g2_a21oi_1 _5118_ (.A1(_0251_),
    .A2(_0266_),
    .Y(_0282_),
    .B1(_0241_));
 sg13g2_or3_1 _5119_ (.A(_0275_),
    .B(_0282_),
    .C(_0260_),
    .X(_0283_));
 sg13g2_nand4_1 _5120_ (.B(net52),
    .C(_0281_),
    .A(_0273_),
    .Y(_0284_),
    .D(_0283_));
 sg13g2_buf_1 _5121_ (.A(_0284_),
    .X(_0285_));
 sg13g2_o21ai_1 _5122_ (.B1(_0285_),
    .Y(_0177_),
    .A1(_4428_),
    .A2(_4429_));
 sg13g2_inv_1 _5123_ (.Y(_0286_),
    .A(_4416_));
 sg13g2_nor2_1 _5124_ (.A(net52),
    .B(_4413_),
    .Y(_0287_));
 sg13g2_buf_1 _5125_ (.A(_0287_),
    .X(_0288_));
 sg13g2_inv_1 _5126_ (.Y(_0289_),
    .A(_4414_));
 sg13g2_inv_1 _5127_ (.Y(_0290_),
    .A(_4415_));
 sg13g2_a21oi_1 _5128_ (.A1(_0289_),
    .A2(_0290_),
    .Y(_0291_),
    .B1(_4418_));
 sg13g2_a221oi_1 _5129_ (.B2(_0291_),
    .C1(net29),
    .B1(net62),
    .A1(_4416_),
    .Y(_0292_),
    .A2(_4427_));
 sg13g2_a22oi_1 _5130_ (.Y(_0178_),
    .B1(_0292_),
    .B2(_0285_),
    .A2(net29),
    .A1(_0286_));
 sg13g2_nand2_1 _5131_ (.Y(_0293_),
    .A(net29),
    .B(_4415_));
 sg13g2_xnor2_1 _5132_ (.Y(_0294_),
    .A(_0290_),
    .B(_4417_));
 sg13g2_nand3_1 _5133_ (.B(_4425_),
    .C(_0294_),
    .A(_4413_),
    .Y(_0295_));
 sg13g2_nand3_1 _5134_ (.B(_0293_),
    .C(_0295_),
    .A(_0285_),
    .Y(_0179_));
 sg13g2_a21oi_1 _5135_ (.A1(_4417_),
    .A2(_0290_),
    .Y(_0296_),
    .B1(_0289_));
 sg13g2_o21ai_1 _5136_ (.B1(_4423_),
    .Y(_0297_),
    .A1(_0296_),
    .A2(_4412_));
 sg13g2_a22oi_1 _5137_ (.Y(_0180_),
    .B1(_0297_),
    .B2(_0285_),
    .A2(net29),
    .A1(_0289_));
 sg13g2_inv_2 _5138_ (.Y(_0298_),
    .A(_4231_));
 sg13g2_a21oi_1 _5139_ (.A1(_4270_),
    .A2(_0298_),
    .Y(_0299_),
    .B1(_4230_));
 sg13g2_inv_2 _5140_ (.Y(_0300_),
    .A(_4230_));
 sg13g2_nor3_1 _5141_ (.A(_0300_),
    .B(_4231_),
    .C(_4271_),
    .Y(_0301_));
 sg13g2_nor3_1 _5142_ (.A(net35),
    .B(_0299_),
    .C(_0301_),
    .Y(_0097_));
 sg13g2_nand2_1 _5143_ (.Y(_0302_),
    .A(_4271_),
    .B(\main.demo._q_th[0] ));
 sg13g2_nand2_1 _5144_ (.Y(_0303_),
    .A(_4270_),
    .B(_0067_));
 sg13g2_nor3_1 _5145_ (.A(_4149_),
    .B(_4361_),
    .C(_4289_),
    .Y(_0304_));
 sg13g2_nor2_1 _5146_ (.A(_4290_),
    .B(_4291_),
    .Y(_0305_));
 sg13g2_nand3_1 _5147_ (.B(_4296_),
    .C(_0305_),
    .A(_0304_),
    .Y(_0306_));
 sg13g2_nor2b_1 _5148_ (.A(_4272_),
    .B_N(_0306_),
    .Y(_0307_));
 sg13g2_inv_1 _5149_ (.Y(_0308_),
    .A(_0307_));
 sg13g2_a21oi_1 _5150_ (.A1(_0302_),
    .A2(_0303_),
    .Y(_0113_),
    .B1(net41));
 sg13g2_a21oi_1 _5151_ (.A1(_4270_),
    .A2(\main.demo._q_th[0] ),
    .Y(_0309_),
    .B1(\main.demo._q_th[1] ));
 sg13g2_nand3_1 _5152_ (.B(\main.demo._q_th[1] ),
    .C(\main.demo._q_th[0] ),
    .A(_4270_),
    .Y(_0310_));
 sg13g2_inv_1 _5153_ (.Y(_0311_),
    .A(_0310_));
 sg13g2_nor3_1 _5154_ (.A(_0309_),
    .B(_0311_),
    .C(net41),
    .Y(_0114_));
 sg13g2_buf_1 _5155_ (.A(\main.demo._q_th[2] ),
    .X(_0312_));
 sg13g2_nor2_1 _5156_ (.A(_0312_),
    .B(_0311_),
    .Y(_0313_));
 sg13g2_inv_1 _5157_ (.Y(_0314_),
    .A(_0312_));
 sg13g2_nor2_1 _5158_ (.A(_0314_),
    .B(_0310_),
    .Y(_0315_));
 sg13g2_nor3_1 _5159_ (.A(_0313_),
    .B(_0315_),
    .C(net41),
    .Y(_0115_));
 sg13g2_buf_1 _5160_ (.A(\main.demo._q_th[3] ),
    .X(_0316_));
 sg13g2_nor2_1 _5161_ (.A(_0316_),
    .B(_0315_),
    .Y(_0317_));
 sg13g2_nand2_1 _5162_ (.Y(_0318_),
    .A(_0315_),
    .B(_0316_));
 sg13g2_inv_1 _5163_ (.Y(_0319_),
    .A(_0318_));
 sg13g2_nor3_1 _5164_ (.A(_0317_),
    .B(_0319_),
    .C(_0308_),
    .Y(_0116_));
 sg13g2_inv_1 _5165_ (.Y(_0320_),
    .A(\main.demo._q_th[4] ));
 sg13g2_nor2_1 _5166_ (.A(_0320_),
    .B(_0318_),
    .Y(_0321_));
 sg13g2_nor2_1 _5167_ (.A(\main.demo._q_th[4] ),
    .B(_0319_),
    .Y(_0322_));
 sg13g2_nor3_1 _5168_ (.A(_0321_),
    .B(net41),
    .C(_0322_),
    .Y(_0117_));
 sg13g2_inv_1 _5169_ (.Y(_0323_),
    .A(\main.demo._q_th[5] ));
 sg13g2_nor3_1 _5170_ (.A(_0323_),
    .B(_0320_),
    .C(_0318_),
    .Y(_0324_));
 sg13g2_nor2_1 _5171_ (.A(\main.demo._q_th[5] ),
    .B(_0321_),
    .Y(_0325_));
 sg13g2_nor3_1 _5172_ (.A(net41),
    .B(_0324_),
    .C(_0325_),
    .Y(_0118_));
 sg13g2_buf_2 _5173_ (.A(\main.demo._q_th[6] ),
    .X(_0326_));
 sg13g2_nor2_1 _5174_ (.A(_0326_),
    .B(_0324_),
    .Y(_0327_));
 sg13g2_nand2_1 _5175_ (.Y(_0328_),
    .A(_0324_),
    .B(_0326_));
 sg13g2_inv_1 _5176_ (.Y(_0329_),
    .A(_0328_));
 sg13g2_nor3_1 _5177_ (.A(net41),
    .B(_0327_),
    .C(_0329_),
    .Y(_0119_));
 sg13g2_buf_1 _5178_ (.A(\main.demo._q_th[7] ),
    .X(_0330_));
 sg13g2_inv_2 _5179_ (.Y(_0331_),
    .A(_0330_));
 sg13g2_nor2_1 _5180_ (.A(_0331_),
    .B(_0328_),
    .Y(_0332_));
 sg13g2_nor2_1 _5181_ (.A(_0330_),
    .B(_0329_),
    .Y(_0333_));
 sg13g2_nor3_1 _5182_ (.A(net41),
    .B(_0332_),
    .C(_0333_),
    .Y(_0120_));
 sg13g2_nor2_1 _5183_ (.A(\main.demo._q_th[8] ),
    .B(_0332_),
    .Y(_0334_));
 sg13g2_and3_1 _5184_ (.X(_0335_),
    .A(_0329_),
    .B(_0330_),
    .C(\main.demo._q_th[8] ));
 sg13g2_nor3_1 _5185_ (.A(net41),
    .B(_0334_),
    .C(_0335_),
    .Y(_0121_));
 sg13g2_inv_1 _5186_ (.Y(_0336_),
    .A(\main.demo.vga._q_xcount[2] ));
 sg13g2_nand2_1 _5187_ (.Y(_0337_),
    .A(\main.demo.vga._q_xcount[1] ),
    .B(\main.demo.vga._q_xcount[0] ));
 sg13g2_nor2_1 _5188_ (.A(_0336_),
    .B(_0337_),
    .Y(_0338_));
 sg13g2_nand2_1 _5189_ (.Y(_0339_),
    .A(_0338_),
    .B(\main.demo.vga._q_xcount[3] ));
 sg13g2_inv_1 _5190_ (.Y(_0340_),
    .A(_0339_));
 sg13g2_buf_1 _5191_ (.A(\main.demo.vga._q_xcount[7] ),
    .X(_0341_));
 sg13g2_inv_1 _5192_ (.Y(_0342_),
    .A(_0341_));
 sg13g2_inv_1 _5193_ (.Y(_0343_),
    .A(\main.demo.vga._q_xcount[6] ));
 sg13g2_buf_1 _5194_ (.A(\main.demo.vga._q_xcount[5] ),
    .X(_0344_));
 sg13g2_nor2_1 _5195_ (.A(_0344_),
    .B(\main.demo.vga._q_xcount[4] ),
    .Y(_0345_));
 sg13g2_inv_1 _5196_ (.Y(_0346_),
    .A(_0345_));
 sg13g2_nor3_1 _5197_ (.A(_0342_),
    .B(_0343_),
    .C(_0346_),
    .Y(_0347_));
 sg13g2_inv_1 _5198_ (.Y(_0348_),
    .A(\main.demo.vga._q_xcount[9] ));
 sg13g2_inv_2 _5199_ (.Y(_0349_),
    .A(\main.demo.vga._q_xcount[8] ));
 sg13g2_inv_1 _5200_ (.Y(_0350_),
    .A(\main.demo.vga._q_xcount[10] ));
 sg13g2_nor3_1 _5201_ (.A(_0348_),
    .B(_0349_),
    .C(_0350_),
    .Y(_0351_));
 sg13g2_nand3_1 _5202_ (.B(_0347_),
    .C(_0351_),
    .A(_0340_),
    .Y(_0352_));
 sg13g2_inv_1 _5203_ (.Y(_0353_),
    .A(\main._w_demo_video_hs ));
 sg13g2_nand2_1 _5204_ (.Y(_0354_),
    .A(_0344_),
    .B(\main.demo.vga._q_xcount[4] ));
 sg13g2_nor2_1 _5205_ (.A(\main.demo.vga._q_xcount[1] ),
    .B(\main.demo.vga._q_xcount[0] ),
    .Y(_0355_));
 sg13g2_inv_1 _5206_ (.Y(_0356_),
    .A(\main.demo.vga._q_xcount[3] ));
 sg13g2_nand3_1 _5207_ (.B(_0356_),
    .C(_0336_),
    .A(_0355_),
    .Y(_0357_));
 sg13g2_nor4_1 _5208_ (.A(_0341_),
    .B(_0343_),
    .C(_0354_),
    .D(_0357_),
    .Y(_0358_));
 sg13g2_a221oi_1 _5209_ (.B2(_0351_),
    .C1(_0012_),
    .B1(_0358_),
    .A1(_0352_),
    .Y(_0124_),
    .A2(_0353_));
 sg13g2_inv_1 _5210_ (.Y(_0359_),
    .A(\main.demo.vga._q_ycount[1] ));
 sg13g2_buf_1 _5211_ (.A(\main.demo.vga._q_ycount[0] ),
    .X(_0360_));
 sg13g2_nand2_1 _5212_ (.Y(_0361_),
    .A(_0359_),
    .B(_0360_));
 sg13g2_buf_1 _5213_ (.A(\main.demo.vga._q_ycount[5] ),
    .X(_0362_));
 sg13g2_inv_1 _5214_ (.Y(_0363_),
    .A(\main.demo.vga._q_ycount[8] ));
 sg13g2_inv_1 _5215_ (.Y(_0364_),
    .A(\main.demo.vga._d_vblank ));
 sg13g2_nor3_1 _5216_ (.A(_0362_),
    .B(_0363_),
    .C(_0364_),
    .Y(_0365_));
 sg13g2_buf_1 _5217_ (.A(\main.demo.vga._q_ycount[2] ),
    .X(_0366_));
 sg13g2_nand2_1 _5218_ (.Y(_0367_),
    .A(\main.demo.vga._q_ycount[3] ),
    .B(_0366_));
 sg13g2_inv_1 _5219_ (.Y(_0368_),
    .A(_0367_));
 sg13g2_buf_1 _5220_ (.A(\main.demo.vga._q_ycount[4] ),
    .X(_0369_));
 sg13g2_inv_1 _5221_ (.Y(_0370_),
    .A(_0369_));
 sg13g2_nand2_1 _5222_ (.Y(_0371_),
    .A(\main.demo.vga._q_ycount[7] ),
    .B(\main.demo.vga._q_ycount[6] ));
 sg13g2_nor2_1 _5223_ (.A(_0370_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_nand3_1 _5224_ (.B(_0368_),
    .C(_0372_),
    .A(_0365_),
    .Y(_0373_));
 sg13g2_inv_1 _5225_ (.Y(_0374_),
    .A(_0012_));
 sg13g2_o21ai_1 _5226_ (.B1(_0374_),
    .Y(_0375_),
    .A1(_0361_),
    .A2(_0373_));
 sg13g2_nor3_1 _5227_ (.A(_0359_),
    .B(_0360_),
    .C(_0373_),
    .Y(_0376_));
 sg13g2_nor2_1 _5228_ (.A(\main._w_demo_video_vs ),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_nor2_1 _5229_ (.A(_0375_),
    .B(_0377_),
    .Y(_0125_));
 sg13g2_inv_1 _5230_ (.Y(_0378_),
    .A(_0360_));
 sg13g2_nor4_2 _5231_ (.A(\main.demo.vga._q_ycount[1] ),
    .B(_0360_),
    .C(\main.demo.vga._q_ycount[3] ),
    .Y(_0379_),
    .D(_0366_));
 sg13g2_nor2_1 _5232_ (.A(_0369_),
    .B(\main.demo.vga._d_vblank ),
    .Y(_0380_));
 sg13g2_inv_1 _5233_ (.Y(_0381_),
    .A(_0362_));
 sg13g2_nor3_1 _5234_ (.A(_0381_),
    .B(_0363_),
    .C(_0371_),
    .Y(_0382_));
 sg13g2_nand3_1 _5235_ (.B(_0380_),
    .C(_0382_),
    .A(_0379_),
    .Y(_0383_));
 sg13g2_nor4_1 _5236_ (.A(_0362_),
    .B(\main.demo.vga._q_ycount[7] ),
    .C(\main.demo.vga._q_ycount[6] ),
    .D(\main.demo.vga._q_ycount[8] ),
    .Y(_0384_));
 sg13g2_and3_1 _5237_ (.X(_0385_),
    .A(_0379_),
    .B(_0384_),
    .C(_0380_));
 sg13g2_a21oi_1 _5238_ (.A1(\main.demo.vga._q_active_v ),
    .A2(_0383_),
    .Y(_0386_),
    .B1(_0385_));
 sg13g2_buf_1 _5239_ (.A(_0386_),
    .X(_0387_));
 sg13g2_nor2_1 _5240_ (.A(_0378_),
    .B(_0387_),
    .Y(_0137_));
 sg13g2_nor2_1 _5241_ (.A(_0359_),
    .B(_0387_),
    .Y(_0138_));
 sg13g2_nor2b_1 _5242_ (.A(net40),
    .B_N(_0366_),
    .Y(_0139_));
 sg13g2_nor2b_1 _5243_ (.A(_0386_),
    .B_N(\main.demo.vga._q_ycount[3] ),
    .Y(_0140_));
 sg13g2_nor2_1 _5244_ (.A(_0370_),
    .B(net40),
    .Y(_0141_));
 sg13g2_nor2_1 _5245_ (.A(_0381_),
    .B(net40),
    .Y(_0142_));
 sg13g2_inv_1 _5246_ (.Y(_0388_),
    .A(\main.demo.vga._q_ycount[6] ));
 sg13g2_nor2_1 _5247_ (.A(_0388_),
    .B(net40),
    .Y(_0143_));
 sg13g2_inv_1 _5248_ (.Y(_0389_),
    .A(\main.demo.vga._q_ycount[7] ));
 sg13g2_nor2_1 _5249_ (.A(_0389_),
    .B(net40),
    .Y(_0144_));
 sg13g2_nor2_1 _5250_ (.A(_0363_),
    .B(net40),
    .Y(_0145_));
 sg13g2_nor2_1 _5251_ (.A(_0364_),
    .B(net40),
    .Y(_0146_));
 sg13g2_inv_1 _5252_ (.Y(_0390_),
    .A(_0337_));
 sg13g2_inv_1 _5253_ (.Y(_0391_),
    .A(_0357_));
 sg13g2_nor3_1 _5254_ (.A(\main.demo.vga._q_xcount[8] ),
    .B(\main.demo.vga._q_xcount[10] ),
    .C(_0348_),
    .Y(_0392_));
 sg13g2_nor2_1 _5255_ (.A(\main.demo.vga._q_xcount[6] ),
    .B(_0342_),
    .Y(_0393_));
 sg13g2_nand4_1 _5256_ (.B(_0345_),
    .C(_0392_),
    .A(_0391_),
    .Y(_0394_),
    .D(_0393_));
 sg13g2_buf_1 _5257_ (.A(_0394_),
    .X(_0395_));
 sg13g2_nand2_2 _5258_ (.Y(_0396_),
    .A(_0395_),
    .B(_0374_));
 sg13g2_nor3_1 _5259_ (.A(_0390_),
    .B(_0355_),
    .C(_0396_),
    .Y(_0149_));
 sg13g2_nor2_1 _5260_ (.A(\main.demo.vga._q_xcount[2] ),
    .B(_0390_),
    .Y(_0397_));
 sg13g2_nor3_1 _5261_ (.A(_0338_),
    .B(_0397_),
    .C(_0396_),
    .Y(_0150_));
 sg13g2_nor2_1 _5262_ (.A(\main.demo.vga._q_xcount[3] ),
    .B(_0338_),
    .Y(_0398_));
 sg13g2_nor3_1 _5263_ (.A(_0340_),
    .B(_0398_),
    .C(_0396_),
    .Y(_0151_));
 sg13g2_nor2_1 _5264_ (.A(\main.demo.vga._q_xcount[4] ),
    .B(_0340_),
    .Y(_0399_));
 sg13g2_inv_1 _5265_ (.Y(_0400_),
    .A(\main.demo.vga._q_xcount[4] ));
 sg13g2_nor2_1 _5266_ (.A(_0400_),
    .B(_0339_),
    .Y(_0401_));
 sg13g2_nor3_1 _5267_ (.A(_0399_),
    .B(_0401_),
    .C(_0396_),
    .Y(_0152_));
 sg13g2_nor3_1 _5268_ (.A(_0343_),
    .B(_0354_),
    .C(_0339_),
    .Y(_0402_));
 sg13g2_nor2_1 _5269_ (.A(_0341_),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_nand2_1 _5270_ (.Y(_0404_),
    .A(_0402_),
    .B(_0341_));
 sg13g2_inv_1 _5271_ (.Y(_0405_),
    .A(_0404_));
 sg13g2_nor3_1 _5272_ (.A(_0403_),
    .B(_0405_),
    .C(_0396_),
    .Y(_0155_));
 sg13g2_inv_2 _5273_ (.Y(_0406_),
    .A(_4411_));
 sg13g2_nand2_1 _5274_ (.Y(_0407_),
    .A(_0406_),
    .B(\main.demo.zic._q_rythm_count[0] ));
 sg13g2_buf_1 _5275_ (.A(net45),
    .X(_0408_));
 sg13g2_nand2_1 _5276_ (.Y(_0409_),
    .A(net39),
    .B(_0068_));
 sg13g2_nor2_1 _5277_ (.A(\main.demo._q_go ),
    .B(_4298_),
    .Y(_0410_));
 sg13g2_buf_2 _5278_ (.A(_0410_),
    .X(_0411_));
 sg13g2_nor2_1 _5279_ (.A(_0012_),
    .B(_0411_),
    .Y(_0412_));
 sg13g2_inv_1 _5280_ (.Y(_0413_),
    .A(_0412_));
 sg13g2_nor2_1 _5281_ (.A(_4424_),
    .B(net28),
    .Y(_0414_));
 sg13g2_inv_1 _5282_ (.Y(_0415_),
    .A(_0414_));
 sg13g2_buf_1 _5283_ (.A(_0415_),
    .X(_0416_));
 sg13g2_a21oi_1 _5284_ (.A1(_0407_),
    .A2(_0409_),
    .Y(_0201_),
    .B1(net27));
 sg13g2_inv_1 _5285_ (.Y(_0417_),
    .A(\main.demo.zic._q_rythm_count[9] ));
 sg13g2_inv_1 _5286_ (.Y(_0418_),
    .A(\main.demo.zic._q_rythm_count[10] ));
 sg13g2_nor3_1 _5287_ (.A(_4395_),
    .B(_4396_),
    .C(_0406_),
    .Y(_0419_));
 sg13g2_nand2_1 _5288_ (.Y(_0420_),
    .A(_0419_),
    .B(\main.demo.zic._q_rythm_count[2] ));
 sg13g2_nor2_1 _5289_ (.A(_4397_),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_nand2_1 _5290_ (.Y(_0422_),
    .A(_0421_),
    .B(\main.demo.zic._q_rythm_count[4] ));
 sg13g2_nor3_1 _5291_ (.A(_4392_),
    .B(_4393_),
    .C(_0422_),
    .Y(_0423_));
 sg13g2_nand3_1 _5292_ (.B(\main.demo.zic._q_rythm_count[8] ),
    .C(\main.demo.zic._q_rythm_count[7] ),
    .A(_0423_),
    .Y(_0424_));
 sg13g2_nor3_1 _5293_ (.A(_0417_),
    .B(_0418_),
    .C(_0424_),
    .Y(_0425_));
 sg13g2_nor2_1 _5294_ (.A(_0417_),
    .B(_0424_),
    .Y(_0426_));
 sg13g2_nor2_1 _5295_ (.A(\main.demo.zic._q_rythm_count[10] ),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_nor3_1 _5296_ (.A(_0415_),
    .B(_0425_),
    .C(_0427_),
    .Y(_0202_));
 sg13g2_inv_1 _5297_ (.Y(_0428_),
    .A(\main.demo.zic._q_rythm_count[7] ));
 sg13g2_nand3_1 _5298_ (.B(\main.demo.zic._q_rythm_count[0] ),
    .C(\main.demo.zic._q_rythm_count[2] ),
    .A(\main.demo.zic._q_rythm_count[1] ),
    .Y(_0429_));
 sg13g2_nand4_1 _5299_ (.B(\main.demo.zic._q_rythm_count[5] ),
    .C(\main.demo.zic._q_rythm_count[4] ),
    .A(\main.demo.zic._q_rythm_count[3] ),
    .Y(_0430_),
    .D(\main.demo.zic._q_rythm_count[6] ));
 sg13g2_nor4_2 _5300_ (.A(_0428_),
    .B(_0429_),
    .C(_0430_),
    .Y(_0431_),
    .D(_0406_));
 sg13g2_nand3_1 _5301_ (.B(\main.demo.zic._q_rythm_count[9] ),
    .C(\main.demo.zic._q_rythm_count[8] ),
    .A(_0431_),
    .Y(_0432_));
 sg13g2_nor3_1 _5302_ (.A(_4421_),
    .B(_0418_),
    .C(_0432_),
    .Y(_0433_));
 sg13g2_nor2_1 _5303_ (.A(\main.demo.zic._q_rythm_count[11] ),
    .B(_0425_),
    .Y(_0434_));
 sg13g2_nor3_1 _5304_ (.A(_0415_),
    .B(_0433_),
    .C(_0434_),
    .Y(_0203_));
 sg13g2_xnor2_1 _5305_ (.Y(_0435_),
    .A(\main.demo.zic._q_rythm_count[12] ),
    .B(_0433_));
 sg13g2_nor2_1 _5306_ (.A(_0435_),
    .B(net27),
    .Y(_0204_));
 sg13g2_buf_1 _5307_ (.A(net45),
    .X(_0436_));
 sg13g2_a21oi_1 _5308_ (.A1(net38),
    .A2(\main.demo.zic._q_rythm_count[0] ),
    .Y(_0437_),
    .B1(\main.demo.zic._q_rythm_count[1] ));
 sg13g2_nor3_1 _5309_ (.A(_0419_),
    .B(_0437_),
    .C(net27),
    .Y(_0205_));
 sg13g2_inv_1 _5310_ (.Y(_0438_),
    .A(_0420_));
 sg13g2_nor2_1 _5311_ (.A(\main.demo.zic._q_rythm_count[2] ),
    .B(_0419_),
    .Y(_0439_));
 sg13g2_nor3_1 _5312_ (.A(_0438_),
    .B(_0439_),
    .C(_0416_),
    .Y(_0206_));
 sg13g2_nor2_1 _5313_ (.A(\main.demo.zic._q_rythm_count[3] ),
    .B(_0438_),
    .Y(_0440_));
 sg13g2_nor3_1 _5314_ (.A(_0421_),
    .B(_0440_),
    .C(net27),
    .Y(_0207_));
 sg13g2_inv_1 _5315_ (.Y(_0441_),
    .A(_0422_));
 sg13g2_nor2_1 _5316_ (.A(\main.demo.zic._q_rythm_count[4] ),
    .B(_0421_),
    .Y(_0442_));
 sg13g2_nor3_1 _5317_ (.A(_0441_),
    .B(_0442_),
    .C(net27),
    .Y(_0208_));
 sg13g2_nor2_1 _5318_ (.A(_4392_),
    .B(_0422_),
    .Y(_0443_));
 sg13g2_nor2_1 _5319_ (.A(\main.demo.zic._q_rythm_count[5] ),
    .B(_0441_),
    .Y(_0444_));
 sg13g2_nor3_1 _5320_ (.A(_0443_),
    .B(_0444_),
    .C(net27),
    .Y(_0209_));
 sg13g2_nor2_1 _5321_ (.A(\main.demo.zic._q_rythm_count[6] ),
    .B(_0443_),
    .Y(_0445_));
 sg13g2_nor3_1 _5322_ (.A(_0423_),
    .B(_0445_),
    .C(net27),
    .Y(_0210_));
 sg13g2_nor2_1 _5323_ (.A(\main.demo.zic._q_rythm_count[7] ),
    .B(_0423_),
    .Y(_0446_));
 sg13g2_nor3_1 _5324_ (.A(_0431_),
    .B(_0446_),
    .C(net27),
    .Y(_0211_));
 sg13g2_nor2_1 _5325_ (.A(\main.demo.zic._q_rythm_count[8] ),
    .B(_0431_),
    .Y(_0447_));
 sg13g2_inv_1 _5326_ (.Y(_0448_),
    .A(_0424_));
 sg13g2_nor3_1 _5327_ (.A(_0447_),
    .B(_0448_),
    .C(_0416_),
    .Y(_0212_));
 sg13g2_nor2_1 _5328_ (.A(\main.demo.zic._q_rythm_count[9] ),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_nor3_1 _5329_ (.A(_0415_),
    .B(_0426_),
    .C(_0449_),
    .Y(_0213_));
 sg13g2_buf_1 _5330_ (.A(\main.demo._d___pip_58_1_4___block_87_atten_l[0] ),
    .X(_0450_));
 sg13g2_buf_1 _5331_ (.A(_0450_),
    .X(_0451_));
 sg13g2_inv_2 _5332_ (.Y(_0452_),
    .A(net70));
 sg13g2_inv_1 _5333_ (.Y(_0453_),
    .A(\main.demo._d_prev_b[5] ));
 sg13g2_buf_1 _5334_ (.A(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ),
    .X(_0454_));
 sg13g2_inv_1 _5335_ (.Y(_0455_),
    .A(net76));
 sg13g2_a21oi_1 _5336_ (.A1(_0452_),
    .A2(_0453_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_o21ai_1 _5337_ (.B1(_0456_),
    .Y(_0457_),
    .A1(_0452_),
    .A2(\main.demo._d_prev_b[3] ));
 sg13g2_inv_1 _5338_ (.Y(_0458_),
    .A(\main.demo._d_prev_b[7] ));
 sg13g2_a21oi_1 _5339_ (.A1(_0458_),
    .A2(net70),
    .Y(_0459_),
    .B1(net76));
 sg13g2_o21ai_1 _5340_ (.B1(_0459_),
    .Y(_0460_),
    .A1(net70),
    .A2(\main.demo._q_prev_b[7] ));
 sg13g2_inv_1 _5341_ (.Y(_0461_),
    .A(\main.demo._w_vga_active ));
 sg13g2_a21oi_1 _5342_ (.A1(_0457_),
    .A2(_0460_),
    .Y(_0072_),
    .B1(_0461_));
 sg13g2_buf_1 _5343_ (.A(\main.demo._w_vga_vga_x[6] ),
    .X(_0462_));
 sg13g2_inv_1 _5344_ (.Y(_0463_),
    .A(_0462_));
 sg13g2_buf_1 _5345_ (.A(\main.demo._w_vga_vga_x[5] ),
    .X(_0464_));
 sg13g2_inv_2 _5346_ (.Y(_0465_),
    .A(net75));
 sg13g2_buf_1 _5347_ (.A(\main.demo._w_vga_vga_y[5] ),
    .X(_0466_));
 sg13g2_buf_1 _5348_ (.A(\main.demo._w_vga_vga_y[6] ),
    .X(_0467_));
 sg13g2_nor2_1 _5349_ (.A(_0466_),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_nor2_1 _5350_ (.A(_0465_),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_buf_2 _5351_ (.A(\main.demo._w_vga_vga_x[7] ),
    .X(_0470_));
 sg13g2_o21ai_1 _5352_ (.B1(_0470_),
    .Y(_0471_),
    .A1(net69),
    .A2(_0469_));
 sg13g2_nand2_1 _5353_ (.Y(_0472_),
    .A(_0466_),
    .B(_0467_));
 sg13g2_buf_2 _5354_ (.A(_0472_),
    .X(_0473_));
 sg13g2_inv_1 _5355_ (.Y(_0474_),
    .A(_0468_));
 sg13g2_nand2_1 _5356_ (.Y(_0475_),
    .A(_0474_),
    .B(_0473_));
 sg13g2_nor2_1 _5357_ (.A(_0465_),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_nor2_1 _5358_ (.A(_0462_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_o21ai_1 _5359_ (.B1(_0477_),
    .Y(_0478_),
    .A1(_0464_),
    .A2(_0473_));
 sg13g2_nand2b_1 _5360_ (.Y(_0479_),
    .B(_0478_),
    .A_N(_0471_));
 sg13g2_nand3b_1 _5361_ (.B(_0474_),
    .C(_0465_),
    .Y(_0480_),
    .A_N(_0003_));
 sg13g2_inv_1 _5362_ (.Y(_0481_),
    .A(_0470_));
 sg13g2_nand2b_1 _5363_ (.Y(_0482_),
    .B(_0481_),
    .A_N(_0480_));
 sg13g2_buf_1 _5364_ (.A(\main.demo._w_vga_vga_x[8] ),
    .X(_0483_));
 sg13g2_a21oi_1 _5365_ (.A1(_0479_),
    .A2(_0482_),
    .Y(_0484_),
    .B1(_0483_));
 sg13g2_inv_1 _5366_ (.Y(_0485_),
    .A(_0483_));
 sg13g2_nor2_1 _5367_ (.A(net69),
    .B(_0476_),
    .Y(_0486_));
 sg13g2_nor2_1 _5368_ (.A(_0470_),
    .B(_0462_),
    .Y(_0487_));
 sg13g2_inv_1 _5369_ (.Y(_0488_),
    .A(_0487_));
 sg13g2_inv_1 _5370_ (.Y(_0489_),
    .A(_0466_));
 sg13g2_a21oi_1 _5371_ (.A1(_0465_),
    .A2(_0489_),
    .Y(_0490_),
    .B1(_0476_));
 sg13g2_inv_1 _5372_ (.Y(_0491_),
    .A(_0490_));
 sg13g2_nor2_1 _5373_ (.A(_0488_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_nor3_1 _5374_ (.A(_0485_),
    .B(_0486_),
    .C(_0492_),
    .Y(_0493_));
 sg13g2_inv_1 _5375_ (.Y(_0494_),
    .A(_0467_));
 sg13g2_nand2_1 _5376_ (.Y(_0495_),
    .A(net69),
    .B(_0470_));
 sg13g2_nor2_1 _5377_ (.A(net75),
    .B(_0489_),
    .Y(_0496_));
 sg13g2_a21oi_1 _5378_ (.A1(net75),
    .A2(_0467_),
    .Y(_0497_),
    .B1(_0496_));
 sg13g2_inv_1 _5379_ (.Y(_0498_),
    .A(_0497_));
 sg13g2_a21oi_1 _5380_ (.A1(net75),
    .A2(_0489_),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_nor2_1 _5381_ (.A(_0495_),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_o21ai_1 _5382_ (.B1(_0500_),
    .Y(_0501_),
    .A1(net75),
    .A2(_0494_));
 sg13g2_buf_1 _5383_ (.A(\main.demo._w_vga_vga_x[9] ),
    .X(_0502_));
 sg13g2_a21o_1 _5384_ (.A2(_0501_),
    .A1(_0493_),
    .B1(_0502_),
    .X(_0503_));
 sg13g2_nand3_1 _5385_ (.B(_0485_),
    .C(_0487_),
    .A(_0499_),
    .Y(_0504_));
 sg13g2_nand2_1 _5386_ (.Y(_0505_),
    .A(_0504_),
    .B(_0502_));
 sg13g2_o21ai_1 _5387_ (.B1(_0505_),
    .Y(_0506_),
    .A1(_0484_),
    .A2(_0503_));
 sg13g2_inv_1 _5388_ (.Y(_0507_),
    .A(_0502_));
 sg13g2_inv_1 _5389_ (.Y(_0508_),
    .A(_0001_));
 sg13g2_nor3_1 _5390_ (.A(_0507_),
    .B(_0508_),
    .C(_0488_),
    .Y(_0509_));
 sg13g2_nand2b_1 _5391_ (.Y(_0510_),
    .B(_0491_),
    .A_N(_0495_));
 sg13g2_nor2b_1 _5392_ (.A(_0466_),
    .B_N(_0004_),
    .Y(_0511_));
 sg13g2_a221oi_1 _5393_ (.B2(_0495_),
    .C1(_0485_),
    .B1(_0469_),
    .A1(_0511_),
    .Y(_0512_),
    .A2(_0487_));
 sg13g2_o21ai_1 _5394_ (.B1(_0469_),
    .Y(_0513_),
    .A1(net69),
    .A2(_0473_));
 sg13g2_nor2_1 _5395_ (.A(_0481_),
    .B(_0513_),
    .Y(_0514_));
 sg13g2_nor4_1 _5396_ (.A(_0470_),
    .B(net69),
    .C(_0465_),
    .D(_0473_),
    .Y(_0515_));
 sg13g2_nor4_1 _5397_ (.A(_0470_),
    .B(net69),
    .C(net75),
    .D(_0475_),
    .Y(_0516_));
 sg13g2_nor3_1 _5398_ (.A(_0514_),
    .B(_0515_),
    .C(_0516_),
    .Y(_0517_));
 sg13g2_a22oi_1 _5399_ (.Y(_0518_),
    .B1(_0485_),
    .B2(_0517_),
    .A2(_0512_),
    .A1(_0510_));
 sg13g2_a22oi_1 _5400_ (.Y(_0519_),
    .B1(_0507_),
    .B2(_0518_),
    .A2(_0509_),
    .A1(_0491_));
 sg13g2_nand2_1 _5401_ (.Y(_0520_),
    .A(_0506_),
    .B(_0519_));
 sg13g2_inv_1 _5402_ (.Y(_0521_),
    .A(_0520_));
 sg13g2_a21oi_1 _5403_ (.A1(_0473_),
    .A2(net75),
    .Y(_0522_),
    .B1(net69));
 sg13g2_nor4_1 _5404_ (.A(_0485_),
    .B(_0522_),
    .C(_0500_),
    .D(_0492_),
    .Y(_0523_));
 sg13g2_nor2_1 _5405_ (.A(_0467_),
    .B(_0465_),
    .Y(_0524_));
 sg13g2_inv_1 _5406_ (.Y(_0525_),
    .A(_0473_));
 sg13g2_nor3_1 _5407_ (.A(_0003_),
    .B(_0524_),
    .C(_0525_),
    .Y(_0526_));
 sg13g2_nor3_1 _5408_ (.A(_0481_),
    .B(_0522_),
    .C(_0477_),
    .Y(_0527_));
 sg13g2_a21oi_1 _5409_ (.A1(_0481_),
    .A2(_0526_),
    .Y(_0528_),
    .B1(_0527_));
 sg13g2_o21ai_1 _5410_ (.B1(_0507_),
    .Y(_0529_),
    .A1(_0483_),
    .A2(_0528_));
 sg13g2_o21ai_1 _5411_ (.B1(_0505_),
    .Y(_0530_),
    .A1(_0523_),
    .A2(_0529_));
 sg13g2_a21oi_1 _5412_ (.A1(_0010_),
    .A2(_0467_),
    .Y(_0531_),
    .B1(_0524_));
 sg13g2_a21oi_1 _5413_ (.A1(_0531_),
    .A2(_0463_),
    .Y(_0532_),
    .B1(_0481_));
 sg13g2_inv_1 _5414_ (.Y(_0533_),
    .A(_0486_));
 sg13g2_a21oi_1 _5415_ (.A1(_0532_),
    .A2(_0533_),
    .Y(_0534_),
    .B1(_0516_));
 sg13g2_a21oi_1 _5416_ (.A1(_0473_),
    .A2(net75),
    .Y(_0535_),
    .B1(_0511_));
 sg13g2_nor3_1 _5417_ (.A(_0466_),
    .B(_0465_),
    .C(_0494_),
    .Y(_0536_));
 sg13g2_nor3_1 _5418_ (.A(_0481_),
    .B(_0496_),
    .C(_0536_),
    .Y(_0537_));
 sg13g2_o21ai_1 _5419_ (.B1(_0533_),
    .Y(_0538_),
    .A1(_0462_),
    .A2(_0537_));
 sg13g2_o21ai_1 _5420_ (.B1(_0538_),
    .Y(_0539_),
    .A1(_0488_),
    .A2(_0535_));
 sg13g2_nand2_1 _5421_ (.Y(_0540_),
    .A(_0539_),
    .B(_0483_));
 sg13g2_o21ai_1 _5422_ (.B1(_0540_),
    .Y(_0541_),
    .A1(_0483_),
    .A2(_0534_));
 sg13g2_a22oi_1 _5423_ (.Y(_0542_),
    .B1(_0507_),
    .B2(_0541_),
    .A2(_0497_),
    .A1(_0509_));
 sg13g2_nor2_1 _5424_ (.A(_0530_),
    .B(_0542_),
    .Y(_0543_));
 sg13g2_inv_1 _5425_ (.Y(_0544_),
    .A(\main.demo._w_vga_vga_x[4] ));
 sg13g2_nand2_1 _5426_ (.Y(_0545_),
    .A(_0530_),
    .B(_0519_));
 sg13g2_buf_2 _5427_ (.A(_0545_),
    .X(_0546_));
 sg13g2_xnor2_1 _5428_ (.Y(_0547_),
    .A(_0544_),
    .B(_0546_));
 sg13g2_inv_1 _5429_ (.Y(_0548_),
    .A(_0547_));
 sg13g2_buf_2 _5430_ (.A(\main.demo._t___stage___block_3_x[1] ),
    .X(_0549_));
 sg13g2_inv_1 _5431_ (.Y(_0550_),
    .A(_0549_));
 sg13g2_xnor2_1 _5432_ (.Y(_0551_),
    .A(_0550_),
    .B(_0546_));
 sg13g2_buf_2 _5433_ (.A(\main.demo._t___stage___block_3_y[0] ),
    .X(_0552_));
 sg13g2_inv_1 _5434_ (.Y(_0553_),
    .A(_0552_));
 sg13g2_a21oi_1 _5435_ (.A1(_0546_),
    .A2(_0016_),
    .Y(_0554_),
    .B1(_0553_));
 sg13g2_o21ai_1 _5436_ (.B1(_0554_),
    .Y(_0555_),
    .A1(_0016_),
    .A2(_0546_));
 sg13g2_o21ai_1 _5437_ (.B1(_0555_),
    .Y(_0556_),
    .A1(_0014_),
    .A2(_0551_));
 sg13g2_nand2_1 _5438_ (.Y(_0557_),
    .A(_0551_),
    .B(_0014_));
 sg13g2_buf_1 _5439_ (.A(\main.demo._t___stage___block_3_x[2] ),
    .X(_0558_));
 sg13g2_inv_2 _5440_ (.Y(_0559_),
    .A(_0558_));
 sg13g2_xnor2_1 _5441_ (.Y(_0560_),
    .A(_0559_),
    .B(_0546_));
 sg13g2_xnor2_1 _5442_ (.Y(_0561_),
    .A(_0015_),
    .B(_0560_));
 sg13g2_a21o_1 _5443_ (.A2(_0557_),
    .A1(_0556_),
    .B1(_0561_),
    .X(_0562_));
 sg13g2_buf_1 _5444_ (.A(\main.demo._t___stage___block_3_y[2] ),
    .X(_0563_));
 sg13g2_inv_1 _5445_ (.Y(_0564_),
    .A(_0563_));
 sg13g2_nand2_1 _5446_ (.Y(_0565_),
    .A(_0560_),
    .B(_0564_));
 sg13g2_nand2_1 _5447_ (.Y(_0566_),
    .A(_0562_),
    .B(_0565_));
 sg13g2_xnor2_1 _5448_ (.Y(_0567_),
    .A(\main.demo._w_vga_vga_x[3] ),
    .B(_0546_));
 sg13g2_xnor2_1 _5449_ (.Y(_0568_),
    .A(_0011_),
    .B(_0567_));
 sg13g2_nor2_1 _5450_ (.A(\main.demo._w_vga_vga_y[3] ),
    .B(_0567_),
    .Y(_0569_));
 sg13g2_a221oi_1 _5451_ (.B2(_0568_),
    .C1(_0569_),
    .B1(_0566_),
    .A1(_4177_),
    .Y(_0570_),
    .A2(_0547_));
 sg13g2_a21oi_1 _5452_ (.A1(_4170_),
    .A2(_0548_),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_nor3_1 _5453_ (.A(_0521_),
    .B(_0543_),
    .C(_0571_),
    .Y(_0572_));
 sg13g2_nand2_1 _5454_ (.Y(_0573_),
    .A(_0571_),
    .B(_0521_));
 sg13g2_buf_2 _5455_ (.A(\main.demo._t___stage___block_3_x[0] ),
    .X(_0574_));
 sg13g2_inv_1 _5456_ (.Y(_0575_),
    .A(_0574_));
 sg13g2_a22oi_1 _5457_ (.Y(_0576_),
    .B1(_0550_),
    .B2(_0312_),
    .A2(\main.demo._q_th[1] ),
    .A1(_0575_));
 sg13g2_a21oi_1 _5458_ (.A1(_0549_),
    .A2(_0314_),
    .Y(_0577_),
    .B1(_0576_));
 sg13g2_o21ai_1 _5459_ (.B1(_0577_),
    .Y(_0578_),
    .A1(_0559_),
    .A2(_0316_));
 sg13g2_nand2b_1 _5460_ (.Y(_0579_),
    .B(\main.demo._q_th[4] ),
    .A_N(\main.demo._w_vga_vga_x[3] ));
 sg13g2_nand2_1 _5461_ (.Y(_0580_),
    .A(_0559_),
    .B(_0316_));
 sg13g2_nand3_1 _5462_ (.B(_0579_),
    .C(_0580_),
    .A(_0578_),
    .Y(_0581_));
 sg13g2_a22oi_1 _5463_ (.Y(_0582_),
    .B1(_0320_),
    .B2(\main.demo._w_vga_vga_x[3] ),
    .A2(\main.demo._w_vga_vga_x[4] ),
    .A1(_0323_));
 sg13g2_nor3_1 _5464_ (.A(_0330_),
    .B(_0326_),
    .C(\main.demo._q_th[8] ),
    .Y(_0583_));
 sg13g2_o21ai_1 _5465_ (.B1(_0583_),
    .Y(_0584_),
    .A1(_0323_),
    .A2(\main.demo._w_vga_vga_x[4] ));
 sg13g2_a21oi_1 _5466_ (.A1(_0581_),
    .A2(_0582_),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_nor2b_1 _5467_ (.A(\main.demo._w_vga_vga_y[7] ),
    .B_N(_0007_),
    .Y(_0586_));
 sg13g2_buf_1 _5468_ (.A(\main.demo._t___stage___block_3_y[1] ),
    .X(_0587_));
 sg13g2_inv_1 _5469_ (.Y(_0588_),
    .A(_0013_));
 sg13g2_nor3_1 _5470_ (.A(net74),
    .B(_0563_),
    .C(_0588_),
    .Y(_0589_));
 sg13g2_nor3_1 _5471_ (.A(\main.demo._w_vga_vga_y[3] ),
    .B(\main.demo._w_vga_vga_y[7] ),
    .C(_0553_),
    .Y(_0590_));
 sg13g2_nor2b_1 _5472_ (.A(_4170_),
    .B_N(_4141_),
    .Y(_0591_));
 sg13g2_nand4_1 _5473_ (.B(_0590_),
    .C(_0468_),
    .A(_0589_),
    .Y(_0592_),
    .D(_0591_));
 sg13g2_o21ai_1 _5474_ (.B1(_0592_),
    .Y(_0593_),
    .A1(_4141_),
    .A2(_0586_));
 sg13g2_nand3b_1 _5475_ (.B(_0593_),
    .C(_4278_),
    .Y(_0594_),
    .A_N(\main.demo._w_vga_vga_y[10] ));
 sg13g2_and3_1 _5476_ (.X(_0595_),
    .A(_0521_),
    .B(_0530_),
    .C(_0542_));
 sg13g2_nor3_1 _5477_ (.A(_0585_),
    .B(_0594_),
    .C(_0595_),
    .Y(_0596_));
 sg13g2_nand3b_1 _5478_ (.B(_0573_),
    .C(_0596_),
    .Y(_0597_),
    .A_N(_0572_));
 sg13g2_xnor2_1 _5479_ (.Y(_0598_),
    .A(_0574_),
    .B(_0552_));
 sg13g2_buf_2 _5480_ (.A(_0598_),
    .X(_0599_));
 sg13g2_inv_1 _5481_ (.Y(_0600_),
    .A(_0599_));
 sg13g2_buf_8 _5482_ (.A(_0600_),
    .X(_0601_));
 sg13g2_inv_1 _5483_ (.Y(_0602_),
    .A(_4159_));
 sg13g2_xnor2_1 _5484_ (.Y(_0603_),
    .A(net74),
    .B(_0549_));
 sg13g2_inv_1 _5485_ (.Y(_0604_),
    .A(_0603_));
 sg13g2_nor2_1 _5486_ (.A(net74),
    .B(_4353_),
    .Y(_0605_));
 sg13g2_nand3_1 _5487_ (.B(_0564_),
    .C(_4164_),
    .A(_0559_),
    .Y(_0606_));
 sg13g2_inv_1 _5488_ (.Y(_0607_),
    .A(_4171_));
 sg13g2_xnor2_1 _5489_ (.Y(_0608_),
    .A(_0558_),
    .B(_0563_));
 sg13g2_a21oi_1 _5490_ (.A1(_4164_),
    .A2(_0564_),
    .Y(_0609_),
    .B1(_0608_));
 sg13g2_a221oi_1 _5491_ (.B2(_0607_),
    .C1(_0609_),
    .B1(_0606_),
    .A1(_4353_),
    .Y(_0610_),
    .A2(net74));
 sg13g2_nand2_1 _5492_ (.Y(_0611_),
    .A(_0604_),
    .B(_0602_));
 sg13g2_o21ai_1 _5493_ (.B1(_0611_),
    .Y(_0612_),
    .A1(_0605_),
    .A2(_0610_));
 sg13g2_o21ai_1 _5494_ (.B1(_0612_),
    .Y(_0613_),
    .A1(_0602_),
    .A2(_0604_));
 sg13g2_o21ai_1 _5495_ (.B1(_0613_),
    .Y(_0614_),
    .A1(_4146_),
    .A2(_0553_));
 sg13g2_buf_8 _5496_ (.A(_0599_),
    .X(_0615_));
 sg13g2_a22oi_1 _5497_ (.Y(_0616_),
    .B1(_4148_),
    .B2(net51),
    .A2(_0553_),
    .A1(_4146_));
 sg13g2_nand4_1 _5498_ (.B(_4140_),
    .C(_4296_),
    .A(_4288_),
    .Y(_0617_),
    .D(\main.demo._q_go ));
 sg13g2_a221oi_1 _5499_ (.B2(_0616_),
    .C1(_0617_),
    .B1(_0614_),
    .A1(_4149_),
    .Y(_0618_),
    .A2(net44));
 sg13g2_nor2_1 _5500_ (.A(\main.demo._d___pip_58_1_4___stage___block_3_cx[5] ),
    .B(_0553_),
    .Y(_0619_));
 sg13g2_nand2b_1 _5501_ (.Y(_0620_),
    .B(_0604_),
    .A_N(\main.demo._d___pip_58_1_4___stage___block_3_cx[4] ));
 sg13g2_inv_1 _5502_ (.Y(_0621_),
    .A(\main.demo._d___pip_58_1_4___stage___block_3_cx[3] ));
 sg13g2_nand2_1 _5503_ (.Y(_0622_),
    .A(_0621_),
    .B(net74));
 sg13g2_nand2_1 _5504_ (.Y(_0623_),
    .A(_0620_),
    .B(_0622_));
 sg13g2_nor2b_1 _5505_ (.A(_0563_),
    .B_N(\main.demo._d___pip_58_1_4___stage___block_3_cx[1] ),
    .Y(_0624_));
 sg13g2_o21ai_1 _5506_ (.B1(_0624_),
    .Y(_0625_),
    .A1(_0559_),
    .A2(\main.demo._d___pip_58_1_4___stage___block_3_cx[2] ));
 sg13g2_o21ai_1 _5507_ (.B1(_0625_),
    .Y(_0626_),
    .A1(_0587_),
    .A2(_0621_));
 sg13g2_a21oi_1 _5508_ (.A1(\main.demo._d___pip_58_1_4___stage___block_3_cx[2] ),
    .A2(_0608_),
    .Y(_0627_),
    .B1(_0626_));
 sg13g2_a22oi_1 _5509_ (.Y(_0628_),
    .B1(\main.demo._d___pip_58_1_4___stage___block_3_cx[4] ),
    .B2(_0603_),
    .A2(\main.demo._d___pip_58_1_4___stage___block_3_cx[5] ),
    .A1(_0553_));
 sg13g2_o21ai_1 _5510_ (.B1(_0628_),
    .Y(_0629_),
    .A1(_0623_),
    .A2(_0627_));
 sg13g2_nor2b_1 _5511_ (.A(_0619_),
    .B_N(_0629_),
    .Y(_0630_));
 sg13g2_o21ai_1 _5512_ (.B1(_0630_),
    .Y(_0631_),
    .A1(\main.demo._d___pip_58_1_4___stage___block_3_cx[6] ),
    .A2(net51));
 sg13g2_a21oi_1 _5513_ (.A1(net51),
    .A2(\main.demo._d___pip_58_1_4___stage___block_3_cx[6] ),
    .Y(_0632_),
    .B1(\main.demo._d___pip_58_1_4___stage___block_3_cx[9] ));
 sg13g2_nand2_1 _5514_ (.Y(_0633_),
    .A(_0631_),
    .B(_0632_));
 sg13g2_buf_2 _5515_ (.A(_0633_),
    .X(_0634_));
 sg13g2_inv_1 _5516_ (.Y(_0635_),
    .A(_0634_));
 sg13g2_buf_1 _5517_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[4] ),
    .X(_0636_));
 sg13g2_buf_1 _5518_ (.A(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ),
    .X(_0637_));
 sg13g2_nand2_1 _5519_ (.Y(_0638_),
    .A(_0636_),
    .B(_0637_));
 sg13g2_buf_1 _5520_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[5] ),
    .X(_0639_));
 sg13g2_buf_1 _5521_ (.A(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ),
    .X(_0640_));
 sg13g2_nand3_1 _5522_ (.B(_0639_),
    .C(_0640_),
    .A(_0638_),
    .Y(_0641_));
 sg13g2_buf_1 _5523_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[3] ),
    .X(_0642_));
 sg13g2_nand2_1 _5524_ (.Y(_0643_),
    .A(_0642_),
    .B(_0637_));
 sg13g2_buf_1 _5525_ (.A(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ),
    .X(_0644_));
 sg13g2_nand2_1 _5526_ (.Y(_0645_),
    .A(_0636_),
    .B(_0644_));
 sg13g2_nand2_1 _5527_ (.Y(_0646_),
    .A(_0643_),
    .B(_0645_));
 sg13g2_buf_1 _5528_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[2] ),
    .X(_0647_));
 sg13g2_nand2_1 _5529_ (.Y(_0648_),
    .A(_0647_),
    .B(_0640_));
 sg13g2_inv_1 _5530_ (.Y(_0649_),
    .A(_0648_));
 sg13g2_nand2_1 _5531_ (.Y(_0650_),
    .A(_0642_),
    .B(_0644_));
 sg13g2_nor2_1 _5532_ (.A(_0650_),
    .B(_0638_),
    .Y(_0651_));
 sg13g2_a21oi_1 _5533_ (.A1(_0646_),
    .A2(_0649_),
    .Y(_0652_),
    .B1(_0651_));
 sg13g2_nand2_1 _5534_ (.Y(_0653_),
    .A(_0642_),
    .B(_0640_));
 sg13g2_nand2_1 _5535_ (.Y(_0654_),
    .A(_0639_),
    .B(_0637_));
 sg13g2_nor2_1 _5536_ (.A(_0645_),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_inv_1 _5537_ (.Y(_0656_),
    .A(_0639_));
 sg13g2_inv_1 _5538_ (.Y(_0657_),
    .A(_0644_));
 sg13g2_o21ai_1 _5539_ (.B1(_0638_),
    .Y(_0658_),
    .A1(_0656_),
    .A2(_0657_));
 sg13g2_nand2b_1 _5540_ (.Y(_0659_),
    .B(_0658_),
    .A_N(_0655_));
 sg13g2_xnor2_1 _5541_ (.Y(_0660_),
    .A(_0653_),
    .B(_0659_));
 sg13g2_nand2_1 _5542_ (.Y(_0661_),
    .A(_0647_),
    .B(_0637_));
 sg13g2_xor2_1 _5543_ (.B(_0661_),
    .A(_0650_),
    .X(_0662_));
 sg13g2_nand2_1 _5544_ (.Y(_0663_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[1] ),
    .B(_0640_));
 sg13g2_inv_1 _5545_ (.Y(_0664_),
    .A(_0663_));
 sg13g2_nand2_1 _5546_ (.Y(_0665_),
    .A(_0647_),
    .B(_0644_));
 sg13g2_nor2_1 _5547_ (.A(_0643_),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_a21oi_1 _5548_ (.A1(_0662_),
    .A2(_0664_),
    .Y(_0667_),
    .B1(_0666_));
 sg13g2_o21ai_1 _5549_ (.B1(_0646_),
    .Y(_0668_),
    .A1(_0650_),
    .A2(_0638_));
 sg13g2_xnor2_1 _5550_ (.Y(_0669_),
    .A(_0648_),
    .B(_0668_));
 sg13g2_nand2_1 _5551_ (.Y(_0670_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[1] ),
    .B(_0637_));
 sg13g2_nand2_1 _5552_ (.Y(_0671_),
    .A(_0665_),
    .B(_0670_));
 sg13g2_nand2_1 _5553_ (.Y(_0672_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[0] ),
    .B(_0640_));
 sg13g2_inv_1 _5554_ (.Y(_0673_),
    .A(_0672_));
 sg13g2_nor2_1 _5555_ (.A(_0665_),
    .B(_0670_),
    .Y(_0674_));
 sg13g2_a21oi_1 _5556_ (.A1(_0671_),
    .A2(_0673_),
    .Y(_0675_),
    .B1(_0674_));
 sg13g2_xnor2_1 _5557_ (.Y(_0676_),
    .A(_0664_),
    .B(_0662_));
 sg13g2_xor2_1 _5558_ (.B(_0676_),
    .A(_0675_),
    .X(_0677_));
 sg13g2_nor2b_1 _5559_ (.A(_0674_),
    .B_N(_0671_),
    .Y(_0678_));
 sg13g2_xnor2_1 _5560_ (.Y(_0679_),
    .A(_0673_),
    .B(_0678_));
 sg13g2_inv_1 _5561_ (.Y(_0680_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[0] ));
 sg13g2_nor3_1 _5562_ (.A(_0680_),
    .B(_0657_),
    .C(_0670_),
    .Y(_0681_));
 sg13g2_nor2b_1 _5563_ (.A(_0679_),
    .B_N(_0681_),
    .Y(_0682_));
 sg13g2_nand2_1 _5564_ (.Y(_0683_),
    .A(_0677_),
    .B(_0682_));
 sg13g2_o21ai_1 _5565_ (.B1(_0683_),
    .Y(_0684_),
    .A1(_0675_),
    .A2(_0676_));
 sg13g2_xor2_1 _5566_ (.B(_0669_),
    .A(_0667_),
    .X(_0685_));
 sg13g2_nand2_1 _5567_ (.Y(_0686_),
    .A(_0684_),
    .B(_0685_));
 sg13g2_o21ai_1 _5568_ (.B1(_0686_),
    .Y(_0687_),
    .A1(_0667_),
    .A2(_0669_));
 sg13g2_xor2_1 _5569_ (.B(_0660_),
    .A(_0652_),
    .X(_0688_));
 sg13g2_nand2_1 _5570_ (.Y(_0689_),
    .A(_0687_),
    .B(_0688_));
 sg13g2_o21ai_1 _5571_ (.B1(_0689_),
    .Y(_0690_),
    .A1(_0652_),
    .A2(_0660_));
 sg13g2_nand2_1 _5572_ (.Y(_0691_),
    .A(_0636_),
    .B(_0640_));
 sg13g2_xnor2_1 _5573_ (.Y(_0692_),
    .A(_0654_),
    .B(_0691_));
 sg13g2_inv_1 _5574_ (.Y(_0693_),
    .A(_0653_));
 sg13g2_a21oi_1 _5575_ (.A1(_0658_),
    .A2(_0693_),
    .Y(_0694_),
    .B1(_0655_));
 sg13g2_xor2_1 _5576_ (.B(_0694_),
    .A(_0692_),
    .X(_0695_));
 sg13g2_nor2_1 _5577_ (.A(_0692_),
    .B(_0694_),
    .Y(_0696_));
 sg13g2_a21oi_1 _5578_ (.A1(_0690_),
    .A2(_0695_),
    .Y(_0697_),
    .B1(_0696_));
 sg13g2_xnor2_1 _5579_ (.Y(_0698_),
    .A(_0641_),
    .B(_0697_));
 sg13g2_nand2_1 _5580_ (.Y(_0699_),
    .A(_0450_),
    .B(_0636_));
 sg13g2_nand2_1 _5581_ (.Y(_0700_),
    .A(net76),
    .B(_0642_));
 sg13g2_nand2_1 _5582_ (.Y(_0701_),
    .A(_0450_),
    .B(_0642_));
 sg13g2_nand2_1 _5583_ (.Y(_0702_),
    .A(net76),
    .B(_0647_));
 sg13g2_xor2_1 _5584_ (.B(_0702_),
    .A(_0701_),
    .X(_0703_));
 sg13g2_nand2_1 _5585_ (.Y(_0704_),
    .A(_0450_),
    .B(_0647_));
 sg13g2_nand2_1 _5586_ (.Y(_0705_),
    .A(_0450_),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[0] ));
 sg13g2_nand2_1 _5587_ (.Y(_0706_),
    .A(net76),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[1] ));
 sg13g2_a21oi_1 _5588_ (.A1(_0704_),
    .A2(_0705_),
    .Y(_0707_),
    .B1(_0706_));
 sg13g2_nor2_1 _5589_ (.A(_0701_),
    .B(_0702_),
    .Y(_0708_));
 sg13g2_a21oi_1 _5590_ (.A1(_0703_),
    .A2(_0707_),
    .Y(_0709_),
    .B1(_0708_));
 sg13g2_xor2_1 _5591_ (.B(_0700_),
    .A(_0699_),
    .X(_0710_));
 sg13g2_nand2b_1 _5592_ (.Y(_0711_),
    .B(_0710_),
    .A_N(_0709_));
 sg13g2_o21ai_1 _5593_ (.B1(_0711_),
    .Y(_0712_),
    .A1(_0699_),
    .A2(_0700_));
 sg13g2_nand2_1 _5594_ (.Y(_0713_),
    .A(_0454_),
    .B(_0636_));
 sg13g2_nand2_1 _5595_ (.Y(_0714_),
    .A(_0450_),
    .B(_0639_));
 sg13g2_xor2_1 _5596_ (.B(_0714_),
    .A(_0713_),
    .X(_0715_));
 sg13g2_nand2_1 _5597_ (.Y(_0716_),
    .A(_0712_),
    .B(_0715_));
 sg13g2_nand2_1 _5598_ (.Y(_0717_),
    .A(_0454_),
    .B(_0639_));
 sg13g2_a21oi_1 _5599_ (.A1(_0716_),
    .A2(_0699_),
    .Y(_0718_),
    .B1(_0717_));
 sg13g2_nand2_1 _5600_ (.Y(_0719_),
    .A(_0635_),
    .B(_0718_));
 sg13g2_o21ai_1 _5601_ (.B1(_0719_),
    .Y(_0720_),
    .A1(_0635_),
    .A2(_0698_));
 sg13g2_xnor2_1 _5602_ (.Y(_0721_),
    .A(_0695_),
    .B(_0690_));
 sg13g2_nand2_1 _5603_ (.Y(_0722_),
    .A(_0721_),
    .B(_0634_));
 sg13g2_nor2b_1 _5604_ (.A(_0634_),
    .B_N(_0716_),
    .Y(_0723_));
 sg13g2_nand2_1 _5605_ (.Y(_0724_),
    .A(_0723_),
    .B(_0717_));
 sg13g2_nand3_1 _5606_ (.B(_0724_),
    .C(_0719_),
    .A(_0722_),
    .Y(_0725_));
 sg13g2_xor2_1 _5607_ (.B(_0703_),
    .A(_0707_),
    .X(_0726_));
 sg13g2_xnor2_1 _5608_ (.Y(_0727_),
    .A(_0682_),
    .B(_0677_));
 sg13g2_nand2_1 _5609_ (.Y(_0728_),
    .A(_0634_),
    .B(_0727_));
 sg13g2_o21ai_1 _5610_ (.B1(_0728_),
    .Y(_0729_),
    .A1(_0634_),
    .A2(_0726_));
 sg13g2_nand2b_1 _5611_ (.Y(_0730_),
    .B(_0603_),
    .A_N(_0729_));
 sg13g2_nand2b_1 _5612_ (.Y(_0731_),
    .B(_0679_),
    .A_N(_0681_));
 sg13g2_nand2b_1 _5613_ (.Y(_0732_),
    .B(_0731_),
    .A_N(_0682_));
 sg13g2_a21oi_1 _5614_ (.A1(net70),
    .A2(\main.demo._d___pip_58_1_4___block_68_frag[0] ),
    .Y(_0733_),
    .B1(_0706_));
 sg13g2_xnor2_1 _5615_ (.Y(_0734_),
    .A(_0704_),
    .B(_0733_));
 sg13g2_nor2_1 _5616_ (.A(_0734_),
    .B(_0634_),
    .Y(_0735_));
 sg13g2_a21oi_1 _5617_ (.A1(_0634_),
    .A2(_0732_),
    .Y(_0736_),
    .B1(_0735_));
 sg13g2_nand2_1 _5618_ (.Y(_0737_),
    .A(_0729_),
    .B(_0604_));
 sg13g2_o21ai_1 _5619_ (.B1(_0737_),
    .Y(_0738_),
    .A1(_0550_),
    .A2(_0736_));
 sg13g2_xnor2_1 _5620_ (.Y(_0739_),
    .A(_0688_),
    .B(_0687_));
 sg13g2_o21ai_1 _5621_ (.B1(_0723_),
    .Y(_0740_),
    .A1(_0715_),
    .A2(_0712_));
 sg13g2_o21ai_1 _5622_ (.B1(_0740_),
    .Y(_0741_),
    .A1(_0635_),
    .A2(_0739_));
 sg13g2_xnor2_1 _5623_ (.Y(_0742_),
    .A(_0601_),
    .B(_0741_));
 sg13g2_inv_1 _5624_ (.Y(_0743_),
    .A(_0016_));
 sg13g2_nor2b_1 _5625_ (.A(_0635_),
    .B_N(_0686_),
    .Y(_0744_));
 sg13g2_o21ai_1 _5626_ (.B1(_0744_),
    .Y(_0745_),
    .A1(_0685_),
    .A2(_0684_));
 sg13g2_nand2b_1 _5627_ (.Y(_0746_),
    .B(_0709_),
    .A_N(_0710_));
 sg13g2_nand3_1 _5628_ (.B(_0711_),
    .C(_0746_),
    .A(_0635_),
    .Y(_0747_));
 sg13g2_nand2_1 _5629_ (.Y(_0748_),
    .A(_0745_),
    .B(_0747_));
 sg13g2_xnor2_1 _5630_ (.Y(_0749_),
    .A(_0743_),
    .B(_0748_));
 sg13g2_nand2_1 _5631_ (.Y(_0750_),
    .A(_0742_),
    .B(_0749_));
 sg13g2_a21oi_1 _5632_ (.A1(_0730_),
    .A2(_0738_),
    .Y(_0751_),
    .B1(_0750_));
 sg13g2_a21oi_1 _5633_ (.A1(_0745_),
    .A2(_0747_),
    .Y(_0752_),
    .B1(_0574_));
 sg13g2_nor2b_1 _5634_ (.A(net44),
    .B_N(_0741_),
    .Y(_0753_));
 sg13g2_a21oi_1 _5635_ (.A1(_0742_),
    .A2(_0752_),
    .Y(_0754_),
    .B1(_0753_));
 sg13g2_nand2b_1 _5636_ (.Y(_0755_),
    .B(_0754_),
    .A_N(_0751_));
 sg13g2_inv_1 _5637_ (.Y(_0756_),
    .A(_0750_));
 sg13g2_xor2_1 _5638_ (.B(_0736_),
    .A(_0017_),
    .X(_0757_));
 sg13g2_nand4_1 _5639_ (.B(_0737_),
    .C(_0730_),
    .A(_0756_),
    .Y(_0758_),
    .D(_0757_));
 sg13g2_nand2_1 _5640_ (.Y(_0759_),
    .A(_0755_),
    .B(_0758_));
 sg13g2_nor2_1 _5641_ (.A(_0725_),
    .B(_0759_),
    .Y(_0760_));
 sg13g2_nor3_1 _5642_ (.A(_0618_),
    .B(_0720_),
    .C(_0760_),
    .Y(_0761_));
 sg13g2_nand2_1 _5643_ (.Y(\main.demo._d_prev_b[1] ),
    .A(_0597_),
    .B(_0761_));
 sg13g2_a21oi_1 _5644_ (.A1(_0597_),
    .A2(_0761_),
    .Y(_0073_),
    .B1(_0461_));
 sg13g2_a21oi_1 _5645_ (.A1(_0452_),
    .A2(_0458_),
    .Y(_0762_),
    .B1(_0455_));
 sg13g2_o21ai_1 _5646_ (.B1(_0762_),
    .Y(_0763_),
    .A1(_0452_),
    .A2(\main.demo._q_prev_b[7] ));
 sg13g2_a21oi_1 _5647_ (.A1(_0453_),
    .A2(net70),
    .Y(_0764_),
    .B1(net76));
 sg13g2_o21ai_1 _5648_ (.B1(_0764_),
    .Y(_0765_),
    .A1(net70),
    .A2(\main.demo._d_prev_b[3] ));
 sg13g2_a21oi_1 _5649_ (.A1(_0763_),
    .A2(_0765_),
    .Y(_0074_),
    .B1(_0461_));
 sg13g2_inv_1 _5650_ (.Y(_0766_),
    .A(\main.demo._d_prev_b[4] ));
 sg13g2_a21oi_1 _5651_ (.A1(_0766_),
    .A2(_0452_),
    .Y(_0767_),
    .B1(_0455_));
 sg13g2_o21ai_1 _5652_ (.B1(_0767_),
    .Y(_0768_),
    .A1(\main.demo._d_prev_b[2] ),
    .A2(_0452_));
 sg13g2_inv_1 _5653_ (.Y(_0769_),
    .A(\main.demo._d_prev_b[6] ));
 sg13g2_a21oi_1 _5654_ (.A1(_0769_),
    .A2(net70),
    .Y(_0770_),
    .B1(net76));
 sg13g2_o21ai_1 _5655_ (.B1(_0770_),
    .Y(_0771_),
    .A1(net70),
    .A2(\main.demo._q_prev_b[6] ));
 sg13g2_a21oi_1 _5656_ (.A1(_0768_),
    .A2(_0771_),
    .Y(_0075_),
    .B1(_0461_));
 sg13g2_nor3_1 _5657_ (.A(_0725_),
    .B(_0720_),
    .C(_0759_),
    .Y(_0772_));
 sg13g2_a21oi_1 _5658_ (.A1(_0759_),
    .A2(_0725_),
    .Y(_0773_),
    .B1(_0772_));
 sg13g2_nor2_1 _5659_ (.A(_0618_),
    .B(_0773_),
    .Y(_0774_));
 sg13g2_inv_1 _5660_ (.Y(\main.demo._d_prev_b[0] ),
    .A(_0774_));
 sg13g2_nor2_1 _5661_ (.A(_0461_),
    .B(_0774_),
    .Y(_0076_));
 sg13g2_a21oi_1 _5662_ (.A1(_0452_),
    .A2(_0769_),
    .Y(_0775_),
    .B1(_0455_));
 sg13g2_o21ai_1 _5663_ (.B1(_0775_),
    .Y(_0776_),
    .A1(_0452_),
    .A2(\main.demo._q_prev_b[6] ));
 sg13g2_a21oi_1 _5664_ (.A1(_0766_),
    .A2(_0451_),
    .Y(_0777_),
    .B1(net76));
 sg13g2_o21ai_1 _5665_ (.B1(_0777_),
    .Y(_0778_),
    .A1(\main.demo._d_prev_b[2] ),
    .A2(_0451_));
 sg13g2_a21oi_1 _5666_ (.A1(_0776_),
    .A2(_0778_),
    .Y(_0077_),
    .B1(_0461_));
 sg13g2_inv_1 _5667_ (.Y(_0779_),
    .A(_4273_));
 sg13g2_nor2_1 _5668_ (.A(_4271_),
    .B(_0306_),
    .Y(_0780_));
 sg13g2_inv_1 _5669_ (.Y(_0781_),
    .A(_0780_));
 sg13g2_buf_1 _5670_ (.A(rst_n_q),
    .X(_0782_));
 sg13g2_nand2_1 _5671_ (.Y(_0783_),
    .A(\main.demo._q_go ),
    .B(_0782_));
 sg13g2_inv_1 _5672_ (.Y(_0784_),
    .A(_0783_));
 sg13g2_o21ai_1 _5673_ (.B1(_0784_),
    .Y(_0785_),
    .A1(_0069_),
    .A2(_0781_));
 sg13g2_a21oi_1 _5674_ (.A1(_0779_),
    .A2(_0781_),
    .Y(_0078_),
    .B1(_0785_));
 sg13g2_buf_1 _5675_ (.A(_4274_),
    .X(_0786_));
 sg13g2_a21oi_1 _5676_ (.A1(_0781_),
    .A2(net68),
    .Y(_0787_),
    .B1(_0783_));
 sg13g2_nand2_1 _5677_ (.Y(_0788_),
    .A(_4274_),
    .B(_4273_));
 sg13g2_buf_1 _5678_ (.A(_0788_),
    .X(_0789_));
 sg13g2_nor2_1 _5679_ (.A(_4274_),
    .B(_4273_),
    .Y(_0790_));
 sg13g2_buf_1 _5680_ (.A(_0790_),
    .X(_0791_));
 sg13g2_inv_1 _5681_ (.Y(_0792_),
    .A(_0791_));
 sg13g2_buf_1 _5682_ (.A(_0792_),
    .X(_0793_));
 sg13g2_nand3_1 _5683_ (.B(_0789_),
    .C(net43),
    .A(_0780_),
    .Y(_0794_));
 sg13g2_nand2_1 _5684_ (.Y(_0079_),
    .A(_0787_),
    .B(_0794_));
 sg13g2_inv_1 _5685_ (.Y(_0795_),
    .A(_0782_));
 sg13g2_buf_1 _5686_ (.A(_0795_),
    .X(_0796_));
 sg13g2_buf_1 _5687_ (.A(net61),
    .X(_0797_));
 sg13g2_nor2_1 _5688_ (.A(net50),
    .B(_4343_),
    .Y(_0080_));
 sg13g2_nor2b_1 _5689_ (.A(net50),
    .B_N(_4308_),
    .Y(_0081_));
 sg13g2_nor2b_1 _5690_ (.A(net50),
    .B_N(_4318_),
    .Y(_0082_));
 sg13g2_nor2b_1 _5691_ (.A(_0797_),
    .B_N(_4325_),
    .Y(_0083_));
 sg13g2_buf_1 _5692_ (.A(net61),
    .X(_0798_));
 sg13g2_nor2_1 _5693_ (.A(net49),
    .B(_4332_),
    .Y(_0084_));
 sg13g2_nor2b_1 _5694_ (.A(_0797_),
    .B_N(_4338_),
    .Y(_0085_));
 sg13g2_buf_1 _5695_ (.A(_0795_),
    .X(_0799_));
 sg13g2_nor3_1 _5696_ (.A(net60),
    .B(_4347_),
    .C(_4348_),
    .Y(_0086_));
 sg13g2_nor2b_1 _5697_ (.A(net50),
    .B_N(_4354_),
    .Y(_0087_));
 sg13g2_nor3_1 _5698_ (.A(net60),
    .B(_4292_),
    .C(_4358_),
    .Y(_0088_));
 sg13g2_nor2_1 _5699_ (.A(net49),
    .B(_4363_),
    .Y(_0089_));
 sg13g2_nor2b_1 _5700_ (.A(net50),
    .B_N(_4370_),
    .Y(_0090_));
 sg13g2_nor2b_1 _5701_ (.A(net50),
    .B_N(_4377_),
    .Y(_0091_));
 sg13g2_buf_1 _5702_ (.A(_0782_),
    .X(_0800_));
 sg13g2_buf_1 _5703_ (.A(net67),
    .X(_0801_));
 sg13g2_and3_1 _5704_ (.X(_0092_),
    .A(_4385_),
    .B(_4295_),
    .C(net59));
 sg13g2_nor2_1 _5705_ (.A(net49),
    .B(_4389_),
    .Y(_0093_));
 sg13g2_nor2b_1 _5706_ (.A(net50),
    .B_N(_4298_),
    .Y(_0094_));
 sg13g2_nor2_1 _5707_ (.A(_0798_),
    .B(_0411_),
    .Y(_0095_));
 sg13g2_inv_1 _5708_ (.Y(_0802_),
    .A(_0789_));
 sg13g2_a21oi_1 _5709_ (.A1(_0780_),
    .A2(_0802_),
    .Y(_0803_),
    .B1(_4325_));
 sg13g2_o21ai_1 _5710_ (.B1(net59),
    .Y(_0804_),
    .A1(_0000_),
    .A2(_0803_));
 sg13g2_a21oi_1 _5711_ (.A1(_4155_),
    .A2(_0803_),
    .Y(_0096_),
    .B1(_0804_));
 sg13g2_nand3_1 _5712_ (.B(_0349_),
    .C(_0350_),
    .A(_0348_),
    .Y(_0805_));
 sg13g2_nor4_1 _5713_ (.A(_0341_),
    .B(\main.demo.vga._q_xcount[6] ),
    .C(_0346_),
    .D(_0805_),
    .Y(_0806_));
 sg13g2_a22oi_1 _5714_ (.Y(_0807_),
    .B1(\main.demo.vga._q_active_h ),
    .B2(_0395_),
    .A2(_0391_),
    .A1(_0806_));
 sg13g2_buf_1 _5715_ (.A(_0807_),
    .X(_0808_));
 sg13g2_buf_1 _5716_ (.A(_0808_),
    .X(_0809_));
 sg13g2_nor2_1 _5717_ (.A(_0798_),
    .B(net33),
    .Y(_0122_));
 sg13g2_nor2_1 _5718_ (.A(net49),
    .B(net40),
    .Y(_0123_));
 sg13g2_nor2b_1 _5719_ (.A(_0808_),
    .B_N(\main.demo.vga._q_xcount[0] ),
    .Y(_0126_));
 sg13g2_nor2_1 _5720_ (.A(_0350_),
    .B(net33),
    .Y(_0127_));
 sg13g2_nor2b_1 _5721_ (.A(_0808_),
    .B_N(\main.demo.vga._q_xcount[1] ),
    .Y(_0128_));
 sg13g2_nor2_1 _5722_ (.A(_0336_),
    .B(net33),
    .Y(_0129_));
 sg13g2_nor2_1 _5723_ (.A(_0356_),
    .B(_0809_),
    .Y(_0130_));
 sg13g2_nor2_1 _5724_ (.A(_0400_),
    .B(_0809_),
    .Y(_0131_));
 sg13g2_nor2b_1 _5725_ (.A(_0808_),
    .B_N(_0344_),
    .Y(_0132_));
 sg13g2_nor2_1 _5726_ (.A(_0343_),
    .B(net33),
    .Y(_0133_));
 sg13g2_nor2_1 _5727_ (.A(_0342_),
    .B(net33),
    .Y(_0134_));
 sg13g2_nor2_1 _5728_ (.A(_0349_),
    .B(net33),
    .Y(_0135_));
 sg13g2_nor2_1 _5729_ (.A(_0348_),
    .B(net33),
    .Y(_0136_));
 sg13g2_nor2_1 _5730_ (.A(\main.demo.vga._q_xcount[0] ),
    .B(net50),
    .Y(_0147_));
 sg13g2_nand4_1 _5731_ (.B(_0345_),
    .C(_0392_),
    .A(_0391_),
    .Y(_0810_),
    .D(_0393_));
 sg13g2_inv_1 _5732_ (.Y(_0811_),
    .A(_0810_));
 sg13g2_nor3_1 _5733_ (.A(_0348_),
    .B(_0349_),
    .C(_0404_),
    .Y(_0812_));
 sg13g2_nor2_1 _5734_ (.A(_0350_),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_nor2_1 _5735_ (.A(_0811_),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_nand2_1 _5736_ (.Y(_0815_),
    .A(_0812_),
    .B(_0350_));
 sg13g2_buf_1 _5737_ (.A(_0795_),
    .X(_0816_));
 sg13g2_a21oi_1 _5738_ (.A1(_0814_),
    .A2(_0815_),
    .Y(_0148_),
    .B1(net58));
 sg13g2_xnor2_1 _5739_ (.Y(_0817_),
    .A(_0344_),
    .B(_0401_));
 sg13g2_a21oi_1 _5740_ (.A1(_0817_),
    .A2(_0395_),
    .Y(_0153_),
    .B1(net58));
 sg13g2_o21ai_1 _5741_ (.B1(_0343_),
    .Y(_0818_),
    .A1(_0354_),
    .A2(_0339_));
 sg13g2_nand2b_1 _5742_ (.Y(_0819_),
    .B(_0818_),
    .A_N(_0402_));
 sg13g2_a21oi_1 _5743_ (.A1(_0819_),
    .A2(_0395_),
    .Y(_0154_),
    .B1(_0816_));
 sg13g2_xnor2_1 _5744_ (.Y(_0820_),
    .A(_0349_),
    .B(_0404_));
 sg13g2_a21oi_1 _5745_ (.A1(_0820_),
    .A2(_0395_),
    .Y(_0156_),
    .B1(_0816_));
 sg13g2_a21oi_1 _5746_ (.A1(_0405_),
    .A2(\main.demo.vga._q_xcount[8] ),
    .Y(_0821_),
    .B1(\main.demo.vga._q_xcount[9] ));
 sg13g2_nor3_1 _5747_ (.A(net60),
    .B(_0812_),
    .C(_0821_),
    .Y(_0157_));
 sg13g2_nand4_1 _5748_ (.B(_0349_),
    .C(_0350_),
    .A(_0343_),
    .Y(_0822_),
    .D(\main.demo.vga._q_xcount[9] ));
 sg13g2_nor4_1 _5749_ (.A(_0342_),
    .B(_0346_),
    .C(_0357_),
    .D(_0822_),
    .Y(_0823_));
 sg13g2_inv_1 _5750_ (.Y(_0824_),
    .A(_0823_));
 sg13g2_nor2_1 _5751_ (.A(_0378_),
    .B(_0824_),
    .Y(_0825_));
 sg13g2_nor2_1 _5752_ (.A(_0360_),
    .B(_0823_),
    .Y(_0826_));
 sg13g2_nor2_1 _5753_ (.A(_0383_),
    .B(_0824_),
    .Y(_0827_));
 sg13g2_nor2_1 _5754_ (.A(_0795_),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_inv_1 _5755_ (.Y(_0829_),
    .A(_0828_));
 sg13g2_nor3_1 _5756_ (.A(_0825_),
    .B(_0826_),
    .C(_0829_),
    .Y(_0158_));
 sg13g2_nor3_2 _5757_ (.A(_0359_),
    .B(_0378_),
    .C(_0824_),
    .Y(_0830_));
 sg13g2_nor2_1 _5758_ (.A(\main.demo.vga._q_ycount[1] ),
    .B(_0825_),
    .Y(_0831_));
 sg13g2_nor3_1 _5759_ (.A(net61),
    .B(_0830_),
    .C(_0831_),
    .Y(_0159_));
 sg13g2_xnor2_1 _5760_ (.Y(_0832_),
    .A(_0366_),
    .B(_0830_));
 sg13g2_inv_1 _5761_ (.Y(_0833_),
    .A(_0827_));
 sg13g2_a21oi_1 _5762_ (.A1(_0832_),
    .A2(_0833_),
    .Y(_0160_),
    .B1(net58));
 sg13g2_nand2_1 _5763_ (.Y(_0834_),
    .A(_0830_),
    .B(_0368_));
 sg13g2_inv_1 _5764_ (.Y(_0835_),
    .A(_0834_));
 sg13g2_a21oi_1 _5765_ (.A1(_0830_),
    .A2(_0366_),
    .Y(_0836_),
    .B1(\main.demo.vga._q_ycount[3] ));
 sg13g2_nor3_1 _5766_ (.A(_0829_),
    .B(_0835_),
    .C(_0836_),
    .Y(_0161_));
 sg13g2_xnor2_1 _5767_ (.Y(_0837_),
    .A(_0370_),
    .B(_0834_));
 sg13g2_a21oi_1 _5768_ (.A1(_0837_),
    .A2(_0833_),
    .Y(_0162_),
    .B1(net58));
 sg13g2_nor3_1 _5769_ (.A(_0359_),
    .B(_0378_),
    .C(_0367_),
    .Y(_0838_));
 sg13g2_nand4_1 _5770_ (.B(_0362_),
    .C(_0369_),
    .A(_0811_),
    .Y(_0839_),
    .D(_0838_));
 sg13g2_inv_1 _5771_ (.Y(_0840_),
    .A(_0839_));
 sg13g2_a21oi_1 _5772_ (.A1(_0835_),
    .A2(_0369_),
    .Y(_0841_),
    .B1(_0362_));
 sg13g2_nor3_1 _5773_ (.A(_0829_),
    .B(_0840_),
    .C(_0841_),
    .Y(_0163_));
 sg13g2_nor2_1 _5774_ (.A(_0388_),
    .B(_0839_),
    .Y(_0842_));
 sg13g2_nor2_1 _5775_ (.A(\main.demo.vga._q_ycount[6] ),
    .B(_0840_),
    .Y(_0843_));
 sg13g2_nor3_1 _5776_ (.A(net61),
    .B(_0842_),
    .C(_0843_),
    .Y(_0164_));
 sg13g2_nor3_1 _5777_ (.A(_0389_),
    .B(_0388_),
    .C(_0839_),
    .Y(_0844_));
 sg13g2_nor2_1 _5778_ (.A(\main.demo.vga._q_ycount[7] ),
    .B(_0842_),
    .Y(_0845_));
 sg13g2_nor3_1 _5779_ (.A(net61),
    .B(_0844_),
    .C(_0845_),
    .Y(_0165_));
 sg13g2_nand4_1 _5780_ (.B(_0362_),
    .C(_0372_),
    .A(_0811_),
    .Y(_0846_),
    .D(_0838_));
 sg13g2_xnor2_1 _5781_ (.Y(_0847_),
    .A(_0363_),
    .B(_0846_));
 sg13g2_nor2_1 _5782_ (.A(net49),
    .B(_0847_),
    .Y(_0166_));
 sg13g2_nand2_1 _5783_ (.Y(_0848_),
    .A(_0844_),
    .B(\main.demo.vga._q_ycount[8] ));
 sg13g2_xnor2_1 _5784_ (.Y(_0849_),
    .A(_0364_),
    .B(_0848_));
 sg13g2_nand4_1 _5785_ (.B(_0379_),
    .C(_0380_),
    .A(_0811_),
    .Y(_0850_),
    .D(_0382_));
 sg13g2_a21oi_1 _5786_ (.A1(_0849_),
    .A2(_0850_),
    .Y(_0167_),
    .B1(net60));
 sg13g2_nor2b_1 _5787_ (.A(net28),
    .B_N(_0066_),
    .Y(_0168_));
 sg13g2_nand2_1 _5788_ (.Y(_0851_),
    .A(\main.demo.zic._q_clock_count[1] ),
    .B(\main.demo.zic._q_clock_count[0] ));
 sg13g2_inv_1 _5789_ (.Y(_0852_),
    .A(_0851_));
 sg13g2_nor3_1 _5790_ (.A(_4401_),
    .B(_0852_),
    .C(net28),
    .Y(_0169_));
 sg13g2_nor2b_1 _5791_ (.A(_0851_),
    .B_N(_4403_),
    .Y(_0853_));
 sg13g2_nor2_1 _5792_ (.A(_4403_),
    .B(_0852_),
    .Y(_0854_));
 sg13g2_nor3_1 _5793_ (.A(_0853_),
    .B(_0854_),
    .C(net28),
    .Y(_0170_));
 sg13g2_nand2_1 _5794_ (.Y(_0855_),
    .A(_0853_),
    .B(_4402_));
 sg13g2_inv_1 _5795_ (.Y(_0856_),
    .A(_0855_));
 sg13g2_nor2_1 _5796_ (.A(_4402_),
    .B(_0853_),
    .Y(_0857_));
 sg13g2_nor3_1 _5797_ (.A(_0856_),
    .B(_0857_),
    .C(net28),
    .Y(_0171_));
 sg13g2_nor2_1 _5798_ (.A(_4406_),
    .B(_0856_),
    .Y(_0858_));
 sg13g2_nor2_1 _5799_ (.A(_4407_),
    .B(_0855_),
    .Y(_0859_));
 sg13g2_nor3_1 _5800_ (.A(_0858_),
    .B(_0859_),
    .C(net28),
    .Y(_0172_));
 sg13g2_nor2_1 _5801_ (.A(\main.demo.zic._q_clock_count[5] ),
    .B(_0859_),
    .Y(_0860_));
 sg13g2_nor3_1 _5802_ (.A(_4405_),
    .B(_4407_),
    .C(_0855_),
    .Y(_0861_));
 sg13g2_nor3_1 _5803_ (.A(_0860_),
    .B(_0861_),
    .C(net28),
    .Y(_0173_));
 sg13g2_nor2_1 _5804_ (.A(\main.demo.zic._q_clock_count[6] ),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_nand2_1 _5805_ (.Y(_0863_),
    .A(_0861_),
    .B(\main.demo.zic._q_clock_count[6] ));
 sg13g2_inv_1 _5806_ (.Y(_0864_),
    .A(_0863_));
 sg13g2_nor3_1 _5807_ (.A(_0862_),
    .B(_0864_),
    .C(net28),
    .Y(_0174_));
 sg13g2_nand2b_1 _5808_ (.Y(_0865_),
    .B(_0863_),
    .A_N(\main.demo.zic._q_clock_count[7] ));
 sg13g2_nand2_1 _5809_ (.Y(_0866_),
    .A(_0864_),
    .B(\main.demo.zic._q_clock_count[7] ));
 sg13g2_and3_1 _5810_ (.X(_0175_),
    .A(_0412_),
    .B(_0865_),
    .C(_0866_));
 sg13g2_xor2_1 _5811_ (.B(_0866_),
    .A(\main.demo.zic._q_clock_count[8] ),
    .X(_0867_));
 sg13g2_nor2_1 _5812_ (.A(_0867_),
    .B(_0413_),
    .Y(_0176_));
 sg13g2_a22oi_1 _5813_ (.Y(_0868_),
    .B1(_0045_),
    .B2(_0249_),
    .A2(net62),
    .A1(_4433_));
 sg13g2_nor2_1 _5814_ (.A(net49),
    .B(_0868_),
    .Y(_0181_));
 sg13g2_nor2_1 _5815_ (.A(net49),
    .B(_0265_),
    .Y(_0182_));
 sg13g2_nor2_1 _5816_ (.A(net49),
    .B(_0241_),
    .Y(_0183_));
 sg13g2_nor2_1 _5817_ (.A(net58),
    .B(_0251_),
    .Y(_0184_));
 sg13g2_nor2_1 _5818_ (.A(net58),
    .B(_4441_),
    .Y(_0185_));
 sg13g2_nor2_1 _5819_ (.A(net58),
    .B(_0236_),
    .Y(_0186_));
 sg13g2_nor2_1 _5820_ (.A(net58),
    .B(_0259_),
    .Y(_0187_));
 sg13g2_nor3_2 _5821_ (.A(_4430_),
    .B(_4443_),
    .C(_0246_),
    .Y(_0869_));
 sg13g2_inv_1 _5822_ (.Y(_0870_),
    .A(_0869_));
 sg13g2_nor2_1 _5823_ (.A(_4436_),
    .B(_0238_),
    .Y(_0871_));
 sg13g2_inv_1 _5824_ (.Y(_0872_),
    .A(_0871_));
 sg13g2_nor2_1 _5825_ (.A(_4435_),
    .B(_0872_),
    .Y(_0873_));
 sg13g2_nor2_1 _5826_ (.A(_4437_),
    .B(_0242_),
    .Y(_0874_));
 sg13g2_inv_1 _5827_ (.Y(_0875_),
    .A(_0874_));
 sg13g2_nor2_1 _5828_ (.A(_4435_),
    .B(_0875_),
    .Y(_0876_));
 sg13g2_inv_1 _5829_ (.Y(_0877_),
    .A(_0262_));
 sg13g2_nor2_1 _5830_ (.A(_0238_),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_nor2_1 _5831_ (.A(_4436_),
    .B(_4437_),
    .Y(_0879_));
 sg13g2_nor2_1 _5832_ (.A(_0877_),
    .B(_0875_),
    .Y(_0880_));
 sg13g2_a21oi_1 _5833_ (.A1(_0263_),
    .A2(_0879_),
    .Y(_0881_),
    .B1(_0880_));
 sg13g2_inv_1 _5834_ (.Y(_0882_),
    .A(_0881_));
 sg13g2_nor4_1 _5835_ (.A(_0873_),
    .B(_0876_),
    .C(_0878_),
    .D(_0882_),
    .Y(_0883_));
 sg13g2_nor2_1 _5836_ (.A(_0870_),
    .B(_0883_),
    .Y(_0884_));
 sg13g2_inv_1 _5837_ (.Y(_0885_),
    .A(_0879_));
 sg13g2_nor2_1 _5838_ (.A(_4435_),
    .B(_0885_),
    .Y(_0886_));
 sg13g2_inv_1 _5839_ (.Y(_0887_),
    .A(_4433_));
 sg13g2_nand2_1 _5840_ (.Y(_0888_),
    .A(_0887_),
    .B(_4432_));
 sg13g2_nor2_1 _5841_ (.A(_0888_),
    .B(_0872_),
    .Y(_0889_));
 sg13g2_nor2_1 _5842_ (.A(_0886_),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_inv_1 _5843_ (.Y(_0891_),
    .A(_0890_));
 sg13g2_a21oi_1 _5844_ (.A1(_4433_),
    .A2(_0874_),
    .Y(_0892_),
    .B1(_0891_));
 sg13g2_inv_1 _5845_ (.Y(_0893_),
    .A(_0892_));
 sg13g2_inv_1 _5846_ (.Y(_0894_),
    .A(_0248_));
 sg13g2_nor2_1 _5847_ (.A(_4438_),
    .B(_0888_),
    .Y(_0895_));
 sg13g2_inv_1 _5848_ (.Y(_0896_),
    .A(_0895_));
 sg13g2_a21oi_1 _5849_ (.A1(_0894_),
    .A2(_0253_),
    .Y(_0897_),
    .B1(_0896_));
 sg13g2_a21oi_1 _5850_ (.A1(_0893_),
    .A2(_0248_),
    .Y(_0898_),
    .B1(_0897_));
 sg13g2_nor2b_1 _5851_ (.A(_0255_),
    .B_N(_0878_),
    .Y(_0899_));
 sg13g2_nor2_1 _5852_ (.A(_4438_),
    .B(_0877_),
    .Y(_0900_));
 sg13g2_nor2_2 _5853_ (.A(_4430_),
    .B(_0253_),
    .Y(_0901_));
 sg13g2_nor2_1 _5854_ (.A(_4432_),
    .B(_0887_),
    .Y(_0902_));
 sg13g2_inv_1 _5855_ (.Y(_0903_),
    .A(_0902_));
 sg13g2_nor2_1 _5856_ (.A(_0903_),
    .B(_0872_),
    .Y(_0904_));
 sg13g2_nor2_1 _5857_ (.A(_0901_),
    .B(_0869_),
    .Y(_0905_));
 sg13g2_inv_1 _5858_ (.Y(_0906_),
    .A(_0905_));
 sg13g2_a22oi_1 _5859_ (.Y(_0907_),
    .B1(_0904_),
    .B2(_0906_),
    .A2(_0901_),
    .A1(_0900_));
 sg13g2_nor2b_1 _5860_ (.A(_0899_),
    .B_N(_0907_),
    .Y(_0908_));
 sg13g2_nand2_1 _5861_ (.Y(_0909_),
    .A(_0898_),
    .B(_0908_));
 sg13g2_nor2_1 _5862_ (.A(_0877_),
    .B(_0885_),
    .Y(_0910_));
 sg13g2_nor3_1 _5863_ (.A(_4439_),
    .B(_0910_),
    .C(_0893_),
    .Y(_0911_));
 sg13g2_a21oi_1 _5864_ (.A1(_0232_),
    .A2(\main.demo.zic._q_idx[6] ),
    .Y(_0912_),
    .B1(_0901_));
 sg13g2_inv_1 _5865_ (.Y(_0913_),
    .A(_0912_));
 sg13g2_nor2_1 _5866_ (.A(_0888_),
    .B(_0885_),
    .Y(_0914_));
 sg13g2_inv_1 _5867_ (.Y(_0915_),
    .A(_0873_));
 sg13g2_nand2_1 _5868_ (.Y(_0916_),
    .A(_0874_),
    .B(_0887_));
 sg13g2_nand3b_1 _5869_ (.B(_0915_),
    .C(_0916_),
    .Y(_0917_),
    .A_N(_0914_));
 sg13g2_a22oi_1 _5870_ (.Y(_0918_),
    .B1(_0248_),
    .B2(_0917_),
    .A2(_4439_),
    .A1(_0913_));
 sg13g2_o21ai_1 _5871_ (.B1(_0918_),
    .Y(_0919_),
    .A1(_0255_),
    .A2(_0911_));
 sg13g2_nor3_1 _5872_ (.A(_0884_),
    .B(_0909_),
    .C(_0919_),
    .Y(_0920_));
 sg13g2_inv_1 _5873_ (.Y(_0921_),
    .A(_0910_));
 sg13g2_nor2_1 _5874_ (.A(_4436_),
    .B(_4435_),
    .Y(_0922_));
 sg13g2_nor2_1 _5875_ (.A(_0903_),
    .B(_0875_),
    .Y(_0923_));
 sg13g2_nor2_1 _5876_ (.A(_0910_),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_inv_1 _5877_ (.Y(_0925_),
    .A(_0924_));
 sg13g2_o21ai_1 _5878_ (.B1(_0901_),
    .Y(_0926_),
    .A1(_0922_),
    .A2(_0925_));
 sg13g2_o21ai_1 _5879_ (.B1(_0926_),
    .Y(_0927_),
    .A1(_0894_),
    .A2(_0921_));
 sg13g2_nor2_1 _5880_ (.A(_0888_),
    .B(_0875_),
    .Y(_0928_));
 sg13g2_inv_1 _5881_ (.Y(_0929_),
    .A(_0928_));
 sg13g2_nor2_1 _5882_ (.A(_4438_),
    .B(_0903_),
    .Y(_0930_));
 sg13g2_inv_1 _5883_ (.Y(_0931_),
    .A(_0930_));
 sg13g2_a21oi_1 _5884_ (.A1(_0929_),
    .A2(_0931_),
    .Y(_0932_),
    .B1(_0905_));
 sg13g2_nor2_1 _5885_ (.A(_0877_),
    .B(_0872_),
    .Y(_0933_));
 sg13g2_o21ai_1 _5886_ (.B1(_0248_),
    .Y(_0934_),
    .A1(_0930_),
    .A2(_0933_));
 sg13g2_inv_1 _5887_ (.Y(_0935_),
    .A(_0934_));
 sg13g2_nor2_1 _5888_ (.A(_0238_),
    .B(_0903_),
    .Y(_0936_));
 sg13g2_inv_1 _5889_ (.Y(_0937_),
    .A(_0904_));
 sg13g2_nand2b_1 _5890_ (.Y(_0938_),
    .B(_0937_),
    .A_N(_0900_));
 sg13g2_a22oi_1 _5891_ (.Y(_0939_),
    .B1(_0248_),
    .B2(_0938_),
    .A2(_0936_),
    .A1(_0254_));
 sg13g2_inv_1 _5892_ (.Y(_0940_),
    .A(_0939_));
 sg13g2_nor2_1 _5893_ (.A(_0935_),
    .B(_0940_),
    .Y(_0941_));
 sg13g2_o21ai_1 _5894_ (.B1(_0941_),
    .Y(_0942_),
    .A1(_4443_),
    .A2(\main.demo.zic._q_idx[6] ));
 sg13g2_nor3_1 _5895_ (.A(_0927_),
    .B(_0932_),
    .C(_0942_),
    .Y(_0943_));
 sg13g2_inv_1 _5896_ (.Y(_0944_),
    .A(_0889_));
 sg13g2_inv_1 _5897_ (.Y(_0945_),
    .A(_0876_));
 sg13g2_nand2_1 _5898_ (.Y(_0946_),
    .A(_0944_),
    .B(_0945_));
 sg13g2_o21ai_1 _5899_ (.B1(_0901_),
    .Y(_0947_),
    .A1(_0946_),
    .A2(_0882_));
 sg13g2_o21ai_1 _5900_ (.B1(_0869_),
    .Y(_0948_),
    .A1(_0891_),
    .A2(_0925_));
 sg13g2_nand3_1 _5901_ (.B(_0902_),
    .C(_0879_),
    .A(_0248_),
    .Y(_0949_));
 sg13g2_nand3_1 _5902_ (.B(_0948_),
    .C(_0949_),
    .A(_0947_),
    .Y(_0950_));
 sg13g2_nand3_1 _5903_ (.B(_0915_),
    .C(_0929_),
    .A(_0881_),
    .Y(_0951_));
 sg13g2_a22oi_1 _5904_ (.Y(_0952_),
    .B1(_0254_),
    .B2(_0951_),
    .A2(_0895_),
    .A1(_0869_));
 sg13g2_nor2b_1 _5905_ (.A(_0950_),
    .B_N(_0952_),
    .Y(_0953_));
 sg13g2_nand3_1 _5906_ (.B(_0943_),
    .C(_0953_),
    .A(_0920_),
    .Y(_0954_));
 sg13g2_inv_1 _5907_ (.Y(_0955_),
    .A(_0898_));
 sg13g2_nor3_1 _5908_ (.A(_0940_),
    .B(_0955_),
    .C(_0950_),
    .Y(_0956_));
 sg13g2_nand3_1 _5909_ (.B(_0907_),
    .C(_0956_),
    .A(_0954_),
    .Y(_0957_));
 sg13g2_a21oi_1 _5910_ (.A1(_0957_),
    .A2(net38),
    .Y(_0958_),
    .B1(\main.demo.zic._q_qpos[0] ));
 sg13g2_and3_1 _5911_ (.X(_0959_),
    .A(_0957_),
    .B(\main.demo.zic._q_qpos[0] ),
    .C(net45));
 sg13g2_nor3_1 _5912_ (.A(net61),
    .B(_0958_),
    .C(_0959_),
    .Y(_0188_));
 sg13g2_nor3_1 _5913_ (.A(_0927_),
    .B(_0940_),
    .C(_0919_),
    .Y(_0960_));
 sg13g2_nand2_1 _5914_ (.Y(_0961_),
    .A(_0954_),
    .B(_0960_));
 sg13g2_nor2_1 _5915_ (.A(\main.demo.zic._q_qpos[4] ),
    .B(_0961_),
    .Y(_0962_));
 sg13g2_nand2_1 _5916_ (.Y(_0963_),
    .A(_0920_),
    .B(_0939_));
 sg13g2_xor2_1 _5917_ (.B(_0963_),
    .A(\main.demo.zic._q_qpos[1] ),
    .X(_0964_));
 sg13g2_inv_1 _5918_ (.Y(_0965_),
    .A(_0964_));
 sg13g2_nand2_1 _5919_ (.Y(_0966_),
    .A(_0957_),
    .B(\main.demo.zic._q_qpos[0] ));
 sg13g2_nand2_1 _5920_ (.Y(_0967_),
    .A(_0963_),
    .B(\main.demo.zic._q_qpos[1] ));
 sg13g2_o21ai_1 _5921_ (.B1(_0967_),
    .Y(_0968_),
    .A1(_0965_),
    .A2(_0966_));
 sg13g2_inv_1 _5922_ (.Y(_0969_),
    .A(_0968_));
 sg13g2_inv_1 _5923_ (.Y(_0970_),
    .A(_0919_));
 sg13g2_o21ai_1 _5924_ (.B1(_0878_),
    .Y(_0971_),
    .A1(_0254_),
    .A2(_0869_));
 sg13g2_nand4_1 _5925_ (.B(_0952_),
    .C(_0941_),
    .A(_0970_),
    .Y(_0972_),
    .D(_0971_));
 sg13g2_nand2_1 _5926_ (.Y(_0973_),
    .A(_0972_),
    .B(\main.demo.zic._q_qpos[2] ));
 sg13g2_nor2_1 _5927_ (.A(\main.demo.zic._q_qpos[2] ),
    .B(_0972_),
    .Y(_0974_));
 sg13g2_a21oi_1 _5928_ (.A1(_0969_),
    .A2(_0973_),
    .Y(_0975_),
    .B1(_0974_));
 sg13g2_inv_1 _5929_ (.Y(_0976_),
    .A(_0975_));
 sg13g2_nor2_1 _5930_ (.A(_0899_),
    .B(_0935_),
    .Y(_0977_));
 sg13g2_nand3_1 _5931_ (.B(_0898_),
    .C(_0977_),
    .A(_0952_),
    .Y(_0978_));
 sg13g2_nand2_1 _5932_ (.Y(_0979_),
    .A(_0978_),
    .B(\main.demo.zic._q_qpos[3] ));
 sg13g2_nor2_1 _5933_ (.A(\main.demo.zic._q_qpos[3] ),
    .B(_0978_),
    .Y(_0980_));
 sg13g2_a21oi_1 _5934_ (.A1(_0976_),
    .A2(_0979_),
    .Y(_0981_),
    .B1(_0980_));
 sg13g2_inv_1 _5935_ (.Y(_0982_),
    .A(_0981_));
 sg13g2_nand2_1 _5936_ (.Y(_0983_),
    .A(_0961_),
    .B(\main.demo.zic._q_qpos[4] ));
 sg13g2_o21ai_1 _5937_ (.B1(_0983_),
    .Y(_0984_),
    .A1(_0962_),
    .A2(_0982_));
 sg13g2_nand2_1 _5938_ (.Y(_0985_),
    .A(_0953_),
    .B(_0908_));
 sg13g2_nor2_1 _5939_ (.A(\main.demo.zic._q_qpos[5] ),
    .B(_0985_),
    .Y(_0986_));
 sg13g2_inv_1 _5940_ (.Y(_0987_),
    .A(_0986_));
 sg13g2_nand2_1 _5941_ (.Y(_0988_),
    .A(_0985_),
    .B(\main.demo.zic._q_qpos[5] ));
 sg13g2_inv_1 _5942_ (.Y(_0989_),
    .A(_0988_));
 sg13g2_a21o_1 _5943_ (.A2(_0987_),
    .A1(_0984_),
    .B1(_0989_),
    .X(_0990_));
 sg13g2_xor2_1 _5944_ (.B(_0884_),
    .A(\main.demo.zic._q_qpos[6] ),
    .X(_0991_));
 sg13g2_nand2_1 _5945_ (.Y(_0992_),
    .A(_0884_),
    .B(\main.demo.zic._q_qpos[6] ));
 sg13g2_inv_1 _5946_ (.Y(_0993_),
    .A(_0992_));
 sg13g2_a21oi_1 _5947_ (.A1(_0990_),
    .A2(_0991_),
    .Y(_0994_),
    .B1(_0993_));
 sg13g2_nor3_1 _5948_ (.A(_0043_),
    .B(_0406_),
    .C(_0994_),
    .Y(_0995_));
 sg13g2_nand2_1 _5949_ (.Y(_0996_),
    .A(_0995_),
    .B(\main.demo.zic._q_qpos[8] ));
 sg13g2_inv_1 _5950_ (.Y(_0997_),
    .A(_0996_));
 sg13g2_buf_1 _5951_ (.A(\main.demo.zic._q_qpos[9] ),
    .X(_0998_));
 sg13g2_a21oi_1 _5952_ (.A1(_0997_),
    .A2(_0998_),
    .Y(_0999_),
    .B1(\main.demo.zic._q_qpos[10] ));
 sg13g2_and3_1 _5953_ (.X(_1000_),
    .A(_0997_),
    .B(_0998_),
    .C(\main.demo.zic._q_qpos[10] ));
 sg13g2_nor3_1 _5954_ (.A(_0796_),
    .B(_0999_),
    .C(_1000_),
    .Y(_0189_));
 sg13g2_inv_1 _5955_ (.Y(_1001_),
    .A(\main.demo.zic._q_qpos[11] ));
 sg13g2_inv_1 _5956_ (.Y(_1002_),
    .A(_0994_));
 sg13g2_nand4_1 _5957_ (.B(\main.demo.zic._q_qpos[8] ),
    .C(\main.demo.zic._q_qpos[7] ),
    .A(_1002_),
    .Y(_1003_),
    .D(net45));
 sg13g2_nand3b_1 _5958_ (.B(_0998_),
    .C(\main.demo.zic._q_qpos[10] ),
    .Y(_1004_),
    .A_N(_1003_));
 sg13g2_o21ai_1 _5959_ (.B1(net59),
    .Y(_1005_),
    .A1(_1001_),
    .A2(_1004_));
 sg13g2_a21oi_1 _5960_ (.A1(_1001_),
    .A2(_1004_),
    .Y(_0190_),
    .B1(_1005_));
 sg13g2_inv_2 _5961_ (.Y(_1006_),
    .A(\main.demo.zic._q_qpos[12] ));
 sg13g2_nand4_1 _5962_ (.B(_0998_),
    .C(\main.demo.zic._q_qpos[10] ),
    .A(\main.demo.zic._q_qpos[8] ),
    .Y(_1007_),
    .D(\main.demo.zic._q_qpos[11] ));
 sg13g2_nand2b_1 _5963_ (.Y(_1008_),
    .B(_0995_),
    .A_N(_1007_));
 sg13g2_o21ai_1 _5964_ (.B1(_0801_),
    .Y(_1009_),
    .A1(_1006_),
    .A2(_1008_));
 sg13g2_a21oi_1 _5965_ (.A1(_1006_),
    .A2(_1008_),
    .Y(_0191_),
    .B1(_1009_));
 sg13g2_xnor2_1 _5966_ (.Y(_1010_),
    .A(_0965_),
    .B(_0966_));
 sg13g2_buf_1 _5967_ (.A(net45),
    .X(_1011_));
 sg13g2_o21ai_1 _5968_ (.B1(net59),
    .Y(_1012_),
    .A1(\main.demo.zic._q_qpos[1] ),
    .A2(net39));
 sg13g2_a21oi_1 _5969_ (.A1(_1010_),
    .A2(net37),
    .Y(_0192_),
    .B1(_1012_));
 sg13g2_nor2b_1 _5970_ (.A(_0974_),
    .B_N(_0973_),
    .Y(_1013_));
 sg13g2_xnor2_1 _5971_ (.Y(_1014_),
    .A(_1013_),
    .B(_0968_));
 sg13g2_o21ai_1 _5972_ (.B1(net59),
    .Y(_1015_),
    .A1(\main.demo.zic._q_qpos[2] ),
    .A2(net39));
 sg13g2_a21oi_1 _5973_ (.A1(_1014_),
    .A2(net37),
    .Y(_0193_),
    .B1(_1015_));
 sg13g2_nor2b_1 _5974_ (.A(_0980_),
    .B_N(_0979_),
    .Y(_1016_));
 sg13g2_xnor2_1 _5975_ (.Y(_1017_),
    .A(_1016_),
    .B(_0975_));
 sg13g2_o21ai_1 _5976_ (.B1(net59),
    .Y(_1018_),
    .A1(\main.demo.zic._q_qpos[3] ),
    .A2(net39));
 sg13g2_a21oi_1 _5977_ (.A1(_1017_),
    .A2(net37),
    .Y(_0194_),
    .B1(_1018_));
 sg13g2_nor2b_1 _5978_ (.A(_0962_),
    .B_N(_0983_),
    .Y(_1019_));
 sg13g2_xnor2_1 _5979_ (.Y(_1020_),
    .A(_1019_),
    .B(_0981_));
 sg13g2_o21ai_1 _5980_ (.B1(net59),
    .Y(_1021_),
    .A1(\main.demo.zic._q_qpos[4] ),
    .A2(net39));
 sg13g2_a21oi_1 _5981_ (.A1(_1020_),
    .A2(net37),
    .Y(_0195_),
    .B1(_1021_));
 sg13g2_nor2_1 _5982_ (.A(_0986_),
    .B(_0989_),
    .Y(_1022_));
 sg13g2_xnor2_1 _5983_ (.Y(_1023_),
    .A(_1022_),
    .B(_0984_));
 sg13g2_o21ai_1 _5984_ (.B1(net59),
    .Y(_1024_),
    .A1(\main.demo.zic._q_qpos[5] ),
    .A2(net39));
 sg13g2_a21oi_1 _5985_ (.A1(_1023_),
    .A2(net37),
    .Y(_0196_),
    .B1(_1024_));
 sg13g2_xnor2_1 _5986_ (.Y(_1025_),
    .A(_0991_),
    .B(_0990_));
 sg13g2_o21ai_1 _5987_ (.B1(net67),
    .Y(_1026_),
    .A1(\main.demo.zic._q_qpos[6] ),
    .A2(net39));
 sg13g2_a21oi_1 _5988_ (.A1(_1025_),
    .A2(net37),
    .Y(_0197_),
    .B1(_1026_));
 sg13g2_xnor2_1 _5989_ (.Y(_1027_),
    .A(_0043_),
    .B(_0994_));
 sg13g2_o21ai_1 _5990_ (.B1(net67),
    .Y(_1028_),
    .A1(\main.demo.zic._q_qpos[7] ),
    .A2(net38));
 sg13g2_a21oi_1 _5991_ (.A1(_1027_),
    .A2(net37),
    .Y(_0198_),
    .B1(_1028_));
 sg13g2_nor2_1 _5992_ (.A(\main.demo.zic._q_qpos[8] ),
    .B(_0995_),
    .Y(_1029_));
 sg13g2_nor3_1 _5993_ (.A(_0796_),
    .B(_1029_),
    .C(_0997_),
    .Y(_0199_));
 sg13g2_inv_1 _5994_ (.Y(_1030_),
    .A(_0998_));
 sg13g2_nor2_1 _5995_ (.A(_1030_),
    .B(_1003_),
    .Y(_1031_));
 sg13g2_a21oi_1 _5996_ (.A1(_1003_),
    .A2(_1030_),
    .Y(_1032_),
    .B1(_0795_));
 sg13g2_nor2b_1 _5997_ (.A(_1031_),
    .B_N(_1032_),
    .Y(_0200_));
 sg13g2_inv_1 _5998_ (.Y(_1033_),
    .A(_0251_));
 sg13g2_nand4_1 _5999_ (.B(_0266_),
    .C(_0868_),
    .A(_1033_),
    .Y(_1034_),
    .D(_0241_));
 sg13g2_nand3b_1 _6000_ (.B(_0252_),
    .C(_0265_),
    .Y(_1035_),
    .A_N(_0868_));
 sg13g2_a22oi_1 _6001_ (.Y(_1036_),
    .B1(_0271_),
    .B2(_0269_),
    .A2(_1035_),
    .A1(_1034_));
 sg13g2_a21oi_1 _6002_ (.A1(_0259_),
    .A2(_0236_),
    .Y(_1037_),
    .B1(_1036_));
 sg13g2_nand2_2 _6003_ (.Y(_1038_),
    .A(_1037_),
    .B(net52));
 sg13g2_buf_1 _6004_ (.A(\main.demo.zic._q_squ_env[4] ),
    .X(_1039_));
 sg13g2_nor2_1 _6005_ (.A(\main.demo.zic._q_squ_env[5] ),
    .B(_1039_),
    .Y(_1040_));
 sg13g2_buf_2 _6006_ (.A(\main.demo.zic._q_squ_env[3] ),
    .X(_1041_));
 sg13g2_nor2_1 _6007_ (.A(\main.demo.zic._q_squ_env[0] ),
    .B(\main.demo.zic._q_squ_env[1] ),
    .Y(_1042_));
 sg13g2_nand2b_1 _6008_ (.Y(_1043_),
    .B(_1042_),
    .A_N(\main.demo.zic._q_squ_env[2] ));
 sg13g2_nor2_1 _6009_ (.A(_1041_),
    .B(_1043_),
    .Y(_1044_));
 sg13g2_a21oi_1 _6010_ (.A1(_1040_),
    .A2(_1044_),
    .Y(_1045_),
    .B1(net52));
 sg13g2_inv_1 _6011_ (.Y(_1046_),
    .A(_1045_));
 sg13g2_nor2_2 _6012_ (.A(_1046_),
    .B(_4412_),
    .Y(_1047_));
 sg13g2_inv_1 _6013_ (.Y(_1048_),
    .A(net29));
 sg13g2_nand2_1 _6014_ (.Y(_1049_),
    .A(_1048_),
    .B(\main.demo.zic._q_squ_env[0] ));
 sg13g2_o21ai_1 _6015_ (.B1(_1049_),
    .Y(_1050_),
    .A1(\main.demo.zic._q_squ_env[0] ),
    .A2(_1047_));
 sg13g2_a21oi_1 _6016_ (.A1(_1038_),
    .A2(_1050_),
    .Y(_0214_),
    .B1(net60));
 sg13g2_nand2b_1 _6017_ (.Y(_1051_),
    .B(_1048_),
    .A_N(\main.demo.zic._q_squ_env[0] ));
 sg13g2_nor2b_1 _6018_ (.A(net29),
    .B_N(_1042_),
    .Y(_1052_));
 sg13g2_a21o_1 _6019_ (.A2(\main.demo.zic._q_squ_env[1] ),
    .A1(_1051_),
    .B1(_1052_),
    .X(_1053_));
 sg13g2_o21ai_1 _6020_ (.B1(_1053_),
    .Y(_1054_),
    .A1(net29),
    .A2(_1045_));
 sg13g2_a21oi_1 _6021_ (.A1(_1038_),
    .A2(_1054_),
    .Y(_0215_),
    .B1(net60));
 sg13g2_a22oi_1 _6022_ (.Y(_1055_),
    .B1(\main.demo.zic._q_squ_env[2] ),
    .B2(_1052_),
    .A2(_1046_),
    .A1(_1048_));
 sg13g2_o21ai_1 _6023_ (.B1(_1055_),
    .Y(_1056_),
    .A1(\main.demo.zic._q_squ_env[2] ),
    .A2(_1052_));
 sg13g2_a21oi_1 _6024_ (.A1(_1038_),
    .A2(_1056_),
    .Y(_0216_),
    .B1(net60));
 sg13g2_xor2_1 _6025_ (.B(_1043_),
    .A(_0038_),
    .X(_1057_));
 sg13g2_a22oi_1 _6026_ (.Y(_1058_),
    .B1(_1041_),
    .B2(net29),
    .A2(_1057_),
    .A1(_1047_));
 sg13g2_a21oi_1 _6027_ (.A1(_1038_),
    .A2(_1058_),
    .Y(_0217_),
    .B1(net60));
 sg13g2_xnor2_1 _6028_ (.Y(_1059_),
    .A(_0039_),
    .B(_1044_));
 sg13g2_a22oi_1 _6029_ (.Y(_1060_),
    .B1(_1039_),
    .B2(_0288_),
    .A2(_1059_),
    .A1(_1047_));
 sg13g2_a21oi_1 _6030_ (.A1(_1038_),
    .A2(_1060_),
    .Y(_0218_),
    .B1(_0799_));
 sg13g2_nor3_1 _6031_ (.A(_1041_),
    .B(_1039_),
    .C(_1043_),
    .Y(_1061_));
 sg13g2_xnor2_1 _6032_ (.Y(_1062_),
    .A(_0040_),
    .B(_1061_));
 sg13g2_a22oi_1 _6033_ (.Y(_1063_),
    .B1(\main.demo.zic._q_squ_env[5] ),
    .B2(_0288_),
    .A2(_1062_),
    .A1(_1047_));
 sg13g2_a21oi_1 _6034_ (.A1(_1038_),
    .A2(_1063_),
    .Y(_0219_),
    .B1(_0799_));
 sg13g2_xor2_1 _6035_ (.B(\main.demo.zic._q_tpos[0] ),
    .A(\main.demo.zic._q_drum_inc[0] ),
    .X(_1064_));
 sg13g2_nand2_1 _6036_ (.Y(_1065_),
    .A(_4430_),
    .B(_0055_));
 sg13g2_inv_1 _6037_ (.Y(_1066_),
    .A(_1065_));
 sg13g2_a21oi_1 _6038_ (.A1(_0944_),
    .A2(_0233_),
    .Y(_1067_),
    .B1(_1066_));
 sg13g2_nand2b_1 _6039_ (.Y(_1068_),
    .B(_4431_),
    .A_N(_0055_));
 sg13g2_nand3_1 _6040_ (.B(_0945_),
    .C(_0931_),
    .A(_0915_),
    .Y(_1069_));
 sg13g2_a221oi_1 _6041_ (.B2(_1065_),
    .C1(_0914_),
    .B1(_1069_),
    .A1(_0933_),
    .Y(_1070_),
    .A2(_1068_));
 sg13g2_a221oi_1 _6042_ (.B2(_1068_),
    .C1(_0886_),
    .B1(_0880_),
    .A1(_0900_),
    .Y(_1071_),
    .A2(_1065_));
 sg13g2_nand2_1 _6043_ (.Y(_1072_),
    .A(_0924_),
    .B(_0896_));
 sg13g2_a221oi_1 _6044_ (.B2(_1065_),
    .C1(_1067_),
    .B1(_1072_),
    .A1(_0904_),
    .Y(_1073_),
    .A2(_1068_));
 sg13g2_buf_1 _6045_ (.A(_1073_),
    .X(_1074_));
 sg13g2_nand3_1 _6046_ (.B(_1071_),
    .C(_1074_),
    .A(_1070_),
    .Y(_1075_));
 sg13g2_nand3b_1 _6047_ (.B(_1075_),
    .C(_1071_),
    .Y(_1076_),
    .A_N(_1067_));
 sg13g2_xnor2_1 _6048_ (.Y(_1077_),
    .A(_1064_),
    .B(_1076_));
 sg13g2_o21ai_1 _6049_ (.B1(net67),
    .Y(_1078_),
    .A1(\main.demo.zic._q_tpos[0] ),
    .A2(net38));
 sg13g2_a21oi_1 _6050_ (.A1(_1077_),
    .A2(_1011_),
    .Y(_0220_),
    .B1(_1078_));
 sg13g2_buf_1 _6051_ (.A(\main.demo.zic._q_tpos[9] ),
    .X(_1079_));
 sg13g2_nand2_1 _6052_ (.Y(_1080_),
    .A(\main.demo.zic._q_tpos[10] ),
    .B(_1079_));
 sg13g2_inv_1 _6053_ (.Y(_1081_),
    .A(\main.demo.zic._q_tpos[6] ));
 sg13g2_and2_1 _6054_ (.A(_1075_),
    .B(_1070_),
    .X(_1082_));
 sg13g2_xor2_1 _6055_ (.B(\main.demo.zic._q_tpos[1] ),
    .A(_4416_),
    .X(_1083_));
 sg13g2_nor2b_1 _6056_ (.A(_1082_),
    .B_N(_1083_),
    .Y(_1084_));
 sg13g2_a21o_1 _6057_ (.A2(\main.demo.zic._q_tpos[1] ),
    .A1(_4416_),
    .B1(_1084_),
    .X(_1085_));
 sg13g2_xor2_1 _6058_ (.B(\main.demo.zic._q_tpos[2] ),
    .A(_4415_),
    .X(_1086_));
 sg13g2_xor2_1 _6059_ (.B(_1074_),
    .A(_1086_),
    .X(_1087_));
 sg13g2_inv_1 _6060_ (.Y(_1088_),
    .A(\main.demo.zic._q_tpos[0] ));
 sg13g2_nand2_1 _6061_ (.Y(_1089_),
    .A(_1076_),
    .B(_1064_));
 sg13g2_o21ai_1 _6062_ (.B1(_1089_),
    .Y(_1090_),
    .A1(_4426_),
    .A2(_1088_));
 sg13g2_xnor2_1 _6063_ (.Y(_1091_),
    .A(_1083_),
    .B(_1082_));
 sg13g2_nand2_1 _6064_ (.Y(_1092_),
    .A(_1090_),
    .B(_1091_));
 sg13g2_xor2_1 _6065_ (.B(_1085_),
    .A(_1087_),
    .X(_1093_));
 sg13g2_nor2b_1 _6066_ (.A(_1092_),
    .B_N(_1093_),
    .Y(_1094_));
 sg13g2_a21o_1 _6067_ (.A2(_1087_),
    .A1(_1085_),
    .B1(_1094_),
    .X(_1095_));
 sg13g2_xor2_1 _6068_ (.B(\main.demo.zic._q_tpos[3] ),
    .A(_4414_),
    .X(_1096_));
 sg13g2_inv_1 _6069_ (.Y(_1097_),
    .A(_1096_));
 sg13g2_xnor2_1 _6070_ (.Y(_1098_),
    .A(_1097_),
    .B(_1074_));
 sg13g2_inv_1 _6071_ (.Y(_1099_),
    .A(\main.demo.zic._q_tpos[2] ));
 sg13g2_nand2_1 _6072_ (.Y(_1100_),
    .A(_1074_),
    .B(_1086_));
 sg13g2_o21ai_1 _6073_ (.B1(_1100_),
    .Y(_1101_),
    .A1(_0290_),
    .A2(_1099_));
 sg13g2_xnor2_1 _6074_ (.Y(_1102_),
    .A(_1098_),
    .B(_1101_));
 sg13g2_nor2b_1 _6075_ (.A(_1098_),
    .B_N(_1101_),
    .Y(_1103_));
 sg13g2_a21o_1 _6076_ (.A2(_1102_),
    .A1(_1095_),
    .B1(_1103_),
    .X(_1104_));
 sg13g2_inv_1 _6077_ (.Y(_1105_),
    .A(\main.demo.zic._q_tpos[4] ));
 sg13g2_nand2_1 _6078_ (.Y(_1106_),
    .A(_4414_),
    .B(\main.demo.zic._q_tpos[3] ));
 sg13g2_o21ai_1 _6079_ (.B1(_1106_),
    .Y(_1107_),
    .A1(_1097_),
    .A2(_1074_));
 sg13g2_xnor2_1 _6080_ (.Y(_1108_),
    .A(_1105_),
    .B(_1107_));
 sg13g2_nand2_1 _6081_ (.Y(_1109_),
    .A(_1104_),
    .B(_1108_));
 sg13g2_nand2_1 _6082_ (.Y(_1110_),
    .A(_1107_),
    .B(\main.demo.zic._q_tpos[4] ));
 sg13g2_nand2_1 _6083_ (.Y(_1111_),
    .A(_1109_),
    .B(_1110_));
 sg13g2_inv_1 _6084_ (.Y(_1112_),
    .A(_1111_));
 sg13g2_nor2_1 _6085_ (.A(_0056_),
    .B(_1112_),
    .Y(_1113_));
 sg13g2_nand2_1 _6086_ (.Y(_1114_),
    .A(_1113_),
    .B(net45));
 sg13g2_nor2_1 _6087_ (.A(_1081_),
    .B(_1114_),
    .Y(_1115_));
 sg13g2_buf_1 _6088_ (.A(\main.demo.zic._q_tpos[7] ),
    .X(_1116_));
 sg13g2_nand2_1 _6089_ (.Y(_1117_),
    .A(\main.demo.zic._q_tpos[8] ),
    .B(_1116_));
 sg13g2_inv_1 _6090_ (.Y(_1118_),
    .A(_1117_));
 sg13g2_nand2_1 _6091_ (.Y(_1119_),
    .A(_1115_),
    .B(_1118_));
 sg13g2_o21ai_1 _6092_ (.B1(_0801_),
    .Y(_1120_),
    .A1(_1080_),
    .A2(_1119_));
 sg13g2_inv_1 _6093_ (.Y(_1121_),
    .A(_1119_));
 sg13g2_a21oi_1 _6094_ (.A1(_1121_),
    .A2(_1079_),
    .Y(_1122_),
    .B1(\main.demo.zic._q_tpos[10] ));
 sg13g2_nor2_1 _6095_ (.A(_1120_),
    .B(_1122_),
    .Y(_0221_));
 sg13g2_inv_1 _6096_ (.Y(_1123_),
    .A(_0042_));
 sg13g2_inv_1 _6097_ (.Y(_1124_),
    .A(\main.demo.zic._q_tpos[5] ));
 sg13g2_nor3_1 _6098_ (.A(_1081_),
    .B(_1124_),
    .C(_1112_),
    .Y(_1125_));
 sg13g2_inv_1 _6099_ (.Y(_1126_),
    .A(_1125_));
 sg13g2_nor3_1 _6100_ (.A(_1117_),
    .B(_1080_),
    .C(_1126_),
    .Y(_1127_));
 sg13g2_xnor2_1 _6101_ (.Y(_1128_),
    .A(_1123_),
    .B(_1127_));
 sg13g2_buf_1 _6102_ (.A(\main.demo.zic._q_tpos[11] ),
    .X(_1129_));
 sg13g2_o21ai_1 _6103_ (.B1(net67),
    .Y(_1130_),
    .A1(_1129_),
    .A2(net38));
 sg13g2_a21oi_1 _6104_ (.A1(_1128_),
    .A2(_1011_),
    .Y(_0222_),
    .B1(_1130_));
 sg13g2_xnor2_1 _6105_ (.Y(_1131_),
    .A(_1091_),
    .B(_1090_));
 sg13g2_o21ai_1 _6106_ (.B1(net67),
    .Y(_1132_),
    .A1(\main.demo.zic._q_tpos[1] ),
    .A2(net38));
 sg13g2_a21oi_1 _6107_ (.A1(_1131_),
    .A2(net37),
    .Y(_0223_),
    .B1(_1132_));
 sg13g2_xor2_1 _6108_ (.B(_1093_),
    .A(_1092_),
    .X(_1133_));
 sg13g2_o21ai_1 _6109_ (.B1(net67),
    .Y(_1134_),
    .A1(\main.demo.zic._q_tpos[2] ),
    .A2(net38));
 sg13g2_a21oi_1 _6110_ (.A1(_1133_),
    .A2(_0408_),
    .Y(_0224_),
    .B1(_1134_));
 sg13g2_xnor2_1 _6111_ (.Y(_1135_),
    .A(_1102_),
    .B(_1095_));
 sg13g2_o21ai_1 _6112_ (.B1(_0800_),
    .Y(_1136_),
    .A1(\main.demo.zic._q_tpos[3] ),
    .A2(_0436_));
 sg13g2_a21oi_1 _6113_ (.A1(_1135_),
    .A2(_0408_),
    .Y(_0225_),
    .B1(_1136_));
 sg13g2_xnor2_1 _6114_ (.Y(_1137_),
    .A(_1108_),
    .B(_1104_));
 sg13g2_o21ai_1 _6115_ (.B1(_0800_),
    .Y(_1138_),
    .A1(\main.demo.zic._q_tpos[4] ),
    .A2(_0436_));
 sg13g2_a21oi_1 _6116_ (.A1(_1137_),
    .A2(net39),
    .Y(_0226_),
    .B1(_1138_));
 sg13g2_nand3_1 _6117_ (.B(_0056_),
    .C(net45),
    .A(_1112_),
    .Y(_1139_));
 sg13g2_a21oi_1 _6118_ (.A1(_0406_),
    .A2(_1124_),
    .Y(_1140_),
    .B1(_0795_));
 sg13g2_and3_1 _6119_ (.X(_0227_),
    .A(_1114_),
    .B(_1139_),
    .C(_1140_));
 sg13g2_a21oi_1 _6120_ (.A1(_1113_),
    .A2(net38),
    .Y(_1141_),
    .B1(\main.demo.zic._q_tpos[6] ));
 sg13g2_nor3_1 _6121_ (.A(net61),
    .B(_1141_),
    .C(_1115_),
    .Y(_0228_));
 sg13g2_nor2_1 _6122_ (.A(_0406_),
    .B(_1126_),
    .Y(_1142_));
 sg13g2_nor2_1 _6123_ (.A(_1116_),
    .B(_1142_),
    .Y(_1143_));
 sg13g2_a21oi_1 _6124_ (.A1(_1142_),
    .A2(_1116_),
    .Y(_1144_),
    .B1(_0795_));
 sg13g2_nor2b_1 _6125_ (.A(_1143_),
    .B_N(_1144_),
    .Y(_0229_));
 sg13g2_a21oi_1 _6126_ (.A1(_1115_),
    .A2(_1116_),
    .Y(_1145_),
    .B1(\main.demo.zic._q_tpos[8] ));
 sg13g2_nor3_1 _6127_ (.A(net61),
    .B(_1121_),
    .C(_1145_),
    .Y(_0230_));
 sg13g2_inv_1 _6128_ (.Y(_1146_),
    .A(_1079_));
 sg13g2_nand2_1 _6129_ (.Y(_1147_),
    .A(_1142_),
    .B(_1118_));
 sg13g2_o21ai_1 _6130_ (.B1(net67),
    .Y(_1148_),
    .A1(_1146_),
    .A2(_1147_));
 sg13g2_a21oi_1 _6131_ (.A1(_1146_),
    .A2(_1147_),
    .Y(_0231_),
    .B1(_1148_));
 sg13g2_inv_1 _6132_ (.Y(_1149_),
    .A(_1129_));
 sg13g2_nor2_1 _6133_ (.A(_1041_),
    .B(_1039_),
    .Y(_1150_));
 sg13g2_inv_1 _6134_ (.Y(_1151_),
    .A(\main.demo.zic._q_squ_env[5] ));
 sg13g2_nand2_1 _6135_ (.Y(_1152_),
    .A(_1150_),
    .B(_1151_));
 sg13g2_nand2_2 _6136_ (.Y(_1153_),
    .A(_1152_),
    .B(_1006_));
 sg13g2_a21oi_1 _6137_ (.A1(_1040_),
    .A2(_0038_),
    .Y(_1154_),
    .B1(\main.demo.zic._q_qpos[12] ));
 sg13g2_inv_1 _6138_ (.Y(_1155_),
    .A(_1154_));
 sg13g2_nand2b_1 _6139_ (.Y(_1156_),
    .B(_1149_),
    .A_N(\main.demo.zic._q_tpos[10] ));
 sg13g2_nand2_1 _6140_ (.Y(_1157_),
    .A(\main.demo.zic._q_tpos[10] ),
    .B(_1129_));
 sg13g2_nand2_1 _6141_ (.Y(_1158_),
    .A(_1156_),
    .B(_1157_));
 sg13g2_buf_2 _6142_ (.A(_1158_),
    .X(_1159_));
 sg13g2_xnor2_1 _6143_ (.Y(_1160_),
    .A(_1079_),
    .B(_1159_));
 sg13g2_inv_1 _6144_ (.Y(_1161_),
    .A(_1160_));
 sg13g2_xnor2_1 _6145_ (.Y(_1162_),
    .A(\main.demo.zic._q_tpos[8] ),
    .B(_1159_));
 sg13g2_nor2b_1 _6146_ (.A(_1153_),
    .B_N(_1162_),
    .Y(_1163_));
 sg13g2_xnor2_1 _6147_ (.Y(_1164_),
    .A(_1116_),
    .B(_1159_));
 sg13g2_xnor2_1 _6148_ (.Y(_1165_),
    .A(_1155_),
    .B(_1164_));
 sg13g2_inv_1 _6149_ (.Y(_1166_),
    .A(_1165_));
 sg13g2_xnor2_1 _6150_ (.Y(_1167_),
    .A(_1081_),
    .B(_1159_));
 sg13g2_inv_1 _6151_ (.Y(_1168_),
    .A(_1153_));
 sg13g2_o21ai_1 _6152_ (.B1(_1168_),
    .Y(_1169_),
    .A1(_1151_),
    .A2(_1150_));
 sg13g2_o21ai_1 _6153_ (.B1(_1169_),
    .Y(_1170_),
    .A1(_0040_),
    .A2(_1006_));
 sg13g2_nor2b_1 _6154_ (.A(_1167_),
    .B_N(_1170_),
    .Y(_1171_));
 sg13g2_xor2_1 _6155_ (.B(_1039_),
    .A(_1041_),
    .X(_1172_));
 sg13g2_nor2_1 _6156_ (.A(_0039_),
    .B(_1006_),
    .Y(_1173_));
 sg13g2_a21oi_1 _6157_ (.A1(_1172_),
    .A2(_1006_),
    .Y(_1174_),
    .B1(_1173_));
 sg13g2_xnor2_1 _6158_ (.Y(_1175_),
    .A(\main.demo.zic._q_tpos[5] ),
    .B(_1159_));
 sg13g2_nor2b_1 _6159_ (.A(_1174_),
    .B_N(_1175_),
    .Y(_1176_));
 sg13g2_nand2_1 _6160_ (.Y(_1177_),
    .A(_1159_),
    .B(_1105_));
 sg13g2_nand3_1 _6161_ (.B(\main.demo.zic._q_tpos[4] ),
    .C(_1157_),
    .A(_1156_),
    .Y(_1178_));
 sg13g2_nand3_1 _6162_ (.B(_1178_),
    .C(_1041_),
    .A(_1177_),
    .Y(_1179_));
 sg13g2_xor2_1 _6163_ (.B(_1175_),
    .A(_1174_),
    .X(_1180_));
 sg13g2_nor2_1 _6164_ (.A(_1179_),
    .B(_1180_),
    .Y(_1181_));
 sg13g2_nor2_1 _6165_ (.A(_1176_),
    .B(_1181_),
    .Y(_1182_));
 sg13g2_xor2_1 _6166_ (.B(_1170_),
    .A(_1167_),
    .X(_1183_));
 sg13g2_nor2_1 _6167_ (.A(_1182_),
    .B(_1183_),
    .Y(_1184_));
 sg13g2_nor2_1 _6168_ (.A(_1171_),
    .B(_1184_),
    .Y(_1185_));
 sg13g2_nor2_1 _6169_ (.A(_1166_),
    .B(_1185_),
    .Y(_1186_));
 sg13g2_a21oi_1 _6170_ (.A1(_1154_),
    .A2(_1164_),
    .Y(_1187_),
    .B1(_1186_));
 sg13g2_inv_1 _6171_ (.Y(_1188_),
    .A(_1187_));
 sg13g2_xnor2_1 _6172_ (.Y(_1189_),
    .A(_1153_),
    .B(_1162_));
 sg13g2_nand2_1 _6173_ (.Y(_1190_),
    .A(_1188_),
    .B(_1189_));
 sg13g2_inv_1 _6174_ (.Y(_1191_),
    .A(_1190_));
 sg13g2_xnor2_1 _6175_ (.Y(_1192_),
    .A(_1155_),
    .B(_1160_));
 sg13g2_o21ai_1 _6176_ (.B1(_1192_),
    .Y(_1193_),
    .A1(_1163_),
    .A2(_1191_));
 sg13g2_o21ai_1 _6177_ (.B1(_1193_),
    .Y(_1194_),
    .A1(_1155_),
    .A2(_1161_));
 sg13g2_xnor2_1 _6178_ (.Y(_1195_),
    .A(_1129_),
    .B(_1153_));
 sg13g2_nand2_1 _6179_ (.Y(_1196_),
    .A(_1194_),
    .B(_1195_));
 sg13g2_o21ai_1 _6180_ (.B1(_1196_),
    .Y(_1197_),
    .A1(_1149_),
    .A2(_1153_));
 sg13g2_xnor2_1 _6181_ (.Y(_1198_),
    .A(_1123_),
    .B(_1154_));
 sg13g2_nand2b_1 _6182_ (.Y(_1199_),
    .B(_1198_),
    .A_N(_1197_));
 sg13g2_inv_1 _6183_ (.Y(_1200_),
    .A(_0411_));
 sg13g2_nand2b_1 _6184_ (.Y(_1201_),
    .B(_1197_),
    .A_N(_1198_));
 sg13g2_nand3_1 _6185_ (.B(_1200_),
    .C(_1201_),
    .A(_1199_),
    .Y(_1202_));
 sg13g2_nor2_1 _6186_ (.A(_0041_),
    .B(_1202_),
    .Y(_1203_));
 sg13g2_a21oi_1 _6187_ (.A1(_1194_),
    .A2(_1195_),
    .Y(_1204_),
    .B1(_0411_));
 sg13g2_o21ai_1 _6188_ (.B1(_1204_),
    .Y(_1205_),
    .A1(_1194_),
    .A2(_1195_));
 sg13g2_nand2_1 _6189_ (.Y(_1206_),
    .A(_1183_),
    .B(_1182_));
 sg13g2_nand3b_1 _6190_ (.B(_1200_),
    .C(_1206_),
    .Y(_1207_),
    .A_N(_1184_));
 sg13g2_nor2_1 _6191_ (.A(\main.demo.zic._q_clock_count[1] ),
    .B(_1207_),
    .Y(_1208_));
 sg13g2_a21oi_1 _6192_ (.A1(_1179_),
    .A2(_1180_),
    .Y(_1209_),
    .B1(_0411_));
 sg13g2_nand2b_1 _6193_ (.Y(_1210_),
    .B(_1209_),
    .A_N(_1181_));
 sg13g2_o21ai_1 _6194_ (.B1(_1210_),
    .Y(_1211_),
    .A1(\main.demo.zic._q_clock_count[0] ),
    .A2(_0066_));
 sg13g2_o21ai_1 _6195_ (.B1(_1211_),
    .Y(_1212_),
    .A1(_0066_),
    .A2(_1210_));
 sg13g2_nand2b_1 _6196_ (.Y(_1213_),
    .B(_1212_),
    .A_N(_1208_));
 sg13g2_nand2_1 _6197_ (.Y(_1214_),
    .A(_1207_),
    .B(\main.demo.zic._q_clock_count[1] ));
 sg13g2_a21oi_1 _6198_ (.A1(_1185_),
    .A2(_1166_),
    .Y(_1215_),
    .B1(_0411_));
 sg13g2_nand2b_1 _6199_ (.Y(_1216_),
    .B(_1215_),
    .A_N(_1186_));
 sg13g2_nor2_1 _6200_ (.A(_4403_),
    .B(_1216_),
    .Y(_1217_));
 sg13g2_a21o_1 _6201_ (.A2(_1214_),
    .A1(_1213_),
    .B1(_1217_),
    .X(_1218_));
 sg13g2_nor2_1 _6202_ (.A(_1189_),
    .B(_1188_),
    .Y(_1219_));
 sg13g2_nor3_1 _6203_ (.A(_0411_),
    .B(_1219_),
    .C(_1191_),
    .Y(_1220_));
 sg13g2_nor2b_1 _6204_ (.A(_1220_),
    .B_N(_4402_),
    .Y(_1221_));
 sg13g2_nand2_1 _6205_ (.Y(_1222_),
    .A(_1216_),
    .B(_4403_));
 sg13g2_nor2b_1 _6206_ (.A(_1221_),
    .B_N(_1222_),
    .Y(_1223_));
 sg13g2_nor2b_1 _6207_ (.A(_4402_),
    .B_N(_1220_),
    .Y(_1224_));
 sg13g2_a21oi_1 _6208_ (.A1(_1218_),
    .A2(_1223_),
    .Y(_1225_),
    .B1(_1224_));
 sg13g2_a22oi_1 _6209_ (.Y(_1226_),
    .B1(_4406_),
    .B2(_1225_),
    .A2(\main.demo.zic._q_clock_count[5] ),
    .A1(_1205_));
 sg13g2_nor3_1 _6210_ (.A(_1192_),
    .B(_1163_),
    .C(_1191_),
    .Y(_1227_));
 sg13g2_nand3b_1 _6211_ (.B(_1193_),
    .C(_1200_),
    .Y(_1228_),
    .A_N(_1227_));
 sg13g2_o21ai_1 _6212_ (.B1(_1228_),
    .Y(_1229_),
    .A1(_4406_),
    .A2(_1225_));
 sg13g2_nor2_1 _6213_ (.A(\main.demo.zic._q_clock_count[5] ),
    .B(_1205_),
    .Y(_1230_));
 sg13g2_a21oi_1 _6214_ (.A1(_1226_),
    .A2(_1229_),
    .Y(_1231_),
    .B1(_1230_));
 sg13g2_nand2_1 _6215_ (.Y(_1232_),
    .A(_1202_),
    .B(_0041_));
 sg13g2_o21ai_1 _6216_ (.B1(_1232_),
    .Y(\main._w_demo_audio1 ),
    .A1(_1203_),
    .A2(_1231_));
 sg13g2_buf_1 _6217_ (.A(_4132_),
    .X(_1233_));
 sg13g2_a21oi_1 _6218_ (.A1(_4124_),
    .A2(_4130_),
    .Y(_1234_),
    .B1(_4116_));
 sg13g2_inv_1 _6219_ (.Y(_1235_),
    .A(_1234_));
 sg13g2_nor2_1 _6220_ (.A(net66),
    .B(_1235_),
    .Y(_1236_));
 sg13g2_a21oi_1 _6221_ (.A1(_4083_),
    .A2(net66),
    .Y(_1237_),
    .B1(_1236_));
 sg13g2_xnor2_1 _6222_ (.Y(_1238_),
    .A(_4087_),
    .B(_1237_));
 sg13g2_xnor2_1 _6223_ (.Y(_1239_),
    .A(_4093_),
    .B(_4089_));
 sg13g2_buf_1 _6224_ (.A(_4031_),
    .X(_1240_));
 sg13g2_buf_1 _6225_ (.A(net65),
    .X(_1241_));
 sg13g2_nand2_1 _6226_ (.Y(_1242_),
    .A(_4086_),
    .B(_4080_));
 sg13g2_nor2_1 _6227_ (.A(_4074_),
    .B(_4068_),
    .Y(_1243_));
 sg13g2_inv_1 _6228_ (.Y(_1244_),
    .A(_1243_));
 sg13g2_inv_1 _6229_ (.Y(_1245_),
    .A(_4056_));
 sg13g2_nor2_1 _6230_ (.A(_4062_),
    .B(_1245_),
    .Y(_1246_));
 sg13g2_nand2_1 _6231_ (.Y(_1247_),
    .A(_4125_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_nand2_1 _6232_ (.Y(_1248_),
    .A(_1246_),
    .B(_1247_));
 sg13g2_nor2_1 _6233_ (.A(_1244_),
    .B(_1248_),
    .Y(_1249_));
 sg13g2_a21oi_1 _6234_ (.A1(_4110_),
    .A2(_4055_),
    .Y(_1250_),
    .B1(_4060_));
 sg13g2_inv_1 _6235_ (.Y(_1251_),
    .A(_1250_));
 sg13g2_a221oi_1 _6236_ (.B2(_1243_),
    .C1(_4072_),
    .B1(_1251_),
    .A1(_4073_),
    .Y(_1252_),
    .A2(_4065_));
 sg13g2_nor2b_1 _6237_ (.A(_1249_),
    .B_N(_1252_),
    .Y(_1253_));
 sg13g2_a21oi_1 _6238_ (.A1(_4086_),
    .A2(_4078_),
    .Y(_1254_),
    .B1(_4085_));
 sg13g2_o21ai_1 _6239_ (.B1(_1254_),
    .Y(_1255_),
    .A1(_1242_),
    .A2(_1253_));
 sg13g2_xnor2_1 _6240_ (.Y(_1256_),
    .A(_4093_),
    .B(_1255_));
 sg13g2_nor2_1 _6241_ (.A(net65),
    .B(_1256_),
    .Y(_1257_));
 sg13g2_a21oi_2 _6242_ (.B1(_1257_),
    .Y(_1258_),
    .A2(net57),
    .A1(_1239_));
 sg13g2_xnor2_1 _6243_ (.Y(_1259_),
    .A(_4080_),
    .B(_4076_));
 sg13g2_nor2_1 _6244_ (.A(_4081_),
    .B(_1253_),
    .Y(_1260_));
 sg13g2_nor2b_1 _6245_ (.A(_4080_),
    .B_N(_1253_),
    .Y(_1261_));
 sg13g2_o21ai_1 _6246_ (.B1(net77),
    .Y(_1262_),
    .A1(_1260_),
    .A2(_1261_));
 sg13g2_o21ai_1 _6247_ (.B1(_1262_),
    .Y(_1263_),
    .A1(net77),
    .A2(_1259_));
 sg13g2_buf_1 _6248_ (.A(_1263_),
    .X(_1264_));
 sg13g2_xor2_1 _6249_ (.B(_4056_),
    .A(_4051_),
    .X(_1265_));
 sg13g2_nor2_1 _6250_ (.A(net77),
    .B(_1265_),
    .Y(_1266_));
 sg13g2_inv_1 _6251_ (.Y(_1267_),
    .A(_1247_));
 sg13g2_nand2_1 _6252_ (.Y(_1268_),
    .A(_1245_),
    .B(_1267_));
 sg13g2_nand2_1 _6253_ (.Y(_1269_),
    .A(_4056_),
    .B(_1247_));
 sg13g2_a21o_1 _6254_ (.A2(_1269_),
    .A1(_1268_),
    .B1(_4031_),
    .X(_1270_));
 sg13g2_nand2b_1 _6255_ (.Y(_1271_),
    .B(_1270_),
    .A_N(_1266_));
 sg13g2_inv_1 _6256_ (.Y(_1272_),
    .A(_1271_));
 sg13g2_xnor2_1 _6257_ (.Y(_1273_),
    .A(_4061_),
    .B(_4058_));
 sg13g2_nor2_1 _6258_ (.A(net77),
    .B(_1273_),
    .Y(_1274_));
 sg13g2_inv_1 _6259_ (.Y(_1275_),
    .A(_4055_));
 sg13g2_nand2_1 _6260_ (.Y(_1276_),
    .A(_1269_),
    .B(_1275_));
 sg13g2_inv_1 _6261_ (.Y(_1277_),
    .A(_1276_));
 sg13g2_nor2_1 _6262_ (.A(_4062_),
    .B(_1277_),
    .Y(_1278_));
 sg13g2_nand2_1 _6263_ (.Y(_1279_),
    .A(_1277_),
    .B(_4062_));
 sg13g2_inv_1 _6264_ (.Y(_1280_),
    .A(_1279_));
 sg13g2_o21ai_1 _6265_ (.B1(_4132_),
    .Y(_1281_),
    .A1(_1278_),
    .A2(_1280_));
 sg13g2_nand2b_1 _6266_ (.Y(_1282_),
    .B(_1281_),
    .A_N(_1274_));
 sg13g2_inv_1 _6267_ (.Y(_1283_),
    .A(_1282_));
 sg13g2_nor2_1 _6268_ (.A(_1272_),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_inv_1 _6269_ (.Y(_1285_),
    .A(_1284_));
 sg13g2_xnor2_1 _6270_ (.Y(_1286_),
    .A(_4067_),
    .B(_4064_));
 sg13g2_a21oi_1 _6271_ (.A1(_1248_),
    .A2(_1250_),
    .Y(_1287_),
    .B1(_4068_));
 sg13g2_and3_1 _6272_ (.X(_1288_),
    .A(_1248_),
    .B(_4068_),
    .C(_1250_));
 sg13g2_o21ai_1 _6273_ (.B1(net77),
    .Y(_1289_),
    .A1(_1287_),
    .A2(_1288_));
 sg13g2_o21ai_1 _6274_ (.B1(_1289_),
    .Y(_1290_),
    .A1(net77),
    .A2(_1286_));
 sg13g2_inv_1 _6275_ (.Y(_1291_),
    .A(_1290_));
 sg13g2_nor2_1 _6276_ (.A(_1285_),
    .B(_1291_),
    .Y(_1292_));
 sg13g2_inv_1 _6277_ (.Y(_1293_),
    .A(_1292_));
 sg13g2_inv_1 _6278_ (.Y(_1294_),
    .A(_4065_));
 sg13g2_inv_1 _6279_ (.Y(_1295_),
    .A(_4060_));
 sg13g2_a21oi_1 _6280_ (.A1(_1294_),
    .A2(_1295_),
    .Y(_1296_),
    .B1(_4066_));
 sg13g2_nor2_1 _6281_ (.A(_4123_),
    .B(_1277_),
    .Y(_1297_));
 sg13g2_nor3_1 _6282_ (.A(_4031_),
    .B(_1296_),
    .C(_1297_),
    .Y(_1298_));
 sg13g2_a21oi_1 _6283_ (.A1(_4070_),
    .A2(net65),
    .Y(_1299_),
    .B1(_1298_));
 sg13g2_xnor2_1 _6284_ (.Y(_1300_),
    .A(_4073_),
    .B(_1299_));
 sg13g2_inv_1 _6285_ (.Y(_1301_),
    .A(_1300_));
 sg13g2_nor2_1 _6286_ (.A(_1293_),
    .B(_1301_),
    .Y(_1302_));
 sg13g2_nand2_1 _6287_ (.Y(_1303_),
    .A(_1264_),
    .B(_1302_));
 sg13g2_inv_1 _6288_ (.Y(_1304_),
    .A(_1296_));
 sg13g2_a21oi_1 _6289_ (.A1(_4080_),
    .A2(_4072_),
    .Y(_1305_),
    .B1(_4078_));
 sg13g2_o21ai_1 _6290_ (.B1(_1305_),
    .Y(_1306_),
    .A1(_1304_),
    .A2(_4114_));
 sg13g2_a21oi_1 _6291_ (.A1(_4124_),
    .A2(_1276_),
    .Y(_1307_),
    .B1(_1306_));
 sg13g2_inv_1 _6292_ (.Y(_1308_),
    .A(_1307_));
 sg13g2_nor2_1 _6293_ (.A(net65),
    .B(_1308_),
    .Y(_1309_));
 sg13g2_a21oi_1 _6294_ (.A1(_4083_),
    .A2(net65),
    .Y(_1310_),
    .B1(_1309_));
 sg13g2_xnor2_1 _6295_ (.Y(_1311_),
    .A(_4086_),
    .B(_1310_));
 sg13g2_inv_1 _6296_ (.Y(_1312_),
    .A(_1311_));
 sg13g2_nor2_1 _6297_ (.A(_1303_),
    .B(_1312_),
    .Y(_1313_));
 sg13g2_inv_1 _6298_ (.Y(_1314_),
    .A(_1313_));
 sg13g2_nand2_1 _6299_ (.Y(_1315_),
    .A(_4138_),
    .B(_1314_));
 sg13g2_xnor2_1 _6300_ (.Y(_1316_),
    .A(_1258_),
    .B(_1315_));
 sg13g2_nor2_1 _6301_ (.A(_1238_),
    .B(_1316_),
    .Y(_1317_));
 sg13g2_nand2_1 _6302_ (.Y(_1318_),
    .A(_1246_),
    .B(_4127_));
 sg13g2_a21oi_1 _6303_ (.A1(_1295_),
    .A2(_4053_),
    .Y(_1319_),
    .B1(_4059_));
 sg13g2_nand3_1 _6304_ (.B(_4067_),
    .C(_1319_),
    .A(_1318_),
    .Y(_1320_));
 sg13g2_a21o_1 _6305_ (.A2(_1319_),
    .A1(_1318_),
    .B1(_4067_),
    .X(_1321_));
 sg13g2_nand3_1 _6306_ (.B(net65),
    .C(_1321_),
    .A(_1320_),
    .Y(_1322_));
 sg13g2_o21ai_1 _6307_ (.B1(_1322_),
    .Y(_1323_),
    .A1(net65),
    .A2(_1286_));
 sg13g2_nand2_1 _6308_ (.Y(_1324_),
    .A(_4138_),
    .B(_1293_));
 sg13g2_xnor2_1 _6309_ (.Y(_1325_),
    .A(_1300_),
    .B(_1324_));
 sg13g2_inv_1 _6310_ (.Y(_1326_),
    .A(_4130_));
 sg13g2_nand2_1 _6311_ (.Y(_1327_),
    .A(_1326_),
    .B(_4061_));
 sg13g2_nand2_1 _6312_ (.Y(_1328_),
    .A(_4130_),
    .B(_4062_));
 sg13g2_nand3_1 _6313_ (.B(net65),
    .C(_1328_),
    .A(_1327_),
    .Y(_1329_));
 sg13g2_o21ai_1 _6314_ (.B1(_1329_),
    .Y(_1330_),
    .A1(_1240_),
    .A2(_1273_));
 sg13g2_nand2_1 _6315_ (.Y(_1331_),
    .A(_4138_),
    .B(_1285_));
 sg13g2_xnor2_1 _6316_ (.Y(_1332_),
    .A(_1290_),
    .B(_1331_));
 sg13g2_nor2_1 _6317_ (.A(_1240_),
    .B(_1265_),
    .Y(_1333_));
 sg13g2_nand2_1 _6318_ (.Y(_1334_),
    .A(_1245_),
    .B(_4126_));
 sg13g2_a21o_1 _6319_ (.A2(_4128_),
    .A1(_1334_),
    .B1(net77),
    .X(_1335_));
 sg13g2_nand2b_1 _6320_ (.Y(_1336_),
    .B(_1335_),
    .A_N(_1333_));
 sg13g2_buf_1 _6321_ (.A(_1336_),
    .X(_1337_));
 sg13g2_nand2_1 _6322_ (.Y(_1338_),
    .A(_4138_),
    .B(_1272_));
 sg13g2_xnor2_1 _6323_ (.Y(_1339_),
    .A(_1282_),
    .B(_1338_));
 sg13g2_nor2_1 _6324_ (.A(_1337_),
    .B(_1339_),
    .Y(_1340_));
 sg13g2_xnor2_1 _6325_ (.Y(_1341_),
    .A(_1337_),
    .B(_1339_));
 sg13g2_nor2_1 _6326_ (.A(_4126_),
    .B(_1267_),
    .Y(_1342_));
 sg13g2_nor2_1 _6327_ (.A(_1342_),
    .B(_1271_),
    .Y(_1343_));
 sg13g2_nor2b_1 _6328_ (.A(_1341_),
    .B_N(_1343_),
    .Y(_1344_));
 sg13g2_inv_1 _6329_ (.Y(_1345_),
    .A(_1330_));
 sg13g2_xnor2_1 _6330_ (.Y(_1346_),
    .A(_1345_),
    .B(_1332_));
 sg13g2_o21ai_1 _6331_ (.B1(_1346_),
    .Y(_1347_),
    .A1(_1340_),
    .A2(_1344_));
 sg13g2_o21ai_1 _6332_ (.B1(_1347_),
    .Y(_1348_),
    .A1(_1330_),
    .A2(_1332_));
 sg13g2_inv_1 _6333_ (.Y(_1349_),
    .A(_1323_));
 sg13g2_xnor2_1 _6334_ (.Y(_1350_),
    .A(_1349_),
    .B(_1325_));
 sg13g2_nand2_1 _6335_ (.Y(_1351_),
    .A(_1348_),
    .B(_1350_));
 sg13g2_o21ai_1 _6336_ (.B1(_1351_),
    .Y(_1352_),
    .A1(_1323_),
    .A2(_1325_));
 sg13g2_a21oi_1 _6337_ (.A1(_4130_),
    .A2(_4122_),
    .Y(_1353_),
    .B1(_4111_));
 sg13g2_mux2_1 _6338_ (.A0(_1353_),
    .A1(_4070_),
    .S(net66),
    .X(_1354_));
 sg13g2_xnor2_1 _6339_ (.Y(_1355_),
    .A(_4074_),
    .B(_1354_));
 sg13g2_inv_1 _6340_ (.Y(_1356_),
    .A(_1355_));
 sg13g2_nor2_1 _6341_ (.A(_1302_),
    .B(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ),
    .Y(_1357_));
 sg13g2_xor2_1 _6342_ (.B(_1357_),
    .A(_1264_),
    .X(_1358_));
 sg13g2_xnor2_1 _6343_ (.Y(_1359_),
    .A(_1356_),
    .B(_1358_));
 sg13g2_nor2_1 _6344_ (.A(_1355_),
    .B(_1358_),
    .Y(_1360_));
 sg13g2_a21oi_1 _6345_ (.A1(_1352_),
    .A2(_1359_),
    .Y(_1361_),
    .B1(_1360_));
 sg13g2_nand2_1 _6346_ (.Y(_1362_),
    .A(_4138_),
    .B(_1303_));
 sg13g2_xnor2_1 _6347_ (.Y(_1363_),
    .A(_1312_),
    .B(_1362_));
 sg13g2_nor2_1 _6348_ (.A(_1244_),
    .B(_1318_),
    .Y(_1364_));
 sg13g2_inv_1 _6349_ (.Y(_1365_),
    .A(_1319_));
 sg13g2_a221oi_1 _6350_ (.B2(_1243_),
    .C1(_4071_),
    .B1(_1365_),
    .A1(_4073_),
    .Y(_1366_),
    .A2(_4066_));
 sg13g2_nor2b_1 _6351_ (.A(_1364_),
    .B_N(_1366_),
    .Y(_1367_));
 sg13g2_nand2b_1 _6352_ (.Y(_1368_),
    .B(_4081_),
    .A_N(_1367_));
 sg13g2_nand2_1 _6353_ (.Y(_1369_),
    .A(_1367_),
    .B(_4080_));
 sg13g2_nand3_1 _6354_ (.B(net57),
    .C(_1369_),
    .A(_1368_),
    .Y(_1370_));
 sg13g2_o21ai_1 _6355_ (.B1(_1370_),
    .Y(_1371_),
    .A1(net57),
    .A2(_1259_));
 sg13g2_nand2b_1 _6356_ (.Y(_1372_),
    .B(_1371_),
    .A_N(_1363_));
 sg13g2_nand2b_1 _6357_ (.Y(_1373_),
    .B(_1372_),
    .A_N(_1361_));
 sg13g2_inv_1 _6358_ (.Y(_1374_),
    .A(_1371_));
 sg13g2_nand2_1 _6359_ (.Y(_1375_),
    .A(_1363_),
    .B(_1374_));
 sg13g2_nand2_1 _6360_ (.Y(_1376_),
    .A(_1373_),
    .B(_1375_));
 sg13g2_inv_1 _6361_ (.Y(_1377_),
    .A(_1376_));
 sg13g2_nand2_1 _6362_ (.Y(_1378_),
    .A(_1316_),
    .B(_1238_));
 sg13g2_o21ai_1 _6363_ (.B1(_1378_),
    .Y(_1379_),
    .A1(_1317_),
    .A2(_1377_));
 sg13g2_xnor2_1 _6364_ (.Y(_1380_),
    .A(_4099_),
    .B(_4095_));
 sg13g2_a21oi_1 _6365_ (.A1(_4092_),
    .A2(_4085_),
    .Y(_1381_),
    .B1(_4091_));
 sg13g2_inv_1 _6366_ (.Y(_1382_),
    .A(_1381_));
 sg13g2_a21oi_1 _6367_ (.A1(_1308_),
    .A2(_4117_),
    .Y(_1383_),
    .B1(_1382_));
 sg13g2_nor2_1 _6368_ (.A(_4100_),
    .B(_1383_),
    .Y(_1384_));
 sg13g2_nor2b_1 _6369_ (.A(_4099_),
    .B_N(_1383_),
    .Y(_1385_));
 sg13g2_o21ai_1 _6370_ (.B1(net66),
    .Y(_1386_),
    .A1(_1384_),
    .A2(_1385_));
 sg13g2_o21ai_1 _6371_ (.B1(_1386_),
    .Y(_1387_),
    .A1(net66),
    .A2(_1380_));
 sg13g2_inv_1 _6372_ (.Y(_1388_),
    .A(_1387_));
 sg13g2_nor2_1 _6373_ (.A(_1314_),
    .B(_1258_),
    .Y(_1389_));
 sg13g2_inv_1 _6374_ (.Y(_1390_),
    .A(_1389_));
 sg13g2_nand2_1 _6375_ (.Y(_1391_),
    .A(net19),
    .B(_1390_));
 sg13g2_xnor2_1 _6376_ (.Y(_1392_),
    .A(_1388_),
    .B(_1391_));
 sg13g2_a21oi_1 _6377_ (.A1(_4086_),
    .A2(_4077_),
    .Y(_1393_),
    .B1(_4084_));
 sg13g2_o21ai_1 _6378_ (.B1(_1393_),
    .Y(_1394_),
    .A1(_1242_),
    .A2(_1367_));
 sg13g2_xnor2_1 _6379_ (.Y(_1395_),
    .A(_4093_),
    .B(_1394_));
 sg13g2_nor2_1 _6380_ (.A(net66),
    .B(_1395_),
    .Y(_1396_));
 sg13g2_a21oi_1 _6381_ (.A1(_1239_),
    .A2(net66),
    .Y(_1397_),
    .B1(_1396_));
 sg13g2_inv_1 _6382_ (.Y(_1398_),
    .A(_1397_));
 sg13g2_nand2b_1 _6383_ (.Y(_1399_),
    .B(_1398_),
    .A_N(_1392_));
 sg13g2_nand2_1 _6384_ (.Y(_1400_),
    .A(_1379_),
    .B(_1399_));
 sg13g2_nand2_1 _6385_ (.Y(_1401_),
    .A(_1392_),
    .B(_1397_));
 sg13g2_nand2_1 _6386_ (.Y(_1402_),
    .A(_1400_),
    .B(_1401_));
 sg13g2_a21oi_1 _6387_ (.A1(_1235_),
    .A2(_4117_),
    .Y(_1403_),
    .B1(_4108_));
 sg13g2_nand2b_1 _6388_ (.Y(_1404_),
    .B(_4100_),
    .A_N(_1403_));
 sg13g2_nand2_1 _6389_ (.Y(_1405_),
    .A(_1403_),
    .B(_4099_));
 sg13g2_nand3_1 _6390_ (.B(net57),
    .C(_1405_),
    .A(_1404_),
    .Y(_1406_));
 sg13g2_o21ai_1 _6391_ (.B1(_1406_),
    .Y(_1407_),
    .A1(net57),
    .A2(_1380_));
 sg13g2_buf_1 _6392_ (.A(_1407_),
    .X(_1408_));
 sg13g2_nand3_1 _6393_ (.B(_4099_),
    .C(_4092_),
    .A(_1255_),
    .Y(_1409_));
 sg13g2_nor2b_1 _6394_ (.A(_4096_),
    .B_N(_4091_),
    .Y(_1410_));
 sg13g2_nor3_1 _6395_ (.A(_1241_),
    .B(_4097_),
    .C(_1410_),
    .Y(_1411_));
 sg13g2_a22oi_1 _6396_ (.Y(_1412_),
    .B1(_1241_),
    .B2(_4102_),
    .A2(_1411_),
    .A1(_1409_));
 sg13g2_xnor2_1 _6397_ (.Y(_1413_),
    .A(_4105_),
    .B(_1412_));
 sg13g2_nor2_1 _6398_ (.A(_1390_),
    .B(_1388_),
    .Y(_1414_));
 sg13g2_inv_1 _6399_ (.Y(_1415_),
    .A(_1414_));
 sg13g2_nand2_1 _6400_ (.Y(_1416_),
    .A(net19),
    .B(_1415_));
 sg13g2_xnor2_1 _6401_ (.Y(_1417_),
    .A(_1413_),
    .B(_1416_));
 sg13g2_nor2b_1 _6402_ (.A(_1408_),
    .B_N(_1417_),
    .Y(_1418_));
 sg13g2_nand2b_1 _6403_ (.Y(_1419_),
    .B(_1408_),
    .A_N(_1417_));
 sg13g2_nor2b_1 _6404_ (.A(_1418_),
    .B_N(_1419_),
    .Y(_1420_));
 sg13g2_nand2_1 _6405_ (.Y(_1421_),
    .A(_1402_),
    .B(_1420_));
 sg13g2_nand3_1 _6406_ (.B(_4124_),
    .C(_1276_),
    .A(_4119_),
    .Y(_1422_));
 sg13g2_nand2b_1 _6407_ (.Y(_1423_),
    .B(_4097_),
    .A_N(_4033_));
 sg13g2_nand3_1 _6408_ (.B(net66),
    .C(_4034_),
    .A(_1423_),
    .Y(_1424_));
 sg13g2_a221oi_1 _6409_ (.B2(_4119_),
    .C1(_1424_),
    .B1(_1306_),
    .A1(_4106_),
    .Y(_1425_),
    .A2(_1382_));
 sg13g2_a22oi_1 _6410_ (.Y(_1426_),
    .B1(net57),
    .B2(_4104_),
    .A2(_1425_),
    .A1(_1422_));
 sg13g2_xnor2_1 _6411_ (.Y(_1427_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ),
    .B(_1426_));
 sg13g2_nor2_1 _6412_ (.A(_1415_),
    .B(_1413_),
    .Y(_1428_));
 sg13g2_inv_1 _6413_ (.Y(_1429_),
    .A(_1428_));
 sg13g2_nand2_1 _6414_ (.Y(_1430_),
    .A(net19),
    .B(_1429_));
 sg13g2_xor2_1 _6415_ (.B(_1430_),
    .A(_1427_),
    .X(_1431_));
 sg13g2_xnor2_1 _6416_ (.Y(_1432_),
    .A(_4105_),
    .B(_4102_));
 sg13g2_inv_1 _6417_ (.Y(_1433_),
    .A(_1432_));
 sg13g2_nand2_1 _6418_ (.Y(_1434_),
    .A(_4099_),
    .B(_4092_));
 sg13g2_nor2_1 _6419_ (.A(_1242_),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_a221oi_1 _6420_ (.B2(_1435_),
    .C1(_4096_),
    .B1(_1364_),
    .A1(_4099_),
    .Y(_1436_),
    .A2(_4090_));
 sg13g2_nand2b_1 _6421_ (.Y(_1437_),
    .B(_1435_),
    .A_N(_1366_));
 sg13g2_or2_1 _6422_ (.X(_1438_),
    .B(_1393_),
    .A(_1434_));
 sg13g2_nand3_1 _6423_ (.B(_1437_),
    .C(_1438_),
    .A(_1436_),
    .Y(_1439_));
 sg13g2_xnor2_1 _6424_ (.Y(_1440_),
    .A(_4036_),
    .B(_1439_));
 sg13g2_nand2_1 _6425_ (.Y(_1441_),
    .A(_1440_),
    .B(net57));
 sg13g2_o21ai_1 _6426_ (.B1(_1441_),
    .Y(_1442_),
    .A1(net57),
    .A2(_1433_));
 sg13g2_inv_1 _6427_ (.Y(_1443_),
    .A(_1442_));
 sg13g2_nand2_1 _6428_ (.Y(_1444_),
    .A(_1431_),
    .B(_1443_));
 sg13g2_nor2b_1 _6429_ (.A(_1418_),
    .B_N(_1444_),
    .Y(_1445_));
 sg13g2_nor2_1 _6430_ (.A(_1443_),
    .B(_1431_),
    .Y(_1446_));
 sg13g2_a21oi_1 _6431_ (.A1(_1421_),
    .A2(_1445_),
    .Y(_1447_),
    .B1(_1446_));
 sg13g2_o21ai_1 _6432_ (.B1(_1427_),
    .Y(_1448_),
    .A1(_1429_),
    .A2(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ));
 sg13g2_nand2b_1 _6433_ (.Y(_1449_),
    .B(_1448_),
    .A_N(_1447_));
 sg13g2_nand2b_1 _6434_ (.Y(_1450_),
    .B(_1447_),
    .A_N(_1448_));
 sg13g2_nand2_1 _6435_ (.Y(_1451_),
    .A(_1449_),
    .B(_1450_));
 sg13g2_buf_2 _6436_ (.A(_1451_),
    .X(_1452_));
 sg13g2_buf_1 _6437_ (.A(_1452_),
    .X(_1453_));
 sg13g2_inv_1 _6438_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ),
    .A(net13));
 sg13g2_inv_1 _6439_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_a[4] ),
    .A(_1453_));
 sg13g2_xnor2_1 _6440_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_a[6] ),
    .A(_1233_),
    .B(_0070_));
 sg13g2_nor2_1 _6441_ (.A(_1233_),
    .B(_0070_),
    .Y(_1454_));
 sg13g2_xor2_1 _6442_ (.B(_1454_),
    .A(_0071_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[7] ));
 sg13g2_xnor2_1 _6443_ (.Y(_1455_),
    .A(_1342_),
    .B(_1337_));
 sg13g2_nor2_1 _6444_ (.A(_1340_),
    .B(_1344_),
    .Y(_1456_));
 sg13g2_xnor2_1 _6445_ (.Y(_1457_),
    .A(_1346_),
    .B(_1456_));
 sg13g2_xnor2_1 _6446_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[0] ),
    .A(_1455_),
    .B(_1457_));
 sg13g2_inv_1 _6447_ (.Y(_1458_),
    .A(_1337_));
 sg13g2_nor2_1 _6448_ (.A(_1458_),
    .B(_1345_),
    .Y(_1459_));
 sg13g2_inv_1 _6449_ (.Y(_1460_),
    .A(_1459_));
 sg13g2_nor2_1 _6450_ (.A(_1460_),
    .B(_1349_),
    .Y(_1461_));
 sg13g2_inv_1 _6451_ (.Y(_1462_),
    .A(_1461_));
 sg13g2_nor2_1 _6452_ (.A(_1462_),
    .B(_1356_),
    .Y(_1463_));
 sg13g2_inv_1 _6453_ (.Y(_1464_),
    .A(_1463_));
 sg13g2_nor2_1 _6454_ (.A(_1464_),
    .B(_1374_),
    .Y(_1465_));
 sg13g2_inv_1 _6455_ (.Y(_1466_),
    .A(_1465_));
 sg13g2_nor2_1 _6456_ (.A(_1466_),
    .B(_1238_),
    .Y(_1467_));
 sg13g2_nand2_1 _6457_ (.Y(_1468_),
    .A(_1398_),
    .B(_1467_));
 sg13g2_nor2b_1 _6458_ (.A(_1468_),
    .B_N(_1408_),
    .Y(_1469_));
 sg13g2_nand3_1 _6459_ (.B(_1442_),
    .C(_1469_),
    .A(net19),
    .Y(_1470_));
 sg13g2_xor2_1 _6460_ (.B(_1470_),
    .A(_1427_),
    .X(_1471_));
 sg13g2_nor2_1 _6461_ (.A(_1469_),
    .B(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ),
    .Y(_1472_));
 sg13g2_xnor2_1 _6462_ (.Y(_1473_),
    .A(_1442_),
    .B(_1472_));
 sg13g2_nor2_1 _6463_ (.A(_1387_),
    .B(_1473_),
    .Y(_1474_));
 sg13g2_xnor2_1 _6464_ (.Y(_1475_),
    .A(_1387_),
    .B(_1473_));
 sg13g2_nand2_1 _6465_ (.Y(_1476_),
    .A(net19),
    .B(_1468_));
 sg13g2_xnor2_1 _6466_ (.Y(_1477_),
    .A(_1408_),
    .B(_1476_));
 sg13g2_nor2_1 _6467_ (.A(_1258_),
    .B(_1477_),
    .Y(_1478_));
 sg13g2_nand2_1 _6468_ (.Y(_1479_),
    .A(net19),
    .B(_1466_));
 sg13g2_xnor2_1 _6469_ (.Y(_1480_),
    .A(_1238_),
    .B(_1479_));
 sg13g2_nor2_1 _6470_ (.A(_1264_),
    .B(_1480_),
    .Y(_1481_));
 sg13g2_nand2_1 _6471_ (.Y(_1482_),
    .A(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .B(_1462_));
 sg13g2_xnor2_1 _6472_ (.Y(_1483_),
    .A(_1355_),
    .B(_1482_));
 sg13g2_nand2_1 _6473_ (.Y(_1484_),
    .A(_1483_),
    .B(_1291_));
 sg13g2_inv_1 _6474_ (.Y(_1485_),
    .A(_1484_));
 sg13g2_nand2_1 _6475_ (.Y(_1486_),
    .A(net19),
    .B(_1460_));
 sg13g2_xnor2_1 _6476_ (.Y(_1487_),
    .A(_1323_),
    .B(_1486_));
 sg13g2_xnor2_1 _6477_ (.Y(_1488_),
    .A(_1282_),
    .B(_1487_));
 sg13g2_inv_1 _6478_ (.Y(_1489_),
    .A(_1488_));
 sg13g2_nand2_1 _6479_ (.Y(_1490_),
    .A(_4138_),
    .B(_1458_));
 sg13g2_xnor2_1 _6480_ (.Y(_1491_),
    .A(_1330_),
    .B(_1490_));
 sg13g2_inv_1 _6481_ (.Y(_1492_),
    .A(_1342_));
 sg13g2_nor2_1 _6482_ (.A(_1492_),
    .B(_1337_),
    .Y(_1493_));
 sg13g2_xnor2_1 _6483_ (.Y(_1494_),
    .A(_1272_),
    .B(_1491_));
 sg13g2_nor2_1 _6484_ (.A(_1493_),
    .B(_1494_),
    .Y(_1495_));
 sg13g2_a21oi_1 _6485_ (.A1(_1272_),
    .A2(_1491_),
    .Y(_1496_),
    .B1(_1495_));
 sg13g2_nand2_1 _6486_ (.Y(_1497_),
    .A(_1487_),
    .B(_1283_));
 sg13g2_o21ai_1 _6487_ (.B1(_1497_),
    .Y(_1498_),
    .A1(_1489_),
    .A2(_1496_));
 sg13g2_nor2_1 _6488_ (.A(_1291_),
    .B(_1483_),
    .Y(_1499_));
 sg13g2_inv_1 _6489_ (.Y(_1500_),
    .A(_1499_));
 sg13g2_o21ai_1 _6490_ (.B1(_1500_),
    .Y(_1501_),
    .A1(_1485_),
    .A2(_1498_));
 sg13g2_nand2_1 _6491_ (.Y(_1502_),
    .A(net19),
    .B(_1464_));
 sg13g2_xnor2_1 _6492_ (.Y(_1503_),
    .A(_1371_),
    .B(_1502_));
 sg13g2_nand2_1 _6493_ (.Y(_1504_),
    .A(_1503_),
    .B(_1301_));
 sg13g2_nor2_1 _6494_ (.A(_1301_),
    .B(_1503_),
    .Y(_1505_));
 sg13g2_a21oi_1 _6495_ (.A1(_1501_),
    .A2(_1504_),
    .Y(_1506_),
    .B1(_1505_));
 sg13g2_nor2_1 _6496_ (.A(_1481_),
    .B(_1506_),
    .Y(_1507_));
 sg13g2_nand2_1 _6497_ (.Y(_1508_),
    .A(_1480_),
    .B(_1264_));
 sg13g2_nor2b_1 _6498_ (.A(_1507_),
    .B_N(_1508_),
    .Y(_1509_));
 sg13g2_nor2_1 _6499_ (.A(_1467_),
    .B(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ),
    .Y(_1510_));
 sg13g2_xnor2_1 _6500_ (.Y(_1511_),
    .A(_1398_),
    .B(_1510_));
 sg13g2_nand2_1 _6501_ (.Y(_1512_),
    .A(_1511_),
    .B(_1311_));
 sg13g2_nor2_1 _6502_ (.A(_1311_),
    .B(_1511_),
    .Y(_1513_));
 sg13g2_a221oi_1 _6503_ (.B2(_1512_),
    .C1(_1513_),
    .B1(_1509_),
    .A1(_1258_),
    .Y(_1514_),
    .A2(_1477_));
 sg13g2_nor2_1 _6504_ (.A(_1478_),
    .B(_1514_),
    .Y(_1515_));
 sg13g2_nand2b_1 _6505_ (.Y(_1516_),
    .B(_1515_),
    .A_N(_1475_));
 sg13g2_nand2b_1 _6506_ (.Y(_1517_),
    .B(_1413_),
    .A_N(_1470_));
 sg13g2_nand3b_1 _6507_ (.B(_1516_),
    .C(_1517_),
    .Y(_1518_),
    .A_N(_1474_));
 sg13g2_nand2b_1 _6508_ (.Y(_1519_),
    .B(_1470_),
    .A_N(_1413_));
 sg13g2_and2_1 _6509_ (.A(_1518_),
    .B(_1519_),
    .X(_1520_));
 sg13g2_xor2_1 _6510_ (.B(_1520_),
    .A(_1471_),
    .X(_1521_));
 sg13g2_inv_1 _6511_ (.Y(_1522_),
    .A(_1521_));
 sg13g2_nand2b_1 _6512_ (.Y(_1523_),
    .B(_1444_),
    .A_N(_1446_));
 sg13g2_o21ai_1 _6513_ (.B1(_1419_),
    .Y(_1524_),
    .A1(_1418_),
    .A2(_1402_));
 sg13g2_xor2_1 _6514_ (.B(_1524_),
    .A(_1523_),
    .X(_1525_));
 sg13g2_inv_1 _6515_ (.Y(_1526_),
    .A(_1525_));
 sg13g2_xor2_1 _6516_ (.B(_1348_),
    .A(_1350_),
    .X(_1527_));
 sg13g2_nor2_1 _6517_ (.A(_1457_),
    .B(_1527_),
    .Y(_1528_));
 sg13g2_inv_1 _6518_ (.Y(_1529_),
    .A(_1528_));
 sg13g2_xor2_1 _6519_ (.B(_1352_),
    .A(_1359_),
    .X(_1530_));
 sg13g2_nor2_1 _6520_ (.A(_1529_),
    .B(_1530_),
    .Y(_1531_));
 sg13g2_inv_1 _6521_ (.Y(_1532_),
    .A(_1531_));
 sg13g2_nand2_1 _6522_ (.Y(_1533_),
    .A(_1372_),
    .B(_1375_));
 sg13g2_xnor2_1 _6523_ (.Y(_1534_),
    .A(_1533_),
    .B(_1361_));
 sg13g2_nor2b_1 _6524_ (.A(_1532_),
    .B_N(_1534_),
    .Y(_1535_));
 sg13g2_inv_1 _6525_ (.Y(_1536_),
    .A(_1535_));
 sg13g2_nand2b_1 _6526_ (.Y(_1537_),
    .B(_1378_),
    .A_N(_1317_));
 sg13g2_xor2_1 _6527_ (.B(_1376_),
    .A(_1537_),
    .X(_1538_));
 sg13g2_nor2b_1 _6528_ (.A(_1536_),
    .B_N(_1538_),
    .Y(_1539_));
 sg13g2_inv_1 _6529_ (.Y(_1540_),
    .A(_1539_));
 sg13g2_nand2_1 _6530_ (.Y(_1541_),
    .A(_1399_),
    .B(_1401_));
 sg13g2_xnor2_1 _6531_ (.Y(_1542_),
    .A(_1541_),
    .B(_1379_));
 sg13g2_nor2_1 _6532_ (.A(_1540_),
    .B(_1542_),
    .Y(_1543_));
 sg13g2_inv_1 _6533_ (.Y(_1544_),
    .A(_1543_));
 sg13g2_xor2_1 _6534_ (.B(_1402_),
    .A(_1420_),
    .X(_1545_));
 sg13g2_nor2_1 _6535_ (.A(_1544_),
    .B(_1545_),
    .Y(_1546_));
 sg13g2_nand3_1 _6536_ (.B(_1526_),
    .C(_1546_),
    .A(net13),
    .Y(_1547_));
 sg13g2_buf_1 _6537_ (.A(_1547_),
    .X(_1548_));
 sg13g2_xnor2_1 _6538_ (.Y(_1549_),
    .A(_1522_),
    .B(_1548_));
 sg13g2_and2_1 _6539_ (.A(_1517_),
    .B(_1519_),
    .X(_1550_));
 sg13g2_xnor2_1 _6540_ (.Y(_1551_),
    .A(_1550_),
    .B(_1518_));
 sg13g2_inv_1 _6541_ (.Y(_1552_),
    .A(_1551_));
 sg13g2_xnor2_1 _6542_ (.Y(_1553_),
    .A(_1552_),
    .B(_1548_));
 sg13g2_xnor2_1 _6543_ (.Y(_1554_),
    .A(_1475_),
    .B(_1515_));
 sg13g2_xnor2_1 _6544_ (.Y(_1555_),
    .A(_1554_),
    .B(_1548_));
 sg13g2_nand2_1 _6545_ (.Y(_1556_),
    .A(_1553_),
    .B(_1555_));
 sg13g2_nor2b_1 _6546_ (.A(_1513_),
    .B_N(_1512_),
    .Y(_1557_));
 sg13g2_xor2_1 _6547_ (.B(_1509_),
    .A(_1557_),
    .X(_1558_));
 sg13g2_inv_1 _6548_ (.Y(_1559_),
    .A(_1558_));
 sg13g2_nand2_1 _6549_ (.Y(_1560_),
    .A(net13),
    .B(_1544_));
 sg13g2_xnor2_1 _6550_ (.Y(_1561_),
    .A(_1545_),
    .B(_1560_));
 sg13g2_nor2_1 _6551_ (.A(_1559_),
    .B(_1561_),
    .Y(_1562_));
 sg13g2_xnor2_1 _6552_ (.Y(_1563_),
    .A(_1488_),
    .B(_1496_));
 sg13g2_buf_1 _6553_ (.A(_1563_),
    .X(_1564_));
 sg13g2_inv_1 _6554_ (.Y(_1565_),
    .A(_1564_));
 sg13g2_inv_1 _6555_ (.Y(_1566_),
    .A(_1530_));
 sg13g2_nand2_1 _6556_ (.Y(_1567_),
    .A(_1452_),
    .B(_1529_));
 sg13g2_xnor2_1 _6557_ (.Y(_1568_),
    .A(_1566_),
    .B(_1567_));
 sg13g2_xnor2_1 _6558_ (.Y(_1569_),
    .A(_1565_),
    .B(_1568_));
 sg13g2_inv_1 _6559_ (.Y(_1570_),
    .A(_1569_));
 sg13g2_xnor2_1 _6560_ (.Y(_1571_),
    .A(_1493_),
    .B(_1494_));
 sg13g2_inv_1 _6561_ (.Y(_1572_),
    .A(_1527_));
 sg13g2_nand2_1 _6562_ (.Y(_1573_),
    .A(_1452_),
    .B(_1457_));
 sg13g2_xnor2_1 _6563_ (.Y(_1574_),
    .A(_1572_),
    .B(_1573_));
 sg13g2_nor2b_1 _6564_ (.A(_1571_),
    .B_N(_1574_),
    .Y(_1575_));
 sg13g2_xor2_1 _6565_ (.B(_1574_),
    .A(_1571_),
    .X(_1576_));
 sg13g2_nand2_1 _6566_ (.Y(_1577_),
    .A(_1457_),
    .B(_1455_));
 sg13g2_nor2b_1 _6567_ (.A(_1576_),
    .B_N(_1577_),
    .Y(_1578_));
 sg13g2_nor2_1 _6568_ (.A(_1575_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_nand2_1 _6569_ (.Y(_1580_),
    .A(_1568_),
    .B(_1564_));
 sg13g2_o21ai_1 _6570_ (.B1(_1580_),
    .Y(_1581_),
    .A1(_1570_),
    .A2(_1579_));
 sg13g2_nand2_1 _6571_ (.Y(_1582_),
    .A(_1452_),
    .B(_1532_));
 sg13g2_xnor2_1 _6572_ (.Y(_1583_),
    .A(_1534_),
    .B(_1582_));
 sg13g2_nor2_1 _6573_ (.A(_1499_),
    .B(_1485_),
    .Y(_1584_));
 sg13g2_xor2_1 _6574_ (.B(_1498_),
    .A(_1584_),
    .X(_1585_));
 sg13g2_inv_1 _6575_ (.Y(_1586_),
    .A(_1585_));
 sg13g2_nand2b_1 _6576_ (.Y(_1587_),
    .B(_1586_),
    .A_N(_1583_));
 sg13g2_nand2_1 _6577_ (.Y(_1588_),
    .A(_1583_),
    .B(_1585_));
 sg13g2_inv_1 _6578_ (.Y(_1589_),
    .A(_1588_));
 sg13g2_a21oi_1 _6579_ (.A1(_1581_),
    .A2(_1587_),
    .Y(_1590_),
    .B1(_1589_));
 sg13g2_nand2_1 _6580_ (.Y(_1591_),
    .A(_1452_),
    .B(_1536_));
 sg13g2_xnor2_1 _6581_ (.Y(_1592_),
    .A(_1538_),
    .B(_1591_));
 sg13g2_nor2b_1 _6582_ (.A(_1505_),
    .B_N(_1504_),
    .Y(_1593_));
 sg13g2_xor2_1 _6583_ (.B(_1501_),
    .A(_1593_),
    .X(_1594_));
 sg13g2_inv_1 _6584_ (.Y(_1595_),
    .A(_1594_));
 sg13g2_nand2_1 _6585_ (.Y(_1596_),
    .A(_1592_),
    .B(_1595_));
 sg13g2_nor2_1 _6586_ (.A(_1595_),
    .B(_1592_),
    .Y(_1597_));
 sg13g2_a21oi_1 _6587_ (.A1(_1590_),
    .A2(_1596_),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_nor2b_1 _6588_ (.A(_1481_),
    .B_N(_1508_),
    .Y(_1599_));
 sg13g2_xor2_1 _6589_ (.B(_1506_),
    .A(_1599_),
    .X(_1600_));
 sg13g2_nand2_1 _6590_ (.Y(_1601_),
    .A(net13),
    .B(_1540_));
 sg13g2_xor2_1 _6591_ (.B(_1601_),
    .A(_1542_),
    .X(_1602_));
 sg13g2_nor2_1 _6592_ (.A(_1600_),
    .B(_1602_),
    .Y(_1603_));
 sg13g2_inv_1 _6593_ (.Y(_1604_),
    .A(_1603_));
 sg13g2_nand2_1 _6594_ (.Y(_1605_),
    .A(_1602_),
    .B(_1600_));
 sg13g2_inv_1 _6595_ (.Y(_1606_),
    .A(_1605_));
 sg13g2_a21oi_1 _6596_ (.A1(_1598_),
    .A2(_1604_),
    .Y(_1607_),
    .B1(_1606_));
 sg13g2_inv_1 _6597_ (.Y(_1608_),
    .A(_1607_));
 sg13g2_nand2_1 _6598_ (.Y(_1609_),
    .A(_1561_),
    .B(_1559_));
 sg13g2_o21ai_1 _6599_ (.B1(_1609_),
    .Y(_1610_),
    .A1(_1562_),
    .A2(_1608_));
 sg13g2_inv_1 _6600_ (.Y(_1611_),
    .A(_1610_));
 sg13g2_nor2_1 _6601_ (.A(_1546_),
    .B(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ),
    .Y(_1612_));
 sg13g2_xnor2_1 _6602_ (.Y(_1613_),
    .A(_1526_),
    .B(_1612_));
 sg13g2_xor2_1 _6603_ (.B(_1477_),
    .A(_1258_),
    .X(_1614_));
 sg13g2_nor2_1 _6604_ (.A(_1481_),
    .B(_1513_),
    .Y(_1615_));
 sg13g2_nand2_1 _6605_ (.Y(_1616_),
    .A(_1506_),
    .B(_1599_));
 sg13g2_a22oi_1 _6606_ (.Y(_1617_),
    .B1(_1615_),
    .B2(_1616_),
    .A2(_1511_),
    .A1(_1311_));
 sg13g2_xor2_1 _6607_ (.B(_1617_),
    .A(_1614_),
    .X(_1618_));
 sg13g2_inv_1 _6608_ (.Y(_1619_),
    .A(_1618_));
 sg13g2_nand2_1 _6609_ (.Y(_1620_),
    .A(_1613_),
    .B(_1619_));
 sg13g2_nor2_1 _6610_ (.A(_1619_),
    .B(_1613_),
    .Y(_1621_));
 sg13g2_a21oi_1 _6611_ (.A1(_1611_),
    .A2(_1620_),
    .Y(_1622_),
    .B1(_1621_));
 sg13g2_inv_1 _6612_ (.Y(_1623_),
    .A(_1554_));
 sg13g2_a21o_1 _6613_ (.A2(_1623_),
    .A1(_1551_),
    .B1(_1548_),
    .X(_1624_));
 sg13g2_o21ai_1 _6614_ (.B1(_1624_),
    .Y(_1625_),
    .A1(_1556_),
    .A2(_1622_));
 sg13g2_xnor2_1 _6615_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[10] ),
    .A(_1549_),
    .B(_1625_));
 sg13g2_xnor2_1 _6616_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[1] ),
    .A(_1577_),
    .B(_1576_));
 sg13g2_xnor2_1 _6617_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[2] ),
    .A(_1569_),
    .B(_1579_));
 sg13g2_nand2_1 _6618_ (.Y(_1626_),
    .A(_1587_),
    .B(_1588_));
 sg13g2_xnor2_1 _6619_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[3] ),
    .A(_1626_),
    .B(_1581_));
 sg13g2_nor2b_1 _6620_ (.A(_1597_),
    .B_N(_1596_),
    .Y(_1627_));
 sg13g2_xnor2_1 _6621_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[4] ),
    .A(_1627_),
    .B(_1590_));
 sg13g2_nand2_1 _6622_ (.Y(_1628_),
    .A(_1604_),
    .B(_1605_));
 sg13g2_xnor2_1 _6623_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[5] ),
    .A(_1628_),
    .B(_1598_));
 sg13g2_nor2b_1 _6624_ (.A(_1562_),
    .B_N(_1609_),
    .Y(_1629_));
 sg13g2_xnor2_1 _6625_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[6] ),
    .A(_1629_),
    .B(_1607_));
 sg13g2_nor2b_1 _6626_ (.A(_1621_),
    .B_N(_1620_),
    .Y(_1630_));
 sg13g2_xnor2_1 _6627_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[7] ),
    .A(_1630_),
    .B(_1610_));
 sg13g2_xnor2_1 _6628_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[8] ),
    .A(_1555_),
    .B(_1622_));
 sg13g2_a21oi_1 _6629_ (.A1(_1548_),
    .A2(_1623_),
    .Y(_1631_),
    .B1(_1622_));
 sg13g2_xor2_1 _6630_ (.B(_1631_),
    .A(_1553_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[9] ));
 sg13g2_xnor2_1 _6631_ (.Y(_1632_),
    .A(_1492_),
    .B(_1271_));
 sg13g2_xor2_1 _6632_ (.B(_1564_),
    .A(_1632_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_nor2_1 _6633_ (.A(_1564_),
    .B(_1585_),
    .Y(_1633_));
 sg13g2_inv_1 _6634_ (.Y(_1634_),
    .A(_1633_));
 sg13g2_nor2_1 _6635_ (.A(_1634_),
    .B(_1595_),
    .Y(_1635_));
 sg13g2_inv_1 _6636_ (.Y(_1636_),
    .A(_1635_));
 sg13g2_nor2_1 _6637_ (.A(_1636_),
    .B(_1600_),
    .Y(_1637_));
 sg13g2_inv_1 _6638_ (.Y(_1638_),
    .A(_1637_));
 sg13g2_nor2_1 _6639_ (.A(_1638_),
    .B(_1558_),
    .Y(_1639_));
 sg13g2_inv_1 _6640_ (.Y(_1640_),
    .A(_1639_));
 sg13g2_nor2_1 _6641_ (.A(_1618_),
    .B(_1640_),
    .Y(_1641_));
 sg13g2_inv_1 _6642_ (.Y(_1642_),
    .A(_1641_));
 sg13g2_nor2_1 _6643_ (.A(_1642_),
    .B(_1554_),
    .Y(_1643_));
 sg13g2_inv_1 _6644_ (.Y(_1644_),
    .A(_1643_));
 sg13g2_nor2_1 _6645_ (.A(_1644_),
    .B(_1552_),
    .Y(_1645_));
 sg13g2_a21oi_1 _6646_ (.A1(_1645_),
    .A2(net13),
    .Y(_1646_),
    .B1(_1521_));
 sg13g2_o21ai_1 _6647_ (.B1(net13),
    .Y(_1647_),
    .A1(_1644_),
    .A2(_1552_));
 sg13g2_nand2_1 _6648_ (.Y(_1648_),
    .A(_1647_),
    .B(_1522_));
 sg13g2_o21ai_1 _6649_ (.B1(_1648_),
    .Y(_1649_),
    .A1(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ),
    .A2(_1522_));
 sg13g2_inv_1 _6650_ (.Y(_1650_),
    .A(_1545_));
 sg13g2_xnor2_1 _6651_ (.Y(_1651_),
    .A(_1522_),
    .B(_1647_));
 sg13g2_nor2_1 _6652_ (.A(_1650_),
    .B(_1651_),
    .Y(_1652_));
 sg13g2_nor2_1 _6653_ (.A(_1526_),
    .B(_1649_),
    .Y(_1653_));
 sg13g2_nor2_1 _6654_ (.A(_1652_),
    .B(_1653_),
    .Y(_1654_));
 sg13g2_inv_1 _6655_ (.Y(_1655_),
    .A(_1652_));
 sg13g2_nand2_1 _6656_ (.Y(_1656_),
    .A(_1651_),
    .B(_1650_));
 sg13g2_nand2_1 _6657_ (.Y(_1657_),
    .A(_1655_),
    .B(_1656_));
 sg13g2_a21oi_1 _6658_ (.A1(_1552_),
    .A2(_1644_),
    .Y(_1658_),
    .B1(_1647_));
 sg13g2_a21o_1 _6659_ (.A2(_1552_),
    .A1(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ),
    .B1(_1658_),
    .X(_1659_));
 sg13g2_nor2_1 _6660_ (.A(_1542_),
    .B(_1659_),
    .Y(_1660_));
 sg13g2_nand2_1 _6661_ (.Y(_1661_),
    .A(net13),
    .B(_1642_));
 sg13g2_xnor2_1 _6662_ (.Y(_1662_),
    .A(_1623_),
    .B(_1661_));
 sg13g2_nor2_1 _6663_ (.A(_1538_),
    .B(_1662_),
    .Y(_1663_));
 sg13g2_nand2_1 _6664_ (.Y(_1664_),
    .A(_1659_),
    .B(_1542_));
 sg13g2_inv_1 _6665_ (.Y(_1665_),
    .A(_1664_));
 sg13g2_nand2_1 _6666_ (.Y(_1666_),
    .A(net13),
    .B(_1638_));
 sg13g2_xnor2_1 _6667_ (.Y(_1667_),
    .A(_1559_),
    .B(_1666_));
 sg13g2_nor2_1 _6668_ (.A(_1566_),
    .B(_1667_),
    .Y(_1668_));
 sg13g2_nand2_1 _6669_ (.Y(_1669_),
    .A(_1452_),
    .B(_1564_));
 sg13g2_xnor2_1 _6670_ (.Y(_1670_),
    .A(_1586_),
    .B(_1669_));
 sg13g2_xnor2_1 _6671_ (.Y(_1671_),
    .A(_1343_),
    .B(_1341_));
 sg13g2_nor2b_1 _6672_ (.A(_1670_),
    .B_N(_1671_),
    .Y(_1672_));
 sg13g2_nand2_1 _6673_ (.Y(_1673_),
    .A(_1564_),
    .B(_1632_));
 sg13g2_xor2_1 _6674_ (.B(_1670_),
    .A(_1671_),
    .X(_1674_));
 sg13g2_nor2_1 _6675_ (.A(_1673_),
    .B(_1674_),
    .Y(_1675_));
 sg13g2_nor2_1 _6676_ (.A(_1672_),
    .B(_1675_),
    .Y(_1676_));
 sg13g2_inv_1 _6677_ (.Y(_1677_),
    .A(_1676_));
 sg13g2_nand2_1 _6678_ (.Y(_1678_),
    .A(_1452_),
    .B(_1634_));
 sg13g2_xnor2_1 _6679_ (.Y(_1679_),
    .A(_1594_),
    .B(_1678_));
 sg13g2_inv_1 _6680_ (.Y(_1680_),
    .A(_1457_));
 sg13g2_nand2_1 _6681_ (.Y(_1681_),
    .A(_1679_),
    .B(_1680_));
 sg13g2_nor2_1 _6682_ (.A(_1680_),
    .B(_1679_),
    .Y(_1682_));
 sg13g2_a21oi_1 _6683_ (.A1(_1677_),
    .A2(_1681_),
    .Y(_1683_),
    .B1(_1682_));
 sg13g2_inv_1 _6684_ (.Y(_1684_),
    .A(_1683_));
 sg13g2_nand2_1 _6685_ (.Y(_1685_),
    .A(_1452_),
    .B(_1636_));
 sg13g2_xor2_1 _6686_ (.B(_1685_),
    .A(_1600_),
    .X(_1686_));
 sg13g2_nand2_1 _6687_ (.Y(_1687_),
    .A(_1686_),
    .B(_1572_));
 sg13g2_nor2_1 _6688_ (.A(_1572_),
    .B(_1686_),
    .Y(_1688_));
 sg13g2_a21oi_1 _6689_ (.A1(_1684_),
    .A2(_1687_),
    .Y(_1689_),
    .B1(_1688_));
 sg13g2_inv_1 _6690_ (.Y(_1690_),
    .A(_1689_));
 sg13g2_nand2_1 _6691_ (.Y(_1691_),
    .A(_1667_),
    .B(_1566_));
 sg13g2_o21ai_1 _6692_ (.B1(_1691_),
    .Y(_1692_),
    .A1(_1668_),
    .A2(_1690_));
 sg13g2_nand2_1 _6693_ (.Y(_1693_),
    .A(_1453_),
    .B(_1640_));
 sg13g2_xnor2_1 _6694_ (.Y(_1694_),
    .A(_1619_),
    .B(_1693_));
 sg13g2_nand2_1 _6695_ (.Y(_1695_),
    .A(_1694_),
    .B(_1534_));
 sg13g2_nand2b_1 _6696_ (.Y(_1696_),
    .B(_1695_),
    .A_N(_1692_));
 sg13g2_nor2_1 _6697_ (.A(_1534_),
    .B(_1694_),
    .Y(_1697_));
 sg13g2_inv_1 _6698_ (.Y(_1698_),
    .A(_1697_));
 sg13g2_nand2_1 _6699_ (.Y(_1699_),
    .A(_1662_),
    .B(_1538_));
 sg13g2_nand2b_1 _6700_ (.Y(_1700_),
    .B(_1699_),
    .A_N(_1663_));
 sg13g2_a21oi_1 _6701_ (.A1(_1696_),
    .A2(_1698_),
    .Y(_1701_),
    .B1(_1700_));
 sg13g2_nor3_1 _6702_ (.A(_1663_),
    .B(_1665_),
    .C(_1701_),
    .Y(_1702_));
 sg13g2_nor2_1 _6703_ (.A(_1660_),
    .B(_1702_),
    .Y(_1703_));
 sg13g2_nand2b_1 _6704_ (.Y(_1704_),
    .B(_1703_),
    .A_N(_1657_));
 sg13g2_a22oi_1 _6705_ (.Y(_1705_),
    .B1(_1654_),
    .B2(_1704_),
    .A2(_1649_),
    .A1(_1526_));
 sg13g2_xor2_1 _6706_ (.B(_1705_),
    .A(_1646_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[10] ));
 sg13g2_xor2_1 _6707_ (.B(_1674_),
    .A(_1673_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[1] ));
 sg13g2_nor2b_1 _6708_ (.A(_1682_),
    .B_N(_1681_),
    .Y(_1706_));
 sg13g2_xnor2_1 _6709_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[2] ),
    .A(_1706_),
    .B(_1676_));
 sg13g2_nor2b_1 _6710_ (.A(_1688_),
    .B_N(_1687_),
    .Y(_1707_));
 sg13g2_xnor2_1 _6711_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[3] ),
    .A(_1707_),
    .B(_1683_));
 sg13g2_nor2b_1 _6712_ (.A(_1668_),
    .B_N(_1691_),
    .Y(_1708_));
 sg13g2_xnor2_1 _6713_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[4] ),
    .A(_1708_),
    .B(_1689_));
 sg13g2_nand2_1 _6714_ (.Y(_1709_),
    .A(_1698_),
    .B(_1695_));
 sg13g2_xor2_1 _6715_ (.B(_1692_),
    .A(_1709_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_nand2_1 _6716_ (.Y(_1710_),
    .A(_1696_),
    .B(_1698_));
 sg13g2_xnor2_1 _6717_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[6] ),
    .A(_1700_),
    .B(_1710_));
 sg13g2_nor2_1 _6718_ (.A(_1660_),
    .B(_1665_),
    .Y(_1711_));
 sg13g2_a21oi_1 _6719_ (.A1(_1710_),
    .A2(_1699_),
    .Y(_1712_),
    .B1(_1663_));
 sg13g2_xnor2_1 _6720_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[7] ),
    .A(_1711_),
    .B(_1712_));
 sg13g2_xnor2_1 _6721_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[8] ),
    .A(_1657_),
    .B(_1703_));
 sg13g2_xnor2_1 _6722_ (.Y(_1713_),
    .A(_1525_),
    .B(_1649_));
 sg13g2_nand2_1 _6723_ (.Y(_1714_),
    .A(_1664_),
    .B(_1655_));
 sg13g2_nor2b_1 _6724_ (.A(_1712_),
    .B_N(_1711_),
    .Y(_1715_));
 sg13g2_o21ai_1 _6725_ (.B1(_1656_),
    .Y(_1716_),
    .A1(_1714_),
    .A2(_1715_));
 sg13g2_xnor2_1 _6726_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[9] ),
    .A(_1713_),
    .B(_1716_));
 sg13g2_buf_1 _6727_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[10] ),
    .X(_1717_));
 sg13g2_buf_1 _6728_ (.A(_1717_),
    .X(_1718_));
 sg13g2_buf_1 _6729_ (.A(_1718_),
    .X(_1719_));
 sg13g2_xor2_1 _6730_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ),
    .A(net56),
    .X(_1720_));
 sg13g2_buf_1 _6731_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .X(_1721_));
 sg13g2_buf_1 _6732_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ),
    .X(_1722_));
 sg13g2_buf_1 _6733_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .X(_1723_));
 sg13g2_nor2_1 _6734_ (.A(_1723_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ),
    .Y(_1724_));
 sg13g2_inv_1 _6735_ (.Y(_1725_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ));
 sg13g2_nand2_1 _6736_ (.Y(_1726_),
    .A(_1724_),
    .B(_1725_));
 sg13g2_nor2_1 _6737_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ),
    .B(_1726_),
    .Y(_1727_));
 sg13g2_inv_1 _6738_ (.Y(_1728_),
    .A(_1727_));
 sg13g2_nor2_1 _6739_ (.A(_1722_),
    .B(_1728_),
    .Y(_1729_));
 sg13g2_inv_1 _6740_ (.Y(_1730_),
    .A(_1729_));
 sg13g2_nor3_1 _6741_ (.A(_1721_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .C(_1730_),
    .Y(_1731_));
 sg13g2_inv_1 _6742_ (.Y(_1732_),
    .A(_1717_));
 sg13g2_buf_1 _6743_ (.A(_1732_),
    .X(_1733_));
 sg13g2_buf_1 _6744_ (.A(_1733_),
    .X(_1734_));
 sg13g2_a21oi_1 _6745_ (.A1(_1731_),
    .A2(net48),
    .Y(_1735_),
    .B1(\main.demo._q___pip_58_1_2___stage___block_3_cx[10] ));
 sg13g2_inv_1 _6746_ (.Y(_1736_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_nand3_1 _6747_ (.B(_1736_),
    .C(_0049_),
    .A(_1725_),
    .Y(_1737_));
 sg13g2_nor2_1 _6748_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ),
    .B(_1737_),
    .Y(_1738_));
 sg13g2_inv_1 _6749_ (.Y(_1739_),
    .A(_1738_));
 sg13g2_nor3_1 _6750_ (.A(_1722_),
    .B(_1721_),
    .C(_1739_),
    .Y(_1740_));
 sg13g2_inv_1 _6751_ (.Y(_1741_),
    .A(_1740_));
 sg13g2_nor2_1 _6752_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .B(_1741_),
    .Y(_1742_));
 sg13g2_inv_1 _6753_ (.Y(_1743_),
    .A(_1742_));
 sg13g2_nor2b_1 _6754_ (.A(net64),
    .B_N(\main.demo._q___pip_58_1_2___stage___block_3_cx[10] ),
    .Y(_1744_));
 sg13g2_a21oi_1 _6755_ (.A1(net64),
    .A2(_0063_),
    .Y(_1745_),
    .B1(_1744_));
 sg13g2_o21ai_1 _6756_ (.B1(_1745_),
    .Y(_1746_),
    .A1(net56),
    .A2(_1743_));
 sg13g2_buf_1 _6757_ (.A(_1746_),
    .X(_1747_));
 sg13g2_inv_1 _6758_ (.Y(_1748_),
    .A(_1731_));
 sg13g2_o21ai_1 _6759_ (.B1(_1745_),
    .Y(_1749_),
    .A1(net56),
    .A2(_1748_));
 sg13g2_inv_1 _6760_ (.Y(_1750_),
    .A(_0054_));
 sg13g2_o21ai_1 _6761_ (.B1(_1721_),
    .Y(_1751_),
    .A1(_1722_),
    .A2(_1739_));
 sg13g2_nor2_1 _6762_ (.A(net64),
    .B(_1740_),
    .Y(_1752_));
 sg13g2_a22oi_1 _6763_ (.Y(_1753_),
    .B1(_1751_),
    .B2(_1752_),
    .A2(_1750_),
    .A1(net64));
 sg13g2_inv_1 _6764_ (.Y(_1754_),
    .A(_0046_));
 sg13g2_nand2_1 _6765_ (.Y(_1755_),
    .A(_1728_),
    .B(_1722_));
 sg13g2_nor2_1 _6766_ (.A(net64),
    .B(_1729_),
    .Y(_1756_));
 sg13g2_a22oi_1 _6767_ (.Y(_1757_),
    .B1(_1755_),
    .B2(_1756_),
    .A2(net64),
    .A1(_1754_));
 sg13g2_nand2_1 _6768_ (.Y(_1758_),
    .A(_1737_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ));
 sg13g2_a21oi_1 _6769_ (.A1(_1739_),
    .A2(_1758_),
    .Y(_1759_),
    .B1(_1717_));
 sg13g2_a21o_1 _6770_ (.A2(_0048_),
    .A1(_1718_),
    .B1(_1759_),
    .X(_1760_));
 sg13g2_inv_1 _6771_ (.Y(_1761_),
    .A(_1724_));
 sg13g2_nand2_1 _6772_ (.Y(_1762_),
    .A(_1761_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ));
 sg13g2_nand3_1 _6773_ (.B(_1733_),
    .C(_1726_),
    .A(_1762_),
    .Y(_1763_));
 sg13g2_o21ai_1 _6774_ (.B1(_1763_),
    .Y(_1764_),
    .A1(net55),
    .A2(_0050_));
 sg13g2_xnor2_1 _6775_ (.Y(_1765_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[2] ),
    .B(_1764_));
 sg13g2_nand2_1 _6776_ (.Y(_1766_),
    .A(_1723_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_nand3_1 _6777_ (.B(_1732_),
    .C(_1766_),
    .A(_1761_),
    .Y(_1767_));
 sg13g2_o21ai_1 _6778_ (.B1(_1767_),
    .Y(_1768_),
    .A1(net55),
    .A2(_0051_));
 sg13g2_nand2_1 _6779_ (.Y(_1769_),
    .A(_1723_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ));
 sg13g2_xor2_1 _6780_ (.B(_1768_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[1] ),
    .X(_1770_));
 sg13g2_nor2b_1 _6781_ (.A(_1769_),
    .B_N(_1770_),
    .Y(_1771_));
 sg13g2_a21oi_1 _6782_ (.A1(\main.demo._q___pip_58_1_2___stage___block_3_cy[1] ),
    .A2(_1768_),
    .Y(_1772_),
    .B1(_1771_));
 sg13g2_nand2_1 _6783_ (.Y(_1773_),
    .A(_1764_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[2] ));
 sg13g2_o21ai_1 _6784_ (.B1(_1773_),
    .Y(_1774_),
    .A1(_1765_),
    .A2(_1772_));
 sg13g2_buf_1 _6785_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .X(_1775_));
 sg13g2_xnor2_1 _6786_ (.Y(_1776_),
    .A(_1775_),
    .B(_1760_));
 sg13g2_nand2_1 _6787_ (.Y(_1777_),
    .A(_1774_),
    .B(_1776_));
 sg13g2_o21ai_1 _6788_ (.B1(_1777_),
    .Y(_1778_),
    .A1(_0047_),
    .A2(_1760_));
 sg13g2_buf_1 _6789_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ),
    .X(_1779_));
 sg13g2_xnor2_1 _6790_ (.Y(_1780_),
    .A(_1779_),
    .B(_1757_));
 sg13g2_nand2_1 _6791_ (.Y(_1781_),
    .A(_1778_),
    .B(_1780_));
 sg13g2_o21ai_1 _6792_ (.B1(_1781_),
    .Y(_1782_),
    .A1(_0062_),
    .A2(_1757_));
 sg13g2_buf_1 _6793_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ),
    .X(_1783_));
 sg13g2_xnor2_1 _6794_ (.Y(_1784_),
    .A(_1783_),
    .B(_1753_));
 sg13g2_nand2_1 _6795_ (.Y(_1785_),
    .A(_1782_),
    .B(_1784_));
 sg13g2_o21ai_1 _6796_ (.B1(_1785_),
    .Y(_1786_),
    .A1(_0061_),
    .A2(_1753_));
 sg13g2_buf_1 _6797_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ),
    .X(_1787_));
 sg13g2_o21ai_1 _6798_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .Y(_1788_),
    .A1(_1721_),
    .A2(_1730_));
 sg13g2_nand3_1 _6799_ (.B(_1748_),
    .C(net48),
    .A(_1788_),
    .Y(_1789_));
 sg13g2_o21ai_1 _6800_ (.B1(_1789_),
    .Y(_1790_),
    .A1(net48),
    .A2(_0052_));
 sg13g2_xor2_1 _6801_ (.B(_1790_),
    .A(_1787_),
    .X(_1791_));
 sg13g2_nor2b_1 _6802_ (.A(_0060_),
    .B_N(_1790_),
    .Y(_1792_));
 sg13g2_a21o_1 _6803_ (.A2(_1791_),
    .A1(_1786_),
    .B1(_1792_),
    .X(_1793_));
 sg13g2_buf_1 _6804_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ),
    .X(_1794_));
 sg13g2_nand2_1 _6805_ (.Y(_1795_),
    .A(_1742_),
    .B(_1744_));
 sg13g2_nand2_1 _6806_ (.Y(_1796_),
    .A(_1747_),
    .B(_1795_));
 sg13g2_xor2_1 _6807_ (.B(_1796_),
    .A(_1794_),
    .X(_1797_));
 sg13g2_a21oi_1 _6808_ (.A1(_1747_),
    .A2(_1795_),
    .Y(_1798_),
    .B1(_0059_));
 sg13g2_a21o_1 _6809_ (.A2(_1797_),
    .A1(_1793_),
    .B1(_1798_),
    .X(_1799_));
 sg13g2_buf_1 _6810_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ),
    .X(_1800_));
 sg13g2_xnor2_1 _6811_ (.Y(_1801_),
    .A(_1800_),
    .B(_1749_));
 sg13g2_nand2_1 _6812_ (.Y(_1802_),
    .A(_1799_),
    .B(_1801_));
 sg13g2_o21ai_1 _6813_ (.B1(_1802_),
    .Y(_1803_),
    .A1(_0058_),
    .A2(_1749_));
 sg13g2_xnor2_1 _6814_ (.Y(_1804_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .B(_1747_));
 sg13g2_nand2_1 _6815_ (.Y(_1805_),
    .A(_1803_),
    .B(_1804_));
 sg13g2_o21ai_1 _6816_ (.B1(_1805_),
    .Y(_1806_),
    .A1(_0057_),
    .A2(_1747_));
 sg13g2_or2_1 _6817_ (.X(_1807_),
    .B(_1806_),
    .A(_1735_));
 sg13g2_nand2_1 _6818_ (.Y(_1808_),
    .A(_1806_),
    .B(_1735_));
 sg13g2_nand2_1 _6819_ (.Y(_1809_),
    .A(_1807_),
    .B(_1808_));
 sg13g2_buf_1 _6820_ (.A(_1809_),
    .X(_1810_));
 sg13g2_buf_1 _6821_ (.A(net21),
    .X(_1811_));
 sg13g2_nor2_1 _6822_ (.A(_0059_),
    .B(net55),
    .Y(_1812_));
 sg13g2_nor2_1 _6823_ (.A(_1775_),
    .B(_1779_),
    .Y(_1813_));
 sg13g2_nand2b_1 _6824_ (.Y(_1814_),
    .B(_1813_),
    .A_N(_1783_));
 sg13g2_nor2_1 _6825_ (.A(_1787_),
    .B(_1814_),
    .Y(_1815_));
 sg13g2_inv_1 _6826_ (.Y(_1816_),
    .A(_1815_));
 sg13g2_nor2_1 _6827_ (.A(_1794_),
    .B(_1816_),
    .Y(_1817_));
 sg13g2_inv_1 _6828_ (.Y(_1818_),
    .A(_1817_));
 sg13g2_nand2_1 _6829_ (.Y(_1819_),
    .A(_1816_),
    .B(_1794_));
 sg13g2_nand3_1 _6830_ (.B(net55),
    .C(_1819_),
    .A(_1818_),
    .Y(_1820_));
 sg13g2_nor2b_1 _6831_ (.A(_1812_),
    .B_N(_1820_),
    .Y(_1821_));
 sg13g2_xnor2_1 _6832_ (.Y(_1822_),
    .A(_0051_),
    .B(_1821_));
 sg13g2_inv_1 _6833_ (.Y(_1823_),
    .A(_0060_));
 sg13g2_inv_1 _6834_ (.Y(_1824_),
    .A(_0047_));
 sg13g2_nor3_1 _6835_ (.A(_1779_),
    .B(_1783_),
    .C(_1824_),
    .Y(_1825_));
 sg13g2_inv_1 _6836_ (.Y(_1826_),
    .A(_1825_));
 sg13g2_nand2_1 _6837_ (.Y(_1827_),
    .A(_1826_),
    .B(_1787_));
 sg13g2_nor2_1 _6838_ (.A(_1787_),
    .B(_1826_),
    .Y(_1828_));
 sg13g2_nor2_1 _6839_ (.A(net64),
    .B(_1828_),
    .Y(_1829_));
 sg13g2_a22oi_1 _6840_ (.Y(_1830_),
    .B1(_1827_),
    .B2(_1829_),
    .A2(_1823_),
    .A1(net64));
 sg13g2_inv_1 _6841_ (.Y(_1831_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[1] ));
 sg13g2_inv_1 _6842_ (.Y(_1832_),
    .A(_1813_));
 sg13g2_nand2_1 _6843_ (.Y(_1833_),
    .A(_1775_),
    .B(_1779_));
 sg13g2_nand3_1 _6844_ (.B(net55),
    .C(_1833_),
    .A(_1832_),
    .Y(_1834_));
 sg13g2_o21ai_1 _6845_ (.B1(_1834_),
    .Y(_1835_),
    .A1(net55),
    .A2(_0062_));
 sg13g2_nor2_1 _6846_ (.A(_1831_),
    .B(_1835_),
    .Y(_1836_));
 sg13g2_nor2b_1 _6847_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[0] ),
    .B_N(_1775_),
    .Y(_1837_));
 sg13g2_xnor2_1 _6848_ (.Y(_1838_),
    .A(_1831_),
    .B(_1835_));
 sg13g2_nor2_1 _6849_ (.A(_1837_),
    .B(_1838_),
    .Y(_1839_));
 sg13g2_nor2_1 _6850_ (.A(_1836_),
    .B(_1839_),
    .Y(_1840_));
 sg13g2_inv_1 _6851_ (.Y(_1841_),
    .A(_1840_));
 sg13g2_nand2_1 _6852_ (.Y(_1842_),
    .A(_1832_),
    .B(_1783_));
 sg13g2_nand3_1 _6853_ (.B(net55),
    .C(_1814_),
    .A(_1842_),
    .Y(_1843_));
 sg13g2_o21ai_1 _6854_ (.B1(_1843_),
    .Y(_1844_),
    .A1(net55),
    .A2(_0061_));
 sg13g2_xnor2_1 _6855_ (.Y(_1845_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[2] ),
    .B(_1844_));
 sg13g2_nor2b_1 _6856_ (.A(_1844_),
    .B_N(\main.demo._q___pip_58_1_2___stage___block_3_cx[2] ),
    .Y(_1846_));
 sg13g2_a21oi_1 _6857_ (.A1(_1841_),
    .A2(_1845_),
    .Y(_1847_),
    .B1(_1846_));
 sg13g2_xnor2_1 _6858_ (.Y(_1848_),
    .A(_0049_),
    .B(_1830_));
 sg13g2_nor2b_1 _6859_ (.A(_1847_),
    .B_N(_1848_),
    .Y(_1849_));
 sg13g2_a21o_1 _6860_ (.A2(_1830_),
    .A1(_1723_),
    .B1(_1849_),
    .X(_1850_));
 sg13g2_xor2_1 _6861_ (.B(_1850_),
    .A(_1822_),
    .X(_1851_));
 sg13g2_inv_1 _6862_ (.Y(_1852_),
    .A(_1828_));
 sg13g2_nor2_1 _6863_ (.A(_1794_),
    .B(_1852_),
    .Y(_1853_));
 sg13g2_xnor2_1 _6864_ (.Y(_1854_),
    .A(_1800_),
    .B(_1853_));
 sg13g2_nor2_1 _6865_ (.A(_0058_),
    .B(net48),
    .Y(_1855_));
 sg13g2_a21oi_1 _6866_ (.A1(_1854_),
    .A2(net48),
    .Y(_1856_),
    .B1(_1855_));
 sg13g2_xnor2_1 _6867_ (.Y(_1857_),
    .A(_0050_),
    .B(_1856_));
 sg13g2_inv_1 _6868_ (.Y(_1858_),
    .A(_1821_));
 sg13g2_nand2_1 _6869_ (.Y(_1859_),
    .A(_1850_),
    .B(_1822_));
 sg13g2_o21ai_1 _6870_ (.B1(_1859_),
    .Y(_1860_),
    .A1(_1736_),
    .A2(_1858_));
 sg13g2_xor2_1 _6871_ (.B(_1860_),
    .A(_1857_),
    .X(_1861_));
 sg13g2_nor2_1 _6872_ (.A(_1851_),
    .B(_1861_),
    .Y(_1862_));
 sg13g2_inv_1 _6873_ (.Y(_1863_),
    .A(_1862_));
 sg13g2_inv_1 _6874_ (.Y(_1864_),
    .A(_0057_));
 sg13g2_nor2_1 _6875_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .B(_1800_),
    .Y(_1865_));
 sg13g2_nor2b_1 _6876_ (.A(_1818_),
    .B_N(_1865_),
    .Y(_1866_));
 sg13g2_nor2_1 _6877_ (.A(net56),
    .B(_1866_),
    .Y(_1867_));
 sg13g2_o21ai_1 _6878_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .Y(_1868_),
    .A1(_1800_),
    .A2(_1818_));
 sg13g2_a22oi_1 _6879_ (.Y(_1869_),
    .B1(_1867_),
    .B2(_1868_),
    .A2(_1864_),
    .A1(net56));
 sg13g2_xnor2_1 _6880_ (.Y(_1870_),
    .A(_0048_),
    .B(_1869_));
 sg13g2_nor2b_1 _6881_ (.A(_1725_),
    .B_N(_1856_),
    .Y(_1871_));
 sg13g2_a21o_1 _6882_ (.A2(_1857_),
    .A1(_1860_),
    .B1(_1871_),
    .X(_1872_));
 sg13g2_xor2_1 _6883_ (.B(_1872_),
    .A(_1870_),
    .X(_1873_));
 sg13g2_nor2_1 _6884_ (.A(_1863_),
    .B(_1873_),
    .Y(_1874_));
 sg13g2_inv_1 _6885_ (.Y(_1875_),
    .A(_1874_));
 sg13g2_nand3_1 _6886_ (.B(_0053_),
    .C(_1865_),
    .A(_1853_),
    .Y(_1876_));
 sg13g2_xor2_1 _6887_ (.B(_1876_),
    .A(_0046_),
    .X(_1877_));
 sg13g2_nand2_1 _6888_ (.Y(_1878_),
    .A(_1872_),
    .B(_1870_));
 sg13g2_nand2_1 _6889_ (.Y(_1879_),
    .A(_1869_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ));
 sg13g2_nand2_1 _6890_ (.Y(_1880_),
    .A(_1878_),
    .B(_1879_));
 sg13g2_xor2_1 _6891_ (.B(_1880_),
    .A(_1877_),
    .X(_1881_));
 sg13g2_nor2_1 _6892_ (.A(_1875_),
    .B(_1881_),
    .Y(_1882_));
 sg13g2_inv_1 _6893_ (.Y(_1883_),
    .A(_1882_));
 sg13g2_nand3_1 _6894_ (.B(net48),
    .C(_0053_),
    .A(_1865_),
    .Y(_1884_));
 sg13g2_nor2_1 _6895_ (.A(_1884_),
    .B(_1818_),
    .Y(_1885_));
 sg13g2_xnor2_1 _6896_ (.Y(_1886_),
    .A(_0054_),
    .B(_1885_));
 sg13g2_inv_1 _6897_ (.Y(_1887_),
    .A(_1722_));
 sg13g2_nand2_1 _6898_ (.Y(_1888_),
    .A(_1880_),
    .B(_1877_));
 sg13g2_o21ai_1 _6899_ (.B1(_1888_),
    .Y(_1889_),
    .A1(_1887_),
    .A2(_1876_));
 sg13g2_xor2_1 _6900_ (.B(_1889_),
    .A(_1886_),
    .X(_1890_));
 sg13g2_nor2_1 _6901_ (.A(_1883_),
    .B(_1890_),
    .Y(_1891_));
 sg13g2_inv_1 _6902_ (.Y(_1892_),
    .A(_1891_));
 sg13g2_xor2_1 _6903_ (.B(_1885_),
    .A(_0052_),
    .X(_1893_));
 sg13g2_nand2_1 _6904_ (.Y(_1894_),
    .A(_1889_),
    .B(_1886_));
 sg13g2_inv_1 _6905_ (.Y(_1895_),
    .A(_1894_));
 sg13g2_a21oi_1 _6906_ (.A1(_1721_),
    .A2(_1885_),
    .Y(_1896_),
    .B1(_1895_));
 sg13g2_nor2_1 _6907_ (.A(_1893_),
    .B(_1896_),
    .Y(_1897_));
 sg13g2_nand2_1 _6908_ (.Y(_1898_),
    .A(_1896_),
    .B(_1893_));
 sg13g2_nor2b_1 _6909_ (.A(_1897_),
    .B_N(_1898_),
    .Y(_1899_));
 sg13g2_buf_1 _6910_ (.A(_1899_),
    .X(_1900_));
 sg13g2_nor2_1 _6911_ (.A(_1892_),
    .B(_1900_),
    .Y(_1901_));
 sg13g2_nand3_1 _6912_ (.B(net48),
    .C(_0053_),
    .A(_1866_),
    .Y(_1902_));
 sg13g2_xor2_1 _6913_ (.B(_1902_),
    .A(_0063_),
    .X(_1903_));
 sg13g2_inv_1 _6914_ (.Y(_1904_),
    .A(_1902_));
 sg13g2_inv_1 _6915_ (.Y(_1905_),
    .A(_1893_));
 sg13g2_and3_1 _6916_ (.X(_1906_),
    .A(_1904_),
    .B(_0052_),
    .C(_1721_));
 sg13g2_a221oi_1 _6917_ (.B2(_1905_),
    .C1(_1906_),
    .B1(_1895_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .Y(_1907_),
    .A2(_1904_));
 sg13g2_xor2_1 _6918_ (.B(_1907_),
    .A(_1903_),
    .X(_1908_));
 sg13g2_inv_1 _6919_ (.Y(_1909_),
    .A(_1908_));
 sg13g2_a21oi_1 _6920_ (.A1(net18),
    .A2(_1901_),
    .Y(_1910_),
    .B1(_1909_));
 sg13g2_nor2_1 _6921_ (.A(_1909_),
    .B(net21),
    .Y(_1911_));
 sg13g2_inv_1 _6922_ (.Y(_1912_),
    .A(_1901_));
 sg13g2_inv_1 _6923_ (.Y(_1913_),
    .A(net21));
 sg13g2_a21oi_1 _6924_ (.A1(_1908_),
    .A2(_1912_),
    .Y(_1914_),
    .B1(net17));
 sg13g2_nor2_1 _6925_ (.A(_1911_),
    .B(_1914_),
    .Y(_1915_));
 sg13g2_buf_1 _6926_ (.A(_1915_),
    .X(_1916_));
 sg13g2_inv_1 _6927_ (.Y(_1917_),
    .A(_1916_));
 sg13g2_xor2_1 _6928_ (.B(_1803_),
    .A(_1804_),
    .X(_1918_));
 sg13g2_inv_1 _6929_ (.Y(_1919_),
    .A(_1918_));
 sg13g2_xor2_1 _6930_ (.B(_1799_),
    .A(_1801_),
    .X(_1920_));
 sg13g2_o21ai_1 _6931_ (.B1(_1916_),
    .Y(_1921_),
    .A1(_1918_),
    .A2(_1920_));
 sg13g2_xor2_1 _6932_ (.B(_1782_),
    .A(_1784_),
    .X(_1922_));
 sg13g2_nand2_1 _6933_ (.Y(_1923_),
    .A(net21),
    .B(_1892_));
 sg13g2_xnor2_1 _6934_ (.Y(_1924_),
    .A(_1900_),
    .B(_1923_));
 sg13g2_nor2_1 _6935_ (.A(_1922_),
    .B(_1924_),
    .Y(_1925_));
 sg13g2_xor2_1 _6936_ (.B(_1778_),
    .A(_1780_),
    .X(_1926_));
 sg13g2_buf_1 _6937_ (.A(_1926_),
    .X(_1927_));
 sg13g2_a21oi_1 _6938_ (.A1(_1890_),
    .A2(_1883_),
    .Y(_1928_),
    .B1(_1923_));
 sg13g2_a21o_1 _6939_ (.A2(_1890_),
    .A1(net17),
    .B1(_1928_),
    .X(_1929_));
 sg13g2_xor2_1 _6940_ (.B(_1774_),
    .A(_1776_),
    .X(_1930_));
 sg13g2_nand2_1 _6941_ (.Y(_1931_),
    .A(net21),
    .B(_1875_));
 sg13g2_xnor2_1 _6942_ (.Y(_1932_),
    .A(_1881_),
    .B(_1931_));
 sg13g2_nor2_1 _6943_ (.A(_1930_),
    .B(_1932_),
    .Y(_1933_));
 sg13g2_inv_1 _6944_ (.Y(_1934_),
    .A(_1873_));
 sg13g2_nand2_1 _6945_ (.Y(_1935_),
    .A(net21),
    .B(_1863_));
 sg13g2_xnor2_1 _6946_ (.Y(_1936_),
    .A(_1934_),
    .B(_1935_));
 sg13g2_xor2_1 _6947_ (.B(_1772_),
    .A(_1765_),
    .X(_1937_));
 sg13g2_nor2b_1 _6948_ (.A(_1936_),
    .B_N(_1937_),
    .Y(_1938_));
 sg13g2_inv_1 _6949_ (.Y(_1939_),
    .A(_1851_));
 sg13g2_nor2b_1 _6950_ (.A(_1939_),
    .B_N(_1769_),
    .Y(_1940_));
 sg13g2_o21ai_1 _6951_ (.B1(_1940_),
    .Y(_1941_),
    .A1(_1723_),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ));
 sg13g2_xnor2_1 _6952_ (.Y(_1942_),
    .A(_1769_),
    .B(_1770_));
 sg13g2_nand2_1 _6953_ (.Y(_1943_),
    .A(_1810_),
    .B(_1851_));
 sg13g2_xnor2_1 _6954_ (.Y(_1944_),
    .A(_1861_),
    .B(_1943_));
 sg13g2_nor2_1 _6955_ (.A(_1942_),
    .B(_1944_),
    .Y(_1945_));
 sg13g2_nand2_1 _6956_ (.Y(_1946_),
    .A(_1944_),
    .B(_1942_));
 sg13g2_o21ai_1 _6957_ (.B1(_1946_),
    .Y(_1947_),
    .A1(_1941_),
    .A2(_1945_));
 sg13g2_nand2b_1 _6958_ (.Y(_1948_),
    .B(_1936_),
    .A_N(_1937_));
 sg13g2_o21ai_1 _6959_ (.B1(_1948_),
    .Y(_1949_),
    .A1(_1938_),
    .A2(_1947_));
 sg13g2_nand2_1 _6960_ (.Y(_1950_),
    .A(_1932_),
    .B(_1930_));
 sg13g2_o21ai_1 _6961_ (.B1(_1950_),
    .Y(_1951_),
    .A1(_1933_),
    .A2(_1949_));
 sg13g2_o21ai_1 _6962_ (.B1(_1951_),
    .Y(_1952_),
    .A1(_1927_),
    .A2(_1929_));
 sg13g2_nand2_1 _6963_ (.Y(_1953_),
    .A(_1929_),
    .B(_1927_));
 sg13g2_nand2_1 _6964_ (.Y(_1954_),
    .A(_1952_),
    .B(_1953_));
 sg13g2_inv_1 _6965_ (.Y(_1955_),
    .A(_1954_));
 sg13g2_nand2_1 _6966_ (.Y(_1956_),
    .A(_1924_),
    .B(_1922_));
 sg13g2_o21ai_1 _6967_ (.B1(_1956_),
    .Y(_1957_),
    .A1(_1925_),
    .A2(_1955_));
 sg13g2_xor2_1 _6968_ (.B(_1786_),
    .A(_1791_),
    .X(_1958_));
 sg13g2_inv_1 _6969_ (.Y(_1959_),
    .A(_1958_));
 sg13g2_a21oi_1 _6970_ (.A1(_1909_),
    .A2(_1901_),
    .Y(_1960_),
    .B1(_1916_));
 sg13g2_nor2_1 _6971_ (.A(_1959_),
    .B(_1960_),
    .Y(_1961_));
 sg13g2_nand2_1 _6972_ (.Y(_1962_),
    .A(_1960_),
    .B(_1959_));
 sg13g2_nor2b_1 _6973_ (.A(_1961_),
    .B_N(_1962_),
    .Y(_1963_));
 sg13g2_nand2_1 _6974_ (.Y(_1964_),
    .A(_1957_),
    .B(_1963_));
 sg13g2_xor2_1 _6975_ (.B(_1793_),
    .A(_1797_),
    .X(_1965_));
 sg13g2_nor2b_1 _6976_ (.A(_1917_),
    .B_N(_1965_),
    .Y(_1966_));
 sg13g2_nor2_1 _6977_ (.A(_1966_),
    .B(_1961_),
    .Y(_1967_));
 sg13g2_nor2_1 _6978_ (.A(_1965_),
    .B(_1916_),
    .Y(_1968_));
 sg13g2_a21oi_1 _6979_ (.A1(_1964_),
    .A2(_1967_),
    .Y(_1969_),
    .B1(_1968_));
 sg13g2_nor2_1 _6980_ (.A(_1920_),
    .B(_1916_),
    .Y(_1970_));
 sg13g2_inv_1 _6981_ (.Y(_1971_),
    .A(_1920_));
 sg13g2_nor2_1 _6982_ (.A(_1971_),
    .B(_1917_),
    .Y(_1972_));
 sg13g2_nor2_1 _6983_ (.A(_1970_),
    .B(_1972_),
    .Y(_1973_));
 sg13g2_nand2_1 _6984_ (.Y(_1974_),
    .A(_1969_),
    .B(_1973_));
 sg13g2_a22oi_1 _6985_ (.Y(_1975_),
    .B1(_1921_),
    .B2(_1974_),
    .A2(_1919_),
    .A1(_1917_));
 sg13g2_xnor2_1 _6986_ (.Y(_1976_),
    .A(_1910_),
    .B(_1975_));
 sg13g2_buf_1 _6987_ (.A(_1976_),
    .X(_1977_));
 sg13g2_xnor2_1 _6988_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[1] ),
    .A(_1720_),
    .B(net15));
 sg13g2_nand2_1 _6989_ (.Y(_1978_),
    .A(net56),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ));
 sg13g2_xnor2_1 _6990_ (.Y(_1979_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_a[2] ),
    .B(_1978_));
 sg13g2_xnor2_1 _6991_ (.Y(_1980_),
    .A(_1979_),
    .B(net18));
 sg13g2_inv_1 _6992_ (.Y(_1981_),
    .A(_1980_));
 sg13g2_inv_1 _6993_ (.Y(_1982_),
    .A(_1720_));
 sg13g2_nor2_1 _6994_ (.A(_1982_),
    .B(net15),
    .Y(_1983_));
 sg13g2_xnor2_1 _6995_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[2] ),
    .A(_1981_),
    .B(_1983_));
 sg13g2_nand2b_1 _6996_ (.Y(_1984_),
    .B(_1978_),
    .A_N(\main.demo._q___pip_58_1_2___stage___block_3_a[2] ));
 sg13g2_inv_1 _6997_ (.Y(_1985_),
    .A(_1984_));
 sg13g2_nor2_1 _6998_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ),
    .B(net48),
    .Y(_1986_));
 sg13g2_inv_1 _6999_ (.Y(_1987_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ));
 sg13g2_nor2_1 _7000_ (.A(net56),
    .B(_1987_),
    .Y(_1988_));
 sg13g2_nor2_2 _7001_ (.A(_1986_),
    .B(_1988_),
    .Y(_1989_));
 sg13g2_xnor2_1 _7002_ (.Y(_1990_),
    .A(_1985_),
    .B(_1989_));
 sg13g2_xor2_1 _7003_ (.B(net18),
    .A(_1990_),
    .X(_1991_));
 sg13g2_nor2_1 _7004_ (.A(_1979_),
    .B(net17),
    .Y(_1992_));
 sg13g2_nor2_1 _7005_ (.A(_1982_),
    .B(_1981_),
    .Y(_1993_));
 sg13g2_nor2_1 _7006_ (.A(_1992_),
    .B(_1993_),
    .Y(_1994_));
 sg13g2_xnor2_1 _7007_ (.Y(_1995_),
    .A(_1991_),
    .B(_1994_));
 sg13g2_nand2_1 _7008_ (.Y(_1996_),
    .A(net15),
    .B(_1993_));
 sg13g2_xnor2_1 _7009_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[3] ),
    .A(_1995_),
    .B(_1996_));
 sg13g2_xnor2_1 _7010_ (.Y(_1997_),
    .A(net56),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_a21oi_1 _7011_ (.A1(_1989_),
    .A2(_1984_),
    .Y(_1998_),
    .B1(_1988_));
 sg13g2_xor2_1 _7012_ (.B(_1998_),
    .A(_1997_),
    .X(_1999_));
 sg13g2_xor2_1 _7013_ (.B(net18),
    .A(_1999_),
    .X(_2000_));
 sg13g2_nand2_1 _7014_ (.Y(_2001_),
    .A(_1993_),
    .B(_1991_));
 sg13g2_nand2_1 _7015_ (.Y(_2002_),
    .A(net18),
    .B(_1990_));
 sg13g2_nand3b_1 _7016_ (.B(_2001_),
    .C(_2002_),
    .Y(_2003_),
    .A_N(_1992_));
 sg13g2_xnor2_1 _7017_ (.Y(_2004_),
    .A(_2000_),
    .B(_2003_));
 sg13g2_o21ai_1 _7018_ (.B1(_2004_),
    .Y(_2005_),
    .A1(_1995_),
    .A2(_1996_));
 sg13g2_nor2_1 _7019_ (.A(_2001_),
    .B(_2004_),
    .Y(_2006_));
 sg13g2_nand2_1 _7020_ (.Y(_2007_),
    .A(_1977_),
    .B(_2006_));
 sg13g2_nand2_1 _7021_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[4] ),
    .A(_2005_),
    .B(_2007_));
 sg13g2_nand3_1 _7022_ (.B(_1984_),
    .C(_1997_),
    .A(_1989_),
    .Y(_2008_));
 sg13g2_o21ai_1 _7023_ (.B1(_1734_),
    .Y(_2009_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_nand2_1 _7024_ (.Y(_2010_),
    .A(_2008_),
    .B(_2009_));
 sg13g2_a21oi_1 _7025_ (.A1(_2010_),
    .A2(_1989_),
    .Y(_2011_),
    .B1(_1986_));
 sg13g2_inv_1 _7026_ (.Y(_2012_),
    .A(_2011_));
 sg13g2_nor2_1 _7027_ (.A(_2012_),
    .B(net17),
    .Y(_2013_));
 sg13g2_inv_1 _7028_ (.Y(_2014_),
    .A(_2000_));
 sg13g2_a21oi_1 _7029_ (.A1(_1999_),
    .A2(_2012_),
    .Y(_2015_),
    .B1(net17));
 sg13g2_a21oi_2 _7030_ (.B1(_2015_),
    .Y(_2016_),
    .A2(_2014_),
    .A1(_2003_));
 sg13g2_nand2_1 _7031_ (.Y(_2017_),
    .A(net17),
    .B(_2012_));
 sg13g2_o21ai_1 _7032_ (.B1(_2017_),
    .Y(_2018_),
    .A1(_2013_),
    .A2(_2016_));
 sg13g2_nand2_1 _7033_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[5] ),
    .A(_2007_),
    .B(_2018_));
 sg13g2_xnor2_1 _7034_ (.Y(_2019_),
    .A(_1719_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ));
 sg13g2_xnor2_1 _7035_ (.Y(_2020_),
    .A(_2019_),
    .B(_2010_));
 sg13g2_xnor2_1 _7036_ (.Y(_2021_),
    .A(_2020_),
    .B(net18));
 sg13g2_xor2_1 _7037_ (.B(_2016_),
    .A(_2021_),
    .X(_2022_));
 sg13g2_xor2_1 _7038_ (.B(_2007_),
    .A(_2022_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_a[6] ));
 sg13g2_xnor2_1 _7039_ (.Y(_2023_),
    .A(_1719_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[7] ));
 sg13g2_a21oi_1 _7040_ (.A1(_2010_),
    .A2(_2019_),
    .Y(_2024_),
    .B1(_1988_));
 sg13g2_inv_1 _7041_ (.Y(_2025_),
    .A(_2024_));
 sg13g2_a21oi_1 _7042_ (.A1(_1734_),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ),
    .Y(_2026_),
    .B1(_2025_));
 sg13g2_xnor2_1 _7043_ (.Y(_2027_),
    .A(_2023_),
    .B(_2026_));
 sg13g2_xor2_1 _7044_ (.B(_1811_),
    .A(_2027_),
    .X(_2028_));
 sg13g2_nand2b_1 _7045_ (.Y(_2029_),
    .B(_2017_),
    .A_N(_2013_));
 sg13g2_nor2_1 _7046_ (.A(_2029_),
    .B(_2016_),
    .Y(_2030_));
 sg13g2_nor2_1 _7047_ (.A(_2020_),
    .B(_1913_),
    .Y(_2031_));
 sg13g2_a221oi_1 _7048_ (.B2(_2021_),
    .C1(_2031_),
    .B1(_2030_),
    .A1(_1811_),
    .Y(_2032_),
    .A2(_2011_));
 sg13g2_xnor2_1 _7049_ (.Y(_2033_),
    .A(_2028_),
    .B(_2032_));
 sg13g2_nand3_1 _7050_ (.B(_2006_),
    .C(_2022_),
    .A(_1977_),
    .Y(_2034_));
 sg13g2_xnor2_1 _7051_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[7] ),
    .A(_2033_),
    .B(_2034_));
 sg13g2_xnor2_1 _7052_ (.Y(_2035_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[0] ),
    .B(_1775_));
 sg13g2_xor2_1 _7053_ (.B(_1927_),
    .A(_2035_),
    .X(_2036_));
 sg13g2_nand2b_1 _7054_ (.Y(_2037_),
    .B(_1956_),
    .A_N(_1925_));
 sg13g2_xor2_1 _7055_ (.B(_1954_),
    .A(_2037_),
    .X(_2038_));
 sg13g2_xor2_1 _7056_ (.B(_2038_),
    .A(_2036_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[0] ));
 sg13g2_xnor2_1 _7057_ (.Y(_2039_),
    .A(_1919_),
    .B(_1916_));
 sg13g2_o21ai_1 _7058_ (.B1(_1956_),
    .Y(_2040_),
    .A1(_1959_),
    .A2(_1960_));
 sg13g2_inv_1 _7059_ (.Y(_2041_),
    .A(_1963_));
 sg13g2_nor3_1 _7060_ (.A(_2041_),
    .B(_2037_),
    .C(_1955_),
    .Y(_2042_));
 sg13g2_a21o_1 _7061_ (.A2(_2040_),
    .A1(_1962_),
    .B1(_2042_),
    .X(_2043_));
 sg13g2_nor2_1 _7062_ (.A(_1968_),
    .B(_1966_),
    .Y(_2044_));
 sg13g2_nand2_1 _7063_ (.Y(_2045_),
    .A(_2043_),
    .B(_2044_));
 sg13g2_nor2_1 _7064_ (.A(_1966_),
    .B(_1972_),
    .Y(_2046_));
 sg13g2_a21oi_1 _7065_ (.A1(_2045_),
    .A2(_2046_),
    .Y(_2047_),
    .B1(_1970_));
 sg13g2_xnor2_1 _7066_ (.Y(_2048_),
    .A(_2039_),
    .B(_2047_));
 sg13g2_xor2_1 _7067_ (.B(_1969_),
    .A(_1973_),
    .X(_2049_));
 sg13g2_inv_1 _7068_ (.Y(_2050_),
    .A(_2038_));
 sg13g2_xnor2_1 _7069_ (.Y(_2051_),
    .A(_2041_),
    .B(_1957_));
 sg13g2_nor2_1 _7070_ (.A(_2050_),
    .B(_2051_),
    .Y(_2052_));
 sg13g2_inv_1 _7071_ (.Y(_2053_),
    .A(_2052_));
 sg13g2_xor2_1 _7072_ (.B(_2043_),
    .A(_2044_),
    .X(_2054_));
 sg13g2_nor2_1 _7073_ (.A(_2053_),
    .B(_2054_),
    .Y(_2055_));
 sg13g2_inv_1 _7074_ (.Y(_2056_),
    .A(_2055_));
 sg13g2_nor2_1 _7075_ (.A(_2049_),
    .B(_2056_),
    .Y(_2057_));
 sg13g2_nand3_1 _7076_ (.B(_2048_),
    .C(_2057_),
    .A(net15),
    .Y(_2058_));
 sg13g2_buf_1 _7077_ (.A(_2058_),
    .X(_2059_));
 sg13g2_nor2_1 _7078_ (.A(_1927_),
    .B(_1922_),
    .Y(_2060_));
 sg13g2_inv_1 _7079_ (.Y(_2061_),
    .A(_2060_));
 sg13g2_nor2_1 _7080_ (.A(_2061_),
    .B(_1958_),
    .Y(_2062_));
 sg13g2_inv_1 _7081_ (.Y(_2063_),
    .A(_2062_));
 sg13g2_nor2_1 _7082_ (.A(_2063_),
    .B(_1965_),
    .Y(_2064_));
 sg13g2_nand2_1 _7083_ (.Y(_2065_),
    .A(_1971_),
    .B(_2064_));
 sg13g2_nor3_1 _7084_ (.A(_1918_),
    .B(_2065_),
    .C(net17),
    .Y(_2066_));
 sg13g2_buf_2 _7085_ (.A(_2066_),
    .X(_2067_));
 sg13g2_xnor2_1 _7086_ (.Y(_2068_),
    .A(_1908_),
    .B(_2067_));
 sg13g2_inv_1 _7087_ (.Y(_2069_),
    .A(_1900_));
 sg13g2_inv_1 _7088_ (.Y(_2070_),
    .A(_2067_));
 sg13g2_nor2b_1 _7089_ (.A(_2070_),
    .B_N(_1881_),
    .Y(_2071_));
 sg13g2_nor2_1 _7090_ (.A(_1873_),
    .B(_2067_),
    .Y(_2072_));
 sg13g2_xor2_1 _7091_ (.B(_1840_),
    .A(_1845_),
    .X(_2073_));
 sg13g2_nand2_1 _7092_ (.Y(_2074_),
    .A(net21),
    .B(_2061_));
 sg13g2_xnor2_1 _7093_ (.Y(_2075_),
    .A(_1959_),
    .B(_2074_));
 sg13g2_nor2b_1 _7094_ (.A(_2073_),
    .B_N(_2075_),
    .Y(_2076_));
 sg13g2_xor2_1 _7095_ (.B(_2075_),
    .A(_2073_),
    .X(_2077_));
 sg13g2_xnor2_1 _7096_ (.Y(_2078_),
    .A(_1837_),
    .B(_1838_));
 sg13g2_nand2_1 _7097_ (.Y(_2079_),
    .A(net21),
    .B(_1927_));
 sg13g2_xor2_1 _7098_ (.B(_2079_),
    .A(_1922_),
    .X(_2080_));
 sg13g2_nor2b_1 _7099_ (.A(_2078_),
    .B_N(_2080_),
    .Y(_2081_));
 sg13g2_xor2_1 _7100_ (.B(_2080_),
    .A(_2078_),
    .X(_2082_));
 sg13g2_nand2_1 _7101_ (.Y(_2083_),
    .A(_1927_),
    .B(_2035_));
 sg13g2_nor2b_1 _7102_ (.A(_2082_),
    .B_N(_2083_),
    .Y(_2084_));
 sg13g2_nor2_1 _7103_ (.A(_2081_),
    .B(_2084_),
    .Y(_2085_));
 sg13g2_nor2_1 _7104_ (.A(_2077_),
    .B(_2085_),
    .Y(_2086_));
 sg13g2_nor2_1 _7105_ (.A(_2076_),
    .B(_2086_),
    .Y(_2087_));
 sg13g2_inv_1 _7106_ (.Y(_2088_),
    .A(_2087_));
 sg13g2_xnor2_1 _7107_ (.Y(_2089_),
    .A(_1848_),
    .B(_1847_));
 sg13g2_nand2_1 _7108_ (.Y(_2090_),
    .A(net18),
    .B(_2063_));
 sg13g2_xnor2_1 _7109_ (.Y(_2091_),
    .A(_1965_),
    .B(_2090_));
 sg13g2_nand2b_1 _7110_ (.Y(_2092_),
    .B(_2091_),
    .A_N(_2089_));
 sg13g2_nor2b_1 _7111_ (.A(_2091_),
    .B_N(_2089_),
    .Y(_2093_));
 sg13g2_a21o_1 _7112_ (.A2(_2092_),
    .A1(_2088_),
    .B1(_2093_),
    .X(_2094_));
 sg13g2_nor2_1 _7113_ (.A(_2064_),
    .B(net17),
    .Y(_2095_));
 sg13g2_xnor2_1 _7114_ (.Y(_2096_),
    .A(_1971_),
    .B(_2095_));
 sg13g2_nand2_1 _7115_ (.Y(_2097_),
    .A(_2096_),
    .B(_1939_));
 sg13g2_nor2_1 _7116_ (.A(_1939_),
    .B(_2096_),
    .Y(_2098_));
 sg13g2_a21o_1 _7117_ (.A2(_2097_),
    .A1(_2094_),
    .B1(_2098_),
    .X(_2099_));
 sg13g2_nand2_1 _7118_ (.Y(_2100_),
    .A(net18),
    .B(_2065_));
 sg13g2_xnor2_1 _7119_ (.Y(_2101_),
    .A(_1918_),
    .B(_2100_));
 sg13g2_inv_1 _7120_ (.Y(_2102_),
    .A(_1861_));
 sg13g2_nand2_1 _7121_ (.Y(_2103_),
    .A(_2101_),
    .B(_2102_));
 sg13g2_nor2_1 _7122_ (.A(_2102_),
    .B(_2101_),
    .Y(_2104_));
 sg13g2_a21o_1 _7123_ (.A2(_2103_),
    .A1(_2099_),
    .B1(_2104_),
    .X(_2105_));
 sg13g2_nor2b_1 _7124_ (.A(_2072_),
    .B_N(_2105_),
    .Y(_2106_));
 sg13g2_nor2_1 _7125_ (.A(_1881_),
    .B(_2067_),
    .Y(_2107_));
 sg13g2_nor2_1 _7126_ (.A(_2107_),
    .B(_2071_),
    .Y(_2108_));
 sg13g2_nand2_1 _7127_ (.Y(_2109_),
    .A(_2106_),
    .B(_2108_));
 sg13g2_inv_1 _7128_ (.Y(_2110_),
    .A(_1890_));
 sg13g2_nor2_1 _7129_ (.A(_2110_),
    .B(_2070_),
    .Y(_2111_));
 sg13g2_inv_1 _7130_ (.Y(_2112_),
    .A(_2111_));
 sg13g2_nand3b_1 _7131_ (.B(_2109_),
    .C(_2112_),
    .Y(_2113_),
    .A_N(_2071_));
 sg13g2_nand2_1 _7132_ (.Y(_2114_),
    .A(_2070_),
    .B(_2110_));
 sg13g2_nand2_1 _7133_ (.Y(_2115_),
    .A(_2113_),
    .B(_2114_));
 sg13g2_a21oi_1 _7134_ (.A1(_2069_),
    .A2(_2070_),
    .Y(_2116_),
    .B1(_2115_));
 sg13g2_xnor2_1 _7135_ (.Y(_2117_),
    .A(_2068_),
    .B(_2116_));
 sg13g2_xnor2_1 _7136_ (.Y(_2118_),
    .A(net14),
    .B(_2117_));
 sg13g2_xnor2_1 _7137_ (.Y(_2119_),
    .A(_1900_),
    .B(_2067_));
 sg13g2_xnor2_1 _7138_ (.Y(_2120_),
    .A(_2119_),
    .B(_2115_));
 sg13g2_nand2_1 _7139_ (.Y(_2121_),
    .A(_2112_),
    .B(_2114_));
 sg13g2_xnor2_1 _7140_ (.Y(_2122_),
    .A(_2121_),
    .B(_2113_));
 sg13g2_inv_1 _7141_ (.Y(_2123_),
    .A(_2122_));
 sg13g2_a21oi_1 _7142_ (.A1(_2120_),
    .A2(_2123_),
    .Y(_2124_),
    .B1(net14));
 sg13g2_xnor2_1 _7143_ (.Y(_2125_),
    .A(_1934_),
    .B(_2067_));
 sg13g2_xnor2_1 _7144_ (.Y(_2126_),
    .A(_2125_),
    .B(_2105_));
 sg13g2_inv_1 _7145_ (.Y(_2127_),
    .A(net14));
 sg13g2_nand2b_1 _7146_ (.Y(_2128_),
    .B(_2103_),
    .A_N(_2104_));
 sg13g2_xnor2_1 _7147_ (.Y(_2129_),
    .A(_2128_),
    .B(_2099_));
 sg13g2_nor2b_1 _7148_ (.A(_2098_),
    .B_N(_2097_),
    .Y(_2130_));
 sg13g2_xor2_1 _7149_ (.B(_2094_),
    .A(_2130_),
    .X(_2131_));
 sg13g2_nand2b_1 _7150_ (.Y(_2132_),
    .B(net15),
    .A_N(_2057_));
 sg13g2_xor2_1 _7151_ (.B(_2132_),
    .A(_2048_),
    .X(_2133_));
 sg13g2_nor2b_1 _7152_ (.A(_2131_),
    .B_N(_2133_),
    .Y(_2134_));
 sg13g2_nor2b_1 _7153_ (.A(_2133_),
    .B_N(_2131_),
    .Y(_2135_));
 sg13g2_xor2_1 _7154_ (.B(_2085_),
    .A(_2077_),
    .X(_2136_));
 sg13g2_nand2_1 _7155_ (.Y(_2137_),
    .A(net15),
    .B(_2053_));
 sg13g2_xor2_1 _7156_ (.B(_2137_),
    .A(_2054_),
    .X(_2138_));
 sg13g2_nor2_1 _7157_ (.A(_2136_),
    .B(_2138_),
    .Y(_2139_));
 sg13g2_xor2_1 _7158_ (.B(_2082_),
    .A(_2083_),
    .X(_2140_));
 sg13g2_nand2_1 _7159_ (.Y(_2141_),
    .A(net15),
    .B(_2050_));
 sg13g2_xor2_1 _7160_ (.B(_2141_),
    .A(_2051_),
    .X(_2142_));
 sg13g2_nor2b_1 _7161_ (.A(_2140_),
    .B_N(_2142_),
    .Y(_2143_));
 sg13g2_xor2_1 _7162_ (.B(_2142_),
    .A(_2140_),
    .X(_2144_));
 sg13g2_nand2_1 _7163_ (.Y(_2145_),
    .A(_2050_),
    .B(_2036_));
 sg13g2_nor2b_1 _7164_ (.A(_2144_),
    .B_N(_2145_),
    .Y(_2146_));
 sg13g2_nor2_1 _7165_ (.A(_2143_),
    .B(_2146_),
    .Y(_2147_));
 sg13g2_nand2_1 _7166_ (.Y(_2148_),
    .A(_2138_),
    .B(_2136_));
 sg13g2_o21ai_1 _7167_ (.B1(_2148_),
    .Y(_2149_),
    .A1(_2139_),
    .A2(_2147_));
 sg13g2_nor2b_1 _7168_ (.A(_2093_),
    .B_N(_2092_),
    .Y(_2150_));
 sg13g2_xnor2_1 _7169_ (.Y(_2151_),
    .A(_2150_),
    .B(_2087_));
 sg13g2_nand2_1 _7170_ (.Y(_2152_),
    .A(net15),
    .B(_2056_));
 sg13g2_xnor2_1 _7171_ (.Y(_2153_),
    .A(_2049_),
    .B(_2152_));
 sg13g2_nand2b_1 _7172_ (.Y(_2154_),
    .B(_2153_),
    .A_N(_2151_));
 sg13g2_nor2b_1 _7173_ (.A(_2153_),
    .B_N(_2151_),
    .Y(_2155_));
 sg13g2_a21o_1 _7174_ (.A2(_2154_),
    .A1(_2149_),
    .B1(_2155_),
    .X(_2156_));
 sg13g2_nor2_1 _7175_ (.A(_2135_),
    .B(_2156_),
    .Y(_2157_));
 sg13g2_nor2_1 _7176_ (.A(_2134_),
    .B(_2157_),
    .Y(_2158_));
 sg13g2_o21ai_1 _7177_ (.B1(_2158_),
    .Y(_2159_),
    .A1(_2127_),
    .A2(_2129_));
 sg13g2_a21oi_1 _7178_ (.A1(net14),
    .A2(_2126_),
    .Y(_2160_),
    .B1(_2159_));
 sg13g2_xnor2_1 _7179_ (.Y(_2161_),
    .A(_2108_),
    .B(_2106_));
 sg13g2_xor2_1 _7180_ (.B(_2059_),
    .A(_2161_),
    .X(_2162_));
 sg13g2_a21oi_1 _7181_ (.A1(_2123_),
    .A2(_2161_),
    .Y(_2163_),
    .B1(_2059_));
 sg13g2_a21o_1 _7182_ (.A2(_2162_),
    .A1(_2160_),
    .B1(_2163_),
    .X(_2164_));
 sg13g2_buf_1 _7183_ (.A(_2164_),
    .X(_2165_));
 sg13g2_xor2_1 _7184_ (.B(net14),
    .A(_2120_),
    .X(_2166_));
 sg13g2_xnor2_1 _7185_ (.Y(_2167_),
    .A(_2122_),
    .B(net14));
 sg13g2_nand3_1 _7186_ (.B(_2166_),
    .C(_2167_),
    .A(_2165_),
    .Y(_2168_));
 sg13g2_nand2b_1 _7187_ (.Y(_2169_),
    .B(_2168_),
    .A_N(_2124_));
 sg13g2_xnor2_1 _7188_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[10] ),
    .A(_2118_),
    .B(_2169_));
 sg13g2_xnor2_1 _7189_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[1] ),
    .A(_2145_),
    .B(_2144_));
 sg13g2_nor2b_1 _7190_ (.A(_2139_),
    .B_N(_2148_),
    .Y(_2170_));
 sg13g2_xnor2_1 _7191_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[2] ),
    .A(_2170_),
    .B(_2147_));
 sg13g2_nor2b_1 _7192_ (.A(_2155_),
    .B_N(_2154_),
    .Y(_2171_));
 sg13g2_xor2_1 _7193_ (.B(_2149_),
    .A(_2171_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[3] ));
 sg13g2_nor2_1 _7194_ (.A(_2135_),
    .B(_2134_),
    .Y(_2172_));
 sg13g2_xor2_1 _7195_ (.B(_2156_),
    .A(_2172_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_xor2_1 _7196_ (.B(net14),
    .A(_2129_),
    .X(_2173_));
 sg13g2_xnor2_1 _7197_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[5] ),
    .A(_2173_),
    .B(_2158_));
 sg13g2_xor2_1 _7198_ (.B(net14),
    .A(_2126_),
    .X(_2174_));
 sg13g2_xnor2_1 _7199_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[6] ),
    .A(_2174_),
    .B(_2159_));
 sg13g2_xor2_1 _7200_ (.B(_2160_),
    .A(_2162_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[7] ));
 sg13g2_xor2_1 _7201_ (.B(_2165_),
    .A(_2167_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[8] ));
 sg13g2_o21ai_1 _7202_ (.B1(_2165_),
    .Y(_2175_),
    .A1(_2127_),
    .A2(_2122_));
 sg13g2_xnor2_1 _7203_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[9] ),
    .A(_2166_),
    .B(_2175_));
 sg13g2_buf_1 _7204_ (.A(_4275_),
    .X(_2176_));
 sg13g2_inv_1 _7205_ (.Y(_2177_),
    .A(_4229_));
 sg13g2_inv_1 _7206_ (.Y(_2178_),
    .A(_4226_));
 sg13g2_inv_1 _7207_ (.Y(_2179_),
    .A(_4223_));
 sg13g2_nor2_2 _7208_ (.A(_2179_),
    .B(_0792_),
    .Y(_2180_));
 sg13g2_inv_1 _7209_ (.Y(_2181_),
    .A(_2180_));
 sg13g2_a21oi_1 _7210_ (.A1(_2177_),
    .A2(_2178_),
    .Y(_2182_),
    .B1(_2181_));
 sg13g2_nor2_1 _7211_ (.A(_2177_),
    .B(net43),
    .Y(_2183_));
 sg13g2_buf_2 _7212_ (.A(_2183_),
    .X(_2184_));
 sg13g2_nor2_2 _7213_ (.A(_2178_),
    .B(_0792_),
    .Y(_2185_));
 sg13g2_nor2_1 _7214_ (.A(_2185_),
    .B(_2180_),
    .Y(_2186_));
 sg13g2_inv_1 _7215_ (.Y(_2187_),
    .A(_2186_));
 sg13g2_nor2_1 _7216_ (.A(_2184_),
    .B(_2187_),
    .Y(_2188_));
 sg13g2_nor2_1 _7217_ (.A(_2182_),
    .B(_2188_),
    .Y(_2189_));
 sg13g2_buf_8 _7218_ (.A(_0018_),
    .X(_2190_));
 sg13g2_buf_8 _7219_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ),
    .X(_2191_));
 sg13g2_nor2_1 _7220_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .B(net72),
    .Y(_2192_));
 sg13g2_buf_8 _7221_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ),
    .X(_2193_));
 sg13g2_nand2_1 _7222_ (.Y(_2194_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .B(_2193_));
 sg13g2_buf_8 _7223_ (.A(_2194_),
    .X(_2195_));
 sg13g2_nand2_1 _7224_ (.Y(_2196_),
    .A(_2192_),
    .B(_2195_));
 sg13g2_nand2_1 _7225_ (.Y(_2197_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[8] ));
 sg13g2_inv_1 _7226_ (.Y(_2198_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ));
 sg13g2_nand2_1 _7227_ (.Y(_2199_),
    .A(_2197_),
    .B(_2198_));
 sg13g2_buf_2 _7228_ (.A(_2199_),
    .X(_2200_));
 sg13g2_nand2_1 _7229_ (.Y(_2201_),
    .A(_2196_),
    .B(_2200_));
 sg13g2_buf_8 _7230_ (.A(_2201_),
    .X(_2202_));
 sg13g2_o21ai_1 _7231_ (.B1(_2202_),
    .Y(_2203_),
    .A1(net73),
    .A2(_2191_));
 sg13g2_buf_1 _7232_ (.A(_2203_),
    .X(_2204_));
 sg13g2_nor2_1 _7233_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .Y(_2205_));
 sg13g2_buf_2 _7234_ (.A(_2205_),
    .X(_2206_));
 sg13g2_inv_2 _7235_ (.Y(_2207_),
    .A(_2206_));
 sg13g2_buf_8 _7236_ (.A(_2207_),
    .X(_2208_));
 sg13g2_inv_4 _7237_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .Y(_2209_));
 sg13g2_nor2_2 _7238_ (.A(_2193_),
    .B(_2209_),
    .Y(_2210_));
 sg13g2_nand2b_1 _7239_ (.Y(_2211_),
    .B(_2202_),
    .A_N(_2210_));
 sg13g2_nand3_1 _7240_ (.B(net47),
    .C(_2211_),
    .A(net32),
    .Y(_2212_));
 sg13g2_buf_1 _7241_ (.A(_2212_),
    .X(_2213_));
 sg13g2_a21oi_1 _7242_ (.A1(_2196_),
    .A2(_2200_),
    .Y(_2214_),
    .B1(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ));
 sg13g2_nand3_1 _7243_ (.B(net47),
    .C(_2214_),
    .A(net32),
    .Y(_2215_));
 sg13g2_nor2_2 _7244_ (.A(_2195_),
    .B(_2200_),
    .Y(_2216_));
 sg13g2_inv_1 _7245_ (.Y(_2217_),
    .A(_2216_));
 sg13g2_inv_1 _7246_ (.Y(_2218_),
    .A(_0018_));
 sg13g2_nand3_1 _7247_ (.B(_2198_),
    .C(net72),
    .A(_2197_),
    .Y(_2219_));
 sg13g2_buf_1 _7248_ (.A(_2219_),
    .X(_2220_));
 sg13g2_nor2_1 _7249_ (.A(_2218_),
    .B(_2220_),
    .Y(_2221_));
 sg13g2_nand2_2 _7250_ (.Y(_2222_),
    .A(_2221_),
    .B(net47));
 sg13g2_nor2_1 _7251_ (.A(_2217_),
    .B(_2222_),
    .Y(_2223_));
 sg13g2_inv_2 _7252_ (.Y(_2224_),
    .A(_2223_));
 sg13g2_nand3_1 _7253_ (.B(_2215_),
    .C(_2224_),
    .A(_2213_),
    .Y(_2225_));
 sg13g2_nand3_1 _7254_ (.B(_2209_),
    .C(_2193_),
    .A(_2202_),
    .Y(_2226_));
 sg13g2_nor2_1 _7255_ (.A(_2222_),
    .B(_2226_),
    .Y(_2227_));
 sg13g2_buf_8 _7256_ (.A(_2206_),
    .X(_2228_));
 sg13g2_a21oi_1 _7257_ (.A1(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .A2(\main.demo._d___pip_58_1_3___stage___block_3_cx[8] ),
    .Y(_2229_),
    .B1(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ));
 sg13g2_nand3_1 _7258_ (.B(net73),
    .C(net72),
    .A(_2229_),
    .Y(_2230_));
 sg13g2_buf_1 _7259_ (.A(_2230_),
    .X(_2231_));
 sg13g2_a21oi_1 _7260_ (.A1(_2196_),
    .A2(_2200_),
    .Y(_2232_),
    .B1(_2210_));
 sg13g2_nor3_1 _7261_ (.A(net53),
    .B(_2231_),
    .C(_2232_),
    .Y(_2233_));
 sg13g2_nor2_1 _7262_ (.A(_2227_),
    .B(_2233_),
    .Y(_2234_));
 sg13g2_nand2_1 _7263_ (.Y(_2235_),
    .A(_2202_),
    .B(net73));
 sg13g2_nand2_1 _7264_ (.Y(_2236_),
    .A(_2216_),
    .B(net72));
 sg13g2_inv_1 _7265_ (.Y(_2237_),
    .A(net72));
 sg13g2_a21oi_1 _7266_ (.A1(_2237_),
    .A2(_2195_),
    .Y(_2238_),
    .B1(_2200_));
 sg13g2_nand2_1 _7267_ (.Y(_2239_),
    .A(_2236_),
    .B(_2238_));
 sg13g2_nor2_1 _7268_ (.A(_2235_),
    .B(_2239_),
    .Y(_2240_));
 sg13g2_inv_1 _7269_ (.Y(_2241_),
    .A(_2193_));
 sg13g2_nand3_1 _7270_ (.B(_2209_),
    .C(_2241_),
    .A(_2202_),
    .Y(_2242_));
 sg13g2_buf_1 _7271_ (.A(_2242_),
    .X(_2243_));
 sg13g2_nor2_1 _7272_ (.A(net53),
    .B(_2243_),
    .Y(_2244_));
 sg13g2_nand2_1 _7273_ (.Y(_2245_),
    .A(_2240_),
    .B(_2244_));
 sg13g2_inv_2 _7274_ (.Y(_2246_),
    .A(_2195_));
 sg13g2_nand4_1 _7275_ (.B(net73),
    .C(_2237_),
    .A(_2229_),
    .Y(_2247_),
    .D(_2246_));
 sg13g2_nor2_2 _7276_ (.A(net53),
    .B(_2247_),
    .Y(_2248_));
 sg13g2_inv_2 _7277_ (.Y(_2249_),
    .A(_2248_));
 sg13g2_nand3_1 _7278_ (.B(_2245_),
    .C(_2249_),
    .A(_2234_),
    .Y(_2250_));
 sg13g2_nor2_1 _7279_ (.A(_2225_),
    .B(_2250_),
    .Y(_2251_));
 sg13g2_nor2_1 _7280_ (.A(net73),
    .B(_2220_),
    .Y(_2252_));
 sg13g2_nand2_1 _7281_ (.Y(_2253_),
    .A(_2252_),
    .B(_2216_));
 sg13g2_nand2_1 _7282_ (.Y(_2254_),
    .A(_2253_),
    .B(net53));
 sg13g2_nand3_1 _7283_ (.B(net47),
    .C(_2216_),
    .A(_2252_),
    .Y(_2255_));
 sg13g2_nand2_1 _7284_ (.Y(_2256_),
    .A(_2254_),
    .B(_2255_));
 sg13g2_nand3_1 _7285_ (.B(net73),
    .C(_2237_),
    .A(_2202_),
    .Y(_2257_));
 sg13g2_buf_1 _7286_ (.A(_2257_),
    .X(_2258_));
 sg13g2_nor2_1 _7287_ (.A(_2243_),
    .B(_2258_),
    .Y(_2259_));
 sg13g2_nand2_1 _7288_ (.Y(_2260_),
    .A(_2256_),
    .B(_2259_));
 sg13g2_buf_2 _7289_ (.A(_2260_),
    .X(_2261_));
 sg13g2_nand2_2 _7290_ (.Y(_2262_),
    .A(_2210_),
    .B(net53));
 sg13g2_inv_1 _7291_ (.Y(_2263_),
    .A(_2262_));
 sg13g2_nand3_1 _7292_ (.B(_2209_),
    .C(_2193_),
    .A(_2206_),
    .Y(_2264_));
 sg13g2_buf_2 _7293_ (.A(_2264_),
    .X(_2265_));
 sg13g2_inv_1 _7294_ (.Y(_2266_),
    .A(_2265_));
 sg13g2_nor2_1 _7295_ (.A(net72),
    .B(_2235_),
    .Y(_2267_));
 sg13g2_o21ai_1 _7296_ (.B1(_2267_),
    .Y(_2268_),
    .A1(_2263_),
    .A2(_2266_));
 sg13g2_buf_1 _7297_ (.A(_2268_),
    .X(_2269_));
 sg13g2_nand2_1 _7298_ (.Y(_2270_),
    .A(_2261_),
    .B(_2269_));
 sg13g2_nand2_1 _7299_ (.Y(_2271_),
    .A(_2235_),
    .B(_2220_));
 sg13g2_a21oi_1 _7300_ (.A1(_2262_),
    .A2(_2265_),
    .Y(_2272_),
    .B1(_2271_));
 sg13g2_nand3_1 _7301_ (.B(_2209_),
    .C(_2241_),
    .A(_2206_),
    .Y(_2273_));
 sg13g2_buf_1 _7302_ (.A(_2273_),
    .X(_2274_));
 sg13g2_inv_1 _7303_ (.Y(_2275_),
    .A(_2274_));
 sg13g2_nand2_1 _7304_ (.Y(_2276_),
    .A(net32),
    .B(_2275_));
 sg13g2_nand2_1 _7305_ (.Y(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ),
    .A(_2228_),
    .B(_2190_));
 sg13g2_nor2_1 _7306_ (.A(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ),
    .B(_2236_),
    .Y(_2277_));
 sg13g2_inv_2 _7307_ (.Y(_2278_),
    .A(_2277_));
 sg13g2_nand2_1 _7308_ (.Y(_2279_),
    .A(_2276_),
    .B(_2278_));
 sg13g2_nor2_1 _7309_ (.A(_2272_),
    .B(_2279_),
    .Y(_2280_));
 sg13g2_nor2_1 _7310_ (.A(_2274_),
    .B(_2231_),
    .Y(_2281_));
 sg13g2_a21oi_2 _7311_ (.B1(_2231_),
    .Y(_2282_),
    .A2(_2265_),
    .A1(_2262_));
 sg13g2_nor2_1 _7312_ (.A(net47),
    .B(_2247_),
    .Y(_2283_));
 sg13g2_nor3_1 _7313_ (.A(_2281_),
    .B(_2282_),
    .C(_2283_),
    .Y(_2284_));
 sg13g2_nand2_1 _7314_ (.Y(_2285_),
    .A(_2280_),
    .B(_2284_));
 sg13g2_nor2_1 _7315_ (.A(_2270_),
    .B(_2285_),
    .Y(_2286_));
 sg13g2_nand4_1 _7316_ (.B(net73),
    .C(_2237_),
    .A(_2202_),
    .Y(_2287_),
    .D(net47));
 sg13g2_buf_2 _7317_ (.A(_2287_),
    .X(_2288_));
 sg13g2_nor2b_1 _7318_ (.A(_2288_),
    .B_N(_2210_),
    .Y(_2289_));
 sg13g2_buf_8 _7319_ (.A(_2289_),
    .X(_2290_));
 sg13g2_nor4_2 _7320_ (.A(net73),
    .B(_2237_),
    .C(_2195_),
    .Y(_2291_),
    .D(_2207_));
 sg13g2_inv_1 _7321_ (.Y(_2292_),
    .A(_2291_));
 sg13g2_nor2b_1 _7322_ (.A(_2290_),
    .B_N(_2292_),
    .Y(_2293_));
 sg13g2_inv_2 _7323_ (.Y(_2294_),
    .A(_2288_));
 sg13g2_nand2_1 _7324_ (.Y(_2295_),
    .A(_2294_),
    .B(_2214_));
 sg13g2_nand2_1 _7325_ (.Y(_2296_),
    .A(_2293_),
    .B(_2295_));
 sg13g2_nand3_1 _7326_ (.B(_2218_),
    .C(net72),
    .A(_2206_),
    .Y(_2297_));
 sg13g2_inv_1 _7327_ (.Y(_2298_),
    .A(_2297_));
 sg13g2_nand3_1 _7328_ (.B(_2241_),
    .C(_2298_),
    .A(_2214_),
    .Y(_2299_));
 sg13g2_nor4_1 _7329_ (.A(_2190_),
    .B(_2191_),
    .C(_2195_),
    .D(_2200_),
    .Y(_2300_));
 sg13g2_nand2_1 _7330_ (.Y(_2301_),
    .A(_2300_),
    .B(_2228_));
 sg13g2_nand2_1 _7331_ (.Y(_2302_),
    .A(_2299_),
    .B(_2301_));
 sg13g2_nand4_1 _7332_ (.B(_2218_),
    .C(net72),
    .A(net53),
    .Y(_2303_),
    .D(_2209_));
 sg13g2_nor2_1 _7333_ (.A(_2241_),
    .B(_2303_),
    .Y(_2304_));
 sg13g2_nor2_1 _7334_ (.A(_2297_),
    .B(_2232_),
    .Y(_2305_));
 sg13g2_nor2_2 _7335_ (.A(_2304_),
    .B(_2305_),
    .Y(_2306_));
 sg13g2_nor2b_1 _7336_ (.A(_2302_),
    .B_N(_2306_),
    .Y(_2307_));
 sg13g2_nor2b_1 _7337_ (.A(_2296_),
    .B_N(_2307_),
    .Y(_2308_));
 sg13g2_nand3_1 _7338_ (.B(_2286_),
    .C(_2308_),
    .A(_2251_),
    .Y(_2309_));
 sg13g2_buf_2 _7339_ (.A(_2309_),
    .X(_2310_));
 sg13g2_nor2_1 _7340_ (.A(_2233_),
    .B(_2290_),
    .Y(_2311_));
 sg13g2_nand2_1 _7341_ (.Y(_2312_),
    .A(_2244_),
    .B(net32));
 sg13g2_inv_2 _7342_ (.Y(_2313_),
    .A(_2282_));
 sg13g2_nand4_1 _7343_ (.B(_2224_),
    .C(_2312_),
    .A(_2311_),
    .Y(_2314_),
    .D(net36));
 sg13g2_nor2b_1 _7344_ (.A(_2239_),
    .B_N(_2235_),
    .Y(_2315_));
 sg13g2_nor2_1 _7345_ (.A(_2274_),
    .B(_2315_),
    .Y(_2316_));
 sg13g2_nor3_1 _7346_ (.A(_2248_),
    .B(_2304_),
    .C(_2316_),
    .Y(_2317_));
 sg13g2_inv_1 _7347_ (.Y(_2318_),
    .A(_2272_));
 sg13g2_nor2_1 _7348_ (.A(_2243_),
    .B(_2288_),
    .Y(_2319_));
 sg13g2_nor2_1 _7349_ (.A(_2291_),
    .B(_2319_),
    .Y(_2320_));
 sg13g2_nand3_1 _7350_ (.B(_2318_),
    .C(_2320_),
    .A(_2317_),
    .Y(_2321_));
 sg13g2_nor2_1 _7351_ (.A(_2314_),
    .B(_2321_),
    .Y(_2322_));
 sg13g2_nand2_1 _7352_ (.Y(_2323_),
    .A(_2310_),
    .B(_2322_));
 sg13g2_nand2_1 _7353_ (.Y(_2324_),
    .A(_2216_),
    .B(net53));
 sg13g2_a21oi_1 _7354_ (.A1(_2265_),
    .A2(_2324_),
    .Y(_2325_),
    .B1(_2258_));
 sg13g2_nand2_1 _7355_ (.Y(_2326_),
    .A(net32),
    .B(_2266_));
 sg13g2_nand2_2 _7356_ (.Y(_2327_),
    .A(_2276_),
    .B(_2326_));
 sg13g2_nor2_1 _7357_ (.A(_2325_),
    .B(_2327_),
    .Y(_2328_));
 sg13g2_nand2_1 _7358_ (.Y(_2329_),
    .A(_2278_),
    .B(_2303_));
 sg13g2_nand2_1 _7359_ (.Y(_2330_),
    .A(_2204_),
    .B(_2263_));
 sg13g2_nand2_1 _7360_ (.Y(_2331_),
    .A(_2301_),
    .B(_2330_));
 sg13g2_nor2_1 _7361_ (.A(_2329_),
    .B(_2331_),
    .Y(_2332_));
 sg13g2_nand2_1 _7362_ (.Y(_2333_),
    .A(_2328_),
    .B(_2332_));
 sg13g2_nor2_1 _7363_ (.A(_2281_),
    .B(_2282_),
    .Y(_2334_));
 sg13g2_nor2_1 _7364_ (.A(_2262_),
    .B(_2258_),
    .Y(_2335_));
 sg13g2_inv_2 _7365_ (.Y(_2336_),
    .A(_2335_));
 sg13g2_nand2_1 _7366_ (.Y(_2337_),
    .A(_2334_),
    .B(_2336_));
 sg13g2_nand2_1 _7367_ (.Y(_2338_),
    .A(net32),
    .B(_2208_));
 sg13g2_nand2_1 _7368_ (.Y(_2339_),
    .A(_2338_),
    .B(_2222_));
 sg13g2_nor2_1 _7369_ (.A(_2291_),
    .B(_2305_),
    .Y(_2340_));
 sg13g2_nand2_1 _7370_ (.Y(_2341_),
    .A(_2340_),
    .B(_2288_));
 sg13g2_nor2_1 _7371_ (.A(_2339_),
    .B(_2341_),
    .Y(_2342_));
 sg13g2_nand2b_1 _7372_ (.Y(_2343_),
    .B(_2342_),
    .A_N(_2337_));
 sg13g2_nor2_1 _7373_ (.A(_2333_),
    .B(_2343_),
    .Y(_2344_));
 sg13g2_nand2_1 _7374_ (.Y(_2345_),
    .A(_2202_),
    .B(_2209_));
 sg13g2_a21oi_1 _7375_ (.A1(_2345_),
    .A2(_2217_),
    .Y(_2346_),
    .B1(_2288_));
 sg13g2_nand2_1 _7376_ (.Y(_2347_),
    .A(_2215_),
    .B(_2224_));
 sg13g2_nor3_1 _7377_ (.A(_2331_),
    .B(_2346_),
    .C(_2347_),
    .Y(_2348_));
 sg13g2_nor2_1 _7378_ (.A(_2265_),
    .B(_2231_),
    .Y(_2349_));
 sg13g2_nor2_1 _7379_ (.A(_2262_),
    .B(_2231_),
    .Y(_2350_));
 sg13g2_nor2_1 _7380_ (.A(_2350_),
    .B(_2277_),
    .Y(_2351_));
 sg13g2_nand2_1 _7381_ (.Y(_2352_),
    .A(_2266_),
    .B(_2220_));
 sg13g2_nand2_1 _7382_ (.Y(_2353_),
    .A(_2351_),
    .B(_2352_));
 sg13g2_nand2_1 _7383_ (.Y(_2354_),
    .A(_2211_),
    .B(_2298_));
 sg13g2_o21ai_1 _7384_ (.B1(_2354_),
    .Y(_2355_),
    .A1(_2222_),
    .A2(_2243_));
 sg13g2_nor3_1 _7385_ (.A(_2349_),
    .B(_2353_),
    .C(_2355_),
    .Y(_2356_));
 sg13g2_nand2_1 _7386_ (.Y(_2357_),
    .A(_2348_),
    .B(_2356_));
 sg13g2_nor2_1 _7387_ (.A(_2344_),
    .B(_2357_),
    .Y(_2358_));
 sg13g2_buf_2 _7388_ (.A(_2358_),
    .X(_2359_));
 sg13g2_nand2_1 _7389_ (.Y(_2360_),
    .A(_2323_),
    .B(_2359_));
 sg13g2_nor2b_1 _7390_ (.A(_2248_),
    .B_N(_2299_),
    .Y(_2361_));
 sg13g2_nor2_1 _7391_ (.A(_2283_),
    .B(_2335_),
    .Y(_2362_));
 sg13g2_nand3_1 _7392_ (.B(_2301_),
    .C(_2362_),
    .A(_2361_),
    .Y(_2363_));
 sg13g2_inv_1 _7393_ (.Y(_2364_),
    .A(_2281_));
 sg13g2_inv_1 _7394_ (.Y(_2365_),
    .A(_2349_));
 sg13g2_nand2_1 _7395_ (.Y(_2366_),
    .A(_2364_),
    .B(_2365_));
 sg13g2_inv_1 _7396_ (.Y(_2367_),
    .A(_2222_));
 sg13g2_nand2_1 _7397_ (.Y(_2368_),
    .A(_2367_),
    .B(_2217_));
 sg13g2_nand2_1 _7398_ (.Y(_2369_),
    .A(_2340_),
    .B(_2368_));
 sg13g2_nor3_1 _7399_ (.A(_2366_),
    .B(_2327_),
    .C(_2369_),
    .Y(_2370_));
 sg13g2_nand2b_1 _7400_ (.Y(_2371_),
    .B(_2370_),
    .A_N(_2363_));
 sg13g2_nor2_1 _7401_ (.A(_2344_),
    .B(_2371_),
    .Y(_2372_));
 sg13g2_inv_1 _7402_ (.Y(_2373_),
    .A(_2372_));
 sg13g2_buf_8 _7403_ (.A(_2310_),
    .X(_2374_));
 sg13g2_nand2_1 _7404_ (.Y(_2375_),
    .A(_2245_),
    .B(_2249_));
 sg13g2_nor2_1 _7405_ (.A(_2227_),
    .B(_2375_),
    .Y(_2376_));
 sg13g2_inv_1 _7406_ (.Y(_2377_),
    .A(_2279_));
 sg13g2_nand2_1 _7407_ (.Y(_2378_),
    .A(_2376_),
    .B(_2377_));
 sg13g2_nor2_1 _7408_ (.A(_2290_),
    .B(_2331_),
    .Y(_2379_));
 sg13g2_inv_1 _7409_ (.Y(_2380_),
    .A(_2283_));
 sg13g2_nand2_1 _7410_ (.Y(_2381_),
    .A(_2380_),
    .B(_2364_));
 sg13g2_inv_1 _7411_ (.Y(_2382_),
    .A(_2381_));
 sg13g2_nand4_1 _7412_ (.B(_2382_),
    .C(_2269_),
    .A(_2379_),
    .Y(_2383_),
    .D(_2306_));
 sg13g2_nor2_1 _7413_ (.A(_2378_),
    .B(_2383_),
    .Y(_2384_));
 sg13g2_nand3_1 _7414_ (.B(net26),
    .C(_2384_),
    .A(_2373_),
    .Y(_2385_));
 sg13g2_nand2_1 _7415_ (.Y(_2386_),
    .A(net26),
    .B(_2384_));
 sg13g2_nand2_1 _7416_ (.Y(_2387_),
    .A(_2386_),
    .B(_2372_));
 sg13g2_nand2_2 _7417_ (.Y(_2388_),
    .A(_2385_),
    .B(_2387_));
 sg13g2_o21ai_1 _7418_ (.B1(_2387_),
    .Y(_2389_),
    .A1(_2360_),
    .A2(_2388_));
 sg13g2_nand2_1 _7419_ (.Y(_2390_),
    .A(_2306_),
    .B(_2299_));
 sg13g2_nor2_1 _7420_ (.A(_2290_),
    .B(_2390_),
    .Y(_2391_));
 sg13g2_nor2_1 _7421_ (.A(_2241_),
    .B(_2345_),
    .Y(_2392_));
 sg13g2_nand3_1 _7422_ (.B(_2208_),
    .C(net32),
    .A(_2392_),
    .Y(_2393_));
 sg13g2_nor2b_1 _7423_ (.A(_2223_),
    .B_N(_2393_),
    .Y(_2394_));
 sg13g2_nand3_1 _7424_ (.B(_2391_),
    .C(_2394_),
    .A(_2376_),
    .Y(_2395_));
 sg13g2_nand3_1 _7425_ (.B(_2276_),
    .C(_2365_),
    .A(_2380_),
    .Y(_2396_));
 sg13g2_nor2_1 _7426_ (.A(_2265_),
    .B(_2258_),
    .Y(_2397_));
 sg13g2_inv_1 _7427_ (.Y(_2398_),
    .A(_2397_));
 sg13g2_nand2_1 _7428_ (.Y(_2399_),
    .A(_2261_),
    .B(_2398_));
 sg13g2_nor2_1 _7429_ (.A(_2396_),
    .B(_2399_),
    .Y(_2400_));
 sg13g2_nor2b_1 _7430_ (.A(_2395_),
    .B_N(_2400_),
    .Y(_2401_));
 sg13g2_nand2_1 _7431_ (.Y(_2402_),
    .A(_2354_),
    .B(_2292_));
 sg13g2_nor3_1 _7432_ (.A(_2304_),
    .B(_2248_),
    .C(_2402_),
    .Y(_2403_));
 sg13g2_inv_1 _7433_ (.Y(_2404_),
    .A(_2403_));
 sg13g2_nor2_1 _7434_ (.A(_2281_),
    .B(_2350_),
    .Y(_2405_));
 sg13g2_nand3_1 _7435_ (.B(_2326_),
    .C(_2405_),
    .A(_2269_),
    .Y(_2406_));
 sg13g2_nand3_1 _7436_ (.B(_2213_),
    .C(_2368_),
    .A(_2312_),
    .Y(_2407_));
 sg13g2_nor3_1 _7437_ (.A(_2404_),
    .B(_2406_),
    .C(_2407_),
    .Y(_2408_));
 sg13g2_nor2_1 _7438_ (.A(_2402_),
    .B(_2294_),
    .Y(_2409_));
 sg13g2_nand2b_1 _7439_ (.Y(_2410_),
    .B(_2409_),
    .A_N(_2339_));
 sg13g2_nor2_1 _7440_ (.A(_2337_),
    .B(_2410_),
    .Y(_2411_));
 sg13g2_inv_1 _7441_ (.Y(_2412_),
    .A(_2333_));
 sg13g2_nand2_1 _7442_ (.Y(_2413_),
    .A(_2411_),
    .B(_2412_));
 sg13g2_buf_8 _7443_ (.A(_2413_),
    .X(_2414_));
 sg13g2_nand2_1 _7444_ (.Y(_2415_),
    .A(_2408_),
    .B(_2414_));
 sg13g2_nand3_1 _7445_ (.B(_2401_),
    .C(_2415_),
    .A(_2310_),
    .Y(_2416_));
 sg13g2_buf_1 _7446_ (.A(_2416_),
    .X(_2417_));
 sg13g2_nand2_1 _7447_ (.Y(_2418_),
    .A(_2380_),
    .B(_2313_));
 sg13g2_nand3_1 _7448_ (.B(_2267_),
    .C(net47),
    .A(_2392_),
    .Y(_2419_));
 sg13g2_nand2_1 _7449_ (.Y(_2420_),
    .A(_2419_),
    .B(_2292_));
 sg13g2_nand3b_1 _7450_ (.B(_2213_),
    .C(_2224_),
    .Y(_2421_),
    .A_N(_2233_));
 sg13g2_nor4_2 _7451_ (.A(_2327_),
    .B(_2418_),
    .C(_2420_),
    .Y(_2422_),
    .D(_2421_));
 sg13g2_nand2_1 _7452_ (.Y(_2423_),
    .A(net26),
    .B(_2422_));
 sg13g2_nand2_1 _7453_ (.Y(_2424_),
    .A(_2224_),
    .B(_2364_));
 sg13g2_nor2_1 _7454_ (.A(_2319_),
    .B(_2424_),
    .Y(_2425_));
 sg13g2_inv_1 _7455_ (.Y(_2426_),
    .A(_2351_));
 sg13g2_a21oi_1 _7456_ (.A1(net32),
    .A2(_2244_),
    .Y(_2427_),
    .B1(_2426_));
 sg13g2_nand2_1 _7457_ (.Y(_2428_),
    .A(_2425_),
    .B(_2427_));
 sg13g2_a21oi_1 _7458_ (.A1(net47),
    .A2(_2300_),
    .Y(_2429_),
    .B1(_2290_));
 sg13g2_nand2_1 _7459_ (.Y(_2430_),
    .A(_2429_),
    .B(_2318_));
 sg13g2_nor2_1 _7460_ (.A(_2428_),
    .B(_2430_),
    .Y(_2431_));
 sg13g2_nand2_2 _7461_ (.Y(_2432_),
    .A(_2414_),
    .B(_2431_));
 sg13g2_inv_2 _7462_ (.Y(_2433_),
    .A(_2432_));
 sg13g2_nand2_1 _7463_ (.Y(_2434_),
    .A(_2423_),
    .B(_2433_));
 sg13g2_nand3_1 _7464_ (.B(_2432_),
    .C(_2422_),
    .A(_2310_),
    .Y(_2435_));
 sg13g2_buf_1 _7465_ (.A(_2435_),
    .X(_2436_));
 sg13g2_nand3_1 _7466_ (.B(_2434_),
    .C(_2436_),
    .A(_2417_),
    .Y(_2437_));
 sg13g2_nor2_1 _7467_ (.A(_2283_),
    .B(_2227_),
    .Y(_2438_));
 sg13g2_nand3_1 _7468_ (.B(_2301_),
    .C(_2213_),
    .A(_2438_),
    .Y(_2439_));
 sg13g2_nand2_1 _7469_ (.Y(_2440_),
    .A(_2425_),
    .B(_2403_));
 sg13g2_nor2_1 _7470_ (.A(_2439_),
    .B(_2440_),
    .Y(_2441_));
 sg13g2_nand2_2 _7471_ (.Y(_2442_),
    .A(_2414_),
    .B(_2441_));
 sg13g2_inv_2 _7472_ (.Y(_2443_),
    .A(_2442_));
 sg13g2_nand2_1 _7473_ (.Y(_2444_),
    .A(_2239_),
    .B(_2263_));
 sg13g2_nand3_1 _7474_ (.B(_2292_),
    .C(_2444_),
    .A(_2245_),
    .Y(_2445_));
 sg13g2_nand3_1 _7475_ (.B(_2380_),
    .C(_2393_),
    .A(_2311_),
    .Y(_2446_));
 sg13g2_nor3_1 _7476_ (.A(_2390_),
    .B(_2445_),
    .C(_2446_),
    .Y(_2447_));
 sg13g2_nand2_1 _7477_ (.Y(_2448_),
    .A(_2310_),
    .B(_2447_));
 sg13g2_a21oi_1 _7478_ (.A1(net26),
    .A2(_2422_),
    .Y(_2449_),
    .B1(_2432_));
 sg13g2_a21oi_1 _7479_ (.A1(_2443_),
    .A2(_2448_),
    .Y(_2450_),
    .B1(_2449_));
 sg13g2_nand2_1 _7480_ (.Y(_2451_),
    .A(_2437_),
    .B(_2450_));
 sg13g2_xnor2_1 _7481_ (.Y(_2452_),
    .A(_2359_),
    .B(_2323_));
 sg13g2_nor2_1 _7482_ (.A(_2452_),
    .B(_2388_),
    .Y(_2453_));
 sg13g2_nand3_1 _7483_ (.B(_2442_),
    .C(_2447_),
    .A(_2310_),
    .Y(_2454_));
 sg13g2_buf_1 _7484_ (.A(_2454_),
    .X(_2455_));
 sg13g2_nand3_1 _7485_ (.B(_2453_),
    .C(_2455_),
    .A(_2451_),
    .Y(_2456_));
 sg13g2_nand2b_1 _7486_ (.Y(_2457_),
    .B(_2456_),
    .A_N(_2389_));
 sg13g2_nand2_1 _7487_ (.Y(_2458_),
    .A(_2414_),
    .B(_2269_));
 sg13g2_nor2_1 _7488_ (.A(_2402_),
    .B(_2290_),
    .Y(_2459_));
 sg13g2_nand3_1 _7489_ (.B(_2278_),
    .C(_2295_),
    .A(_2459_),
    .Y(_2460_));
 sg13g2_nor3_1 _7490_ (.A(_2366_),
    .B(_2272_),
    .C(_2460_),
    .Y(_2461_));
 sg13g2_nor2b_1 _7491_ (.A(_2458_),
    .B_N(_2461_),
    .Y(_2462_));
 sg13g2_buf_8 _7492_ (.A(_2462_),
    .X(_2463_));
 sg13g2_nand2b_1 _7493_ (.Y(_2464_),
    .B(_2382_),
    .A_N(_2350_));
 sg13g2_nand3_1 _7494_ (.B(_2419_),
    .C(_2306_),
    .A(_2320_),
    .Y(_2465_));
 sg13g2_nor4_1 _7495_ (.A(_2327_),
    .B(_2399_),
    .C(_2464_),
    .D(_2465_),
    .Y(_2466_));
 sg13g2_nand2_1 _7496_ (.Y(_2467_),
    .A(_2466_),
    .B(net26));
 sg13g2_nor2_1 _7497_ (.A(_2463_),
    .B(_2467_),
    .Y(_2468_));
 sg13g2_nand2_1 _7498_ (.Y(_2469_),
    .A(_2467_),
    .B(_2463_));
 sg13g2_nand2b_1 _7499_ (.Y(_2470_),
    .B(_2469_),
    .A_N(_2468_));
 sg13g2_inv_1 _7500_ (.Y(_2471_),
    .A(_2470_));
 sg13g2_nand2_1 _7501_ (.Y(_2472_),
    .A(_2457_),
    .B(_2471_));
 sg13g2_buf_2 _7502_ (.A(_2472_),
    .X(_2473_));
 sg13g2_inv_1 _7503_ (.Y(_2474_),
    .A(_0022_));
 sg13g2_inv_1 _7504_ (.Y(_2475_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ));
 sg13g2_a21oi_1 _7505_ (.A1(_2434_),
    .A2(_2436_),
    .Y(_2476_),
    .B1(_2417_));
 sg13g2_nand2b_1 _7506_ (.Y(_2477_),
    .B(_2437_),
    .A_N(_2476_));
 sg13g2_buf_2 _7507_ (.A(_2477_),
    .X(_2478_));
 sg13g2_nor2_2 _7508_ (.A(_2475_),
    .B(_2478_),
    .Y(_2479_));
 sg13g2_nand4_1 _7509_ (.B(_2474_),
    .C(net36),
    .A(_2473_),
    .Y(_2480_),
    .D(_2479_));
 sg13g2_inv_1 _7510_ (.Y(_2481_),
    .A(_2480_));
 sg13g2_buf_2 _7511_ (.A(_0020_),
    .X(_2482_));
 sg13g2_nand2_1 _7512_ (.Y(_2483_),
    .A(_2448_),
    .B(_2443_));
 sg13g2_nand2_1 _7513_ (.Y(_2484_),
    .A(_2483_),
    .B(_2455_));
 sg13g2_a21oi_2 _7514_ (.B1(_2449_),
    .Y(_2485_),
    .A2(_2436_),
    .A1(_2417_));
 sg13g2_xnor2_1 _7515_ (.Y(_2486_),
    .A(_2484_),
    .B(_2485_));
 sg13g2_buf_2 _7516_ (.A(_2486_),
    .X(_2487_));
 sg13g2_nor2_2 _7517_ (.A(_2482_),
    .B(_2487_),
    .Y(_2488_));
 sg13g2_inv_2 _7518_ (.Y(_2489_),
    .A(_2485_));
 sg13g2_nor2_1 _7519_ (.A(_2484_),
    .B(_2452_),
    .Y(_2490_));
 sg13g2_nand2_1 _7520_ (.Y(_2491_),
    .A(_2489_),
    .B(_2490_));
 sg13g2_nor2_1 _7521_ (.A(_2359_),
    .B(_2323_),
    .Y(_2492_));
 sg13g2_a21oi_1 _7522_ (.A1(_2360_),
    .A2(_2483_),
    .Y(_2493_),
    .B1(_2492_));
 sg13g2_inv_1 _7523_ (.Y(_2494_),
    .A(_2493_));
 sg13g2_nand2_1 _7524_ (.Y(_2495_),
    .A(_2491_),
    .B(_2494_));
 sg13g2_nor2_1 _7525_ (.A(_2388_),
    .B(_2470_),
    .Y(_2496_));
 sg13g2_nand2_1 _7526_ (.Y(_2497_),
    .A(_2495_),
    .B(_2496_));
 sg13g2_a21oi_1 _7527_ (.A1(_2467_),
    .A2(_2463_),
    .Y(_2498_),
    .B1(_2397_));
 sg13g2_nand2_1 _7528_ (.Y(_2499_),
    .A(_2497_),
    .B(_2498_));
 sg13g2_nand3_1 _7529_ (.B(_2362_),
    .C(_2364_),
    .A(_2377_),
    .Y(_2500_));
 sg13g2_nor2_1 _7530_ (.A(_2410_),
    .B(_2500_),
    .Y(_2501_));
 sg13g2_nand2_2 _7531_ (.Y(_2502_),
    .A(_2414_),
    .B(_2501_));
 sg13g2_nand3_1 _7532_ (.B(_2380_),
    .C(_2306_),
    .A(_2269_),
    .Y(_2503_));
 sg13g2_nor3_1 _7533_ (.A(_2426_),
    .B(_2503_),
    .C(_2296_),
    .Y(_2504_));
 sg13g2_nand3_1 _7534_ (.B(_2504_),
    .C(_2251_),
    .A(_2374_),
    .Y(_2505_));
 sg13g2_xnor2_1 _7535_ (.Y(_2506_),
    .A(_2502_),
    .B(_2505_));
 sg13g2_nand2_2 _7536_ (.Y(_2507_),
    .A(_2499_),
    .B(_2506_));
 sg13g2_buf_2 _7537_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ),
    .X(_2508_));
 sg13g2_nand3_1 _7538_ (.B(_2508_),
    .C(_2261_),
    .A(_2507_),
    .Y(_2509_));
 sg13g2_nand2b_1 _7539_ (.Y(_2510_),
    .B(_2509_),
    .A_N(_2488_));
 sg13g2_nand4_1 _7540_ (.B(_2508_),
    .C(_2261_),
    .A(_2507_),
    .Y(_2511_),
    .D(_2488_));
 sg13g2_buf_1 _7541_ (.A(_2511_),
    .X(_2512_));
 sg13g2_nand2_1 _7542_ (.Y(_2513_),
    .A(_2510_),
    .B(_2512_));
 sg13g2_xnor2_1 _7543_ (.Y(_2514_),
    .A(_2481_),
    .B(_2513_));
 sg13g2_buf_2 _7544_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ),
    .X(_2515_));
 sg13g2_inv_4 _7545_ (.A(_2515_),
    .Y(_2516_));
 sg13g2_nand2_1 _7546_ (.Y(_2517_),
    .A(_2451_),
    .B(_2455_));
 sg13g2_xnor2_1 _7547_ (.Y(_2518_),
    .A(_2452_),
    .B(_2517_));
 sg13g2_nor2_2 _7548_ (.A(net63),
    .B(_2518_),
    .Y(_2519_));
 sg13g2_inv_1 _7549_ (.Y(_2520_),
    .A(_2388_));
 sg13g2_nand2_1 _7550_ (.Y(_2521_),
    .A(_2495_),
    .B(_2520_));
 sg13g2_nand3_1 _7551_ (.B(_2388_),
    .C(_2494_),
    .A(_2491_),
    .Y(_2522_));
 sg13g2_buf_2 _7552_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .X(_2523_));
 sg13g2_nand3_1 _7553_ (.B(_2522_),
    .C(_2523_),
    .A(_2521_),
    .Y(_2524_));
 sg13g2_buf_1 _7554_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .X(_2525_));
 sg13g2_inv_2 _7555_ (.Y(_2526_),
    .A(net71));
 sg13g2_nand2_1 _7556_ (.Y(_2527_),
    .A(_2473_),
    .B(net36));
 sg13g2_nor2_1 _7557_ (.A(_2526_),
    .B(_2527_),
    .Y(_2528_));
 sg13g2_nand2b_1 _7558_ (.Y(_2529_),
    .B(_2528_),
    .A_N(_2524_));
 sg13g2_xnor2_1 _7559_ (.Y(_2530_),
    .A(_2442_),
    .B(_2448_));
 sg13g2_inv_1 _7560_ (.Y(_2531_),
    .A(_2359_));
 sg13g2_nand2_1 _7561_ (.Y(_2532_),
    .A(_2323_),
    .B(_2531_));
 sg13g2_nand3_1 _7562_ (.B(_2322_),
    .C(_2359_),
    .A(_2374_),
    .Y(_2533_));
 sg13g2_nand2_1 _7563_ (.Y(_2534_),
    .A(_2532_),
    .B(_2533_));
 sg13g2_nand2_1 _7564_ (.Y(_2535_),
    .A(_2530_),
    .B(_2534_));
 sg13g2_nor2_1 _7565_ (.A(_2485_),
    .B(_2535_),
    .Y(_2536_));
 sg13g2_nor3_1 _7566_ (.A(_2520_),
    .B(_2493_),
    .C(_2536_),
    .Y(_2537_));
 sg13g2_a21oi_1 _7567_ (.A1(_2491_),
    .A2(_2494_),
    .Y(_2538_),
    .B1(_2388_));
 sg13g2_nor3_1 _7568_ (.A(_2526_),
    .B(_2537_),
    .C(_2538_),
    .Y(_2539_));
 sg13g2_nand3_1 _7569_ (.B(_2523_),
    .C(net36),
    .A(_2473_),
    .Y(_2540_));
 sg13g2_nand2b_1 _7570_ (.Y(_2541_),
    .B(_2540_),
    .A_N(_2539_));
 sg13g2_buf_1 _7571_ (.A(_2541_),
    .X(_2542_));
 sg13g2_nand2_1 _7572_ (.Y(_2543_),
    .A(_2529_),
    .B(_2542_));
 sg13g2_xor2_1 _7573_ (.B(_2543_),
    .A(_2519_),
    .X(_2544_));
 sg13g2_nand2_1 _7574_ (.Y(_2545_),
    .A(_2514_),
    .B(_2544_));
 sg13g2_nand2_1 _7575_ (.Y(_2546_),
    .A(_2513_),
    .B(_2480_));
 sg13g2_nand3_1 _7576_ (.B(_2512_),
    .C(_2481_),
    .A(_2510_),
    .Y(_2547_));
 sg13g2_nand2_1 _7577_ (.Y(_2548_),
    .A(_2546_),
    .B(_2547_));
 sg13g2_xnor2_1 _7578_ (.Y(_2549_),
    .A(_2519_),
    .B(_2543_));
 sg13g2_nand2_1 _7579_ (.Y(_2550_),
    .A(_2548_),
    .B(_2549_));
 sg13g2_nand3_1 _7580_ (.B(_2474_),
    .C(net36),
    .A(_2473_),
    .Y(_2551_));
 sg13g2_nand2b_1 _7581_ (.Y(_2552_),
    .B(_2551_),
    .A_N(_2479_));
 sg13g2_nand2_1 _7582_ (.Y(_2553_),
    .A(_2552_),
    .B(_2480_));
 sg13g2_inv_2 _7583_ (.Y(_2554_),
    .A(_2508_));
 sg13g2_nand2_1 _7584_ (.Y(_2555_),
    .A(_2521_),
    .B(_2522_));
 sg13g2_nor2_1 _7585_ (.A(_2554_),
    .B(_2555_),
    .Y(_2556_));
 sg13g2_a21oi_1 _7586_ (.A1(net26),
    .A2(_2401_),
    .Y(_2557_),
    .B1(_2415_));
 sg13g2_nor2b_1 _7587_ (.A(_2557_),
    .B_N(_2417_),
    .Y(_2558_));
 sg13g2_nor2_1 _7588_ (.A(_2482_),
    .B(_2558_),
    .Y(_2559_));
 sg13g2_nand2_1 _7589_ (.Y(_2560_),
    .A(_2556_),
    .B(_2559_));
 sg13g2_nand2_1 _7590_ (.Y(_2561_),
    .A(_2553_),
    .B(_2560_));
 sg13g2_nor2_2 _7591_ (.A(net63),
    .B(_2487_),
    .Y(_2562_));
 sg13g2_inv_1 _7592_ (.Y(_2563_),
    .A(_2523_));
 sg13g2_nor2_1 _7593_ (.A(_2563_),
    .B(_2518_),
    .Y(_2564_));
 sg13g2_nand2_1 _7594_ (.Y(_2565_),
    .A(_2539_),
    .B(_2564_));
 sg13g2_nand2_1 _7595_ (.Y(_2566_),
    .A(_2517_),
    .B(_2534_));
 sg13g2_nand3_1 _7596_ (.B(_2455_),
    .C(_2452_),
    .A(_2451_),
    .Y(_2567_));
 sg13g2_nand2_2 _7597_ (.Y(_2568_),
    .A(_2566_),
    .B(_2567_));
 sg13g2_nand2_1 _7598_ (.Y(_2569_),
    .A(_2568_),
    .B(net71));
 sg13g2_nand2_1 _7599_ (.Y(_2570_),
    .A(_2524_),
    .B(_2569_));
 sg13g2_nand2_1 _7600_ (.Y(_2571_),
    .A(_2565_),
    .B(_2570_));
 sg13g2_xnor2_1 _7601_ (.Y(_2572_),
    .A(_2562_),
    .B(_2571_));
 sg13g2_nor2_1 _7602_ (.A(_2560_),
    .B(_2553_),
    .Y(_2573_));
 sg13g2_a21oi_1 _7603_ (.A1(_2561_),
    .A2(_2572_),
    .Y(_2574_),
    .B1(_2573_));
 sg13g2_nand3_1 _7604_ (.B(_2550_),
    .C(_2574_),
    .A(_2545_),
    .Y(_2575_));
 sg13g2_buf_1 _7605_ (.A(_2575_),
    .X(_2576_));
 sg13g2_inv_1 _7606_ (.Y(_2577_),
    .A(_2565_));
 sg13g2_a21oi_1 _7607_ (.A1(_2570_),
    .A2(_2562_),
    .Y(_2578_),
    .B1(_2577_));
 sg13g2_inv_1 _7608_ (.Y(_2579_),
    .A(_2578_));
 sg13g2_nand2_1 _7609_ (.Y(_2580_),
    .A(_2545_),
    .B(_2550_));
 sg13g2_nand2b_1 _7610_ (.Y(_2581_),
    .B(_2580_),
    .A_N(_2574_));
 sg13g2_inv_1 _7611_ (.Y(_2582_),
    .A(_2581_));
 sg13g2_a21oi_2 _7612_ (.B1(_2582_),
    .Y(_2583_),
    .A2(_2579_),
    .A1(_2576_));
 sg13g2_inv_1 _7613_ (.Y(_2584_),
    .A(_2547_));
 sg13g2_a21oi_1 _7614_ (.A1(_2549_),
    .A2(_2546_),
    .Y(_2585_),
    .B1(_2584_));
 sg13g2_inv_1 _7615_ (.Y(_2586_),
    .A(_2482_));
 sg13g2_nand2_2 _7616_ (.Y(_2587_),
    .A(_2568_),
    .B(_2586_));
 sg13g2_nand3_1 _7617_ (.B(_2489_),
    .C(_2490_),
    .A(_2496_),
    .Y(_2588_));
 sg13g2_buf_8 _7618_ (.A(_2588_),
    .X(_2589_));
 sg13g2_nand2_2 _7619_ (.Y(_2590_),
    .A(_2589_),
    .B(_2336_));
 sg13g2_nor2_2 _7620_ (.A(_2554_),
    .B(_2590_),
    .Y(_2591_));
 sg13g2_xnor2_1 _7621_ (.Y(_2592_),
    .A(_2587_),
    .B(_2591_));
 sg13g2_xor2_1 _7622_ (.B(_2512_),
    .A(_2592_),
    .X(_2593_));
 sg13g2_nand2_2 _7623_ (.Y(_2594_),
    .A(_2507_),
    .B(_2261_));
 sg13g2_nor2_1 _7624_ (.A(_2563_),
    .B(_2594_),
    .Y(_2595_));
 sg13g2_nand2_1 _7625_ (.Y(_2596_),
    .A(_2595_),
    .B(_2528_));
 sg13g2_nand3_1 _7626_ (.B(_2523_),
    .C(_2261_),
    .A(_2507_),
    .Y(_2597_));
 sg13g2_nand3_1 _7627_ (.B(net71),
    .C(net36),
    .A(_2473_),
    .Y(_2598_));
 sg13g2_nand2_1 _7628_ (.Y(_2599_),
    .A(_2597_),
    .B(_2598_));
 sg13g2_nand2_1 _7629_ (.Y(_2600_),
    .A(_2596_),
    .B(_2599_));
 sg13g2_nor2_2 _7630_ (.A(net63),
    .B(_2555_),
    .Y(_2601_));
 sg13g2_nand2_1 _7631_ (.Y(_2602_),
    .A(_2600_),
    .B(_2601_));
 sg13g2_inv_1 _7632_ (.Y(_2603_),
    .A(_2601_));
 sg13g2_nand3_1 _7633_ (.B(_2599_),
    .C(_2603_),
    .A(_2596_),
    .Y(_2604_));
 sg13g2_nand2_1 _7634_ (.Y(_2605_),
    .A(_2602_),
    .B(_2604_));
 sg13g2_xnor2_1 _7635_ (.Y(_2606_),
    .A(_2593_),
    .B(_2605_));
 sg13g2_nand2b_1 _7636_ (.Y(_2607_),
    .B(_2606_),
    .A_N(_2585_));
 sg13g2_xor2_1 _7637_ (.B(_2605_),
    .A(_2593_),
    .X(_2608_));
 sg13g2_nand2_1 _7638_ (.Y(_2609_),
    .A(_2608_),
    .B(_2585_));
 sg13g2_nand2_1 _7639_ (.Y(_2610_),
    .A(_2607_),
    .B(_2609_));
 sg13g2_inv_1 _7640_ (.Y(_2611_),
    .A(_2529_));
 sg13g2_a21oi_1 _7641_ (.A1(_2519_),
    .A2(_2542_),
    .Y(_2612_),
    .B1(_2611_));
 sg13g2_nand2_1 _7642_ (.Y(_2613_),
    .A(_2610_),
    .B(_2612_));
 sg13g2_inv_1 _7643_ (.Y(_2614_),
    .A(_2612_));
 sg13g2_nand3_1 _7644_ (.B(_2609_),
    .C(_2614_),
    .A(_2607_),
    .Y(_2615_));
 sg13g2_buf_1 _7645_ (.A(_2615_),
    .X(_2616_));
 sg13g2_nand2_1 _7646_ (.Y(_2617_),
    .A(_2613_),
    .B(_2616_));
 sg13g2_nand2b_1 _7647_ (.Y(_2618_),
    .B(_2617_),
    .A_N(_2583_));
 sg13g2_nand3_1 _7648_ (.B(_2616_),
    .C(_2583_),
    .A(_2613_),
    .Y(_2619_));
 sg13g2_nand2_1 _7649_ (.Y(_2620_),
    .A(_2618_),
    .B(_2619_));
 sg13g2_nor2b_1 _7650_ (.A(_2573_),
    .B_N(_2561_),
    .Y(_2621_));
 sg13g2_xnor2_1 _7651_ (.Y(_2622_),
    .A(_2572_),
    .B(_2621_));
 sg13g2_nand2_1 _7652_ (.Y(_2623_),
    .A(_2568_),
    .B(_2523_));
 sg13g2_inv_1 _7653_ (.Y(_2624_),
    .A(_2487_));
 sg13g2_nand2_1 _7654_ (.Y(_2625_),
    .A(_2624_),
    .B(_2525_));
 sg13g2_nand2_1 _7655_ (.Y(_2626_),
    .A(_2623_),
    .B(_2625_));
 sg13g2_nor2_1 _7656_ (.A(_2526_),
    .B(_2487_),
    .Y(_2627_));
 sg13g2_nand3_1 _7657_ (.B(_2523_),
    .C(_2627_),
    .A(_2568_),
    .Y(_2628_));
 sg13g2_nor2_2 _7658_ (.A(_2516_),
    .B(_2478_),
    .Y(_2629_));
 sg13g2_inv_1 _7659_ (.Y(_2630_),
    .A(_2629_));
 sg13g2_nand3_1 _7660_ (.B(_2628_),
    .C(_2630_),
    .A(_2626_),
    .Y(_2631_));
 sg13g2_nand2_1 _7661_ (.Y(_2632_),
    .A(_2623_),
    .B(_2627_));
 sg13g2_nand3_1 _7662_ (.B(_2625_),
    .C(_2523_),
    .A(_2568_),
    .Y(_2633_));
 sg13g2_nand3_1 _7663_ (.B(_2633_),
    .C(_2629_),
    .A(_2632_),
    .Y(_2634_));
 sg13g2_nand2_1 _7664_ (.Y(_2635_),
    .A(_2631_),
    .B(_2634_));
 sg13g2_inv_1 _7665_ (.Y(_2636_),
    .A(_2559_));
 sg13g2_xnor2_1 _7666_ (.Y(_2637_),
    .A(_2636_),
    .B(_2556_));
 sg13g2_nand2_1 _7667_ (.Y(_2638_),
    .A(_2635_),
    .B(_2637_));
 sg13g2_nand2_1 _7668_ (.Y(_2639_),
    .A(_2622_),
    .B(_2638_));
 sg13g2_inv_1 _7669_ (.Y(_2640_),
    .A(_2628_));
 sg13g2_a21oi_1 _7670_ (.A1(_2626_),
    .A2(_2629_),
    .Y(_2641_),
    .B1(_2640_));
 sg13g2_inv_1 _7671_ (.Y(_2642_),
    .A(_2641_));
 sg13g2_nor2_1 _7672_ (.A(_2638_),
    .B(_2622_),
    .Y(_2643_));
 sg13g2_a21oi_1 _7673_ (.A1(_2639_),
    .A2(_2642_),
    .Y(_2644_),
    .B1(_2643_));
 sg13g2_nand2_1 _7674_ (.Y(_2645_),
    .A(_2581_),
    .B(_2576_));
 sg13g2_nand2_1 _7675_ (.Y(_2646_),
    .A(_2645_),
    .B(_2578_));
 sg13g2_nand3_1 _7676_ (.B(_2576_),
    .C(_2579_),
    .A(_2581_),
    .Y(_2647_));
 sg13g2_nand2_1 _7677_ (.Y(_2648_),
    .A(_2646_),
    .B(_2647_));
 sg13g2_nor2_1 _7678_ (.A(_2644_),
    .B(_2648_),
    .Y(_2649_));
 sg13g2_inv_1 _7679_ (.Y(_2650_),
    .A(_2649_));
 sg13g2_nor2_1 _7680_ (.A(_2537_),
    .B(_2538_),
    .Y(_2651_));
 sg13g2_nand2_1 _7681_ (.Y(_2652_),
    .A(_2651_),
    .B(_2508_));
 sg13g2_nand2_1 _7682_ (.Y(_2653_),
    .A(_2626_),
    .B(_2628_));
 sg13g2_xnor2_1 _7683_ (.Y(_2654_),
    .A(_2652_),
    .B(_2653_));
 sg13g2_xnor2_1 _7684_ (.Y(_2655_),
    .A(_2636_),
    .B(_2629_));
 sg13g2_nor2b_1 _7685_ (.A(_2654_),
    .B_N(_2655_),
    .Y(_2656_));
 sg13g2_nor2_1 _7686_ (.A(_2636_),
    .B(_2630_),
    .Y(_2657_));
 sg13g2_xnor2_1 _7687_ (.Y(_2658_),
    .A(_2479_),
    .B(_2562_));
 sg13g2_xor2_1 _7688_ (.B(_2658_),
    .A(_2657_),
    .X(_2659_));
 sg13g2_nand3_1 _7689_ (.B(_2565_),
    .C(_2570_),
    .A(_2551_),
    .Y(_2660_));
 sg13g2_inv_1 _7690_ (.Y(_2661_),
    .A(_2551_));
 sg13g2_nand2_1 _7691_ (.Y(_2662_),
    .A(_2571_),
    .B(_2661_));
 sg13g2_nand2_1 _7692_ (.Y(_2663_),
    .A(_2660_),
    .B(_2662_));
 sg13g2_nand2b_1 _7693_ (.Y(_2664_),
    .B(_2663_),
    .A_N(_2659_));
 sg13g2_nand3_1 _7694_ (.B(_2662_),
    .C(_2659_),
    .A(_2660_),
    .Y(_2665_));
 sg13g2_nand2_1 _7695_ (.Y(_2666_),
    .A(_2664_),
    .B(_2665_));
 sg13g2_nand2b_1 _7696_ (.Y(_2667_),
    .B(_2666_),
    .A_N(_2656_));
 sg13g2_nand3_1 _7697_ (.B(_2665_),
    .C(_2656_),
    .A(_2664_),
    .Y(_2668_));
 sg13g2_nand2_1 _7698_ (.Y(_2669_),
    .A(_2667_),
    .B(_2668_));
 sg13g2_a21oi_1 _7699_ (.A1(_2626_),
    .A2(_2556_),
    .Y(_2670_),
    .B1(_2640_));
 sg13g2_nand2_1 _7700_ (.Y(_2671_),
    .A(_2669_),
    .B(_2670_));
 sg13g2_inv_1 _7701_ (.Y(_2672_),
    .A(_2670_));
 sg13g2_nand3_1 _7702_ (.B(_2668_),
    .C(_2672_),
    .A(_2667_),
    .Y(_2673_));
 sg13g2_nand2_1 _7703_ (.Y(_2674_),
    .A(_2671_),
    .B(_2673_));
 sg13g2_nand2_1 _7704_ (.Y(_2675_),
    .A(_2652_),
    .B(_2636_));
 sg13g2_nand2_1 _7705_ (.Y(_2676_),
    .A(_2675_),
    .B(_2560_));
 sg13g2_nand3_1 _7706_ (.B(_2634_),
    .C(_2676_),
    .A(_2631_),
    .Y(_2677_));
 sg13g2_nand2_1 _7707_ (.Y(_2678_),
    .A(_2638_),
    .B(_2677_));
 sg13g2_nor2_1 _7708_ (.A(net63),
    .B(_2558_),
    .Y(_2679_));
 sg13g2_inv_1 _7709_ (.Y(_2680_),
    .A(_2679_));
 sg13g2_nand2_1 _7710_ (.Y(_2681_),
    .A(_2624_),
    .B(_2523_));
 sg13g2_nand2b_1 _7711_ (.Y(_2682_),
    .B(_2525_),
    .A_N(_2478_));
 sg13g2_nand2_1 _7712_ (.Y(_2683_),
    .A(_2681_),
    .B(_2682_));
 sg13g2_nor2_1 _7713_ (.A(_2563_),
    .B(_2478_),
    .Y(_2684_));
 sg13g2_nand2_1 _7714_ (.Y(_2685_),
    .A(_2627_),
    .B(_2684_));
 sg13g2_nand2_2 _7715_ (.Y(_2686_),
    .A(_2683_),
    .B(_2685_));
 sg13g2_xnor2_1 _7716_ (.Y(_2687_),
    .A(_2680_),
    .B(_2686_));
 sg13g2_nor2_2 _7717_ (.A(_2554_),
    .B(_2518_),
    .Y(_2688_));
 sg13g2_nand2b_1 _7718_ (.Y(_2689_),
    .B(_2688_),
    .A_N(_2687_));
 sg13g2_nand2_1 _7719_ (.Y(_2690_),
    .A(_2678_),
    .B(_2689_));
 sg13g2_o21ai_1 _7720_ (.B1(_2685_),
    .Y(_2691_),
    .A1(_2680_),
    .A2(_2686_));
 sg13g2_nor2_1 _7721_ (.A(_2689_),
    .B(_2678_),
    .Y(_2692_));
 sg13g2_a21oi_1 _7722_ (.A1(_2690_),
    .A2(_2691_),
    .Y(_2693_),
    .B1(_2692_));
 sg13g2_nand2_1 _7723_ (.Y(_2694_),
    .A(_2674_),
    .B(_2693_));
 sg13g2_xor2_1 _7724_ (.B(_2686_),
    .A(_2688_),
    .X(_2695_));
 sg13g2_nor2_1 _7725_ (.A(_2680_),
    .B(_2695_),
    .Y(_2696_));
 sg13g2_nand2b_1 _7726_ (.Y(_2697_),
    .B(_2678_),
    .A_N(_2696_));
 sg13g2_nand3_1 _7727_ (.B(_2677_),
    .C(_2696_),
    .A(_2638_),
    .Y(_2698_));
 sg13g2_inv_1 _7728_ (.Y(_2699_),
    .A(_2688_));
 sg13g2_o21ai_1 _7729_ (.B1(_2685_),
    .Y(_2700_),
    .A1(_2686_),
    .A2(_2699_));
 sg13g2_a21oi_1 _7730_ (.A1(_2697_),
    .A2(_2698_),
    .Y(_2701_),
    .B1(_2700_));
 sg13g2_nand3_1 _7731_ (.B(_2698_),
    .C(_2700_),
    .A(_2697_),
    .Y(_2702_));
 sg13g2_nor2_1 _7732_ (.A(_2526_),
    .B(_2558_),
    .Y(_2703_));
 sg13g2_xnor2_1 _7733_ (.Y(_2704_),
    .A(_2703_),
    .B(_2684_));
 sg13g2_nor2_1 _7734_ (.A(_2554_),
    .B(_2487_),
    .Y(_2705_));
 sg13g2_nand2b_1 _7735_ (.Y(_2706_),
    .B(_2705_),
    .A_N(_2704_));
 sg13g2_nand2b_1 _7736_ (.Y(_2707_),
    .B(_2704_),
    .A_N(_2705_));
 sg13g2_buf_1 _7737_ (.A(_0021_),
    .X(_2708_));
 sg13g2_nor4_1 _7738_ (.A(_2708_),
    .B(_0022_),
    .C(_2558_),
    .D(_2478_),
    .Y(_2709_));
 sg13g2_nand3_1 _7739_ (.B(_2707_),
    .C(_2709_),
    .A(_2706_),
    .Y(_2710_));
 sg13g2_nand2_1 _7740_ (.Y(_2711_),
    .A(_2684_),
    .B(_2703_));
 sg13g2_nand2_1 _7741_ (.Y(_2712_),
    .A(_2706_),
    .B(_2711_));
 sg13g2_xnor2_1 _7742_ (.Y(_2713_),
    .A(_2688_),
    .B(_2687_));
 sg13g2_nor2_1 _7743_ (.A(_2712_),
    .B(_2713_),
    .Y(_2714_));
 sg13g2_nand2_1 _7744_ (.Y(_2715_),
    .A(_2713_),
    .B(_2712_));
 sg13g2_o21ai_1 _7745_ (.B1(_2715_),
    .Y(_2716_),
    .A1(_2710_),
    .A2(_2714_));
 sg13g2_nand2_1 _7746_ (.Y(_2717_),
    .A(_2702_),
    .B(_2716_));
 sg13g2_nor2_1 _7747_ (.A(_2701_),
    .B(_2717_),
    .Y(_2718_));
 sg13g2_nand2_1 _7748_ (.Y(_2719_),
    .A(_2694_),
    .B(_2718_));
 sg13g2_inv_1 _7749_ (.Y(_2720_),
    .A(_2693_));
 sg13g2_nand3_1 _7750_ (.B(_2673_),
    .C(_2720_),
    .A(_2671_),
    .Y(_2721_));
 sg13g2_buf_1 _7751_ (.A(_2721_),
    .X(_2722_));
 sg13g2_nand2_2 _7752_ (.Y(_2723_),
    .A(_2719_),
    .B(_2722_));
 sg13g2_nand2_1 _7753_ (.Y(_2724_),
    .A(_2648_),
    .B(_2644_));
 sg13g2_nand2_1 _7754_ (.Y(_2725_),
    .A(_2723_),
    .B(_2724_));
 sg13g2_nand3_1 _7755_ (.B(_2650_),
    .C(_2725_),
    .A(_2620_),
    .Y(_2726_));
 sg13g2_nand2_1 _7756_ (.Y(_2727_),
    .A(_2725_),
    .B(_2650_));
 sg13g2_inv_2 _7757_ (.Y(_2728_),
    .A(_2620_));
 sg13g2_nand2_1 _7758_ (.Y(_2729_),
    .A(_2727_),
    .B(_2728_));
 sg13g2_nand3_1 _7759_ (.B(_2729_),
    .C(_2443_),
    .A(_2726_),
    .Y(_2730_));
 sg13g2_nand2_1 _7760_ (.Y(_2731_),
    .A(_2694_),
    .B(_2722_));
 sg13g2_nand2b_1 _7761_ (.Y(_2732_),
    .B(_2731_),
    .A_N(_2718_));
 sg13g2_nand3_1 _7762_ (.B(_2722_),
    .C(_2718_),
    .A(_2694_),
    .Y(_2733_));
 sg13g2_nand3_1 _7763_ (.B(_2733_),
    .C(_2415_),
    .A(_2732_),
    .Y(_2734_));
 sg13g2_buf_2 _7764_ (.A(_2734_),
    .X(_2735_));
 sg13g2_nand2_1 _7765_ (.Y(_2736_),
    .A(_2735_),
    .B(_2433_));
 sg13g2_nand2b_1 _7766_ (.Y(_2737_),
    .B(_2657_),
    .A_N(_2658_));
 sg13g2_nand2_1 _7767_ (.Y(_2738_),
    .A(_2664_),
    .B(_2737_));
 sg13g2_nand2_1 _7768_ (.Y(_2739_),
    .A(_2543_),
    .B(_2509_));
 sg13g2_inv_1 _7769_ (.Y(_2740_),
    .A(_2509_));
 sg13g2_nand3_1 _7770_ (.B(_2542_),
    .C(_2740_),
    .A(_2529_),
    .Y(_2741_));
 sg13g2_nand2_1 _7771_ (.Y(_2742_),
    .A(_2739_),
    .B(_2741_));
 sg13g2_nand2_1 _7772_ (.Y(_2743_),
    .A(_2562_),
    .B(_2479_));
 sg13g2_xnor2_1 _7773_ (.Y(_2744_),
    .A(_2488_),
    .B(_2519_));
 sg13g2_xor2_1 _7774_ (.B(_2744_),
    .A(_2743_),
    .X(_2745_));
 sg13g2_inv_1 _7775_ (.Y(_2746_),
    .A(_2745_));
 sg13g2_nand2_1 _7776_ (.Y(_2747_),
    .A(_2742_),
    .B(_2746_));
 sg13g2_nand3_1 _7777_ (.B(_2745_),
    .C(_2741_),
    .A(_2739_),
    .Y(_2748_));
 sg13g2_nand2_1 _7778_ (.Y(_2749_),
    .A(_2747_),
    .B(_2748_));
 sg13g2_nand2b_1 _7779_ (.Y(_2750_),
    .B(_2749_),
    .A_N(_2738_));
 sg13g2_nand3_1 _7780_ (.B(_2748_),
    .C(_2738_),
    .A(_2747_),
    .Y(_2751_));
 sg13g2_nand2_1 _7781_ (.Y(_2752_),
    .A(_2750_),
    .B(_2751_));
 sg13g2_a21oi_1 _7782_ (.A1(_2661_),
    .A2(_2570_),
    .Y(_2753_),
    .B1(_2577_));
 sg13g2_nand2_1 _7783_ (.Y(_2754_),
    .A(_2752_),
    .B(_2753_));
 sg13g2_inv_1 _7784_ (.Y(_2755_),
    .A(_2753_));
 sg13g2_nand3_1 _7785_ (.B(_2751_),
    .C(_2755_),
    .A(_2750_),
    .Y(_2756_));
 sg13g2_nand2_1 _7786_ (.Y(_2757_),
    .A(_2754_),
    .B(_2756_));
 sg13g2_inv_1 _7787_ (.Y(_2758_),
    .A(_2668_));
 sg13g2_a21oi_1 _7788_ (.A1(_2667_),
    .A2(_2672_),
    .Y(_2759_),
    .B1(_2758_));
 sg13g2_nand2_1 _7789_ (.Y(_2760_),
    .A(_2757_),
    .B(_2759_));
 sg13g2_inv_1 _7790_ (.Y(_2761_),
    .A(_2759_));
 sg13g2_nand3_1 _7791_ (.B(_2756_),
    .C(_2761_),
    .A(_2754_),
    .Y(_2762_));
 sg13g2_nand2_1 _7792_ (.Y(_2763_),
    .A(_2760_),
    .B(_2762_));
 sg13g2_xnor2_1 _7793_ (.Y(_2764_),
    .A(_2723_),
    .B(_2763_));
 sg13g2_nand2_1 _7794_ (.Y(_2765_),
    .A(_2736_),
    .B(_2764_));
 sg13g2_nand2b_1 _7795_ (.Y(_2766_),
    .B(_2432_),
    .A_N(_2735_));
 sg13g2_nand2_1 _7796_ (.Y(_2767_),
    .A(_2765_),
    .B(_2766_));
 sg13g2_nand2_1 _7797_ (.Y(_2768_),
    .A(_2730_),
    .B(_2767_));
 sg13g2_nand2_1 _7798_ (.Y(_2769_),
    .A(_2726_),
    .B(_2729_));
 sg13g2_nand2_1 _7799_ (.Y(_2770_),
    .A(_2769_),
    .B(_2442_));
 sg13g2_nand2_1 _7800_ (.Y(_2771_),
    .A(_2768_),
    .B(_2770_));
 sg13g2_xnor2_1 _7801_ (.Y(_2772_),
    .A(_2761_),
    .B(_2757_));
 sg13g2_nand2_1 _7802_ (.Y(_2773_),
    .A(_2772_),
    .B(_2723_));
 sg13g2_nor2_1 _7803_ (.A(_2583_),
    .B(_2617_),
    .Y(_2774_));
 sg13g2_nor2_1 _7804_ (.A(_2649_),
    .B(_2774_),
    .Y(_2775_));
 sg13g2_nand2_1 _7805_ (.Y(_2776_),
    .A(_2773_),
    .B(_2775_));
 sg13g2_nand2_1 _7806_ (.Y(_2777_),
    .A(_2617_),
    .B(_2583_));
 sg13g2_nand2_1 _7807_ (.Y(_2778_),
    .A(_2776_),
    .B(_2777_));
 sg13g2_nand2_2 _7808_ (.Y(_2779_),
    .A(_2616_),
    .B(_2607_));
 sg13g2_nor2b_1 _7809_ (.A(_2512_),
    .B_N(_2592_),
    .Y(_2780_));
 sg13g2_nand2b_1 _7810_ (.Y(_2781_),
    .B(_2605_),
    .A_N(_2593_));
 sg13g2_nand2b_1 _7811_ (.Y(_2782_),
    .B(_2781_),
    .A_N(_2780_));
 sg13g2_nor2_2 _7812_ (.A(_2482_),
    .B(_2590_),
    .Y(_2783_));
 sg13g2_nand2_1 _7813_ (.Y(_2784_),
    .A(_2783_),
    .B(_2688_));
 sg13g2_nand2_2 _7814_ (.Y(_2785_),
    .A(_2589_),
    .B(_2398_));
 sg13g2_nor2_2 _7815_ (.A(_2554_),
    .B(_2785_),
    .Y(_2786_));
 sg13g2_nand2_1 _7816_ (.Y(_2787_),
    .A(_2651_),
    .B(_2586_));
 sg13g2_xor2_1 _7817_ (.B(_2787_),
    .A(_2786_),
    .X(_2788_));
 sg13g2_xnor2_1 _7818_ (.Y(_2789_),
    .A(_2784_),
    .B(_2788_));
 sg13g2_nor2_1 _7819_ (.A(net63),
    .B(_2527_),
    .Y(_2790_));
 sg13g2_buf_2 _7820_ (.A(_2790_),
    .X(_2791_));
 sg13g2_nor2_1 _7821_ (.A(_2708_),
    .B(_2590_),
    .Y(_2792_));
 sg13g2_inv_1 _7822_ (.Y(_2793_),
    .A(_2792_));
 sg13g2_o21ai_1 _7823_ (.B1(_2793_),
    .Y(_2794_),
    .A1(_2526_),
    .A2(_2594_));
 sg13g2_buf_1 _7824_ (.A(_2794_),
    .X(_2795_));
 sg13g2_inv_2 _7825_ (.Y(_2796_),
    .A(_2594_));
 sg13g2_nand3_1 _7826_ (.B(net71),
    .C(_2792_),
    .A(_2796_),
    .Y(_2797_));
 sg13g2_nand2_1 _7827_ (.Y(_2798_),
    .A(_2795_),
    .B(_2797_));
 sg13g2_nand2b_1 _7828_ (.Y(_2799_),
    .B(_2798_),
    .A_N(_2791_));
 sg13g2_nand3_1 _7829_ (.B(_2797_),
    .C(_2791_),
    .A(_2795_),
    .Y(_2800_));
 sg13g2_nand3b_1 _7830_ (.B(_2799_),
    .C(_2800_),
    .Y(_2801_),
    .A_N(_2789_));
 sg13g2_buf_1 _7831_ (.A(_2801_),
    .X(_2802_));
 sg13g2_nand2_1 _7832_ (.Y(_2803_),
    .A(_2799_),
    .B(_2800_));
 sg13g2_nand2_1 _7833_ (.Y(_2804_),
    .A(_2803_),
    .B(_2789_));
 sg13g2_nand3_1 _7834_ (.B(_2802_),
    .C(_2804_),
    .A(_2782_),
    .Y(_2805_));
 sg13g2_nand2_1 _7835_ (.Y(_2806_),
    .A(_2802_),
    .B(_2804_));
 sg13g2_nand2b_1 _7836_ (.Y(_2807_),
    .B(_2806_),
    .A_N(_2782_));
 sg13g2_nand2_1 _7837_ (.Y(_2808_),
    .A(_2805_),
    .B(_2807_));
 sg13g2_inv_1 _7838_ (.Y(_2809_),
    .A(_2596_));
 sg13g2_a21oi_1 _7839_ (.A1(_2601_),
    .A2(_2599_),
    .Y(_2810_),
    .B1(_2809_));
 sg13g2_nand2_1 _7840_ (.Y(_2811_),
    .A(_2808_),
    .B(_2810_));
 sg13g2_inv_1 _7841_ (.Y(_2812_),
    .A(_2810_));
 sg13g2_nand3_1 _7842_ (.B(_2807_),
    .C(_2812_),
    .A(_2805_),
    .Y(_2813_));
 sg13g2_nand2_2 _7843_ (.Y(_2814_),
    .A(_2811_),
    .B(_2813_));
 sg13g2_xor2_1 _7844_ (.B(_2814_),
    .A(_2779_),
    .X(_2815_));
 sg13g2_nand2_1 _7845_ (.Y(_2816_),
    .A(_2778_),
    .B(_2815_));
 sg13g2_xnor2_1 _7846_ (.Y(_2817_),
    .A(_2779_),
    .B(_2814_));
 sg13g2_nand3_1 _7847_ (.B(_2777_),
    .C(_2817_),
    .A(_2776_),
    .Y(_2818_));
 sg13g2_nand2_1 _7848_ (.Y(_2819_),
    .A(_2816_),
    .B(_2818_));
 sg13g2_nand2_1 _7849_ (.Y(_2820_),
    .A(_2819_),
    .B(_2359_));
 sg13g2_nand2_1 _7850_ (.Y(_2821_),
    .A(_2771_),
    .B(_2820_));
 sg13g2_nor2_1 _7851_ (.A(_2728_),
    .B(_2815_),
    .Y(_2822_));
 sg13g2_nand2_1 _7852_ (.Y(_2823_),
    .A(_2822_),
    .B(_2727_));
 sg13g2_nor2b_1 _7853_ (.A(_2814_),
    .B_N(_2779_),
    .Y(_2824_));
 sg13g2_nand2b_1 _7854_ (.Y(_2825_),
    .B(_2814_),
    .A_N(_2779_));
 sg13g2_o21ai_1 _7855_ (.B1(_2825_),
    .Y(_2826_),
    .A1(_2774_),
    .A2(_2824_));
 sg13g2_nand2_1 _7856_ (.Y(_2827_),
    .A(_2823_),
    .B(_2826_));
 sg13g2_inv_1 _7857_ (.Y(_2828_),
    .A(_2805_));
 sg13g2_a21oi_2 _7858_ (.B1(_2828_),
    .Y(_2829_),
    .A2(_2812_),
    .A1(_2807_));
 sg13g2_nand2_2 _7859_ (.Y(_2830_),
    .A(_2796_),
    .B(_2515_));
 sg13g2_nor2_1 _7860_ (.A(_2526_),
    .B(_2590_),
    .Y(_2831_));
 sg13g2_inv_2 _7861_ (.Y(_2832_),
    .A(_2785_));
 sg13g2_inv_1 _7862_ (.Y(_2833_),
    .A(_2708_));
 sg13g2_nand2_1 _7863_ (.Y(_2834_),
    .A(_2832_),
    .B(_2833_));
 sg13g2_xnor2_1 _7864_ (.Y(_2835_),
    .A(_2831_),
    .B(_2834_));
 sg13g2_xnor2_1 _7865_ (.Y(_2836_),
    .A(_2830_),
    .B(_2835_));
 sg13g2_nor2b_1 _7866_ (.A(_2787_),
    .B_N(_2786_),
    .Y(_2837_));
 sg13g2_nand3_1 _7867_ (.B(_2586_),
    .C(net36),
    .A(_2473_),
    .Y(_2838_));
 sg13g2_inv_1 _7868_ (.Y(_2839_),
    .A(_2589_));
 sg13g2_nor2_1 _7869_ (.A(_2554_),
    .B(_2839_),
    .Y(_2840_));
 sg13g2_inv_1 _7870_ (.Y(_2841_),
    .A(_2840_));
 sg13g2_nand2_1 _7871_ (.Y(_2842_),
    .A(_2838_),
    .B(_2841_));
 sg13g2_nand4_1 _7872_ (.B(_2586_),
    .C(_2508_),
    .A(_2473_),
    .Y(_2843_),
    .D(net36));
 sg13g2_buf_1 _7873_ (.A(_2843_),
    .X(_2844_));
 sg13g2_nand2_1 _7874_ (.Y(_2845_),
    .A(_2842_),
    .B(_2844_));
 sg13g2_xor2_1 _7875_ (.B(_2845_),
    .A(_2837_),
    .X(_2846_));
 sg13g2_xnor2_1 _7876_ (.Y(_2847_),
    .A(_2836_),
    .B(_2846_));
 sg13g2_inv_1 _7877_ (.Y(_2848_),
    .A(_2847_));
 sg13g2_or2_1 _7878_ (.X(_2849_),
    .B(_2788_),
    .A(_2784_));
 sg13g2_nand3_1 _7879_ (.B(_2849_),
    .C(_2802_),
    .A(_2848_),
    .Y(_2850_));
 sg13g2_nand2_1 _7880_ (.Y(_2851_),
    .A(_2802_),
    .B(_2849_));
 sg13g2_nand2_1 _7881_ (.Y(_2852_),
    .A(_2851_),
    .B(_2847_));
 sg13g2_nand2_1 _7882_ (.Y(_2853_),
    .A(_2850_),
    .B(_2852_));
 sg13g2_inv_1 _7883_ (.Y(_2854_),
    .A(_2797_));
 sg13g2_a21oi_1 _7884_ (.A1(_2795_),
    .A2(_2791_),
    .Y(_2855_),
    .B1(_2854_));
 sg13g2_nand2_1 _7885_ (.Y(_2856_),
    .A(_2853_),
    .B(_2855_));
 sg13g2_inv_1 _7886_ (.Y(_2857_),
    .A(_2855_));
 sg13g2_nand3_1 _7887_ (.B(_2852_),
    .C(_2857_),
    .A(_2850_),
    .Y(_2858_));
 sg13g2_nand2_1 _7888_ (.Y(_2859_),
    .A(_2856_),
    .B(_2858_));
 sg13g2_xnor2_1 _7889_ (.Y(_2860_),
    .A(_2829_),
    .B(_2859_));
 sg13g2_inv_4 _7890_ (.A(_2860_),
    .Y(_2861_));
 sg13g2_nand2_1 _7891_ (.Y(_2862_),
    .A(_2827_),
    .B(_2861_));
 sg13g2_nand3_1 _7892_ (.B(_2860_),
    .C(_2826_),
    .A(_2823_),
    .Y(_2863_));
 sg13g2_nand3_1 _7893_ (.B(_2863_),
    .C(_2373_),
    .A(_2862_),
    .Y(_2864_));
 sg13g2_nand3_1 _7894_ (.B(_2818_),
    .C(_2531_),
    .A(_2816_),
    .Y(_2865_));
 sg13g2_buf_1 _7895_ (.A(_2865_),
    .X(_2866_));
 sg13g2_nand3_1 _7896_ (.B(_2864_),
    .C(_2866_),
    .A(_2821_),
    .Y(_2867_));
 sg13g2_nand2_1 _7897_ (.Y(_2868_),
    .A(_2862_),
    .B(_2863_));
 sg13g2_nand2_1 _7898_ (.Y(_2869_),
    .A(_2868_),
    .B(_2372_));
 sg13g2_nand2_1 _7899_ (.Y(_2870_),
    .A(_2867_),
    .B(_2869_));
 sg13g2_nand2_1 _7900_ (.Y(_2871_),
    .A(_2589_),
    .B(net71));
 sg13g2_nor2_1 _7901_ (.A(_2871_),
    .B(_2834_),
    .Y(_2872_));
 sg13g2_nor2_1 _7902_ (.A(net63),
    .B(_2590_),
    .Y(_2873_));
 sg13g2_inv_1 _7903_ (.Y(_2874_),
    .A(_2873_));
 sg13g2_a22oi_1 _7904_ (.Y(_2875_),
    .B1(net71),
    .B2(_2832_),
    .A2(_2589_),
    .A1(_2833_));
 sg13g2_or2_1 _7905_ (.X(_2876_),
    .B(_2875_),
    .A(_2872_));
 sg13g2_buf_1 _7906_ (.A(_2876_),
    .X(_2877_));
 sg13g2_nor2_1 _7907_ (.A(_2874_),
    .B(_2877_),
    .Y(_2878_));
 sg13g2_nor2_1 _7908_ (.A(_2872_),
    .B(_2878_),
    .Y(_2879_));
 sg13g2_nor2_1 _7909_ (.A(net63),
    .B(_2785_),
    .Y(_2880_));
 sg13g2_inv_1 _7910_ (.Y(_2881_),
    .A(_2880_));
 sg13g2_inv_1 _7911_ (.Y(_2882_),
    .A(net26));
 sg13g2_o21ai_1 _7912_ (.B1(_2871_),
    .Y(_2883_),
    .A1(_2708_),
    .A2(_2882_));
 sg13g2_nand3_1 _7913_ (.B(_2833_),
    .C(net71),
    .A(net26),
    .Y(_2884_));
 sg13g2_nand2_1 _7914_ (.Y(_2885_),
    .A(_2883_),
    .B(_2884_));
 sg13g2_xnor2_1 _7915_ (.Y(_2886_),
    .A(_2881_),
    .B(_2885_));
 sg13g2_nor2_1 _7916_ (.A(_2554_),
    .B(_2882_),
    .Y(_2887_));
 sg13g2_buf_2 _7917_ (.A(_2887_),
    .X(_2888_));
 sg13g2_inv_1 _7918_ (.Y(_2889_),
    .A(_2888_));
 sg13g2_nor2_2 _7919_ (.A(_2482_),
    .B(_2594_),
    .Y(_2890_));
 sg13g2_nor2_1 _7920_ (.A(_2889_),
    .B(_2890_),
    .Y(_2891_));
 sg13g2_xnor2_1 _7921_ (.Y(_2892_),
    .A(_2783_),
    .B(_2891_));
 sg13g2_xnor2_1 _7922_ (.Y(_2893_),
    .A(_2886_),
    .B(_2892_));
 sg13g2_xnor2_1 _7923_ (.Y(_2894_),
    .A(_2873_),
    .B(_2877_));
 sg13g2_xnor2_1 _7924_ (.Y(_2895_),
    .A(_2888_),
    .B(_2890_));
 sg13g2_nand2_1 _7925_ (.Y(_2896_),
    .A(_2895_),
    .B(_2844_));
 sg13g2_nor2_1 _7926_ (.A(_2844_),
    .B(_2895_),
    .Y(_2897_));
 sg13g2_a21oi_1 _7927_ (.A1(_2894_),
    .A2(_2896_),
    .Y(_2898_),
    .B1(_2897_));
 sg13g2_xnor2_1 _7928_ (.Y(_2899_),
    .A(_2893_),
    .B(_2898_));
 sg13g2_xor2_1 _7929_ (.B(_2899_),
    .A(_2879_),
    .X(_2900_));
 sg13g2_inv_1 _7930_ (.Y(_2901_),
    .A(_2836_));
 sg13g2_nand3_1 _7931_ (.B(_2844_),
    .C(_2837_),
    .A(_2842_),
    .Y(_2902_));
 sg13g2_o21ai_1 _7932_ (.B1(_2902_),
    .Y(_2903_),
    .A1(_2901_),
    .A2(_2846_));
 sg13g2_xnor2_1 _7933_ (.Y(_2904_),
    .A(_2844_),
    .B(_2895_));
 sg13g2_xor2_1 _7934_ (.B(_2904_),
    .A(_2894_),
    .X(_2905_));
 sg13g2_nand2b_1 _7935_ (.Y(_2906_),
    .B(_2905_),
    .A_N(_2903_));
 sg13g2_inv_1 _7936_ (.Y(_2907_),
    .A(_2835_));
 sg13g2_nand3_1 _7937_ (.B(net71),
    .C(_2832_),
    .A(_2792_),
    .Y(_2908_));
 sg13g2_o21ai_1 _7938_ (.B1(_2908_),
    .Y(_2909_),
    .A1(_2830_),
    .A2(_2907_));
 sg13g2_nand2b_1 _7939_ (.Y(_2910_),
    .B(_2903_),
    .A_N(_2905_));
 sg13g2_inv_1 _7940_ (.Y(_2911_),
    .A(_2910_));
 sg13g2_a21oi_1 _7941_ (.A1(_2906_),
    .A2(_2909_),
    .Y(_2912_),
    .B1(_2911_));
 sg13g2_xnor2_1 _7942_ (.Y(_2913_),
    .A(_2900_),
    .B(_2912_));
 sg13g2_nand2_1 _7943_ (.Y(_2914_),
    .A(_2858_),
    .B(_2852_));
 sg13g2_nand2_1 _7944_ (.Y(_2915_),
    .A(_2910_),
    .B(_2906_));
 sg13g2_nand2b_1 _7945_ (.Y(_2916_),
    .B(_2915_),
    .A_N(_2909_));
 sg13g2_nand3_1 _7946_ (.B(_2906_),
    .C(_2909_),
    .A(_2910_),
    .Y(_2917_));
 sg13g2_nand2_1 _7947_ (.Y(_2918_),
    .A(_2916_),
    .B(_2917_));
 sg13g2_xnor2_1 _7948_ (.Y(_2919_),
    .A(_2914_),
    .B(_2918_));
 sg13g2_nand4_1 _7949_ (.B(_2727_),
    .C(_2919_),
    .A(_2822_),
    .Y(_2920_),
    .D(_2861_));
 sg13g2_nand2_1 _7950_ (.Y(_2921_),
    .A(_2919_),
    .B(_2861_));
 sg13g2_nor2_1 _7951_ (.A(_2826_),
    .B(_2921_),
    .Y(_2922_));
 sg13g2_nand2b_1 _7952_ (.Y(_2923_),
    .B(_2918_),
    .A_N(_2914_));
 sg13g2_nor2_1 _7953_ (.A(_2829_),
    .B(_2859_),
    .Y(_2924_));
 sg13g2_nor2b_1 _7954_ (.A(_2918_),
    .B_N(_2914_),
    .Y(_2925_));
 sg13g2_a21oi_1 _7955_ (.A1(_2923_),
    .A2(_2924_),
    .Y(_2926_),
    .B1(_2925_));
 sg13g2_nor2b_1 _7956_ (.A(_2922_),
    .B_N(_2926_),
    .Y(_2927_));
 sg13g2_nand2_1 _7957_ (.Y(_2928_),
    .A(_2920_),
    .B(_2927_));
 sg13g2_xnor2_1 _7958_ (.Y(_2929_),
    .A(_2913_),
    .B(_2928_));
 sg13g2_xnor2_1 _7959_ (.Y(_2930_),
    .A(_2502_),
    .B(_2929_));
 sg13g2_nor2_1 _7960_ (.A(_2860_),
    .B(_2815_),
    .Y(_2931_));
 sg13g2_nor2b_1 _7961_ (.A(_2775_),
    .B_N(_2777_),
    .Y(_2932_));
 sg13g2_nand2_1 _7962_ (.Y(_2933_),
    .A(_2859_),
    .B(_2829_));
 sg13g2_a21oi_1 _7963_ (.A1(_2824_),
    .A2(_2933_),
    .Y(_2934_),
    .B1(_2924_));
 sg13g2_inv_1 _7964_ (.Y(_2935_),
    .A(_2934_));
 sg13g2_a21oi_1 _7965_ (.A1(_2931_),
    .A2(_2932_),
    .Y(_2936_),
    .B1(_2935_));
 sg13g2_nor2_1 _7966_ (.A(_2763_),
    .B(_2728_),
    .Y(_2937_));
 sg13g2_nand3_1 _7967_ (.B(_2723_),
    .C(_2937_),
    .A(_2931_),
    .Y(_2938_));
 sg13g2_nand3b_1 _7968_ (.B(_2936_),
    .C(_2938_),
    .Y(_2939_),
    .A_N(_2919_));
 sg13g2_nand2_1 _7969_ (.Y(_2940_),
    .A(_2936_),
    .B(_2938_));
 sg13g2_nand2_1 _7970_ (.Y(_2941_),
    .A(_2940_),
    .B(_2919_));
 sg13g2_nand2_1 _7971_ (.Y(_2942_),
    .A(_2939_),
    .B(_2941_));
 sg13g2_nand2b_1 _7972_ (.Y(_2943_),
    .B(_2942_),
    .A_N(_2463_));
 sg13g2_nand3_1 _7973_ (.B(_2941_),
    .C(_2463_),
    .A(_2939_),
    .Y(_2944_));
 sg13g2_nand2_1 _7974_ (.Y(_2945_),
    .A(_2943_),
    .B(_2944_));
 sg13g2_nand3b_1 _7975_ (.B(_2930_),
    .C(_2945_),
    .Y(_2946_),
    .A_N(_2870_));
 sg13g2_a21oi_1 _7976_ (.A1(_2708_),
    .A2(_2526_),
    .Y(_2947_),
    .B1(_2882_));
 sg13g2_nand2_1 _7977_ (.Y(_2948_),
    .A(_2947_),
    .B(_2884_));
 sg13g2_o21ai_1 _7978_ (.B1(_2884_),
    .Y(_2949_),
    .A1(_2889_),
    .A2(_2948_));
 sg13g2_buf_2 _7979_ (.A(_2949_),
    .X(_2950_));
 sg13g2_nor3_1 _7980_ (.A(_2482_),
    .B(_2874_),
    .C(_2594_),
    .Y(_2951_));
 sg13g2_xnor2_1 _7981_ (.Y(_2952_),
    .A(_2888_),
    .B(_2885_));
 sg13g2_nand2_1 _7982_ (.Y(_2953_),
    .A(_2830_),
    .B(_2783_));
 sg13g2_xnor2_1 _7983_ (.Y(_2954_),
    .A(_2880_),
    .B(_2953_));
 sg13g2_a22oi_1 _7984_ (.Y(_2955_),
    .B1(_2952_),
    .B2(_2954_),
    .A2(_2951_),
    .A1(_2785_));
 sg13g2_xnor2_1 _7985_ (.Y(_2956_),
    .A(_2888_),
    .B(_2948_));
 sg13g2_nand2_1 _7986_ (.Y(_2957_),
    .A(_2783_),
    .B(_2880_));
 sg13g2_a22oi_1 _7987_ (.Y(_2958_),
    .B1(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .B2(_2832_),
    .A2(_2589_),
    .A1(_2515_));
 sg13g2_nor2_1 _7988_ (.A(_2475_),
    .B(_2839_),
    .Y(_2959_));
 sg13g2_inv_1 _7989_ (.Y(_2960_),
    .A(_2959_));
 sg13g2_nor2_1 _7990_ (.A(_2960_),
    .B(_2881_),
    .Y(_2961_));
 sg13g2_inv_1 _7991_ (.Y(_2962_),
    .A(_2961_));
 sg13g2_nand2b_1 _7992_ (.Y(_2963_),
    .B(_2962_),
    .A_N(_2958_));
 sg13g2_nor2_1 _7993_ (.A(_2957_),
    .B(_2963_),
    .Y(_2964_));
 sg13g2_nand2_1 _7994_ (.Y(_2965_),
    .A(_2963_),
    .B(_2957_));
 sg13g2_nand2b_1 _7995_ (.Y(_2966_),
    .B(_2965_),
    .A_N(_2964_));
 sg13g2_xnor2_1 _7996_ (.Y(_2967_),
    .A(_2956_),
    .B(_2966_));
 sg13g2_xnor2_1 _7997_ (.Y(_2968_),
    .A(_2955_),
    .B(_2967_));
 sg13g2_xnor2_1 _7998_ (.Y(_2969_),
    .A(_2950_),
    .B(_2968_));
 sg13g2_xnor2_1 _7999_ (.Y(_2970_),
    .A(_2952_),
    .B(_2954_));
 sg13g2_xnor2_1 _8000_ (.Y(_2971_),
    .A(_2888_),
    .B(_2877_));
 sg13g2_nor2_1 _8001_ (.A(_2873_),
    .B(_2890_),
    .Y(_2972_));
 sg13g2_nand2_1 _8002_ (.Y(_2973_),
    .A(_2890_),
    .B(_2791_));
 sg13g2_o21ai_1 _8003_ (.B1(_2973_),
    .Y(_2974_),
    .A1(_2951_),
    .A2(_2972_));
 sg13g2_nand3_1 _8004_ (.B(_2791_),
    .C(_2874_),
    .A(_2890_),
    .Y(_2975_));
 sg13g2_nand3_1 _8005_ (.B(_2974_),
    .C(_2975_),
    .A(_2971_),
    .Y(_2976_));
 sg13g2_and2_1 _8006_ (.A(_2976_),
    .B(_2975_),
    .X(_2977_));
 sg13g2_nor2_1 _8007_ (.A(_2970_),
    .B(_2977_),
    .Y(_2978_));
 sg13g2_nor2_1 _8008_ (.A(_2889_),
    .B(_2877_),
    .Y(_2979_));
 sg13g2_nor2_1 _8009_ (.A(_2872_),
    .B(_2979_),
    .Y(_2980_));
 sg13g2_xnor2_1 _8010_ (.Y(_2981_),
    .A(_2970_),
    .B(_2977_));
 sg13g2_nor2_1 _8011_ (.A(_2980_),
    .B(_2981_),
    .Y(_2982_));
 sg13g2_nor2_1 _8012_ (.A(_2978_),
    .B(_2982_),
    .Y(_2983_));
 sg13g2_nor2_1 _8013_ (.A(_2969_),
    .B(_2983_),
    .Y(_2984_));
 sg13g2_nand2_1 _8014_ (.Y(_2985_),
    .A(_2983_),
    .B(_2969_));
 sg13g2_nor2b_2 _8015_ (.A(_2984_),
    .B_N(_2985_),
    .Y(_2986_));
 sg13g2_a21oi_1 _8016_ (.A1(_2740_),
    .A2(_2542_),
    .Y(_2987_),
    .B1(_2611_));
 sg13g2_o21ai_1 _8017_ (.B1(_2748_),
    .Y(_2988_),
    .A1(_2743_),
    .A2(_2744_));
 sg13g2_nand2_1 _8018_ (.Y(_2989_),
    .A(_2519_),
    .B(_2488_));
 sg13g2_xnor2_1 _8019_ (.Y(_2990_),
    .A(_2587_),
    .B(_2601_));
 sg13g2_xnor2_1 _8020_ (.Y(_2991_),
    .A(_2989_),
    .B(_2990_));
 sg13g2_xnor2_1 _8021_ (.Y(_2992_),
    .A(_2591_),
    .B(_2600_));
 sg13g2_xnor2_1 _8022_ (.Y(_2993_),
    .A(_2991_),
    .B(_2992_));
 sg13g2_xor2_1 _8023_ (.B(_2993_),
    .A(_2988_),
    .X(_2994_));
 sg13g2_xnor2_1 _8024_ (.Y(_2995_),
    .A(_2987_),
    .B(_2994_));
 sg13g2_and2_1 _8025_ (.A(_2756_),
    .B(_2751_),
    .X(_2996_));
 sg13g2_nand2_1 _8026_ (.Y(_2997_),
    .A(_2995_),
    .B(_2996_));
 sg13g2_inv_1 _8027_ (.Y(_2998_),
    .A(_2762_));
 sg13g2_nor2_1 _8028_ (.A(_2996_),
    .B(_2995_),
    .Y(_2999_));
 sg13g2_a21oi_1 _8029_ (.A1(_2997_),
    .A2(_2998_),
    .Y(_3000_),
    .B1(_2999_));
 sg13g2_nand2b_1 _8030_ (.Y(_3001_),
    .B(_2988_),
    .A_N(_2993_));
 sg13g2_o21ai_1 _8031_ (.B1(_3001_),
    .Y(_3002_),
    .A1(_2987_),
    .A2(_2994_));
 sg13g2_nand2_1 _8032_ (.Y(_3003_),
    .A(_2992_),
    .B(_2991_));
 sg13g2_inv_1 _8033_ (.Y(_3004_),
    .A(_2587_));
 sg13g2_nand3_1 _8034_ (.B(_2562_),
    .C(_3004_),
    .A(_2603_),
    .Y(_3005_));
 sg13g2_nand2_1 _8035_ (.Y(_3006_),
    .A(_3003_),
    .B(_3005_));
 sg13g2_nand2_1 _8036_ (.Y(_3007_),
    .A(_2601_),
    .B(_3004_));
 sg13g2_inv_1 _8037_ (.Y(_3008_),
    .A(_2787_));
 sg13g2_xnor2_1 _8038_ (.Y(_3009_),
    .A(_3008_),
    .B(_2791_));
 sg13g2_nor2_1 _8039_ (.A(_3007_),
    .B(_3009_),
    .Y(_3010_));
 sg13g2_inv_1 _8040_ (.Y(_3011_),
    .A(_3010_));
 sg13g2_nand2_1 _8041_ (.Y(_3012_),
    .A(_3009_),
    .B(_3007_));
 sg13g2_nand2_1 _8042_ (.Y(_3013_),
    .A(_3011_),
    .B(_3012_));
 sg13g2_xnor2_1 _8043_ (.Y(_3014_),
    .A(_2786_),
    .B(_2798_));
 sg13g2_xnor2_1 _8044_ (.Y(_3015_),
    .A(_3013_),
    .B(_3014_));
 sg13g2_or2_1 _8045_ (.X(_3016_),
    .B(_3015_),
    .A(_3006_));
 sg13g2_buf_1 _8046_ (.A(_3016_),
    .X(_3017_));
 sg13g2_nand2_1 _8047_ (.Y(_3018_),
    .A(_3015_),
    .B(_3006_));
 sg13g2_nand2_1 _8048_ (.Y(_3019_),
    .A(_3017_),
    .B(_3018_));
 sg13g2_a21oi_1 _8049_ (.A1(_2591_),
    .A2(_2599_),
    .Y(_3020_),
    .B1(_2809_));
 sg13g2_nand2_1 _8050_ (.Y(_3021_),
    .A(_3019_),
    .B(_3020_));
 sg13g2_inv_1 _8051_ (.Y(_3022_),
    .A(_3020_));
 sg13g2_nand3_1 _8052_ (.B(_3018_),
    .C(_3022_),
    .A(_3017_),
    .Y(_3023_));
 sg13g2_nand2_1 _8053_ (.Y(_3024_),
    .A(_3021_),
    .B(_3023_));
 sg13g2_xnor2_1 _8054_ (.Y(_3025_),
    .A(_3002_),
    .B(_3024_));
 sg13g2_inv_1 _8055_ (.Y(_3026_),
    .A(_3018_));
 sg13g2_a21oi_2 _8056_ (.B1(_3026_),
    .Y(_3027_),
    .A2(_3022_),
    .A1(_3017_));
 sg13g2_xnor2_1 _8057_ (.Y(_3028_),
    .A(_2841_),
    .B(_2835_));
 sg13g2_nand2_1 _8058_ (.Y(_3029_),
    .A(_2791_),
    .B(_3008_));
 sg13g2_nand2_1 _8059_ (.Y(_3030_),
    .A(_2830_),
    .B(_2838_));
 sg13g2_nand2_1 _8060_ (.Y(_3031_),
    .A(_3030_),
    .B(_2973_));
 sg13g2_nor2_1 _8061_ (.A(_3029_),
    .B(_3031_),
    .Y(_3032_));
 sg13g2_inv_1 _8062_ (.Y(_3033_),
    .A(_3032_));
 sg13g2_nand2_1 _8063_ (.Y(_3034_),
    .A(_3031_),
    .B(_3029_));
 sg13g2_nand2_1 _8064_ (.Y(_3035_),
    .A(_3033_),
    .B(_3034_));
 sg13g2_xor2_1 _8065_ (.B(_3035_),
    .A(_3028_),
    .X(_3036_));
 sg13g2_a21oi_1 _8066_ (.A1(_3014_),
    .A2(_3012_),
    .Y(_3037_),
    .B1(_3010_));
 sg13g2_nand2_1 _8067_ (.Y(_3038_),
    .A(_3036_),
    .B(_3037_));
 sg13g2_xnor2_1 _8068_ (.Y(_3039_),
    .A(_3028_),
    .B(_3035_));
 sg13g2_inv_1 _8069_ (.Y(_3040_),
    .A(_3037_));
 sg13g2_nand2_1 _8070_ (.Y(_3041_),
    .A(_3039_),
    .B(_3040_));
 sg13g2_nand2_1 _8071_ (.Y(_3042_),
    .A(_3038_),
    .B(_3041_));
 sg13g2_a21oi_1 _8072_ (.A1(_2795_),
    .A2(_2786_),
    .Y(_3043_),
    .B1(_2854_));
 sg13g2_nand2_1 _8073_ (.Y(_3044_),
    .A(_3042_),
    .B(_3043_));
 sg13g2_inv_1 _8074_ (.Y(_3045_),
    .A(_3043_));
 sg13g2_nand3_1 _8075_ (.B(_3041_),
    .C(_3045_),
    .A(_3038_),
    .Y(_3046_));
 sg13g2_nand2_1 _8076_ (.Y(_3047_),
    .A(_3044_),
    .B(_3046_));
 sg13g2_xor2_1 _8077_ (.B(_3047_),
    .A(_3027_),
    .X(_3048_));
 sg13g2_nand2_1 _8078_ (.Y(_3049_),
    .A(_3025_),
    .B(_3048_));
 sg13g2_nor2_1 _8079_ (.A(_3000_),
    .B(_3049_),
    .Y(_3050_));
 sg13g2_nor2b_1 _8080_ (.A(_3024_),
    .B_N(_3002_),
    .Y(_3051_));
 sg13g2_nand2_1 _8081_ (.Y(_3052_),
    .A(_3047_),
    .B(_3027_));
 sg13g2_nor2_1 _8082_ (.A(_3027_),
    .B(_3047_),
    .Y(_3053_));
 sg13g2_a21oi_1 _8083_ (.A1(_3051_),
    .A2(_3052_),
    .Y(_3054_),
    .B1(_3053_));
 sg13g2_nor2b_1 _8084_ (.A(_3050_),
    .B_N(_3054_),
    .Y(_3055_));
 sg13g2_nand2_1 _8085_ (.Y(_3056_),
    .A(_3055_),
    .B(_2938_));
 sg13g2_inv_1 _8086_ (.Y(_3057_),
    .A(_2908_));
 sg13g2_a21oi_1 _8087_ (.A1(_2835_),
    .A2(_2840_),
    .Y(_3058_),
    .B1(_3057_));
 sg13g2_a21oi_1 _8088_ (.A1(_3034_),
    .A2(_3028_),
    .Y(_3059_),
    .B1(_3032_));
 sg13g2_a21oi_1 _8089_ (.A1(_2974_),
    .A2(_2975_),
    .Y(_3060_),
    .B1(_2971_));
 sg13g2_nand2b_1 _8090_ (.Y(_3061_),
    .B(_2976_),
    .A_N(_3060_));
 sg13g2_xnor2_1 _8091_ (.Y(_3062_),
    .A(_3059_),
    .B(_3061_));
 sg13g2_xnor2_1 _8092_ (.Y(_3063_),
    .A(_3058_),
    .B(_3062_));
 sg13g2_nand2_1 _8093_ (.Y(_3064_),
    .A(_3046_),
    .B(_3041_));
 sg13g2_nor2b_1 _8094_ (.A(_3063_),
    .B_N(_3064_),
    .Y(_3065_));
 sg13g2_nor2b_1 _8095_ (.A(_3064_),
    .B_N(_3063_),
    .Y(_3066_));
 sg13g2_nor2_1 _8096_ (.A(_3059_),
    .B(_3061_),
    .Y(_3067_));
 sg13g2_nor2_1 _8097_ (.A(_3058_),
    .B(_3062_),
    .Y(_3068_));
 sg13g2_nor2_1 _8098_ (.A(_3067_),
    .B(_3068_),
    .Y(_3069_));
 sg13g2_xnor2_1 _8099_ (.Y(_3070_),
    .A(_2980_),
    .B(_2981_));
 sg13g2_xnor2_1 _8100_ (.Y(_3071_),
    .A(_3069_),
    .B(_3070_));
 sg13g2_nor3_1 _8101_ (.A(_3065_),
    .B(_3066_),
    .C(_3071_),
    .Y(_3072_));
 sg13g2_inv_1 _8102_ (.Y(_3073_),
    .A(_3065_));
 sg13g2_or2_1 _8103_ (.X(_3074_),
    .B(_3070_),
    .A(_3069_));
 sg13g2_o21ai_1 _8104_ (.B1(_3074_),
    .Y(_3075_),
    .A1(_3073_),
    .A2(_3071_));
 sg13g2_a21oi_2 _8105_ (.B1(_3075_),
    .Y(_3076_),
    .A2(_3072_),
    .A1(_3056_));
 sg13g2_xor2_1 _8106_ (.B(_3076_),
    .A(_2986_),
    .X(_3077_));
 sg13g2_nand2_1 _8107_ (.Y(_3078_),
    .A(_3077_),
    .B(_2343_));
 sg13g2_xnor2_1 _8108_ (.Y(_3079_),
    .A(_2986_),
    .B(_3076_));
 sg13g2_nand2_1 _8109_ (.Y(_3080_),
    .A(_3079_),
    .B(_2411_));
 sg13g2_nand2_1 _8110_ (.Y(_3081_),
    .A(_3078_),
    .B(_3080_));
 sg13g2_nor2_1 _8111_ (.A(_2463_),
    .B(_2942_),
    .Y(_3082_));
 sg13g2_inv_1 _8112_ (.Y(_3083_),
    .A(_2502_));
 sg13g2_nor2_1 _8113_ (.A(_3083_),
    .B(_2929_),
    .Y(_3084_));
 sg13g2_nand2_1 _8114_ (.Y(_3085_),
    .A(_2929_),
    .B(_3083_));
 sg13g2_o21ai_1 _8115_ (.B1(_3085_),
    .Y(_3086_),
    .A1(_3082_),
    .A2(_3084_));
 sg13g2_nand3_1 _8116_ (.B(_3081_),
    .C(_3086_),
    .A(_2946_),
    .Y(_3087_));
 sg13g2_nand3_1 _8117_ (.B(_2869_),
    .C(_2867_),
    .A(_2945_),
    .Y(_3088_));
 sg13g2_nor2_1 _8118_ (.A(_3082_),
    .B(_3084_),
    .Y(_3089_));
 sg13g2_nand2_1 _8119_ (.Y(_3090_),
    .A(_3088_),
    .B(_3089_));
 sg13g2_xnor2_1 _8120_ (.Y(_3091_),
    .A(_2343_),
    .B(_3079_));
 sg13g2_nand3_1 _8121_ (.B(_3091_),
    .C(_3085_),
    .A(_3090_),
    .Y(_3092_));
 sg13g2_nand3_1 _8122_ (.B(_3092_),
    .C(_4247_),
    .A(_3087_),
    .Y(_3093_));
 sg13g2_nand3_1 _8123_ (.B(_3091_),
    .C(_3086_),
    .A(_2946_),
    .Y(_3094_));
 sg13g2_nand3_1 _8124_ (.B(_3081_),
    .C(_3085_),
    .A(_3090_),
    .Y(_3095_));
 sg13g2_inv_1 _8125_ (.Y(_3096_),
    .A(_4247_));
 sg13g2_nand3_1 _8126_ (.B(_3095_),
    .C(_3096_),
    .A(_3094_),
    .Y(_3097_));
 sg13g2_nand2_1 _8127_ (.Y(_3098_),
    .A(_3093_),
    .B(_3097_));
 sg13g2_nand2_1 _8128_ (.Y(_3099_),
    .A(_2819_),
    .B(_2531_));
 sg13g2_nand3_1 _8129_ (.B(_2818_),
    .C(_2359_),
    .A(_2816_),
    .Y(_3100_));
 sg13g2_nand2_1 _8130_ (.Y(_3101_),
    .A(_3099_),
    .B(_3100_));
 sg13g2_nand2b_1 _8131_ (.Y(_3102_),
    .B(_3101_),
    .A_N(_2771_));
 sg13g2_nand2_1 _8132_ (.Y(_3103_),
    .A(_2820_),
    .B(_2866_));
 sg13g2_nand2_1 _8133_ (.Y(_3104_),
    .A(_3103_),
    .B(_2771_));
 sg13g2_nand2_1 _8134_ (.Y(_3105_),
    .A(_3102_),
    .B(_3104_));
 sg13g2_nand2_1 _8135_ (.Y(_3106_),
    .A(_3105_),
    .B(_4229_));
 sg13g2_nand3_1 _8136_ (.B(_3104_),
    .C(_2177_),
    .A(_3102_),
    .Y(_3107_));
 sg13g2_nand2_1 _8137_ (.Y(_3108_),
    .A(_2770_),
    .B(_2730_));
 sg13g2_nand2b_1 _8138_ (.Y(_3109_),
    .B(_3108_),
    .A_N(_2767_));
 sg13g2_nand3_1 _8139_ (.B(_2730_),
    .C(_2767_),
    .A(_2770_),
    .Y(_3110_));
 sg13g2_nand2_1 _8140_ (.Y(_3111_),
    .A(_3109_),
    .B(_3110_));
 sg13g2_nor2_1 _8141_ (.A(_0300_),
    .B(_3111_),
    .Y(_3112_));
 sg13g2_nand3_1 _8142_ (.B(_3107_),
    .C(_3112_),
    .A(_3106_),
    .Y(_3113_));
 sg13g2_inv_1 _8143_ (.Y(_3114_),
    .A(_0026_));
 sg13g2_nand2_1 _8144_ (.Y(_3115_),
    .A(_3105_),
    .B(_3114_));
 sg13g2_nand2_1 _8145_ (.Y(_3116_),
    .A(_3113_),
    .B(_3115_));
 sg13g2_nand2_1 _8146_ (.Y(_3117_),
    .A(_2821_),
    .B(_2866_));
 sg13g2_nand2_1 _8147_ (.Y(_3118_),
    .A(_2869_),
    .B(_2864_));
 sg13g2_xor2_1 _8148_ (.B(_3118_),
    .A(_3117_),
    .X(_3119_));
 sg13g2_nand2_1 _8149_ (.Y(_3120_),
    .A(_3119_),
    .B(_4226_));
 sg13g2_xnor2_1 _8150_ (.Y(_3121_),
    .A(_3117_),
    .B(_3118_));
 sg13g2_nand2_1 _8151_ (.Y(_3122_),
    .A(_3121_),
    .B(_2178_));
 sg13g2_nand2_1 _8152_ (.Y(_3123_),
    .A(_3120_),
    .B(_3122_));
 sg13g2_nand2_1 _8153_ (.Y(_3124_),
    .A(_3116_),
    .B(_3123_));
 sg13g2_inv_1 _8154_ (.Y(_3125_),
    .A(_0025_));
 sg13g2_nand2_1 _8155_ (.Y(_3126_),
    .A(_3121_),
    .B(_3125_));
 sg13g2_nand2_1 _8156_ (.Y(_3127_),
    .A(_3124_),
    .B(_3126_));
 sg13g2_inv_1 _8157_ (.Y(_3128_),
    .A(_2945_));
 sg13g2_nand2_1 _8158_ (.Y(_3129_),
    .A(_2870_),
    .B(_3128_));
 sg13g2_nand2_1 _8159_ (.Y(_3130_),
    .A(_3088_),
    .B(_3129_));
 sg13g2_xnor2_1 _8160_ (.Y(_3131_),
    .A(_4223_),
    .B(_3130_));
 sg13g2_nand2_1 _8161_ (.Y(_3132_),
    .A(_3127_),
    .B(_3131_));
 sg13g2_inv_1 _8162_ (.Y(_3133_),
    .A(_3130_));
 sg13g2_inv_1 _8163_ (.Y(_3134_),
    .A(_0024_));
 sg13g2_nand2_1 _8164_ (.Y(_3135_),
    .A(_3133_),
    .B(_3134_));
 sg13g2_nand2_1 _8165_ (.Y(_3136_),
    .A(_3132_),
    .B(_3135_));
 sg13g2_inv_1 _8166_ (.Y(_3137_),
    .A(_0023_));
 sg13g2_inv_1 _8167_ (.Y(_3138_),
    .A(_3118_));
 sg13g2_nand2_1 _8168_ (.Y(_3139_),
    .A(_3138_),
    .B(_3117_));
 sg13g2_nor2b_1 _8169_ (.A(_3082_),
    .B_N(_2864_),
    .Y(_3140_));
 sg13g2_nand2_1 _8170_ (.Y(_3141_),
    .A(_3139_),
    .B(_3140_));
 sg13g2_nand2_1 _8171_ (.Y(_3142_),
    .A(_2942_),
    .B(_2463_));
 sg13g2_nand2_1 _8172_ (.Y(_3143_),
    .A(_3141_),
    .B(_3142_));
 sg13g2_inv_1 _8173_ (.Y(_3144_),
    .A(_2930_));
 sg13g2_nand2_1 _8174_ (.Y(_3145_),
    .A(_3143_),
    .B(_3144_));
 sg13g2_nand3_1 _8175_ (.B(_2930_),
    .C(_3142_),
    .A(_3141_),
    .Y(_3146_));
 sg13g2_nand2_1 _8176_ (.Y(_3147_),
    .A(_3145_),
    .B(_3146_));
 sg13g2_xnor2_1 _8177_ (.Y(_3148_),
    .A(_3137_),
    .B(_3147_));
 sg13g2_nand2_1 _8178_ (.Y(_3149_),
    .A(_3136_),
    .B(_3148_));
 sg13g2_inv_1 _8179_ (.Y(_3150_),
    .A(_3147_));
 sg13g2_nand2_1 _8180_ (.Y(_3151_),
    .A(_3150_),
    .B(_3137_));
 sg13g2_nand2_1 _8181_ (.Y(_3152_),
    .A(_3149_),
    .B(_3151_));
 sg13g2_xnor2_1 _8182_ (.Y(_3153_),
    .A(_3098_),
    .B(_3152_));
 sg13g2_nand2b_1 _8183_ (.Y(_3154_),
    .B(_3153_),
    .A_N(_2189_));
 sg13g2_inv_1 _8184_ (.Y(_3155_),
    .A(_3098_));
 sg13g2_nand2_2 _8185_ (.Y(_3156_),
    .A(_3152_),
    .B(_3155_));
 sg13g2_nand3_1 _8186_ (.B(_3151_),
    .C(_3098_),
    .A(_3149_),
    .Y(_3157_));
 sg13g2_buf_1 _8187_ (.A(_3157_),
    .X(_3158_));
 sg13g2_nand2_1 _8188_ (.Y(_3159_),
    .A(_3156_),
    .B(_3158_));
 sg13g2_buf_8 _8189_ (.A(_3159_),
    .X(_3160_));
 sg13g2_nand2_1 _8190_ (.Y(_3161_),
    .A(net12),
    .B(_2181_));
 sg13g2_nand3_1 _8191_ (.B(\main.demo._d___pip_58_1_3___stage___block_3_a[2] ),
    .C(_3161_),
    .A(_3154_),
    .Y(_3162_));
 sg13g2_buf_1 _8192_ (.A(_3162_),
    .X(_3163_));
 sg13g2_nand2_1 _8193_ (.Y(_3164_),
    .A(net12),
    .B(_2180_));
 sg13g2_nand3_1 _8194_ (.B(_3158_),
    .C(_2189_),
    .A(_3156_),
    .Y(_3165_));
 sg13g2_inv_1 _8195_ (.Y(_3166_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[2] ));
 sg13g2_nand3_1 _8196_ (.B(_3165_),
    .C(_3166_),
    .A(_3164_),
    .Y(_3167_));
 sg13g2_nand2_1 _8197_ (.Y(_3168_),
    .A(_3163_),
    .B(_3167_));
 sg13g2_inv_1 _8198_ (.Y(_3169_),
    .A(_2185_));
 sg13g2_nand2_1 _8199_ (.Y(_3170_),
    .A(net12),
    .B(_3169_));
 sg13g2_xnor2_1 _8200_ (.Y(_3171_),
    .A(_2184_),
    .B(_2185_));
 sg13g2_nand3_1 _8201_ (.B(_3158_),
    .C(_3171_),
    .A(_3156_),
    .Y(_3172_));
 sg13g2_nand2_1 _8202_ (.Y(_3173_),
    .A(_3170_),
    .B(_3172_));
 sg13g2_nor2_1 _8203_ (.A(_0030_),
    .B(_3173_),
    .Y(_3174_));
 sg13g2_xnor2_1 _8204_ (.Y(_3175_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ),
    .B(_3173_));
 sg13g2_nand2_1 _8205_ (.Y(_3176_),
    .A(_3175_),
    .B(_2184_));
 sg13g2_nand2b_1 _8206_ (.Y(_3177_),
    .B(_3176_),
    .A_N(_3174_));
 sg13g2_xnor2_1 _8207_ (.Y(_3178_),
    .A(_3168_),
    .B(_3177_));
 sg13g2_inv_1 _8208_ (.Y(_3179_),
    .A(_3178_));
 sg13g2_nor2_1 _8209_ (.A(net43),
    .B(_3179_),
    .Y(_3180_));
 sg13g2_nor2_1 _8210_ (.A(_4274_),
    .B(_0779_),
    .Y(_3181_));
 sg13g2_buf_2 _8211_ (.A(_3181_),
    .X(_3182_));
 sg13g2_inv_1 _8212_ (.Y(_3183_),
    .A(_3182_));
 sg13g2_inv_1 _8213_ (.Y(_3184_),
    .A(_3111_));
 sg13g2_nor2_1 _8214_ (.A(_4230_),
    .B(_3184_),
    .Y(_3185_));
 sg13g2_nor3_1 _8215_ (.A(_3183_),
    .B(_3112_),
    .C(_3185_),
    .Y(_3186_));
 sg13g2_inv_1 _8216_ (.Y(_3187_),
    .A(_3186_));
 sg13g2_a21o_1 _8217_ (.A2(_3107_),
    .A1(_3106_),
    .B1(_3112_),
    .X(_3188_));
 sg13g2_and2_1 _8218_ (.A(_3188_),
    .B(_3113_),
    .X(_3189_));
 sg13g2_nand3_1 _8219_ (.B(_3110_),
    .C(_0599_),
    .A(_3109_),
    .Y(_3190_));
 sg13g2_xnor2_1 _8220_ (.Y(_3191_),
    .A(_2433_),
    .B(_2764_));
 sg13g2_xnor2_1 _8221_ (.Y(_3192_),
    .A(_2735_),
    .B(_3191_));
 sg13g2_nand2_1 _8222_ (.Y(_3193_),
    .A(_3192_),
    .B(_0600_));
 sg13g2_nand2_1 _8223_ (.Y(_3194_),
    .A(_3190_),
    .B(_3193_));
 sg13g2_nand2_1 _8224_ (.Y(_3195_),
    .A(_3194_),
    .B(_4229_));
 sg13g2_nand3_1 _8225_ (.B(_2177_),
    .C(_3193_),
    .A(_3190_),
    .Y(_3196_));
 sg13g2_nand2_1 _8226_ (.Y(_3197_),
    .A(_3192_),
    .B(_0599_));
 sg13g2_a21oi_1 _8227_ (.A1(_2732_),
    .A2(_2733_),
    .Y(_3198_),
    .B1(_2415_));
 sg13g2_nand3b_1 _8228_ (.B(_0600_),
    .C(_2735_),
    .Y(_3199_),
    .A_N(_3198_));
 sg13g2_a21oi_1 _8229_ (.A1(_3197_),
    .A2(_3199_),
    .Y(_3200_),
    .B1(_0300_));
 sg13g2_nand3_1 _8230_ (.B(_3196_),
    .C(_3200_),
    .A(_3195_),
    .Y(_3201_));
 sg13g2_nand2_1 _8231_ (.Y(_3202_),
    .A(_3194_),
    .B(_3114_));
 sg13g2_nand2_1 _8232_ (.Y(_3203_),
    .A(_3201_),
    .B(_3202_));
 sg13g2_nand2_1 _8233_ (.Y(_3204_),
    .A(_3105_),
    .B(net51));
 sg13g2_nand2_1 _8234_ (.Y(_3205_),
    .A(_3184_),
    .B(net44));
 sg13g2_nand2_1 _8235_ (.Y(_3206_),
    .A(_3204_),
    .B(_3205_));
 sg13g2_nand2_1 _8236_ (.Y(_3207_),
    .A(_3206_),
    .B(_2178_));
 sg13g2_nand3_1 _8237_ (.B(_4226_),
    .C(_3205_),
    .A(_3204_),
    .Y(_3208_));
 sg13g2_nand2_1 _8238_ (.Y(_3209_),
    .A(_3207_),
    .B(_3208_));
 sg13g2_nand2_1 _8239_ (.Y(_3210_),
    .A(_3203_),
    .B(_3209_));
 sg13g2_nand2_1 _8240_ (.Y(_3211_),
    .A(_3206_),
    .B(_3125_));
 sg13g2_nand2_1 _8241_ (.Y(_3212_),
    .A(_3210_),
    .B(_3211_));
 sg13g2_nand2_1 _8242_ (.Y(_3213_),
    .A(_3121_),
    .B(net51));
 sg13g2_nand2_1 _8243_ (.Y(_3214_),
    .A(_3105_),
    .B(net44));
 sg13g2_nand2_1 _8244_ (.Y(_3215_),
    .A(_3213_),
    .B(_3214_));
 sg13g2_xnor2_1 _8245_ (.Y(_3216_),
    .A(_2179_),
    .B(_3215_));
 sg13g2_nand2_1 _8246_ (.Y(_3217_),
    .A(_3212_),
    .B(_3216_));
 sg13g2_nand2_1 _8247_ (.Y(_3218_),
    .A(_3130_),
    .B(net51));
 sg13g2_nand2_1 _8248_ (.Y(_3219_),
    .A(_3119_),
    .B(net44));
 sg13g2_nand3_1 _8249_ (.B(_3137_),
    .C(_3219_),
    .A(_3218_),
    .Y(_3220_));
 sg13g2_nand2_1 _8250_ (.Y(_3221_),
    .A(_3215_),
    .B(_3134_));
 sg13g2_nand3_1 _8251_ (.B(_3220_),
    .C(_3221_),
    .A(_3217_),
    .Y(_3222_));
 sg13g2_a21o_1 _8252_ (.A2(_3219_),
    .A1(_3218_),
    .B1(_3137_),
    .X(_3223_));
 sg13g2_nand2_1 _8253_ (.Y(_3224_),
    .A(_3222_),
    .B(_3223_));
 sg13g2_nand3_1 _8254_ (.B(_3146_),
    .C(net51),
    .A(_3145_),
    .Y(_3225_));
 sg13g2_nand2_1 _8255_ (.Y(_3226_),
    .A(_3133_),
    .B(net44));
 sg13g2_nand2_1 _8256_ (.Y(_3227_),
    .A(_3225_),
    .B(_3226_));
 sg13g2_nand2_1 _8257_ (.Y(_3228_),
    .A(_3227_),
    .B(_3096_));
 sg13g2_nand3_1 _8258_ (.B(_3226_),
    .C(_4247_),
    .A(_3225_),
    .Y(_3229_));
 sg13g2_nand2_1 _8259_ (.Y(_3230_),
    .A(_3228_),
    .B(_3229_));
 sg13g2_inv_1 _8260_ (.Y(_3231_),
    .A(_3230_));
 sg13g2_nand2_1 _8261_ (.Y(_3232_),
    .A(_3224_),
    .B(_3231_));
 sg13g2_nand3_1 _8262_ (.B(_3230_),
    .C(_3223_),
    .A(_3222_),
    .Y(_3233_));
 sg13g2_buf_2 _8263_ (.A(_3233_),
    .X(_3234_));
 sg13g2_nand2_1 _8264_ (.Y(_3235_),
    .A(_3232_),
    .B(_3234_));
 sg13g2_buf_8 _8265_ (.A(_3235_),
    .X(_3236_));
 sg13g2_nand2_1 _8266_ (.Y(_3237_),
    .A(_3236_),
    .B(_2181_));
 sg13g2_xnor2_1 _8267_ (.Y(_3238_),
    .A(_2185_),
    .B(_2180_));
 sg13g2_nand3_1 _8268_ (.B(_3234_),
    .C(_3238_),
    .A(_3232_),
    .Y(_3239_));
 sg13g2_nand2_1 _8269_ (.Y(_3240_),
    .A(_3237_),
    .B(_3239_));
 sg13g2_inv_1 _8270_ (.Y(_3241_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ));
 sg13g2_nand2_1 _8271_ (.Y(_3242_),
    .A(_3240_),
    .B(_3241_));
 sg13g2_nand3_1 _8272_ (.B(_3239_),
    .C(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ),
    .A(_3237_),
    .Y(_3243_));
 sg13g2_nand2_2 _8273_ (.Y(_3244_),
    .A(_3242_),
    .B(_3243_));
 sg13g2_nor2_2 _8274_ (.A(_3183_),
    .B(_3244_),
    .Y(_3245_));
 sg13g2_xnor2_1 _8275_ (.Y(_3246_),
    .A(_3189_),
    .B(_3245_));
 sg13g2_nor2_1 _8276_ (.A(_3187_),
    .B(_3246_),
    .Y(_3247_));
 sg13g2_nand2_2 _8277_ (.Y(_3248_),
    .A(_3178_),
    .B(_3182_));
 sg13g2_xnor2_1 _8278_ (.Y(_3249_),
    .A(_3123_),
    .B(_3116_));
 sg13g2_a21oi_1 _8279_ (.A1(_3248_),
    .A2(_0789_),
    .Y(_3250_),
    .B1(_3249_));
 sg13g2_nand3_1 _8280_ (.B(_0789_),
    .C(_3249_),
    .A(_3248_),
    .Y(_3251_));
 sg13g2_nand2b_1 _8281_ (.Y(_3252_),
    .B(_3251_),
    .A_N(_3250_));
 sg13g2_and2_1 _8282_ (.A(_3245_),
    .B(_3189_),
    .X(_3253_));
 sg13g2_buf_1 _8283_ (.A(_3253_),
    .X(_3254_));
 sg13g2_nand2b_1 _8284_ (.Y(_3255_),
    .B(_3254_),
    .A_N(_3252_));
 sg13g2_nand2b_1 _8285_ (.Y(_3256_),
    .B(_3252_),
    .A_N(_3254_));
 sg13g2_nand2_1 _8286_ (.Y(_3257_),
    .A(_3255_),
    .B(_3256_));
 sg13g2_nand2b_1 _8287_ (.Y(_3258_),
    .B(_3257_),
    .A_N(_3247_));
 sg13g2_nand3_1 _8288_ (.B(_3247_),
    .C(_3256_),
    .A(_3255_),
    .Y(_3259_));
 sg13g2_nand2_1 _8289_ (.Y(_3260_),
    .A(_3258_),
    .B(_3259_));
 sg13g2_xnor2_1 _8290_ (.Y(_3261_),
    .A(_3180_),
    .B(_3260_));
 sg13g2_nor2_1 _8291_ (.A(net54),
    .B(_3261_),
    .Y(_3262_));
 sg13g2_xnor2_1 _8292_ (.Y(_3263_),
    .A(_3241_),
    .B(_3173_));
 sg13g2_inv_1 _8293_ (.Y(_3264_),
    .A(_2184_));
 sg13g2_nand2_1 _8294_ (.Y(_3265_),
    .A(_3263_),
    .B(_3264_));
 sg13g2_buf_1 _8295_ (.A(_0791_),
    .X(_3266_));
 sg13g2_nand3_1 _8296_ (.B(_3265_),
    .C(net46),
    .A(_3176_),
    .Y(_3267_));
 sg13g2_xnor2_1 _8297_ (.Y(_3268_),
    .A(_3186_),
    .B(_3246_));
 sg13g2_xnor2_1 _8298_ (.Y(_3269_),
    .A(_3267_),
    .B(_3268_));
 sg13g2_nor2_2 _8299_ (.A(_3096_),
    .B(net43),
    .Y(_3270_));
 sg13g2_inv_2 _8300_ (.Y(_3271_),
    .A(_3270_));
 sg13g2_nand2_1 _8301_ (.Y(_3272_),
    .A(net12),
    .B(_3271_));
 sg13g2_nand2_1 _8302_ (.Y(_3273_),
    .A(_0791_),
    .B(_4220_));
 sg13g2_buf_8 _8303_ (.A(_3273_),
    .X(_3274_));
 sg13g2_nand2_1 _8304_ (.Y(_3275_),
    .A(_2188_),
    .B(_3274_));
 sg13g2_xnor2_1 _8305_ (.Y(_3276_),
    .A(_3270_),
    .B(_3275_));
 sg13g2_nand3_1 _8306_ (.B(_3158_),
    .C(_3276_),
    .A(_3156_),
    .Y(_3277_));
 sg13g2_nand2_1 _8307_ (.Y(_3278_),
    .A(_3272_),
    .B(_3277_));
 sg13g2_xnor2_1 _8308_ (.Y(_3279_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[4] ),
    .B(_3278_));
 sg13g2_nor2_1 _8309_ (.A(_3168_),
    .B(_3263_),
    .Y(_3280_));
 sg13g2_nand2_1 _8310_ (.Y(_3281_),
    .A(_3280_),
    .B(_2184_));
 sg13g2_inv_1 _8311_ (.Y(_3282_),
    .A(_3163_));
 sg13g2_a21oi_1 _8312_ (.A1(_3174_),
    .A2(_3167_),
    .Y(_3283_),
    .B1(_3282_));
 sg13g2_nand2_1 _8313_ (.Y(_3284_),
    .A(_3281_),
    .B(_3283_));
 sg13g2_nand2_1 _8314_ (.Y(_3285_),
    .A(net12),
    .B(_3274_));
 sg13g2_xnor2_1 _8315_ (.Y(_3286_),
    .A(_3274_),
    .B(_2188_));
 sg13g2_nand3_1 _8316_ (.B(_3158_),
    .C(_3286_),
    .A(_3156_),
    .Y(_3287_));
 sg13g2_nand2_1 _8317_ (.Y(_3288_),
    .A(_3285_),
    .B(_3287_));
 sg13g2_inv_1 _8318_ (.Y(_3289_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[3] ));
 sg13g2_nand2_1 _8319_ (.Y(_3290_),
    .A(_3288_),
    .B(_3289_));
 sg13g2_nand3_1 _8320_ (.B(_3287_),
    .C(\main.demo._d___pip_58_1_3___stage___block_3_a[3] ),
    .A(_3285_),
    .Y(_3291_));
 sg13g2_nand2_2 _8321_ (.Y(_3292_),
    .A(_3290_),
    .B(_3291_));
 sg13g2_inv_2 _8322_ (.Y(_3293_),
    .A(_3292_));
 sg13g2_nand2_1 _8323_ (.Y(_3294_),
    .A(_3284_),
    .B(_3293_));
 sg13g2_nor2_1 _8324_ (.A(_0028_),
    .B(_3288_),
    .Y(_3295_));
 sg13g2_inv_1 _8325_ (.Y(_3296_),
    .A(_3295_));
 sg13g2_nand2_1 _8326_ (.Y(_3297_),
    .A(_3294_),
    .B(_3296_));
 sg13g2_xnor2_1 _8327_ (.Y(_3298_),
    .A(_3279_),
    .B(_3297_));
 sg13g2_nor2_1 _8328_ (.A(net43),
    .B(_3298_),
    .Y(_3299_));
 sg13g2_xnor2_1 _8329_ (.Y(_3300_),
    .A(_3131_),
    .B(_3127_));
 sg13g2_nand3_1 _8330_ (.B(_3283_),
    .C(_3292_),
    .A(_3281_),
    .Y(_3301_));
 sg13g2_nand3_1 _8331_ (.B(_3301_),
    .C(_3182_),
    .A(_3294_),
    .Y(_3302_));
 sg13g2_o21ai_1 _8332_ (.B1(_3302_),
    .Y(_3303_),
    .A1(_0789_),
    .A2(_3263_));
 sg13g2_xor2_1 _8333_ (.B(_3303_),
    .A(_3300_),
    .X(_3304_));
 sg13g2_inv_1 _8334_ (.Y(_3305_),
    .A(_3304_));
 sg13g2_nand2_1 _8335_ (.Y(_3306_),
    .A(_3305_),
    .B(_3250_));
 sg13g2_nand2b_1 _8336_ (.Y(_3307_),
    .B(_3303_),
    .A_N(_3300_));
 sg13g2_inv_1 _8337_ (.Y(_3308_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[4] ));
 sg13g2_xnor2_1 _8338_ (.Y(_3309_),
    .A(_3308_),
    .B(_3278_));
 sg13g2_xnor2_1 _8339_ (.Y(_3310_),
    .A(_3309_),
    .B(_3297_));
 sg13g2_nand2_1 _8340_ (.Y(_3311_),
    .A(_3310_),
    .B(_3182_));
 sg13g2_a21oi_1 _8341_ (.A1(_3178_),
    .A2(_4274_),
    .Y(_3312_),
    .B1(_4276_));
 sg13g2_nand2_1 _8342_ (.Y(_3313_),
    .A(_3311_),
    .B(_3312_));
 sg13g2_nand2b_1 _8343_ (.Y(_3314_),
    .B(_3313_),
    .A_N(_3307_));
 sg13g2_nor2_1 _8344_ (.A(_3183_),
    .B(_3298_),
    .Y(_3315_));
 sg13g2_nor2b_1 _8345_ (.A(_3315_),
    .B_N(_3312_),
    .Y(_3316_));
 sg13g2_nand2_1 _8346_ (.Y(_3317_),
    .A(_3316_),
    .B(_3307_));
 sg13g2_nand2_1 _8347_ (.Y(_3318_),
    .A(_3314_),
    .B(_3317_));
 sg13g2_xor2_1 _8348_ (.B(_3136_),
    .A(_3148_),
    .X(_3319_));
 sg13g2_nand2_1 _8349_ (.Y(_3320_),
    .A(_3318_),
    .B(_3319_));
 sg13g2_inv_1 _8350_ (.Y(_3321_),
    .A(_3319_));
 sg13g2_nand3_1 _8351_ (.B(_3317_),
    .C(_3321_),
    .A(_3314_),
    .Y(_3322_));
 sg13g2_nand2_1 _8352_ (.Y(_3323_),
    .A(_3320_),
    .B(_3322_));
 sg13g2_xnor2_1 _8353_ (.Y(_3324_),
    .A(_3306_),
    .B(_3323_));
 sg13g2_inv_2 _8354_ (.Y(_3325_),
    .A(_3259_));
 sg13g2_a21oi_1 _8355_ (.A1(_3251_),
    .A2(_3254_),
    .Y(_3326_),
    .B1(_3250_));
 sg13g2_xor2_1 _8356_ (.B(_3304_),
    .A(_3326_),
    .X(_3327_));
 sg13g2_nor2_1 _8357_ (.A(_3304_),
    .B(_3255_),
    .Y(_3328_));
 sg13g2_a21oi_2 _8358_ (.B1(_3328_),
    .Y(_3329_),
    .A2(_3327_),
    .A1(_3325_));
 sg13g2_inv_4 _8359_ (.A(_3329_),
    .Y(_3330_));
 sg13g2_nand2_1 _8360_ (.Y(_3331_),
    .A(_3324_),
    .B(_3330_));
 sg13g2_nand2b_1 _8361_ (.Y(_3332_),
    .B(_3323_),
    .A_N(_3306_));
 sg13g2_nand3_1 _8362_ (.B(_3322_),
    .C(_3306_),
    .A(_3320_),
    .Y(_3333_));
 sg13g2_nand2_1 _8363_ (.Y(_3334_),
    .A(_3332_),
    .B(_3333_));
 sg13g2_nand2_1 _8364_ (.Y(_3335_),
    .A(_3334_),
    .B(_3329_));
 sg13g2_nand3b_1 _8365_ (.B(_3331_),
    .C(_3335_),
    .Y(_3336_),
    .A_N(_3299_));
 sg13g2_nand2_1 _8366_ (.Y(_3337_),
    .A(_3331_),
    .B(_3335_));
 sg13g2_nand2_1 _8367_ (.Y(_3338_),
    .A(_3337_),
    .B(_3299_));
 sg13g2_nand2_1 _8368_ (.Y(_3339_),
    .A(_3336_),
    .B(_3338_));
 sg13g2_inv_1 _8369_ (.Y(_3340_),
    .A(_3180_));
 sg13g2_xnor2_1 _8370_ (.Y(_3341_),
    .A(_3340_),
    .B(_3260_));
 sg13g2_nand3_1 _8371_ (.B(_0316_),
    .C(_0312_),
    .A(_3341_),
    .Y(_3342_));
 sg13g2_nand2_1 _8372_ (.Y(_3343_),
    .A(_3294_),
    .B(_3301_));
 sg13g2_nor2_1 _8373_ (.A(net43),
    .B(_3343_),
    .Y(_3344_));
 sg13g2_xor2_1 _8374_ (.B(_3259_),
    .A(_3327_),
    .X(_3345_));
 sg13g2_xnor2_1 _8375_ (.Y(_3346_),
    .A(_3344_),
    .B(_3345_));
 sg13g2_nand2_1 _8376_ (.Y(_3347_),
    .A(_3342_),
    .B(_3346_));
 sg13g2_inv_1 _8377_ (.Y(_3348_),
    .A(_0316_));
 sg13g2_o21ai_1 _8378_ (.B1(_3348_),
    .Y(_3349_),
    .A1(_0314_),
    .A2(_3261_));
 sg13g2_nand2_1 _8379_ (.Y(_3350_),
    .A(_3347_),
    .B(_3349_));
 sg13g2_inv_1 _8380_ (.Y(_3351_),
    .A(_0037_));
 sg13g2_nand3_1 _8381_ (.B(_3350_),
    .C(_3351_),
    .A(_3339_),
    .Y(_3352_));
 sg13g2_nand2_1 _8382_ (.Y(_3353_),
    .A(_3352_),
    .B(\main.demo._q_th[5] ));
 sg13g2_nand2_1 _8383_ (.Y(_3354_),
    .A(_3279_),
    .B(_3295_));
 sg13g2_nor2_1 _8384_ (.A(_0027_),
    .B(_3278_),
    .Y(_3355_));
 sg13g2_inv_1 _8385_ (.Y(_3356_),
    .A(_3355_));
 sg13g2_nand2_1 _8386_ (.Y(_3357_),
    .A(_3354_),
    .B(_3356_));
 sg13g2_nand2_1 _8387_ (.Y(_3358_),
    .A(_3293_),
    .B(_3279_));
 sg13g2_nor2_1 _8388_ (.A(_3283_),
    .B(_3358_),
    .Y(_3359_));
 sg13g2_nor2_1 _8389_ (.A(_3357_),
    .B(_3359_),
    .Y(_3360_));
 sg13g2_nor2_1 _8390_ (.A(_3292_),
    .B(_3309_),
    .Y(_3361_));
 sg13g2_nand3_1 _8391_ (.B(_3361_),
    .C(_2184_),
    .A(_3280_),
    .Y(_3362_));
 sg13g2_nand2_1 _8392_ (.Y(_3363_),
    .A(_3360_),
    .B(_3362_));
 sg13g2_inv_1 _8393_ (.Y(_3364_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[5] ));
 sg13g2_nor2_2 _8394_ (.A(_0298_),
    .B(net43),
    .Y(_3365_));
 sg13g2_inv_1 _8395_ (.Y(_3366_),
    .A(_3274_));
 sg13g2_nor2_1 _8396_ (.A(_3366_),
    .B(_2187_),
    .Y(_3367_));
 sg13g2_inv_1 _8397_ (.Y(_3368_),
    .A(_3367_));
 sg13g2_nor2_1 _8398_ (.A(_3270_),
    .B(_3368_),
    .Y(_3369_));
 sg13g2_nand2_1 _8399_ (.Y(_3370_),
    .A(_3369_),
    .B(_3264_));
 sg13g2_xnor2_1 _8400_ (.Y(_3371_),
    .A(_3365_),
    .B(_3370_));
 sg13g2_nand2_1 _8401_ (.Y(_3372_),
    .A(_3153_),
    .B(_3371_));
 sg13g2_inv_1 _8402_ (.Y(_3373_),
    .A(_3365_));
 sg13g2_nand2_1 _8403_ (.Y(_3374_),
    .A(net12),
    .B(_3373_));
 sg13g2_nand2_1 _8404_ (.Y(_3375_),
    .A(_3372_),
    .B(_3374_));
 sg13g2_xnor2_1 _8405_ (.Y(_3376_),
    .A(_3364_),
    .B(_3375_));
 sg13g2_inv_1 _8406_ (.Y(_3377_),
    .A(_3376_));
 sg13g2_nand2_1 _8407_ (.Y(_3378_),
    .A(_3363_),
    .B(_3377_));
 sg13g2_nand3_1 _8408_ (.B(_3362_),
    .C(_3376_),
    .A(_3360_),
    .Y(_3379_));
 sg13g2_and3_1 _8409_ (.X(_3380_),
    .A(_3378_),
    .B(_3379_),
    .C(net46));
 sg13g2_nand3_1 _8410_ (.B(_3379_),
    .C(_3182_),
    .A(_3378_),
    .Y(_3381_));
 sg13g2_inv_1 _8411_ (.Y(_3382_),
    .A(_3343_));
 sg13g2_nand2_1 _8412_ (.Y(_3383_),
    .A(_3382_),
    .B(_0802_));
 sg13g2_nor2_1 _8413_ (.A(_4277_),
    .B(_3244_),
    .Y(_3384_));
 sg13g2_inv_1 _8414_ (.Y(_3385_),
    .A(_3384_));
 sg13g2_nand3_1 _8415_ (.B(_3383_),
    .C(_3385_),
    .A(_3381_),
    .Y(_3386_));
 sg13g2_xnor2_1 _8416_ (.Y(_3387_),
    .A(_3160_),
    .B(_3386_));
 sg13g2_inv_1 _8417_ (.Y(_3388_),
    .A(_3314_));
 sg13g2_a21oi_1 _8418_ (.A1(_3317_),
    .A2(_3319_),
    .Y(_3389_),
    .B1(_3388_));
 sg13g2_xnor2_1 _8419_ (.Y(_3390_),
    .A(_3387_),
    .B(_3389_));
 sg13g2_inv_2 _8420_ (.Y(_3391_),
    .A(_3332_));
 sg13g2_a21oi_1 _8421_ (.A1(_3330_),
    .A2(_3333_),
    .Y(_3392_),
    .B1(_3391_));
 sg13g2_xnor2_1 _8422_ (.Y(_3393_),
    .A(_3390_),
    .B(_3392_));
 sg13g2_xor2_1 _8423_ (.B(_3393_),
    .A(_3380_),
    .X(_3394_));
 sg13g2_nand2_1 _8424_ (.Y(_3395_),
    .A(_3353_),
    .B(_3394_));
 sg13g2_nand3_1 _8425_ (.B(_3350_),
    .C(_0037_),
    .A(_3339_),
    .Y(_3396_));
 sg13g2_inv_2 _8426_ (.Y(_3397_),
    .A(_3394_));
 sg13g2_nand2b_1 _8427_ (.Y(_3398_),
    .B(_3397_),
    .A_N(_3396_));
 sg13g2_nand2_1 _8428_ (.Y(_3399_),
    .A(_3395_),
    .B(_3398_));
 sg13g2_nand2_2 _8429_ (.Y(_3400_),
    .A(_0791_),
    .B(_4217_));
 sg13g2_nor2_1 _8430_ (.A(_3365_),
    .B(_3370_),
    .Y(_3401_));
 sg13g2_nor2_1 _8431_ (.A(_3401_),
    .B(net12),
    .Y(_3402_));
 sg13g2_xnor2_1 _8432_ (.Y(_3403_),
    .A(_3400_),
    .B(_3402_));
 sg13g2_xnor2_1 _8433_ (.Y(_3404_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[6] ),
    .B(_3403_));
 sg13g2_o21ai_1 _8434_ (.B1(_3296_),
    .Y(_3405_),
    .A1(_3163_),
    .A2(_3292_));
 sg13g2_nor2_1 _8435_ (.A(_3309_),
    .B(_3376_),
    .Y(_3406_));
 sg13g2_nor2_1 _8436_ (.A(_0032_),
    .B(_3375_),
    .Y(_3407_));
 sg13g2_inv_1 _8437_ (.Y(_3408_),
    .A(_3407_));
 sg13g2_o21ai_1 _8438_ (.B1(_3408_),
    .Y(_3409_),
    .A1(_3356_),
    .A2(_3376_));
 sg13g2_a21oi_1 _8439_ (.A1(_3405_),
    .A2(_3406_),
    .Y(_3410_),
    .B1(_3409_));
 sg13g2_nor2_1 _8440_ (.A(_3292_),
    .B(_3168_),
    .Y(_3411_));
 sg13g2_nand3_1 _8441_ (.B(_3411_),
    .C(_3406_),
    .A(_3177_),
    .Y(_3412_));
 sg13g2_nand2_1 _8442_ (.Y(_3413_),
    .A(_3410_),
    .B(_3412_));
 sg13g2_nand2b_1 _8443_ (.Y(_3414_),
    .B(_3413_),
    .A_N(_3404_));
 sg13g2_nand3_1 _8444_ (.B(_3404_),
    .C(_3412_),
    .A(_3410_),
    .Y(_3415_));
 sg13g2_nand3_1 _8445_ (.B(_3415_),
    .C(net46),
    .A(_3414_),
    .Y(_3416_));
 sg13g2_nand2_1 _8446_ (.Y(_3417_),
    .A(_3386_),
    .B(_3153_));
 sg13g2_nor4_1 _8447_ (.A(_2325_),
    .B(_2366_),
    .C(_2350_),
    .D(_2344_),
    .Y(_3418_));
 sg13g2_nor2b_1 _8448_ (.A(_2955_),
    .B_N(_2967_),
    .Y(_3419_));
 sg13g2_a21oi_1 _8449_ (.A1(_2968_),
    .A2(_2950_),
    .Y(_3420_),
    .B1(_3419_));
 sg13g2_nor2_1 _8450_ (.A(net63),
    .B(_2882_),
    .Y(_3421_));
 sg13g2_xnor2_1 _8451_ (.Y(_3422_),
    .A(_3421_),
    .B(_2959_));
 sg13g2_xor2_1 _8452_ (.B(_3422_),
    .A(_2961_),
    .X(_3423_));
 sg13g2_xor2_1 _8453_ (.B(_3423_),
    .A(_2956_),
    .X(_3424_));
 sg13g2_a21oi_1 _8454_ (.A1(_2965_),
    .A2(_2956_),
    .Y(_3425_),
    .B1(_2964_));
 sg13g2_nor2_1 _8455_ (.A(_3424_),
    .B(_3425_),
    .Y(_3426_));
 sg13g2_nand2_1 _8456_ (.Y(_3427_),
    .A(_3425_),
    .B(_3424_));
 sg13g2_nand2b_1 _8457_ (.Y(_3428_),
    .B(_3427_),
    .A_N(_3426_));
 sg13g2_xnor2_1 _8458_ (.Y(_3429_),
    .A(_2950_),
    .B(_3428_));
 sg13g2_nand2b_1 _8459_ (.Y(_3430_),
    .B(_3429_),
    .A_N(_3420_));
 sg13g2_nand2b_1 _8460_ (.Y(_3431_),
    .B(_3420_),
    .A_N(_3429_));
 sg13g2_nand2_1 _8461_ (.Y(_3432_),
    .A(_3430_),
    .B(_3431_));
 sg13g2_nor2b_1 _8462_ (.A(_2984_),
    .B_N(_3074_),
    .Y(_3433_));
 sg13g2_nand2_1 _8463_ (.Y(_3434_),
    .A(_2928_),
    .B(_2913_));
 sg13g2_a22oi_1 _8464_ (.Y(_3435_),
    .B1(_3433_),
    .B2(_3434_),
    .A2(_2969_),
    .A1(_2983_));
 sg13g2_xor2_1 _8465_ (.B(_3435_),
    .A(_3432_),
    .X(_3436_));
 sg13g2_nor2_1 _8466_ (.A(_3418_),
    .B(_3436_),
    .Y(_3437_));
 sg13g2_nand2_1 _8467_ (.Y(_3438_),
    .A(_3436_),
    .B(_3418_));
 sg13g2_nand2b_1 _8468_ (.Y(_3439_),
    .B(_3438_),
    .A_N(_3437_));
 sg13g2_nand3_1 _8469_ (.B(_3085_),
    .C(_3078_),
    .A(_3090_),
    .Y(_3440_));
 sg13g2_nand2_1 _8470_ (.Y(_3441_),
    .A(_3440_),
    .B(_3080_));
 sg13g2_xor2_1 _8471_ (.B(_3441_),
    .A(_3439_),
    .X(_3442_));
 sg13g2_xnor2_1 _8472_ (.Y(_3443_),
    .A(_0298_),
    .B(_3442_));
 sg13g2_nand2_1 _8473_ (.Y(_3444_),
    .A(_3087_),
    .B(_3092_));
 sg13g2_o21ai_1 _8474_ (.B1(_3156_),
    .Y(_3445_),
    .A1(_0035_),
    .A2(_3444_));
 sg13g2_xnor2_1 _8475_ (.Y(_3446_),
    .A(_3443_),
    .B(_3445_));
 sg13g2_nand2_1 _8476_ (.Y(_3447_),
    .A(_3236_),
    .B(_3274_));
 sg13g2_xnor2_1 _8477_ (.Y(_3448_),
    .A(_3274_),
    .B(_2186_));
 sg13g2_nand3_1 _8478_ (.B(_3234_),
    .C(_3448_),
    .A(_3232_),
    .Y(_3449_));
 sg13g2_nand2_1 _8479_ (.Y(_3450_),
    .A(_3447_),
    .B(_3449_));
 sg13g2_xnor2_1 _8480_ (.Y(_3451_),
    .A(_3166_),
    .B(_3450_));
 sg13g2_nand3_1 _8481_ (.B(_3243_),
    .C(_2185_),
    .A(_3242_),
    .Y(_3452_));
 sg13g2_or2_1 _8482_ (.X(_3453_),
    .B(_3240_),
    .A(_0030_));
 sg13g2_nand2_1 _8483_ (.Y(_3454_),
    .A(_3452_),
    .B(_3453_));
 sg13g2_xor2_1 _8484_ (.B(_3454_),
    .A(_3451_),
    .X(_3455_));
 sg13g2_nor2_1 _8485_ (.A(_4277_),
    .B(_3455_),
    .Y(_3456_));
 sg13g2_nand2_1 _8486_ (.Y(_3457_),
    .A(_3310_),
    .B(_0802_));
 sg13g2_nand3_1 _8487_ (.B(_3415_),
    .C(_3182_),
    .A(_3414_),
    .Y(_3458_));
 sg13g2_nand3b_1 _8488_ (.B(_3457_),
    .C(_3458_),
    .Y(_3459_),
    .A_N(_3456_));
 sg13g2_xnor2_1 _8489_ (.Y(_3460_),
    .A(_3446_),
    .B(_3459_));
 sg13g2_nor2_1 _8490_ (.A(_3417_),
    .B(_3460_),
    .Y(_3461_));
 sg13g2_nand2_1 _8491_ (.Y(_3462_),
    .A(_3460_),
    .B(_3417_));
 sg13g2_nand2b_1 _8492_ (.Y(_3463_),
    .B(_3462_),
    .A_N(_3461_));
 sg13g2_nand3_1 _8493_ (.B(_3390_),
    .C(_3330_),
    .A(_3324_),
    .Y(_3464_));
 sg13g2_nor2b_1 _8494_ (.A(_3389_),
    .B_N(_3387_),
    .Y(_3465_));
 sg13g2_a21oi_1 _8495_ (.A1(_3391_),
    .A2(_3390_),
    .Y(_3466_),
    .B1(_3465_));
 sg13g2_nand2_1 _8496_ (.Y(_3467_),
    .A(_3464_),
    .B(_3466_));
 sg13g2_nand2b_1 _8497_ (.Y(_3468_),
    .B(_3467_),
    .A_N(_3463_));
 sg13g2_nand3_1 _8498_ (.B(_3463_),
    .C(_3466_),
    .A(_3464_),
    .Y(_3469_));
 sg13g2_nand2_1 _8499_ (.Y(_3470_),
    .A(_3468_),
    .B(_3469_));
 sg13g2_inv_2 _8500_ (.Y(_3471_),
    .A(_3470_));
 sg13g2_nand2b_1 _8501_ (.Y(_3472_),
    .B(_3471_),
    .A_N(_3416_));
 sg13g2_nand2_1 _8502_ (.Y(_3473_),
    .A(_3470_),
    .B(_3416_));
 sg13g2_nand2_1 _8503_ (.Y(_3474_),
    .A(_3472_),
    .B(_3473_));
 sg13g2_nand2b_1 _8504_ (.Y(_3475_),
    .B(_3474_),
    .A_N(_0036_));
 sg13g2_nand3_1 _8505_ (.B(_0036_),
    .C(_3473_),
    .A(_3472_),
    .Y(_3476_));
 sg13g2_nand3_1 _8506_ (.B(_3475_),
    .C(_3476_),
    .A(_3399_),
    .Y(_3477_));
 sg13g2_inv_1 _8507_ (.Y(_3478_),
    .A(_0031_));
 sg13g2_nand2_1 _8508_ (.Y(_3479_),
    .A(_3403_),
    .B(_3478_));
 sg13g2_nand2_1 _8509_ (.Y(_3480_),
    .A(_3414_),
    .B(_3479_));
 sg13g2_nand2_1 _8510_ (.Y(_3481_),
    .A(net46),
    .B(_4214_));
 sg13g2_xnor2_1 _8511_ (.Y(_3482_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[7] ),
    .B(_3481_));
 sg13g2_a21o_1 _8512_ (.A2(_3400_),
    .A1(_3401_),
    .B1(net12),
    .X(_3483_));
 sg13g2_xnor2_1 _8513_ (.Y(_3484_),
    .A(_3482_),
    .B(_3483_));
 sg13g2_nand2_1 _8514_ (.Y(_3485_),
    .A(_3480_),
    .B(_3484_));
 sg13g2_inv_1 _8515_ (.Y(_3486_),
    .A(_3484_));
 sg13g2_nand3_1 _8516_ (.B(_3479_),
    .C(_3486_),
    .A(_3414_),
    .Y(_3487_));
 sg13g2_nand3_1 _8517_ (.B(_3487_),
    .C(net46),
    .A(_3485_),
    .Y(_3488_));
 sg13g2_nand2_1 _8518_ (.Y(_3489_),
    .A(_3459_),
    .B(_3446_));
 sg13g2_a21oi_1 _8519_ (.A1(_3427_),
    .A2(_2950_),
    .Y(_3490_),
    .B1(_3426_));
 sg13g2_xor2_1 _8520_ (.B(_2458_),
    .A(_0033_),
    .X(_3491_));
 sg13g2_a22oi_1 _8521_ (.Y(_3492_),
    .B1(_2956_),
    .B2(_3423_),
    .A2(_2961_),
    .A1(_2882_));
 sg13g2_nand2_1 _8522_ (.Y(_3493_),
    .A(_2960_),
    .B(_3421_));
 sg13g2_o21ai_1 _8523_ (.B1(_3493_),
    .Y(_3494_),
    .A1(_2482_),
    .A2(_2882_));
 sg13g2_o21ai_1 _8524_ (.B1(_3494_),
    .Y(_3495_),
    .A1(_2482_),
    .A2(_3493_));
 sg13g2_xnor2_1 _8525_ (.Y(_3496_),
    .A(_2950_),
    .B(_3495_));
 sg13g2_xnor2_1 _8526_ (.Y(_3497_),
    .A(_3492_),
    .B(_3496_));
 sg13g2_xnor2_1 _8527_ (.Y(_3498_),
    .A(_3491_),
    .B(_3497_));
 sg13g2_xnor2_1 _8528_ (.Y(_3499_),
    .A(_3490_),
    .B(_3498_));
 sg13g2_nand2b_1 _8529_ (.Y(_3500_),
    .B(_2986_),
    .A_N(_3076_));
 sg13g2_nor2b_1 _8530_ (.A(_2984_),
    .B_N(_3430_),
    .Y(_3501_));
 sg13g2_inv_1 _8531_ (.Y(_3502_),
    .A(_3431_));
 sg13g2_a21oi_1 _8532_ (.A1(_3500_),
    .A2(_3501_),
    .Y(_3503_),
    .B1(_3502_));
 sg13g2_xor2_1 _8533_ (.B(_3503_),
    .A(_3499_),
    .X(_3504_));
 sg13g2_o21ai_1 _8534_ (.B1(_3438_),
    .Y(_3505_),
    .A1(_3437_),
    .A2(_3441_));
 sg13g2_xnor2_1 _8535_ (.Y(_3506_),
    .A(_3504_),
    .B(_3505_));
 sg13g2_inv_1 _8536_ (.Y(_3507_),
    .A(_0034_));
 sg13g2_inv_1 _8537_ (.Y(_3508_),
    .A(_3442_));
 sg13g2_inv_1 _8538_ (.Y(_3509_),
    .A(_3443_));
 sg13g2_a22oi_1 _8539_ (.Y(_3510_),
    .B1(_3509_),
    .B2(_3445_),
    .A2(_3508_),
    .A1(_3507_));
 sg13g2_xnor2_1 _8540_ (.Y(_3511_),
    .A(_3506_),
    .B(_3510_));
 sg13g2_nand3_1 _8541_ (.B(_3487_),
    .C(_3182_),
    .A(_3485_),
    .Y(_3512_));
 sg13g2_nand2_1 _8542_ (.Y(_3513_),
    .A(_3382_),
    .B(_4276_));
 sg13g2_nand3_1 _8543_ (.B(_3379_),
    .C(_0802_),
    .A(_3378_),
    .Y(_3514_));
 sg13g2_nand3_1 _8544_ (.B(_3513_),
    .C(_3514_),
    .A(_3512_),
    .Y(_3515_));
 sg13g2_xnor2_1 _8545_ (.Y(_3516_),
    .A(_3511_),
    .B(_3515_));
 sg13g2_xnor2_1 _8546_ (.Y(_3517_),
    .A(_3489_),
    .B(_3516_));
 sg13g2_a21oi_1 _8547_ (.A1(_3333_),
    .A2(_3328_),
    .Y(_3518_),
    .B1(_3391_));
 sg13g2_nor2b_1 _8548_ (.A(_3463_),
    .B_N(_3390_),
    .Y(_3519_));
 sg13g2_nor2b_1 _8549_ (.A(_3518_),
    .B_N(_3519_),
    .Y(_3520_));
 sg13g2_a21oi_1 _8550_ (.A1(_3465_),
    .A2(_3462_),
    .Y(_3521_),
    .B1(_3461_));
 sg13g2_nor2b_1 _8551_ (.A(_3520_),
    .B_N(_3521_),
    .Y(_3522_));
 sg13g2_nand4_1 _8552_ (.B(_3325_),
    .C(_3324_),
    .A(_3519_),
    .Y(_3523_),
    .D(_3327_));
 sg13g2_nand2_1 _8553_ (.Y(_3524_),
    .A(_3522_),
    .B(_3523_));
 sg13g2_nand2b_1 _8554_ (.Y(_3525_),
    .B(_3524_),
    .A_N(_3517_));
 sg13g2_nand3_1 _8555_ (.B(_3523_),
    .C(_3517_),
    .A(_3522_),
    .Y(_3526_));
 sg13g2_nand2_1 _8556_ (.Y(_3527_),
    .A(_3525_),
    .B(_3526_));
 sg13g2_nand2b_1 _8557_ (.Y(_3528_),
    .B(_3527_),
    .A_N(_3488_));
 sg13g2_nand3_1 _8558_ (.B(_3526_),
    .C(_3488_),
    .A(_3525_),
    .Y(_3529_));
 sg13g2_nand2_1 _8559_ (.Y(_3530_),
    .A(_3528_),
    .B(_3529_));
 sg13g2_nor2_1 _8560_ (.A(_0326_),
    .B(_3474_),
    .Y(_3531_));
 sg13g2_a21oi_1 _8561_ (.A1(_3530_),
    .A2(_0331_),
    .Y(_3532_),
    .B1(_3531_));
 sg13g2_nand2_2 _8562_ (.Y(_3533_),
    .A(_3477_),
    .B(_3532_));
 sg13g2_nor2_1 _8563_ (.A(_0331_),
    .B(_3530_),
    .Y(_3534_));
 sg13g2_nor2_2 _8564_ (.A(net54),
    .B(_3534_),
    .Y(_3535_));
 sg13g2_nand2_1 _8565_ (.Y(_3536_),
    .A(_3533_),
    .B(_3535_));
 sg13g2_o21ai_1 _8566_ (.B1(_3536_),
    .Y(_3537_),
    .A1(net68),
    .A2(_3269_));
 sg13g2_or2_1 _8567_ (.X(_3538_),
    .B(_3537_),
    .A(_3262_));
 sg13g2_inv_2 _8568_ (.Y(_3539_),
    .A(_3236_));
 sg13g2_nor2_1 _8569_ (.A(_0789_),
    .B(_0601_),
    .Y(_3540_));
 sg13g2_inv_1 _8570_ (.Y(_3541_),
    .A(_3540_));
 sg13g2_nor2_1 _8571_ (.A(_3541_),
    .B(_3455_),
    .Y(_3542_));
 sg13g2_nor2_1 _8572_ (.A(_4276_),
    .B(_3542_),
    .Y(_3543_));
 sg13g2_nand2_1 _8573_ (.Y(_3544_),
    .A(_3381_),
    .B(_3543_));
 sg13g2_nand2_1 _8574_ (.Y(_3545_),
    .A(_3236_),
    .B(_3271_));
 sg13g2_xnor2_1 _8575_ (.Y(_3546_),
    .A(_3271_),
    .B(_3367_));
 sg13g2_nand3_1 _8576_ (.B(_3234_),
    .C(_3546_),
    .A(_3232_),
    .Y(_3547_));
 sg13g2_nand2_1 _8577_ (.Y(_3548_),
    .A(_3545_),
    .B(_3547_));
 sg13g2_xnor2_1 _8578_ (.Y(_3549_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[3] ),
    .B(_3548_));
 sg13g2_inv_1 _8579_ (.Y(_3550_),
    .A(_3549_));
 sg13g2_nor2_1 _8580_ (.A(_3451_),
    .B(_3550_),
    .Y(_3551_));
 sg13g2_nand2_1 _8581_ (.Y(_3552_),
    .A(_3454_),
    .B(_3551_));
 sg13g2_nor2_1 _8582_ (.A(_0029_),
    .B(_3450_),
    .Y(_3553_));
 sg13g2_nor2_1 _8583_ (.A(_0028_),
    .B(_3548_),
    .Y(_3554_));
 sg13g2_a21oi_1 _8584_ (.A1(_3549_),
    .A2(_3553_),
    .Y(_3555_),
    .B1(_3554_));
 sg13g2_nand2_1 _8585_ (.Y(_3556_),
    .A(_3552_),
    .B(_3555_));
 sg13g2_nor2_1 _8586_ (.A(_3369_),
    .B(_3236_),
    .Y(_3557_));
 sg13g2_xnor2_1 _8587_ (.Y(_3558_),
    .A(_3365_),
    .B(_3557_));
 sg13g2_nor2_1 _8588_ (.A(_0027_),
    .B(_3558_),
    .Y(_3559_));
 sg13g2_inv_1 _8589_ (.Y(_3560_),
    .A(_3559_));
 sg13g2_nand2_1 _8590_ (.Y(_3561_),
    .A(_3558_),
    .B(_0027_));
 sg13g2_nand2_1 _8591_ (.Y(_3562_),
    .A(_3560_),
    .B(_3561_));
 sg13g2_inv_1 _8592_ (.Y(_3563_),
    .A(_3562_));
 sg13g2_nand2_1 _8593_ (.Y(_3564_),
    .A(_3556_),
    .B(_3563_));
 sg13g2_nand3_1 _8594_ (.B(_3562_),
    .C(_3555_),
    .A(_3552_),
    .Y(_3565_));
 sg13g2_nand3_1 _8595_ (.B(_3565_),
    .C(_3182_),
    .A(_3564_),
    .Y(_3566_));
 sg13g2_nand2_1 _8596_ (.Y(_3567_),
    .A(_3244_),
    .B(_3169_));
 sg13g2_and2_1 _8597_ (.A(_3567_),
    .B(_3452_),
    .X(_3568_));
 sg13g2_nand2_1 _8598_ (.Y(_3569_),
    .A(_3568_),
    .B(_3540_));
 sg13g2_nand2_1 _8599_ (.Y(_3570_),
    .A(_3566_),
    .B(_3569_));
 sg13g2_nand2_1 _8600_ (.Y(_3571_),
    .A(_3217_),
    .B(_3221_));
 sg13g2_nand2_1 _8601_ (.Y(_3572_),
    .A(_3223_),
    .B(_3220_));
 sg13g2_xor2_1 _8602_ (.B(_3572_),
    .A(_3571_),
    .X(_3573_));
 sg13g2_inv_1 _8603_ (.Y(_3574_),
    .A(_3573_));
 sg13g2_nand3_1 _8604_ (.B(_3570_),
    .C(_3574_),
    .A(_3544_),
    .Y(_3575_));
 sg13g2_nand2_1 _8605_ (.Y(_3576_),
    .A(_3570_),
    .B(_3574_));
 sg13g2_inv_1 _8606_ (.Y(_3577_),
    .A(_3544_));
 sg13g2_nand2_1 _8607_ (.Y(_3578_),
    .A(_3576_),
    .B(_3577_));
 sg13g2_nand2_1 _8608_ (.Y(_3579_),
    .A(_3575_),
    .B(_3578_));
 sg13g2_xnor2_1 _8609_ (.Y(_3580_),
    .A(_3539_),
    .B(_3579_));
 sg13g2_nand2_1 _8610_ (.Y(_3581_),
    .A(_3570_),
    .B(_3573_));
 sg13g2_nand3_1 _8611_ (.B(_3569_),
    .C(_3574_),
    .A(_3566_),
    .Y(_3582_));
 sg13g2_nand2_1 _8612_ (.Y(_3583_),
    .A(_3302_),
    .B(_3541_));
 sg13g2_xor2_1 _8613_ (.B(_3212_),
    .A(_3216_),
    .X(_3584_));
 sg13g2_nand2_1 _8614_ (.Y(_3585_),
    .A(_3583_),
    .B(_3584_));
 sg13g2_nand3_1 _8615_ (.B(_3582_),
    .C(_3585_),
    .A(_3581_),
    .Y(_3586_));
 sg13g2_nor2_1 _8616_ (.A(_4275_),
    .B(_0615_),
    .Y(_3587_));
 sg13g2_buf_2 _8617_ (.A(_3587_),
    .X(_3588_));
 sg13g2_a21oi_1 _8618_ (.A1(_3581_),
    .A2(_3582_),
    .Y(_3589_),
    .B1(_3585_));
 sg13g2_a21oi_1 _8619_ (.A1(_3586_),
    .A2(_3588_),
    .Y(_3590_),
    .B1(_3589_));
 sg13g2_inv_1 _8620_ (.Y(_3591_),
    .A(_3590_));
 sg13g2_nand2_1 _8621_ (.Y(_3592_),
    .A(_3580_),
    .B(_3591_));
 sg13g2_nand2_1 _8622_ (.Y(_3593_),
    .A(_3579_),
    .B(_3236_));
 sg13g2_nand3_1 _8623_ (.B(_3578_),
    .C(_3539_),
    .A(_3575_),
    .Y(_3594_));
 sg13g2_nand2_1 _8624_ (.Y(_3595_),
    .A(_3593_),
    .B(_3594_));
 sg13g2_nand2_1 _8625_ (.Y(_3596_),
    .A(_3595_),
    .B(_3590_));
 sg13g2_nand2_1 _8626_ (.Y(_3597_),
    .A(_3592_),
    .B(_3596_));
 sg13g2_inv_4 _8627_ (.A(_3588_),
    .Y(_3598_));
 sg13g2_inv_1 _8628_ (.Y(_3599_),
    .A(_3568_));
 sg13g2_nor2_1 _8629_ (.A(net34),
    .B(_3599_),
    .Y(_3600_));
 sg13g2_inv_1 _8630_ (.Y(_3601_),
    .A(_3600_));
 sg13g2_nand2_1 _8631_ (.Y(_3602_),
    .A(_3597_),
    .B(_3601_));
 sg13g2_nand3_1 _8632_ (.B(_3596_),
    .C(_3600_),
    .A(_3592_),
    .Y(_3603_));
 sg13g2_nand2_1 _8633_ (.Y(_3604_),
    .A(_3602_),
    .B(_3603_));
 sg13g2_nand3_1 _8634_ (.B(_3569_),
    .C(_3573_),
    .A(_3566_),
    .Y(_3605_));
 sg13g2_nand3b_1 _8635_ (.B(_3576_),
    .C(_3605_),
    .Y(_3606_),
    .A_N(_3585_));
 sg13g2_nand2_1 _8636_ (.Y(_3607_),
    .A(_3606_),
    .B(_3586_));
 sg13g2_nand2_1 _8637_ (.Y(_3608_),
    .A(_3607_),
    .B(net34));
 sg13g2_nand3_1 _8638_ (.B(_3586_),
    .C(_3588_),
    .A(_3606_),
    .Y(_3609_));
 sg13g2_nand2_1 _8639_ (.Y(_3610_),
    .A(_3608_),
    .B(_3609_));
 sg13g2_inv_1 _8640_ (.Y(_3611_),
    .A(_3610_));
 sg13g2_xor2_1 _8641_ (.B(_3203_),
    .A(_3209_),
    .X(_3612_));
 sg13g2_nor2b_1 _8642_ (.A(_3248_),
    .B_N(_3612_),
    .Y(_3613_));
 sg13g2_inv_1 _8643_ (.Y(_3614_),
    .A(_3613_));
 sg13g2_xor2_1 _8644_ (.B(_3583_),
    .A(_3584_),
    .X(_3615_));
 sg13g2_inv_1 _8645_ (.Y(_3616_),
    .A(_3615_));
 sg13g2_nor2_1 _8646_ (.A(_3614_),
    .B(_3616_),
    .Y(_3617_));
 sg13g2_nand2_1 _8647_ (.Y(_3618_),
    .A(_3611_),
    .B(_3617_));
 sg13g2_inv_1 _8648_ (.Y(_3619_),
    .A(_3618_));
 sg13g2_nand2_1 _8649_ (.Y(_3620_),
    .A(_3604_),
    .B(_3619_));
 sg13g2_nand3_1 _8650_ (.B(_3603_),
    .C(_3618_),
    .A(_3602_),
    .Y(_3621_));
 sg13g2_nand2_1 _8651_ (.Y(_3622_),
    .A(_3620_),
    .B(_3621_));
 sg13g2_nand2_1 _8652_ (.Y(_3623_),
    .A(_3610_),
    .B(_3617_));
 sg13g2_inv_1 _8653_ (.Y(_3624_),
    .A(_3617_));
 sg13g2_nand3_1 _8654_ (.B(_3609_),
    .C(_3624_),
    .A(_3608_),
    .Y(_3625_));
 sg13g2_xnor2_1 _8655_ (.Y(_3626_),
    .A(_3614_),
    .B(_3615_));
 sg13g2_a21oi_1 _8656_ (.A1(_3195_),
    .A2(_3196_),
    .Y(_3627_),
    .B1(_3200_));
 sg13g2_nor2b_1 _8657_ (.A(_3627_),
    .B_N(_3201_),
    .Y(_3628_));
 sg13g2_nand2_1 _8658_ (.Y(_3629_),
    .A(_3245_),
    .B(_3628_));
 sg13g2_xor2_1 _8659_ (.B(_3248_),
    .A(_3612_),
    .X(_3630_));
 sg13g2_nor2_1 _8660_ (.A(_3629_),
    .B(_3630_),
    .Y(_3631_));
 sg13g2_nand2_1 _8661_ (.Y(_3632_),
    .A(_3626_),
    .B(_3631_));
 sg13g2_nand3_1 _8662_ (.B(_3625_),
    .C(_3632_),
    .A(_3623_),
    .Y(_3633_));
 sg13g2_xnor2_1 _8663_ (.Y(_3634_),
    .A(_3629_),
    .B(_3630_));
 sg13g2_xnor2_1 _8664_ (.Y(_3635_),
    .A(_3628_),
    .B(_3245_));
 sg13g2_nand3_1 _8665_ (.B(_0300_),
    .C(_3199_),
    .A(_3197_),
    .Y(_3636_));
 sg13g2_nand2b_1 _8666_ (.Y(_3637_),
    .B(_3636_),
    .A_N(_3200_));
 sg13g2_nor2_1 _8667_ (.A(_3183_),
    .B(_3637_),
    .Y(_3638_));
 sg13g2_nor2b_1 _8668_ (.A(_3635_),
    .B_N(_3638_),
    .Y(_3639_));
 sg13g2_nor2b_1 _8669_ (.A(_3634_),
    .B_N(_3639_),
    .Y(_3640_));
 sg13g2_nand2_1 _8670_ (.Y(_3641_),
    .A(_3626_),
    .B(_3640_));
 sg13g2_inv_1 _8671_ (.Y(_3642_),
    .A(_3641_));
 sg13g2_a21oi_1 _8672_ (.A1(_3623_),
    .A2(_3625_),
    .Y(_3643_),
    .B1(_3632_));
 sg13g2_a21oi_1 _8673_ (.A1(_3633_),
    .A2(_3642_),
    .Y(_3644_),
    .B1(_3643_));
 sg13g2_inv_4 _8674_ (.A(_3644_),
    .Y(_3645_));
 sg13g2_inv_1 _8675_ (.Y(_3646_),
    .A(_3592_));
 sg13g2_a21oi_2 _8676_ (.B1(_3646_),
    .Y(_3647_),
    .A2(_3600_),
    .A1(_3596_));
 sg13g2_nor2_1 _8677_ (.A(net34),
    .B(_3455_),
    .Y(_3648_));
 sg13g2_inv_1 _8678_ (.Y(_3649_),
    .A(_3575_));
 sg13g2_a21oi_2 _8679_ (.B1(_3649_),
    .Y(_3650_),
    .A2(_3539_),
    .A1(_3578_));
 sg13g2_nor2_1 _8680_ (.A(net51),
    .B(_3150_),
    .Y(_3651_));
 sg13g2_a21oi_1 _8681_ (.A1(_3444_),
    .A2(_0615_),
    .Y(_3652_),
    .B1(_3651_));
 sg13g2_xnor2_1 _8682_ (.Y(_3653_),
    .A(_0298_),
    .B(_3652_));
 sg13g2_nand2b_1 _8683_ (.Y(_3654_),
    .B(_3227_),
    .A_N(_0035_));
 sg13g2_nand2_1 _8684_ (.Y(_3655_),
    .A(_3234_),
    .B(_3654_));
 sg13g2_xor2_1 _8685_ (.B(_3655_),
    .A(_3653_),
    .X(_3656_));
 sg13g2_nor2_1 _8686_ (.A(_3453_),
    .B(_3451_),
    .Y(_3657_));
 sg13g2_nor3_1 _8687_ (.A(_3169_),
    .B(_3244_),
    .C(_3451_),
    .Y(_3658_));
 sg13g2_nor3_1 _8688_ (.A(_3553_),
    .B(_3657_),
    .C(_3658_),
    .Y(_3659_));
 sg13g2_xnor2_1 _8689_ (.Y(_3660_),
    .A(_3549_),
    .B(_3659_));
 sg13g2_nand2_1 _8690_ (.Y(_3661_),
    .A(_3660_),
    .B(_3540_));
 sg13g2_nand3_1 _8691_ (.B(_3385_),
    .C(_3661_),
    .A(_3458_),
    .Y(_3662_));
 sg13g2_xnor2_1 _8692_ (.Y(_3663_),
    .A(_3656_),
    .B(_3662_));
 sg13g2_xnor2_1 _8693_ (.Y(_3664_),
    .A(_3650_),
    .B(_3663_));
 sg13g2_xnor2_1 _8694_ (.Y(_3665_),
    .A(_3648_),
    .B(_3664_));
 sg13g2_xnor2_1 _8695_ (.Y(_3666_),
    .A(_3647_),
    .B(_3665_));
 sg13g2_nand3_1 _8696_ (.B(_3645_),
    .C(_3666_),
    .A(_3622_),
    .Y(_3667_));
 sg13g2_nand2b_1 _8697_ (.Y(_3668_),
    .B(_3647_),
    .A_N(_3665_));
 sg13g2_nor2_1 _8698_ (.A(_3618_),
    .B(_3604_),
    .Y(_3669_));
 sg13g2_nor2b_1 _8699_ (.A(_3647_),
    .B_N(_3665_),
    .Y(_3670_));
 sg13g2_a21oi_1 _8700_ (.A1(_3668_),
    .A2(_3669_),
    .Y(_3671_),
    .B1(_3670_));
 sg13g2_nand2_1 _8701_ (.Y(_3672_),
    .A(_3667_),
    .B(_3671_));
 sg13g2_nand2_1 _8702_ (.Y(_3673_),
    .A(_3663_),
    .B(_3650_));
 sg13g2_nor2_1 _8703_ (.A(_3650_),
    .B(_3663_),
    .Y(_3674_));
 sg13g2_a21oi_1 _8704_ (.A1(_3673_),
    .A2(_3648_),
    .Y(_3675_),
    .B1(_3674_));
 sg13g2_inv_1 _8705_ (.Y(_3676_),
    .A(_3660_));
 sg13g2_nor2_1 _8706_ (.A(net34),
    .B(_3676_),
    .Y(_3677_));
 sg13g2_nand2_1 _8707_ (.Y(_3678_),
    .A(_3662_),
    .B(_3656_));
 sg13g2_nor2_1 _8708_ (.A(net44),
    .B(_3508_),
    .Y(_3679_));
 sg13g2_a21oi_1 _8709_ (.A1(net44),
    .A2(_3444_),
    .Y(_3680_),
    .B1(_3679_));
 sg13g2_xnor2_1 _8710_ (.Y(_3681_),
    .A(_0033_),
    .B(_3680_));
 sg13g2_a22oi_1 _8711_ (.Y(_3682_),
    .B1(_3653_),
    .B2(_3655_),
    .A2(_3652_),
    .A1(_3507_));
 sg13g2_xnor2_1 _8712_ (.Y(_3683_),
    .A(_3681_),
    .B(_3682_));
 sg13g2_nand2_1 _8713_ (.Y(_3684_),
    .A(_3564_),
    .B(_3565_));
 sg13g2_inv_1 _8714_ (.Y(_3685_),
    .A(_3684_));
 sg13g2_a21oi_1 _8715_ (.A1(_3685_),
    .A2(_3540_),
    .Y(_3686_),
    .B1(_3456_));
 sg13g2_nand2_1 _8716_ (.Y(_3687_),
    .A(_3512_),
    .B(_3686_));
 sg13g2_xnor2_1 _8717_ (.Y(_3688_),
    .A(_3683_),
    .B(_3687_));
 sg13g2_xnor2_1 _8718_ (.Y(_3689_),
    .A(_3678_),
    .B(_3688_));
 sg13g2_xor2_1 _8719_ (.B(_3689_),
    .A(_3677_),
    .X(_3690_));
 sg13g2_xor2_1 _8720_ (.B(_3690_),
    .A(_3675_),
    .X(_3691_));
 sg13g2_inv_1 _8721_ (.Y(_3692_),
    .A(_3691_));
 sg13g2_nand2_1 _8722_ (.Y(_3693_),
    .A(_3672_),
    .B(_3692_));
 sg13g2_nand3_1 _8723_ (.B(_3671_),
    .C(_3691_),
    .A(_3667_),
    .Y(_3694_));
 sg13g2_nand2_1 _8724_ (.Y(_3695_),
    .A(_3693_),
    .B(_3694_));
 sg13g2_nand2_1 _8725_ (.Y(_3696_),
    .A(net46),
    .B(_4210_));
 sg13g2_xor2_1 _8726_ (.B(_3696_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[7] ),
    .X(_3697_));
 sg13g2_inv_1 _8727_ (.Y(_3698_),
    .A(_3369_));
 sg13g2_nor2_1 _8728_ (.A(_3365_),
    .B(_3698_),
    .Y(_3699_));
 sg13g2_nand3_1 _8729_ (.B(_3400_),
    .C(_3481_),
    .A(_3699_),
    .Y(_3700_));
 sg13g2_nand2_1 _8730_ (.Y(_3701_),
    .A(_3539_),
    .B(_3700_));
 sg13g2_xnor2_1 _8731_ (.Y(_3702_),
    .A(_3697_),
    .B(_3701_));
 sg13g2_a21o_1 _8732_ (.A2(_3400_),
    .A1(_3699_),
    .B1(_3236_),
    .X(_3703_));
 sg13g2_xnor2_1 _8733_ (.Y(_3704_),
    .A(_3481_),
    .B(_3703_));
 sg13g2_nor2_1 _8734_ (.A(_3699_),
    .B(_3236_),
    .Y(_3705_));
 sg13g2_xor2_1 _8735_ (.B(_3705_),
    .A(_3400_),
    .X(_3706_));
 sg13g2_nor2_1 _8736_ (.A(_0032_),
    .B(_3706_),
    .Y(_3707_));
 sg13g2_xnor2_1 _8737_ (.Y(_3708_),
    .A(_3364_),
    .B(_3706_));
 sg13g2_xnor2_1 _8738_ (.Y(_3709_),
    .A(_3308_),
    .B(_3558_));
 sg13g2_nand2b_1 _8739_ (.Y(_3710_),
    .B(_3549_),
    .A_N(_3709_));
 sg13g2_o21ai_1 _8740_ (.B1(_3561_),
    .Y(_3711_),
    .A1(_3554_),
    .A2(_3559_));
 sg13g2_o21ai_1 _8741_ (.B1(_3711_),
    .Y(_3712_),
    .A1(_3710_),
    .A2(_3659_));
 sg13g2_nor2b_1 _8742_ (.A(_3708_),
    .B_N(_3712_),
    .Y(_3713_));
 sg13g2_xnor2_1 _8743_ (.Y(_3714_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[6] ),
    .B(_3704_));
 sg13g2_o21ai_1 _8744_ (.B1(_3714_),
    .Y(_3715_),
    .A1(_3707_),
    .A2(_3713_));
 sg13g2_o21ai_1 _8745_ (.B1(_3715_),
    .Y(_3716_),
    .A1(_0031_),
    .A2(_3704_));
 sg13g2_xor2_1 _8746_ (.B(_3716_),
    .A(_3702_),
    .X(_3717_));
 sg13g2_nand2_1 _8747_ (.Y(_3718_),
    .A(_3717_),
    .B(net46));
 sg13g2_inv_1 _8748_ (.Y(_3719_),
    .A(_3718_));
 sg13g2_nand2_1 _8749_ (.Y(_3720_),
    .A(_3695_),
    .B(_3719_));
 sg13g2_nand3_1 _8750_ (.B(_3694_),
    .C(_3718_),
    .A(_3693_),
    .Y(_3721_));
 sg13g2_nand2_1 _8751_ (.Y(_3722_),
    .A(_3720_),
    .B(_3721_));
 sg13g2_inv_1 _8752_ (.Y(_3723_),
    .A(_3708_));
 sg13g2_nor2_1 _8753_ (.A(_3709_),
    .B(_3708_),
    .Y(_3724_));
 sg13g2_a221oi_1 _8754_ (.B2(_3724_),
    .C1(_3707_),
    .B1(_3556_),
    .A1(_3559_),
    .Y(_3725_),
    .A2(_3723_));
 sg13g2_xnor2_1 _8755_ (.Y(_3726_),
    .A(_3714_),
    .B(_3725_));
 sg13g2_nor2_1 _8756_ (.A(net43),
    .B(_3726_),
    .Y(_3727_));
 sg13g2_xor2_1 _8757_ (.B(_3666_),
    .A(_3727_),
    .X(_3728_));
 sg13g2_a21oi_1 _8758_ (.A1(_3622_),
    .A2(_3645_),
    .Y(_3729_),
    .B1(_3669_));
 sg13g2_xnor2_1 _8759_ (.Y(_3730_),
    .A(_3728_),
    .B(_3729_));
 sg13g2_nor2_1 _8760_ (.A(_0326_),
    .B(_3730_),
    .Y(_3731_));
 sg13g2_a21oi_1 _8761_ (.A1(_3722_),
    .A2(_0331_),
    .Y(_3732_),
    .B1(_3731_));
 sg13g2_nor2_1 _8762_ (.A(_0793_),
    .B(_3685_),
    .Y(_3733_));
 sg13g2_nand2_1 _8763_ (.Y(_3734_),
    .A(_3623_),
    .B(_3625_));
 sg13g2_inv_1 _8764_ (.Y(_3735_),
    .A(_3632_));
 sg13g2_nand2_1 _8765_ (.Y(_3736_),
    .A(_3734_),
    .B(_3735_));
 sg13g2_nand2_1 _8766_ (.Y(_3737_),
    .A(_3736_),
    .B(_3633_));
 sg13g2_nand2_1 _8767_ (.Y(_3738_),
    .A(_3737_),
    .B(_3641_));
 sg13g2_nand3_1 _8768_ (.B(_3633_),
    .C(_3642_),
    .A(_3736_),
    .Y(_3739_));
 sg13g2_nand2_1 _8769_ (.Y(_3740_),
    .A(_3738_),
    .B(_3739_));
 sg13g2_nand2b_1 _8770_ (.Y(_3741_),
    .B(_3740_),
    .A_N(_3733_));
 sg13g2_nand3_1 _8771_ (.B(_3739_),
    .C(_3733_),
    .A(_3738_),
    .Y(_3742_));
 sg13g2_nand2_1 _8772_ (.Y(_3743_),
    .A(_3741_),
    .B(_3742_));
 sg13g2_nand2_1 _8773_ (.Y(_3744_),
    .A(_3676_),
    .B(net46));
 sg13g2_nor2_1 _8774_ (.A(_3631_),
    .B(_3640_),
    .Y(_3745_));
 sg13g2_xor2_1 _8775_ (.B(_3745_),
    .A(_3626_),
    .X(_3746_));
 sg13g2_xor2_1 _8776_ (.B(_3746_),
    .A(_3744_),
    .X(_3747_));
 sg13g2_nand2_1 _8777_ (.Y(_3748_),
    .A(_3455_),
    .B(_3266_));
 sg13g2_xnor2_1 _8778_ (.Y(_3749_),
    .A(_3639_),
    .B(_3634_));
 sg13g2_xnor2_1 _8779_ (.Y(_3750_),
    .A(_3748_),
    .B(_3749_));
 sg13g2_nand2_1 _8780_ (.Y(_3751_),
    .A(_3750_),
    .B(_0312_));
 sg13g2_nand2_1 _8781_ (.Y(_3752_),
    .A(_3751_),
    .B(_3348_));
 sg13g2_nor2_1 _8782_ (.A(_3348_),
    .B(_3751_),
    .Y(_3753_));
 sg13g2_a21oi_1 _8783_ (.A1(_3747_),
    .A2(_3752_),
    .Y(_3754_),
    .B1(_3753_));
 sg13g2_nand3_1 _8784_ (.B(_3351_),
    .C(_3754_),
    .A(_3743_),
    .Y(_3755_));
 sg13g2_nand2_1 _8785_ (.Y(_3756_),
    .A(_3755_),
    .B(\main.demo._q_th[5] ));
 sg13g2_xnor2_1 _8786_ (.Y(_3757_),
    .A(_3708_),
    .B(_3712_));
 sg13g2_nor2_1 _8787_ (.A(_0793_),
    .B(_3757_),
    .Y(_3758_));
 sg13g2_xnor2_1 _8788_ (.Y(_3759_),
    .A(_3645_),
    .B(_3622_));
 sg13g2_xnor2_1 _8789_ (.Y(_3760_),
    .A(_3758_),
    .B(_3759_));
 sg13g2_inv_2 _8790_ (.Y(_3761_),
    .A(_3760_));
 sg13g2_nand2_1 _8791_ (.Y(_3762_),
    .A(_3756_),
    .B(_3761_));
 sg13g2_inv_2 _8792_ (.Y(_3763_),
    .A(_3743_));
 sg13g2_nor2b_1 _8793_ (.A(_3763_),
    .B_N(_3754_),
    .Y(_3764_));
 sg13g2_nand3_1 _8794_ (.B(_3764_),
    .C(_0037_),
    .A(_3760_),
    .Y(_3765_));
 sg13g2_nand2_1 _8795_ (.Y(_3766_),
    .A(_3762_),
    .B(_3765_));
 sg13g2_xnor2_1 _8796_ (.Y(_3767_),
    .A(_0036_),
    .B(_3730_));
 sg13g2_nand2_1 _8797_ (.Y(_3768_),
    .A(_3766_),
    .B(_3767_));
 sg13g2_nand2_1 _8798_ (.Y(_3769_),
    .A(_3732_),
    .B(_3768_));
 sg13g2_nor2_1 _8799_ (.A(_0331_),
    .B(_3722_),
    .Y(_3770_));
 sg13g2_nor2_1 _8800_ (.A(net54),
    .B(_3770_),
    .Y(_3771_));
 sg13g2_nand2_1 _8801_ (.Y(_3772_),
    .A(_3769_),
    .B(_3771_));
 sg13g2_buf_8 _8802_ (.A(_3772_),
    .X(_3773_));
 sg13g2_nand2_1 _8803_ (.Y(_3774_),
    .A(_3599_),
    .B(_3266_));
 sg13g2_xnor2_1 _8804_ (.Y(_3775_),
    .A(_3638_),
    .B(_3635_));
 sg13g2_xnor2_1 _8805_ (.Y(_3776_),
    .A(_3774_),
    .B(_3775_));
 sg13g2_nand2_1 _8806_ (.Y(_3777_),
    .A(_3637_),
    .B(_3588_));
 sg13g2_o21ai_1 _8807_ (.B1(_3777_),
    .Y(_3778_),
    .A1(_3588_),
    .A2(_3776_));
 sg13g2_nand2_1 _8808_ (.Y(_3779_),
    .A(net11),
    .B(_3778_));
 sg13g2_a21oi_1 _8809_ (.A1(_3538_),
    .A2(_3779_),
    .Y(_3780_),
    .B1(net54));
 sg13g2_nor2_1 _8810_ (.A(_3779_),
    .B(_3538_),
    .Y(_3781_));
 sg13g2_inv_1 _8811_ (.Y(_3782_),
    .A(_3781_));
 sg13g2_nor2_1 _8812_ (.A(net68),
    .B(_3394_),
    .Y(_3783_));
 sg13g2_nand2_1 _8813_ (.Y(_3784_),
    .A(_3761_),
    .B(_3783_));
 sg13g2_nor2b_1 _8814_ (.A(net34),
    .B_N(_3776_),
    .Y(_3785_));
 sg13g2_a21oi_1 _8815_ (.A1(_3750_),
    .A2(net34),
    .Y(_3786_),
    .B1(_3785_));
 sg13g2_nand2_1 _8816_ (.Y(_3787_),
    .A(net11),
    .B(_3786_));
 sg13g2_nor2_1 _8817_ (.A(_4274_),
    .B(_3397_),
    .Y(_3788_));
 sg13g2_buf_2 _8818_ (.A(_3788_),
    .X(_3789_));
 sg13g2_nand2b_1 _8819_ (.Y(_3790_),
    .B(_3789_),
    .A_N(_3537_));
 sg13g2_o21ai_1 _8820_ (.B1(_3790_),
    .Y(_3791_),
    .A1(_3784_),
    .A2(_3787_));
 sg13g2_a21o_1 _8821_ (.A2(_3782_),
    .A1(_3780_),
    .B1(_3791_),
    .X(\main.demo._t___block_68_frag[0] ));
 sg13g2_inv_1 _8822_ (.Y(_3792_),
    .A(_3747_));
 sg13g2_nor2_1 _8823_ (.A(_3588_),
    .B(_3792_),
    .Y(_3793_));
 sg13g2_a21oi_1 _8824_ (.A1(_3588_),
    .A2(_3750_),
    .Y(_3794_),
    .B1(_3793_));
 sg13g2_nand2_1 _8825_ (.Y(_3795_),
    .A(net11),
    .B(_3794_));
 sg13g2_nor2_1 _8826_ (.A(net54),
    .B(_3345_),
    .Y(_3796_));
 sg13g2_a21oi_1 _8827_ (.A1(_3261_),
    .A2(net54),
    .Y(_3797_),
    .B1(_3796_));
 sg13g2_a21oi_2 _8828_ (.B1(_3797_),
    .Y(_3798_),
    .A2(_3535_),
    .A1(_3533_));
 sg13g2_nand2_1 _8829_ (.Y(_3799_),
    .A(_3798_),
    .B(_3789_));
 sg13g2_o21ai_1 _8830_ (.B1(_3799_),
    .Y(_3800_),
    .A1(_3784_),
    .A2(_3795_));
 sg13g2_nand2b_1 _8831_ (.Y(_3801_),
    .B(_3787_),
    .A_N(_3798_));
 sg13g2_nand3_1 _8832_ (.B(_3786_),
    .C(_3798_),
    .A(net11),
    .Y(_3802_));
 sg13g2_nand2_1 _8833_ (.Y(_3803_),
    .A(_3801_),
    .B(_3802_));
 sg13g2_nand2_1 _8834_ (.Y(_3804_),
    .A(_3782_),
    .B(_3803_));
 sg13g2_xnor2_1 _8835_ (.Y(_3805_),
    .A(_3798_),
    .B(_3787_));
 sg13g2_nand2_1 _8836_ (.Y(_3806_),
    .A(_3781_),
    .B(_3805_));
 sg13g2_nand3_1 _8837_ (.B(net68),
    .C(_3806_),
    .A(_3804_),
    .Y(_3807_));
 sg13g2_nand2b_1 _8838_ (.Y(\main.demo._t___block_68_frag[1] ),
    .B(_3807_),
    .A_N(_3800_));
 sg13g2_inv_1 _8839_ (.Y(_3808_),
    .A(_3337_));
 sg13g2_nor2b_1 _8840_ (.A(_4274_),
    .B_N(_3346_),
    .Y(_3809_));
 sg13g2_a21o_1 _8841_ (.A2(net68),
    .A1(_3808_),
    .B1(_3809_),
    .X(_3810_));
 sg13g2_inv_1 _8842_ (.Y(_3811_),
    .A(_3810_));
 sg13g2_a21oi_1 _8843_ (.A1(_3533_),
    .A2(_3535_),
    .Y(_3812_),
    .B1(_3811_));
 sg13g2_nand2b_1 _8844_ (.Y(_3813_),
    .B(_3795_),
    .A_N(_3812_));
 sg13g2_nand3_1 _8845_ (.B(_3794_),
    .C(_3812_),
    .A(net11),
    .Y(_3814_));
 sg13g2_buf_8 _8846_ (.A(_3814_),
    .X(_3815_));
 sg13g2_nand2_1 _8847_ (.Y(_3816_),
    .A(_3813_),
    .B(_3815_));
 sg13g2_nand2_1 _8848_ (.Y(_3817_),
    .A(_3806_),
    .B(_3802_));
 sg13g2_xor2_1 _8849_ (.B(_3817_),
    .A(_3816_),
    .X(_3818_));
 sg13g2_nor2_1 _8850_ (.A(net34),
    .B(_3792_),
    .Y(_3819_));
 sg13g2_a21oi_1 _8851_ (.A1(_3763_),
    .A2(net34),
    .Y(_3820_),
    .B1(_3819_));
 sg13g2_nand2_1 _8852_ (.Y(_3821_),
    .A(net11),
    .B(_3820_));
 sg13g2_nor2_1 _8853_ (.A(_3784_),
    .B(_3821_),
    .Y(_3822_));
 sg13g2_a21oi_1 _8854_ (.A1(_3789_),
    .A2(_3812_),
    .Y(_3823_),
    .B1(_3822_));
 sg13g2_o21ai_1 _8855_ (.B1(_3823_),
    .Y(\main.demo._t___block_68_frag[2] ),
    .A1(_2176_),
    .A2(_3818_));
 sg13g2_nand2_1 _8856_ (.Y(_3824_),
    .A(_3397_),
    .B(_0786_));
 sg13g2_o21ai_1 _8857_ (.B1(_3824_),
    .Y(_3825_),
    .A1(_0786_),
    .A2(_3339_));
 sg13g2_a21oi_1 _8858_ (.A1(_3533_),
    .A2(_3535_),
    .Y(_3826_),
    .B1(_3825_));
 sg13g2_inv_1 _8859_ (.Y(_3827_),
    .A(_3826_));
 sg13g2_nand2_1 _8860_ (.Y(_3828_),
    .A(_3821_),
    .B(_3827_));
 sg13g2_nand3_1 _8861_ (.B(_3820_),
    .C(_3826_),
    .A(net11),
    .Y(_3829_));
 sg13g2_nand2_1 _8862_ (.Y(_3830_),
    .A(_3828_),
    .B(_3829_));
 sg13g2_nor2_1 _8863_ (.A(_3803_),
    .B(_3816_),
    .Y(_3831_));
 sg13g2_inv_1 _8864_ (.Y(_3832_),
    .A(_3813_));
 sg13g2_a21oi_1 _8865_ (.A1(_3802_),
    .A2(_3815_),
    .Y(_3833_),
    .B1(_3832_));
 sg13g2_a21oi_1 _8866_ (.A1(_3831_),
    .A2(_3781_),
    .Y(_3834_),
    .B1(_3833_));
 sg13g2_xnor2_1 _8867_ (.Y(_3835_),
    .A(_3830_),
    .B(_3834_));
 sg13g2_a22oi_1 _8868_ (.Y(_3836_),
    .B1(_3789_),
    .B2(_3826_),
    .A2(_3783_),
    .A1(_3761_));
 sg13g2_o21ai_1 _8869_ (.B1(_3836_),
    .Y(\main.demo._t___block_68_frag[3] ),
    .A1(_2176_),
    .A2(_3835_));
 sg13g2_a21oi_1 _8870_ (.A1(_3471_),
    .A2(net68),
    .Y(_3837_),
    .B1(_3789_));
 sg13g2_a21oi_1 _8871_ (.A1(_3533_),
    .A2(_3535_),
    .Y(_3838_),
    .B1(_3837_));
 sg13g2_o21ai_1 _8872_ (.B1(_3609_),
    .Y(_3839_),
    .A1(_3588_),
    .A2(_3760_));
 sg13g2_nand2_1 _8873_ (.Y(_3840_),
    .A(_3773_),
    .B(_3839_));
 sg13g2_nand2b_1 _8874_ (.Y(_3841_),
    .B(_3840_),
    .A_N(_3838_));
 sg13g2_nand3_1 _8875_ (.B(_3839_),
    .C(_3838_),
    .A(_3773_),
    .Y(_3842_));
 sg13g2_nand2_1 _8876_ (.Y(_3843_),
    .A(_3841_),
    .B(_3842_));
 sg13g2_nor2_1 _8877_ (.A(_3830_),
    .B(_3816_),
    .Y(_3844_));
 sg13g2_nand2_1 _8878_ (.Y(_3845_),
    .A(_3817_),
    .B(_3844_));
 sg13g2_inv_1 _8879_ (.Y(_3846_),
    .A(_3815_));
 sg13g2_inv_1 _8880_ (.Y(_3847_),
    .A(_3829_));
 sg13g2_o21ai_1 _8881_ (.B1(_3828_),
    .Y(_3848_),
    .A1(_3846_),
    .A2(_3847_));
 sg13g2_nand2_1 _8882_ (.Y(_3849_),
    .A(_3845_),
    .B(_3848_));
 sg13g2_nand2b_1 _8883_ (.Y(_3850_),
    .B(_3849_),
    .A_N(_3843_));
 sg13g2_nand3_1 _8884_ (.B(_3843_),
    .C(_3848_),
    .A(_3845_),
    .Y(_3851_));
 sg13g2_nand3_1 _8885_ (.B(_3851_),
    .C(net68),
    .A(_3850_),
    .Y(_3852_));
 sg13g2_nor2_1 _8886_ (.A(_3598_),
    .B(_3761_),
    .Y(_3853_));
 sg13g2_a21oi_1 _8887_ (.A1(_3730_),
    .A2(_3598_),
    .Y(_3854_),
    .B1(_3853_));
 sg13g2_nand2_1 _8888_ (.Y(_3855_),
    .A(net11),
    .B(_3854_));
 sg13g2_nor2_1 _8889_ (.A(_3784_),
    .B(_3855_),
    .Y(_3856_));
 sg13g2_nor2_1 _8890_ (.A(_3789_),
    .B(_3856_),
    .Y(_3857_));
 sg13g2_nand2_1 _8891_ (.Y(\main.demo._t___block_68_frag[4] ),
    .A(_3852_),
    .B(_3857_));
 sg13g2_nor2_1 _8892_ (.A(_3830_),
    .B(_3843_),
    .Y(_3858_));
 sg13g2_nand2_1 _8893_ (.Y(_3859_),
    .A(_3847_),
    .B(_3841_));
 sg13g2_nand2_1 _8894_ (.Y(_3860_),
    .A(_3859_),
    .B(_3842_));
 sg13g2_a21oi_1 _8895_ (.A1(_3858_),
    .A2(_3833_),
    .Y(_3861_),
    .B1(_3860_));
 sg13g2_nand3_1 _8896_ (.B(_3858_),
    .C(_3781_),
    .A(_3831_),
    .Y(_3862_));
 sg13g2_nand2_1 _8897_ (.Y(_3863_),
    .A(_3861_),
    .B(_3862_));
 sg13g2_nor2_1 _8898_ (.A(net54),
    .B(_3530_),
    .Y(_3864_));
 sg13g2_a21oi_1 _8899_ (.A1(_3474_),
    .A2(net54),
    .Y(_3865_),
    .B1(_3864_));
 sg13g2_nand2_1 _8900_ (.Y(_3866_),
    .A(_3536_),
    .B(_3865_));
 sg13g2_xor2_1 _8901_ (.B(_3855_),
    .A(_3866_),
    .X(_3867_));
 sg13g2_nand2_1 _8902_ (.Y(_3868_),
    .A(_3863_),
    .B(_3867_));
 sg13g2_inv_1 _8903_ (.Y(_3869_),
    .A(_3867_));
 sg13g2_nand3_1 _8904_ (.B(_3862_),
    .C(_3869_),
    .A(_3861_),
    .Y(_3870_));
 sg13g2_nand3_1 _8905_ (.B(_3870_),
    .C(net68),
    .A(_3868_),
    .Y(_3871_));
 sg13g2_nand3_1 _8906_ (.B(_3789_),
    .C(_3865_),
    .A(_3536_),
    .Y(_3872_));
 sg13g2_nand2_1 _8907_ (.Y(\main.demo._t___block_68_frag[5] ),
    .A(_3871_),
    .B(_3872_));
 sg13g2_a21oi_1 _8908_ (.A1(_4139_),
    .A2(_4288_),
    .Y(_3873_),
    .B1(_0065_));
 sg13g2_xnor2_1 _8909_ (.Y(_3874_),
    .A(\main.demo._w_vga_vga_x[10] ),
    .B(_3873_));
 sg13g2_nand2_1 _8910_ (.Y(_3875_),
    .A(_4384_),
    .B(_4147_));
 sg13g2_nand2_1 _8911_ (.Y(_3876_),
    .A(_3875_),
    .B(_4289_));
 sg13g2_buf_2 _8912_ (.A(_3876_),
    .X(_3877_));
 sg13g2_o21ai_1 _8913_ (.B1(_4139_),
    .Y(_3878_),
    .A1(_0602_),
    .A2(_3877_));
 sg13g2_a21oi_1 _8914_ (.A1(_0602_),
    .A2(_3877_),
    .Y(_3879_),
    .B1(_3878_));
 sg13g2_nor2b_1 _8915_ (.A(_0004_),
    .B_N(_3879_),
    .Y(_3880_));
 sg13g2_inv_1 _8916_ (.Y(_3881_),
    .A(_0005_));
 sg13g2_o21ai_1 _8917_ (.B1(_4139_),
    .Y(_3882_),
    .A1(_4353_),
    .A2(_3877_));
 sg13g2_a21oi_1 _8918_ (.A1(_4353_),
    .A2(_3877_),
    .Y(_3883_),
    .B1(_3882_));
 sg13g2_o21ai_1 _8919_ (.B1(_4139_),
    .Y(_3884_),
    .A1(_0607_),
    .A2(_3877_));
 sg13g2_a21oi_1 _8920_ (.A1(_0607_),
    .A2(_3877_),
    .Y(_3885_),
    .B1(_3884_));
 sg13g2_inv_1 _8921_ (.Y(_3886_),
    .A(_3885_));
 sg13g2_nor2_1 _8922_ (.A(_0006_),
    .B(_3886_),
    .Y(_3887_));
 sg13g2_inv_1 _8923_ (.Y(_3888_),
    .A(_3887_));
 sg13g2_xnor2_1 _8924_ (.Y(_3889_),
    .A(_3881_),
    .B(_3883_));
 sg13g2_nor2_1 _8925_ (.A(_3888_),
    .B(_3889_),
    .Y(_3890_));
 sg13g2_a21oi_1 _8926_ (.A1(_3881_),
    .A2(_3883_),
    .Y(_3891_),
    .B1(_3890_));
 sg13g2_xnor2_1 _8927_ (.Y(_3892_),
    .A(_0004_),
    .B(_3879_));
 sg13g2_nor2b_1 _8928_ (.A(_3891_),
    .B_N(_3892_),
    .Y(_3893_));
 sg13g2_nor2_1 _8929_ (.A(_3880_),
    .B(_3893_),
    .Y(_3894_));
 sg13g2_inv_1 _8930_ (.Y(_3895_),
    .A(_3877_));
 sg13g2_a21oi_1 _8931_ (.A1(_3895_),
    .A2(_4146_),
    .Y(_3896_),
    .B1(_4155_));
 sg13g2_o21ai_1 _8932_ (.B1(_3896_),
    .Y(_3897_),
    .A1(_4146_),
    .A2(_3895_));
 sg13g2_xnor2_1 _8933_ (.Y(_3898_),
    .A(net69),
    .B(_3897_));
 sg13g2_nor2b_1 _8934_ (.A(_3894_),
    .B_N(_3898_),
    .Y(_3899_));
 sg13g2_nand2_1 _8935_ (.Y(_3900_),
    .A(_3897_),
    .B(_0003_));
 sg13g2_a21oi_1 _8936_ (.A1(_4154_),
    .A2(_4288_),
    .Y(_3901_),
    .B1(_4155_));
 sg13g2_o21ai_1 _8937_ (.B1(_3901_),
    .Y(_3902_),
    .A1(_4288_),
    .A2(_4154_));
 sg13g2_xnor2_1 _8938_ (.Y(_3903_),
    .A(_0470_),
    .B(_3902_));
 sg13g2_xnor2_1 _8939_ (.Y(_3904_),
    .A(_3900_),
    .B(_3903_));
 sg13g2_nor2b_1 _8940_ (.A(_3903_),
    .B_N(_3900_),
    .Y(_3905_));
 sg13g2_a21o_1 _8941_ (.A2(_3904_),
    .A1(_3899_),
    .B1(_3905_),
    .X(_3906_));
 sg13g2_nand2_1 _8942_ (.Y(_3907_),
    .A(_4139_),
    .B(_4288_));
 sg13g2_xnor2_1 _8943_ (.Y(_3908_),
    .A(_0508_),
    .B(_3907_));
 sg13g2_nand2_1 _8944_ (.Y(_3909_),
    .A(_3902_),
    .B(_0002_));
 sg13g2_xor2_1 _8945_ (.B(_3909_),
    .A(_3908_),
    .X(_3910_));
 sg13g2_nand2_1 _8946_ (.Y(_3911_),
    .A(_3906_),
    .B(_3910_));
 sg13g2_nand2_1 _8947_ (.Y(_3912_),
    .A(_3909_),
    .B(_3908_));
 sg13g2_nand2_1 _8948_ (.Y(_3913_),
    .A(_3911_),
    .B(_3912_));
 sg13g2_nor2_1 _8949_ (.A(_0508_),
    .B(_3907_),
    .Y(_3914_));
 sg13g2_xnor2_1 _8950_ (.Y(_3915_),
    .A(_0502_),
    .B(_3914_));
 sg13g2_nor3_1 _8951_ (.A(_0507_),
    .B(_0001_),
    .C(_3907_),
    .Y(_3916_));
 sg13g2_a21o_1 _8952_ (.A2(_3915_),
    .A1(_3913_),
    .B1(_3916_),
    .X(_3917_));
 sg13g2_xor2_1 _8953_ (.B(_3917_),
    .A(_3874_),
    .X(_3918_));
 sg13g2_nor2_1 _8954_ (.A(_3918_),
    .B(_4207_),
    .Y(_3919_));
 sg13g2_buf_1 _8955_ (.A(_3919_),
    .X(_3920_));
 sg13g2_inv_1 _8956_ (.Y(_3921_),
    .A(_3920_));
 sg13g2_buf_1 _8957_ (.A(_3921_),
    .X(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ));
 sg13g2_inv_1 _8958_ (.Y(_3922_),
    .A(_3918_));
 sg13g2_nor2_1 _8959_ (.A(_3922_),
    .B(_4207_),
    .Y(_3923_));
 sg13g2_buf_1 _8960_ (.A(_3923_),
    .X(_3924_));
 sg13g2_inv_1 _8961_ (.Y(_3925_),
    .A(net22));
 sg13g2_buf_1 _8962_ (.A(_4207_),
    .X(_3926_));
 sg13g2_a22oi_1 _8963_ (.Y(_3927_),
    .B1(_0743_),
    .B2(net23),
    .A2(_3926_),
    .A1(_0552_));
 sg13g2_o21ai_1 _8964_ (.B1(_3927_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[0] ),
    .A1(_0575_),
    .A2(_3925_));
 sg13g2_xor2_1 _8965_ (.B(_3906_),
    .A(_3910_),
    .X(_3928_));
 sg13g2_xor2_1 _8966_ (.B(_3899_),
    .A(_3904_),
    .X(_3929_));
 sg13g2_inv_1 _8967_ (.Y(_3930_),
    .A(_3929_));
 sg13g2_xor2_1 _8968_ (.B(_3885_),
    .A(_0006_),
    .X(_3931_));
 sg13g2_nor2_1 _8969_ (.A(_0574_),
    .B(_0549_),
    .Y(_3932_));
 sg13g2_nand3_1 _8970_ (.B(_0559_),
    .C(_3932_),
    .A(_3931_),
    .Y(_3933_));
 sg13g2_nand2_1 _8971_ (.Y(_3934_),
    .A(_3889_),
    .B(_3888_));
 sg13g2_nor2b_1 _8972_ (.A(_3890_),
    .B_N(_3934_),
    .Y(_3935_));
 sg13g2_nor2_1 _8973_ (.A(_3933_),
    .B(_3935_),
    .Y(_3936_));
 sg13g2_xnor2_1 _8974_ (.Y(_3937_),
    .A(_3892_),
    .B(_3891_));
 sg13g2_xor2_1 _8975_ (.B(_3898_),
    .A(_3880_),
    .X(_3938_));
 sg13g2_xor2_1 _8976_ (.B(_3893_),
    .A(_3938_),
    .X(_3939_));
 sg13g2_nor2_1 _8977_ (.A(_3937_),
    .B(_3939_),
    .Y(_3940_));
 sg13g2_nand3_1 _8978_ (.B(_3936_),
    .C(_3940_),
    .A(_3930_),
    .Y(_3941_));
 sg13g2_xor2_1 _8979_ (.B(_3913_),
    .A(_3915_),
    .X(_3942_));
 sg13g2_nor3_1 _8980_ (.A(_3928_),
    .B(_3941_),
    .C(_3942_),
    .Y(_3943_));
 sg13g2_and3_1 _8981_ (.X(\main.demo._t___pip_58_1_0___stage___block_3_cx[10] ),
    .A(_4206_),
    .B(_3918_),
    .C(_3943_));
 sg13g2_xor2_1 _8982_ (.B(_0549_),
    .A(_0574_),
    .X(_3944_));
 sg13g2_buf_1 _8983_ (.A(net22),
    .X(_3945_));
 sg13g2_a22oi_1 _8984_ (.Y(_3946_),
    .B1(_3944_),
    .B2(net20),
    .A2(net24),
    .A1(net74));
 sg13g2_o21ai_1 _8985_ (.B1(_3946_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[1] ),
    .A1(_0017_),
    .A2(net16));
 sg13g2_xnor2_1 _8986_ (.Y(_3947_),
    .A(_0558_),
    .B(_3932_));
 sg13g2_a22oi_1 _8987_ (.Y(_3948_),
    .B1(_3947_),
    .B2(_3945_),
    .A2(net24),
    .A1(_0563_));
 sg13g2_o21ai_1 _8988_ (.B1(_3948_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[2] ),
    .A1(_0559_),
    .A2(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ));
 sg13g2_xnor2_1 _8989_ (.Y(_3949_),
    .A(_0011_),
    .B(_4167_));
 sg13g2_nor3_1 _8990_ (.A(_0549_),
    .B(_0558_),
    .C(_0743_),
    .Y(_3950_));
 sg13g2_xor2_1 _8991_ (.B(_3931_),
    .A(_3950_),
    .X(_3951_));
 sg13g2_a22oi_1 _8992_ (.Y(_3952_),
    .B1(_3951_),
    .B2(_3945_),
    .A2(_3949_),
    .A1(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ));
 sg13g2_o21ai_1 _8993_ (.B1(_3952_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[3] ),
    .A1(net16),
    .A2(_3931_));
 sg13g2_inv_1 _8994_ (.Y(_3953_),
    .A(_3935_));
 sg13g2_nand2_1 _8995_ (.Y(_3954_),
    .A(_4174_),
    .B(_4169_));
 sg13g2_nand2_1 _8996_ (.Y(_3955_),
    .A(_4176_),
    .B(_3954_));
 sg13g2_inv_1 _8997_ (.Y(_3956_),
    .A(_3955_));
 sg13g2_xor2_1 _8998_ (.B(_3935_),
    .A(_3933_),
    .X(_3957_));
 sg13g2_a22oi_1 _8999_ (.Y(_3958_),
    .B1(_3957_),
    .B2(net20),
    .A2(_3956_),
    .A1(net25));
 sg13g2_o21ai_1 _9000_ (.B1(_3958_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[4] ),
    .A1(net16),
    .A2(_3953_));
 sg13g2_inv_1 _9001_ (.Y(_3959_),
    .A(_3937_));
 sg13g2_xnor2_1 _9002_ (.Y(_3960_),
    .A(_4175_),
    .B(_4183_));
 sg13g2_buf_1 _9003_ (.A(_3960_),
    .X(_3961_));
 sg13g2_xnor2_1 _9004_ (.Y(_3962_),
    .A(_3936_),
    .B(_3937_));
 sg13g2_a22oi_1 _9005_ (.Y(_3963_),
    .B1(_3962_),
    .B2(net20),
    .A2(_3961_),
    .A1(net25));
 sg13g2_o21ai_1 _9006_ (.B1(_3963_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[5] ),
    .A1(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .A2(_3959_));
 sg13g2_inv_1 _9007_ (.Y(_3964_),
    .A(_3939_));
 sg13g2_nand2b_1 _9008_ (.Y(_3965_),
    .B(_4189_),
    .A_N(_4190_));
 sg13g2_xnor2_1 _9009_ (.Y(_3966_),
    .A(_3965_),
    .B(_4185_));
 sg13g2_nand2_1 _9010_ (.Y(_3967_),
    .A(_3959_),
    .B(_3936_));
 sg13g2_xor2_1 _9011_ (.B(_3967_),
    .A(_3939_),
    .X(_3968_));
 sg13g2_a22oi_1 _9012_ (.Y(_3969_),
    .B1(_3968_),
    .B2(net20),
    .A2(_3966_),
    .A1(net25));
 sg13g2_o21ai_1 _9013_ (.B1(_3969_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[6] ),
    .A1(net16),
    .A2(_3964_));
 sg13g2_xor2_1 _9014_ (.B(_4191_),
    .A(_4192_),
    .X(_3970_));
 sg13g2_nand4_1 _9015_ (.B(_3931_),
    .C(_3953_),
    .A(_3940_),
    .Y(_3971_),
    .D(_3950_));
 sg13g2_xnor2_1 _9016_ (.Y(_3972_),
    .A(_3930_),
    .B(_3971_));
 sg13g2_a22oi_1 _9017_ (.Y(_3973_),
    .B1(_3972_),
    .B2(net22),
    .A2(_3970_),
    .A1(net25));
 sg13g2_o21ai_1 _9018_ (.B1(_3973_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[7] ),
    .A1(net16),
    .A2(_3930_));
 sg13g2_inv_1 _9019_ (.Y(_3974_),
    .A(_3928_));
 sg13g2_xor2_1 _9020_ (.B(_4194_),
    .A(_4197_),
    .X(_3975_));
 sg13g2_xor2_1 _9021_ (.B(_3928_),
    .A(_3941_),
    .X(_3976_));
 sg13g2_a22oi_1 _9022_ (.Y(_3977_),
    .B1(_3976_),
    .B2(net22),
    .A2(_3975_),
    .A1(net24));
 sg13g2_o21ai_1 _9023_ (.B1(_3977_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[8] ),
    .A1(_3921_),
    .A2(_3974_));
 sg13g2_nand2b_1 _9024_ (.Y(_3978_),
    .B(_4201_),
    .A_N(_4145_));
 sg13g2_xnor2_1 _9025_ (.Y(_3979_),
    .A(_3978_),
    .B(_4199_));
 sg13g2_nor3_1 _9026_ (.A(_3929_),
    .B(_3971_),
    .C(_3928_),
    .Y(_3980_));
 sg13g2_xnor2_1 _9027_ (.Y(_3981_),
    .A(_3980_),
    .B(_3942_));
 sg13g2_a22oi_1 _9028_ (.Y(_3982_),
    .B1(net22),
    .B2(_3981_),
    .A2(_3942_),
    .A1(net23));
 sg13g2_o21ai_1 _9029_ (.B1(_3982_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[9] ),
    .A1(_4206_),
    .A2(_3979_));
 sg13g2_a22oi_1 _9030_ (.Y(_3983_),
    .B1(_0552_),
    .B2(net22),
    .A2(net24),
    .A1(_0574_));
 sg13g2_o21ai_1 _9031_ (.B1(_3983_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[0] ),
    .A1(_0013_),
    .A2(net16));
 sg13g2_inv_1 _9032_ (.Y(_3984_),
    .A(_0015_));
 sg13g2_nor2_1 _9033_ (.A(net74),
    .B(_0552_),
    .Y(_3985_));
 sg13g2_inv_1 _9034_ (.Y(_3986_),
    .A(_3985_));
 sg13g2_nor3_1 _9035_ (.A(_3984_),
    .B(_3986_),
    .C(_3949_),
    .Y(_3987_));
 sg13g2_nand2_1 _9036_ (.Y(_3988_),
    .A(_3955_),
    .B(_3987_));
 sg13g2_nor4_1 _9037_ (.A(_3961_),
    .B(_3966_),
    .C(_3988_),
    .D(_3970_),
    .Y(_3989_));
 sg13g2_inv_1 _9038_ (.Y(_3990_),
    .A(_3989_));
 sg13g2_nor2_1 _9039_ (.A(_3975_),
    .B(_3990_),
    .Y(_3991_));
 sg13g2_nand2_1 _9040_ (.Y(_3992_),
    .A(_3979_),
    .B(_3991_));
 sg13g2_nand2b_1 _9041_ (.Y(_3993_),
    .B(_3922_),
    .A_N(_3943_));
 sg13g2_a21oi_1 _9042_ (.A1(_3918_),
    .A2(_3943_),
    .Y(_3994_),
    .B1(_4206_));
 sg13g2_a22oi_1 _9043_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[10] ),
    .B1(_3993_),
    .B2(_3994_),
    .A2(_3992_),
    .A1(net20));
 sg13g2_nand2_1 _9044_ (.Y(_3995_),
    .A(net74),
    .B(_0552_));
 sg13g2_nand3_1 _9045_ (.B(_3986_),
    .C(_3995_),
    .A(net22),
    .Y(_3996_));
 sg13g2_nand2_1 _9046_ (.Y(_3997_),
    .A(net25),
    .B(_3944_));
 sg13g2_nand2b_1 _9047_ (.Y(_3998_),
    .B(_3920_),
    .A_N(_0014_));
 sg13g2_nand3_1 _9048_ (.B(_3997_),
    .C(_3998_),
    .A(_3996_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[1] ));
 sg13g2_xnor2_1 _9049_ (.Y(_3999_),
    .A(_3984_),
    .B(_3985_));
 sg13g2_a22oi_1 _9050_ (.Y(_4000_),
    .B1(_3999_),
    .B2(net22),
    .A2(_3947_),
    .A1(net24));
 sg13g2_o21ai_1 _9051_ (.B1(_4000_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[2] ),
    .A1(_0015_),
    .A2(net16));
 sg13g2_a22oi_1 _9052_ (.Y(_4001_),
    .B1(_3949_),
    .B2(net23),
    .A2(_3951_),
    .A1(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ));
 sg13g2_inv_1 _9053_ (.Y(_4002_),
    .A(_0589_));
 sg13g2_nand2_1 _9054_ (.Y(_4003_),
    .A(_3949_),
    .B(_4002_));
 sg13g2_nor2_1 _9055_ (.A(_4002_),
    .B(_3949_),
    .Y(_4004_));
 sg13g2_inv_1 _9056_ (.Y(_4005_),
    .A(_4004_));
 sg13g2_nand3_1 _9057_ (.B(_4003_),
    .C(_4005_),
    .A(net20),
    .Y(_4006_));
 sg13g2_nand2_1 _9058_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[3] ),
    .A(_4001_),
    .B(_4006_));
 sg13g2_xnor2_1 _9059_ (.Y(_4007_),
    .A(_3987_),
    .B(_3955_));
 sg13g2_a22oi_1 _9060_ (.Y(_4008_),
    .B1(_3956_),
    .B2(net23),
    .A2(_3957_),
    .A1(net24));
 sg13g2_o21ai_1 _9061_ (.B1(_4008_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[4] ),
    .A1(_3925_),
    .A2(_4007_));
 sg13g2_a22oi_1 _9062_ (.Y(_4009_),
    .B1(_3961_),
    .B2(net23),
    .A2(_3962_),
    .A1(net25));
 sg13g2_nor2_1 _9063_ (.A(_4005_),
    .B(_3956_),
    .Y(_4010_));
 sg13g2_inv_1 _9064_ (.Y(_4011_),
    .A(_4010_));
 sg13g2_nor2_1 _9065_ (.A(_4011_),
    .B(_3961_),
    .Y(_4012_));
 sg13g2_inv_1 _9066_ (.Y(_4013_),
    .A(_4012_));
 sg13g2_nand2_1 _9067_ (.Y(_4014_),
    .A(_3961_),
    .B(_4011_));
 sg13g2_nand3_1 _9068_ (.B(_4013_),
    .C(_4014_),
    .A(net20),
    .Y(_4015_));
 sg13g2_nand2_1 _9069_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[5] ),
    .A(_4009_),
    .B(_4015_));
 sg13g2_nor2_1 _9070_ (.A(_3988_),
    .B(_3961_),
    .Y(_4016_));
 sg13g2_xor2_1 _9071_ (.B(_3966_),
    .A(_4016_),
    .X(_4017_));
 sg13g2_a22oi_1 _9072_ (.Y(_4018_),
    .B1(_3966_),
    .B2(net23),
    .A2(_3968_),
    .A1(net24));
 sg13g2_o21ai_1 _9073_ (.B1(_4018_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[6] ),
    .A1(_3925_),
    .A2(_4017_));
 sg13g2_a22oi_1 _9074_ (.Y(_4019_),
    .B1(_3970_),
    .B2(net23),
    .A2(_3972_),
    .A1(net25));
 sg13g2_nor2_1 _9075_ (.A(_4013_),
    .B(_3966_),
    .Y(_4020_));
 sg13g2_nand2b_1 _9076_ (.Y(_4021_),
    .B(_3970_),
    .A_N(_4020_));
 sg13g2_nand2b_1 _9077_ (.Y(_4022_),
    .B(_4020_),
    .A_N(_3970_));
 sg13g2_nand3_1 _9078_ (.B(_4021_),
    .C(_4022_),
    .A(net20),
    .Y(_4023_));
 sg13g2_nand2_1 _9079_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[7] ),
    .A(_4019_),
    .B(_4023_));
 sg13g2_nand2_1 _9080_ (.Y(_4024_),
    .A(_3990_),
    .B(_3975_));
 sg13g2_nand2b_1 _9081_ (.Y(_4025_),
    .B(_4024_),
    .A_N(_3991_));
 sg13g2_a22oi_1 _9082_ (.Y(_4026_),
    .B1(_3975_),
    .B2(net23),
    .A2(_3976_),
    .A1(net24));
 sg13g2_o21ai_1 _9083_ (.B1(_4026_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[8] ),
    .A1(_3925_),
    .A2(_4025_));
 sg13g2_nor2_1 _9084_ (.A(_4022_),
    .B(_3975_),
    .Y(_4027_));
 sg13g2_xor2_1 _9085_ (.B(_3979_),
    .A(_4027_),
    .X(_4028_));
 sg13g2_a22oi_1 _9086_ (.Y(_4029_),
    .B1(_4028_),
    .B2(_3924_),
    .A2(_3981_),
    .A1(_3926_));
 sg13g2_o21ai_1 _9087_ (.B1(_4029_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[9] ),
    .A1(_3921_),
    .A2(_3979_));
 sg13g2_nand2_1 _9088_ (.Y(\main.demo._t___pip_58_1_3___block_87_atten_l[0] ),
    .A(net53),
    .B(_0064_));
 sg13g2_inv_1 _9089_ (.Y(\main.demo._t___pip_58_1_3___block_87_atten_h[0] ),
    .A(\main.demo._t___pip_58_1_3___block_87_atten_l[0] ));
 sg13g2_inv_1 _9090_ (.Y(_4030_),
    .A(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ));
 sg13g2_nor2_1 _9091_ (.A(_4030_),
    .B(\main.demo._t___pip_58_1_3___block_87_atten_h[0] ),
    .Y(\main.demo._t___pip_58_1_3___block_87_atten_h[2] ));
 sg13g2_a21oi_1 _9092_ (.A1(_4030_),
    .A2(_0064_),
    .Y(\main.demo._t___pip_58_1_3___block_87_atten_h[1] ),
    .B1(\main.demo._t___pip_58_1_3___block_87_atten_h[2] ));
 sg13g2_nor2_1 _9093_ (.A(_0386_),
    .B(net33),
    .Y(\main.demo.vga._d_active ));
 sg13g2_dfrbp_1 _9094_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net92),
    .D(net25),
    .Q_N(_4562_),
    .Q(_0070_));
 sg13g2_dfrbp_1 _9095_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net93),
    .D(net16),
    .Q_N(_4563_),
    .Q(_0071_));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _9094__92 (.L_HI(net92));
 sg13g2_buf_1 _9098_ (.A(net78),
    .X(uio_oe[0]));
 sg13g2_buf_1 _9099_ (.A(net79),
    .X(uio_oe[1]));
 sg13g2_buf_1 _9100_ (.A(net80),
    .X(uio_oe[2]));
 sg13g2_buf_1 _9101_ (.A(net81),
    .X(uio_oe[3]));
 sg13g2_buf_1 _9102_ (.A(net82),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9103_ (.A(net83),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9104_ (.A(net84),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9105_ (.A(net94),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9106_ (.A(net85),
    .X(uio_out[0]));
 sg13g2_buf_1 _9107_ (.A(net86),
    .X(uio_out[1]));
 sg13g2_buf_1 _9108_ (.A(net87),
    .X(uio_out[2]));
 sg13g2_buf_1 _9109_ (.A(net88),
    .X(uio_out[3]));
 sg13g2_buf_1 _9110_ (.A(net89),
    .X(uio_out[4]));
 sg13g2_buf_1 _9111_ (.A(net90),
    .X(uio_out[5]));
 sg13g2_buf_1 _9112_ (.A(net91),
    .X(uio_out[6]));
 sg13g2_buf_1 _9113_ (.A(\main.demo._q_prev_vs ),
    .X(net6));
 sg13g2_dfrbp_1 \main._q_uio_o[7]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net95),
    .D(\main._w_demo_audio1 ),
    .Q_N(_4561_),
    .Q(net2));
 sg13g2_dfrbp_1 \main._q_uo[0]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net96),
    .D(_0072_),
    .Q_N(_4560_),
    .Q(net3));
 sg13g2_dfrbp_1 \main._q_uo[1]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net97),
    .D(_0073_),
    .Q_N(_4559_),
    .Q(net4));
 sg13g2_dfrbp_1 \main._q_uo[2]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net98),
    .D(_0074_),
    .Q_N(_4564_),
    .Q(net5));
 sg13g2_dfrbp_1 \main._q_uo[3]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net99),
    .D(\main._w_demo_video_vs ),
    .Q_N(_4558_),
    .Q(\main.demo._q_prev_vs ));
 sg13g2_dfrbp_1 \main._q_uo[4]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net100),
    .D(_0075_),
    .Q_N(_4557_),
    .Q(net7));
 sg13g2_dfrbp_1 \main._q_uo[5]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net101),
    .D(_0076_),
    .Q_N(_4556_),
    .Q(net8));
 sg13g2_dfrbp_1 \main._q_uo[6]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net102),
    .D(_0077_),
    .Q_N(_4565_),
    .Q(net9));
 sg13g2_dfrbp_1 \main._q_uo[7]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net103),
    .D(\main._w_demo_video_hs ),
    .Q_N(_4566_),
    .Q(net10));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[0]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net104),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[0] ),
    .Q_N(_4567_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[10]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net105),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[10] ),
    .Q_N(_4568_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[1]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net106),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[1] ),
    .Q_N(_4569_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[2]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net107),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[2] ),
    .Q_N(_4570_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[3]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net108),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[3] ),
    .Q_N(_4571_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[4]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net109),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[4] ),
    .Q_N(_4572_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[5]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net110),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[5] ),
    .Q_N(_4573_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[6]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net111),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[6] ),
    .Q_N(_4574_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[7]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net112),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[7] ),
    .Q_N(_4575_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[8]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net113),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[8] ),
    .Q_N(_4576_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cx[9]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[9] ),
    .Q_N(_4577_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[0]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net115),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[0] ),
    .Q_N(_4578_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[10]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net116),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[10] ),
    .Q_N(_4579_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[10] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[1]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net117),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[1] ),
    .Q_N(_4580_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[2]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net118),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[2] ),
    .Q_N(_4581_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[3]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net119),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[3] ),
    .Q_N(_4582_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[4]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net120),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[4] ),
    .Q_N(_4583_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[5]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net121),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[5] ),
    .Q_N(_4584_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[6]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net122),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[6] ),
    .Q_N(_4585_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[7]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net123),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[7] ),
    .Q_N(_4586_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[8]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net124),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[8] ),
    .Q_N(_4587_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_1___stage___block_3_cy[9]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net125),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[9] ),
    .Q_N(_4588_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_a[1]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net126),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ),
    .Q_N(_4589_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_a[2]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net127),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .Q_N(_4590_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_a[3]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net128),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ),
    .Q_N(_4591_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_a[4]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net129),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[4] ),
    .Q_N(_4592_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_a[6]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net130),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[6] ),
    .Q_N(_4593_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_a[7]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net131),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[7] ),
    .Q_N(_4594_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[7] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[0]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net132),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[0] ),
    .Q_N(_4595_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[10]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net133),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[10] ),
    .Q_N(_0063_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[10] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[1]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net134),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[1] ),
    .Q_N(_4596_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[2]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net135),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[2] ),
    .Q_N(_4597_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[3]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net136),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[3] ),
    .Q_N(_0049_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[4]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net137),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[4] ),
    .Q_N(_0051_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[5]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net138),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[5] ),
    .Q_N(_0050_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[6]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net139),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[6] ),
    .Q_N(_0048_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[7]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net140),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[7] ),
    .Q_N(_0046_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[8]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net141),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[8] ),
    .Q_N(_0054_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cx[9]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net142),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[9] ),
    .Q_N(_0052_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[0]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net143),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[0] ),
    .Q_N(_4598_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[10]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net144),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[10] ),
    .Q_N(_0053_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[10] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[1]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net145),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[1] ),
    .Q_N(_4599_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[2]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net146),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[2] ),
    .Q_N(_4600_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[3]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net147),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[3] ),
    .Q_N(_0047_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[4]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net148),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[4] ),
    .Q_N(_0062_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[5]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net149),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[5] ),
    .Q_N(_0061_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[6]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net150),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[6] ),
    .Q_N(_0060_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[7]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net151),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[7] ),
    .Q_N(_0059_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[8]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net152),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[8] ),
    .Q_N(_0058_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_2___stage___block_3_cy[9]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net153),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[9] ),
    .Q_N(_0057_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_a[1]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net154),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[1] ),
    .Q_N(_0030_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_a[2]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net155),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[2] ),
    .Q_N(_0029_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_a[3]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net156),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[3] ),
    .Q_N(_0028_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_a[4]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net157),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[4] ),
    .Q_N(_0027_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_a[5]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net158),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[5] ),
    .Q_N(_0032_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_a[6]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net159),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[6] ),
    .Q_N(_0031_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_a[7]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net160),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[7] ),
    .Q_N(_4601_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[7] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[0]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net161),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[0] ),
    .Q_N(_0022_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[10]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net162),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[10] ),
    .Q_N(_4602_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[1]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net163),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[1] ),
    .Q_N(_0021_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[2]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net164),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[2] ),
    .Q_N(_4603_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[3]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net165),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[3] ),
    .Q_N(_4604_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[4]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net166),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[4] ),
    .Q_N(_0020_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[5]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net167),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[5] ),
    .Q_N(_4605_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[6]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net168),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[6] ),
    .Q_N(_4606_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[7]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net169),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[7] ),
    .Q_N(_0064_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[8]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net170),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[8] ),
    .Q_N(_0018_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[8] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_3___stage___block_3_cx[9]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net171),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[9] ),
    .Q_N(_4607_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_68_frag[0]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net172),
    .D(\main.demo._t___block_68_frag[0] ),
    .Q_N(_4608_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_68_frag[1]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net173),
    .D(\main.demo._t___block_68_frag[1] ),
    .Q_N(_4609_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_68_frag[2]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net174),
    .D(\main.demo._t___block_68_frag[2] ),
    .Q_N(_4610_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_68_frag[3]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net175),
    .D(\main.demo._t___block_68_frag[3] ),
    .Q_N(_4611_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_68_frag[4]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net176),
    .D(\main.demo._t___block_68_frag[4] ),
    .Q_N(_4612_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_68_frag[5]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net177),
    .D(\main.demo._t___block_68_frag[5] ),
    .Q_N(_4613_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_87_atten_h[0]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net178),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_h[0] ),
    .Q_N(_4614_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_87_atten_h[1]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net179),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_h[1] ),
    .Q_N(_4615_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_87_atten_h[2]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net180),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_h[2] ),
    .Q_N(_4616_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_87_atten_l[0]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net181),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_l[0] ),
    .Q_N(_4617_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_l[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___block_87_atten_l[1]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net182),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ),
    .Q_N(_4618_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___stage___block_3_cx[1]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net183),
    .D(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .Q_N(_4619_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___stage___block_3_cx[2]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net184),
    .D(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .Q_N(_4620_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___stage___block_3_cx[3]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net185),
    .D(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ),
    .Q_N(_4621_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___stage___block_3_cx[4]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net186),
    .D(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .Q_N(_4622_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___stage___block_3_cx[5]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net187),
    .D(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ),
    .Q_N(_4623_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___stage___block_3_cx[6]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net188),
    .D(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .Q_N(_4624_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_58_1_4___stage___block_3_cx[9]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net189),
    .D(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .Q_N(_4555_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 \main.demo._q_effect[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net190),
    .D(_0078_),
    .Q_N(_0069_),
    .Q(\main.demo._q_effect[0] ));
 sg13g2_dfrbp_1 \main.demo._q_effect[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net191),
    .D(_0079_),
    .Q_N(_4554_),
    .Q(\main.demo._q_effect[1] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[0]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net192),
    .D(_0080_),
    .Q_N(_4553_),
    .Q(\main.demo._q_frame[0] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[10]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net193),
    .D(_0081_),
    .Q_N(_4552_),
    .Q(\main.demo._q_frame[10] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[11]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net194),
    .D(_0082_),
    .Q_N(_4551_),
    .Q(\main.demo._q_frame[11] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[12]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net195),
    .D(_0083_),
    .Q_N(_4550_),
    .Q(\main.demo._q_frame[12] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[13]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net196),
    .D(_0084_),
    .Q_N(_4549_),
    .Q(\main.demo._q_frame[13] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[14]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net197),
    .D(_0085_),
    .Q_N(_4548_),
    .Q(\main.demo._q_frame[14] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[1]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net198),
    .D(_0086_),
    .Q_N(_4547_),
    .Q(\main.demo._q_frame[1] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[2]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net199),
    .D(_0087_),
    .Q_N(_4546_),
    .Q(\main.demo._q_frame[2] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[3]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net200),
    .D(_0088_),
    .Q_N(_4545_),
    .Q(\main.demo._q_frame[3] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[4]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net201),
    .D(_0089_),
    .Q_N(_4544_),
    .Q(\main.demo._q_frame[4] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[5]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net202),
    .D(_0090_),
    .Q_N(_4543_),
    .Q(\main.demo._q_frame[5] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[6]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net203),
    .D(_0091_),
    .Q_N(_4542_),
    .Q(\main.demo._q_frame[6] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[7]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net204),
    .D(_0092_),
    .Q_N(_4541_),
    .Q(\main.demo._q_frame[7] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[8]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net205),
    .D(_0093_),
    .Q_N(_4540_),
    .Q(\main.demo._q_frame[8] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[9]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net206),
    .D(_0094_),
    .Q_N(_4539_),
    .Q(\main.demo._q_frame[9] ));
 sg13g2_dfrbp_1 \main.demo._q_go$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net207),
    .D(_0095_),
    .Q_N(_4625_),
    .Q(\main.demo._q_go ));
 sg13g2_dfrbp_1 \main.demo._q_prev_b[0]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net208),
    .D(\main.demo._d_prev_b[0] ),
    .Q_N(_4626_),
    .Q(\main.demo._d_prev_b[2] ));
 sg13g2_dfrbp_1 \main.demo._q_prev_b[1]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net209),
    .D(\main.demo._d_prev_b[1] ),
    .Q_N(_4627_),
    .Q(\main.demo._d_prev_b[3] ));
 sg13g2_dfrbp_1 \main.demo._q_prev_b[2]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net210),
    .D(\main.demo._d_prev_b[2] ),
    .Q_N(_4628_),
    .Q(\main.demo._d_prev_b[4] ));
 sg13g2_dfrbp_1 \main.demo._q_prev_b[3]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net211),
    .D(\main.demo._d_prev_b[3] ),
    .Q_N(_4629_),
    .Q(\main.demo._d_prev_b[5] ));
 sg13g2_dfrbp_1 \main.demo._q_prev_b[4]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net212),
    .D(\main.demo._d_prev_b[4] ),
    .Q_N(_4630_),
    .Q(\main.demo._d_prev_b[6] ));
 sg13g2_dfrbp_1 \main.demo._q_prev_b[5]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net213),
    .D(\main.demo._d_prev_b[5] ),
    .Q_N(_4631_),
    .Q(\main.demo._d_prev_b[7] ));
 sg13g2_dfrbp_1 \main.demo._q_prev_b[6]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net214),
    .D(\main.demo._d_prev_b[6] ),
    .Q_N(_4632_),
    .Q(\main.demo._q_prev_b[6] ));
 sg13g2_dfrbp_1 \main.demo._q_prev_b[7]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net215),
    .D(\main.demo._d_prev_b[7] ),
    .Q_N(_4538_),
    .Q(\main.demo._q_prev_b[7] ));
 sg13g2_dfrbp_1 \main.demo._q_rot_en$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net216),
    .D(_0096_),
    .Q_N(_0000_),
    .Q(\main.demo._q_rot_en ));
 sg13g2_dfrbp_1 \main.demo._q_speed[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net217),
    .D(_0097_),
    .Q_N(_4537_),
    .Q(\main.demo._q_speed[0] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[10]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net218),
    .D(_0098_),
    .Q_N(_0019_),
    .Q(\main.demo._q_speed[10] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[11]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net219),
    .D(_0099_),
    .Q_N(_4536_),
    .Q(\main.demo._q_speed[11] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[12]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net220),
    .D(_0100_),
    .Q_N(_4535_),
    .Q(\main.demo._q_speed[12] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[13]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net221),
    .D(_0101_),
    .Q_N(_4534_),
    .Q(\main.demo._q_speed[13] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[14]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net222),
    .D(_0102_),
    .Q_N(_4533_),
    .Q(\main.demo._q_speed[14] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[15]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net223),
    .D(_0103_),
    .Q_N(_4532_),
    .Q(\main.demo._q_speed[15] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[1]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net224),
    .D(_0104_),
    .Q_N(_0026_),
    .Q(\main.demo._q_speed[1] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[2]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net225),
    .D(_0105_),
    .Q_N(_0025_),
    .Q(\main.demo._q_speed[2] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[3]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net226),
    .D(_0106_),
    .Q_N(_0024_),
    .Q(\main.demo._q_speed[3] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[4]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net227),
    .D(_0107_),
    .Q_N(_0023_),
    .Q(\main.demo._q_speed[4] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net228),
    .D(_0108_),
    .Q_N(_0035_),
    .Q(\main.demo._q_speed[5] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net229),
    .D(_0109_),
    .Q_N(_0034_),
    .Q(\main.demo._q_speed[6] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[7]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net230),
    .D(_0110_),
    .Q_N(_0033_),
    .Q(\main.demo._q_speed[7] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[8]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net231),
    .D(_0111_),
    .Q_N(_4531_),
    .Q(\main.demo._q_speed[8] ));
 sg13g2_dfrbp_1 \main.demo._q_speed[9]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net232),
    .D(_0112_),
    .Q_N(_4530_),
    .Q(\main.demo._q_speed[9] ));
 sg13g2_dfrbp_1 \main.demo._q_th[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net233),
    .D(_0113_),
    .Q_N(_0067_),
    .Q(\main.demo._q_th[0] ));
 sg13g2_dfrbp_1 \main.demo._q_th[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net234),
    .D(_0114_),
    .Q_N(_4529_),
    .Q(\main.demo._q_th[1] ));
 sg13g2_dfrbp_1 \main.demo._q_th[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net235),
    .D(_0115_),
    .Q_N(_4528_),
    .Q(\main.demo._q_th[2] ));
 sg13g2_dfrbp_1 \main.demo._q_th[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net236),
    .D(_0116_),
    .Q_N(_4527_),
    .Q(\main.demo._q_th[3] ));
 sg13g2_dfrbp_1 \main.demo._q_th[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net237),
    .D(_0117_),
    .Q_N(_4526_),
    .Q(\main.demo._q_th[4] ));
 sg13g2_dfrbp_1 \main.demo._q_th[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net238),
    .D(_0118_),
    .Q_N(_0037_),
    .Q(\main.demo._q_th[5] ));
 sg13g2_dfrbp_1 \main.demo._q_th[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net239),
    .D(_0119_),
    .Q_N(_0036_),
    .Q(\main.demo._q_th[6] ));
 sg13g2_dfrbp_1 \main.demo._q_th[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net240),
    .D(_0120_),
    .Q_N(_4525_),
    .Q(\main.demo._q_th[7] ));
 sg13g2_dfrbp_1 \main.demo._q_th[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net241),
    .D(_0121_),
    .Q_N(_4633_),
    .Q(\main.demo._q_th[8] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_active$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net242),
    .D(\main.demo.vga._d_active ),
    .Q_N(_4524_),
    .Q(\main.demo._w_vga_active ));
 sg13g2_dfrbp_1 \main.demo.vga._q_active_h$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net243),
    .D(_0122_),
    .Q_N(_4523_),
    .Q(\main.demo.vga._q_active_h ));
 sg13g2_dfrbp_1 \main.demo.vga._q_active_v$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net244),
    .D(_0123_),
    .Q_N(_4522_),
    .Q(\main.demo.vga._q_active_v ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_hs$_SDFFE_PP0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net245),
    .D(_0124_),
    .Q_N(_4521_),
    .Q(\main._w_demo_video_hs ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_vs$_SDFFE_PP0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net246),
    .D(_0125_),
    .Q_N(_4520_),
    .Q(\main._w_demo_video_vs ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[0]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net247),
    .D(_0126_),
    .Q_N(_0016_),
    .Q(\main.demo._t___stage___block_3_x[0] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[10]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net248),
    .D(_0127_),
    .Q_N(_4519_),
    .Q(\main.demo._w_vga_vga_x[10] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[1]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net249),
    .D(_0128_),
    .Q_N(_0017_),
    .Q(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[2]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net250),
    .D(_0129_),
    .Q_N(_4518_),
    .Q(\main.demo._t___stage___block_3_x[2] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[3]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net251),
    .D(_0130_),
    .Q_N(_0006_),
    .Q(\main.demo._w_vga_vga_x[3] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[4]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net252),
    .D(_0131_),
    .Q_N(_0005_),
    .Q(\main.demo._w_vga_vga_x[4] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[5]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net253),
    .D(_0132_),
    .Q_N(_0004_),
    .Q(\main.demo._w_vga_vga_x[5] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[6]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net254),
    .D(_0133_),
    .Q_N(_0003_),
    .Q(\main.demo._w_vga_vga_x[6] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[7]$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net255),
    .D(_0134_),
    .Q_N(_0002_),
    .Q(\main.demo._w_vga_vga_x[7] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[8]$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net256),
    .D(_0135_),
    .Q_N(_0001_),
    .Q(\main.demo._w_vga_vga_x[8] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_x[9]$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net257),
    .D(_0136_),
    .Q_N(_0065_),
    .Q(\main.demo._w_vga_vga_x[9] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[0]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net258),
    .D(_0137_),
    .Q_N(_0013_),
    .Q(\main.demo._t___stage___block_3_y[0] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[1]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net259),
    .D(_0138_),
    .Q_N(_0014_),
    .Q(\main.demo._t___stage___block_3_y[1] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[2]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net260),
    .D(_0139_),
    .Q_N(_0015_),
    .Q(\main.demo._t___stage___block_3_y[2] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[3]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net261),
    .D(_0140_),
    .Q_N(_0011_),
    .Q(\main.demo._w_vga_vga_y[3] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[4]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net262),
    .D(_0141_),
    .Q_N(_4517_),
    .Q(\main.demo._w_vga_vga_y[4] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[5]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net263),
    .D(_0142_),
    .Q_N(_0010_),
    .Q(\main.demo._w_vga_vga_y[5] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[6]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net264),
    .D(_0143_),
    .Q_N(_0009_),
    .Q(\main.demo._w_vga_vga_y[6] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[7]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net265),
    .D(_0144_),
    .Q_N(_0008_),
    .Q(\main.demo._w_vga_vga_y[7] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[8]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net266),
    .D(_0145_),
    .Q_N(_4516_),
    .Q(\main.demo._w_vga_vga_y[8] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[9]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net267),
    .D(_0146_),
    .Q_N(_0007_),
    .Q(\main.demo._w_vga_vga_y[10] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[0]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net268),
    .D(_0147_),
    .Q_N(_4515_),
    .Q(\main.demo.vga._q_xcount[0] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[10]$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net269),
    .D(_0148_),
    .Q_N(_4514_),
    .Q(\main.demo.vga._q_xcount[10] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[1]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net270),
    .D(_0149_),
    .Q_N(_4513_),
    .Q(\main.demo.vga._q_xcount[1] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[2]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net271),
    .D(_0150_),
    .Q_N(_4512_),
    .Q(\main.demo.vga._q_xcount[2] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[3]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net272),
    .D(_0151_),
    .Q_N(_4511_),
    .Q(\main.demo.vga._q_xcount[3] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[4]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net273),
    .D(_0152_),
    .Q_N(_4510_),
    .Q(\main.demo.vga._q_xcount[4] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[5]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net274),
    .D(_0153_),
    .Q_N(_4509_),
    .Q(\main.demo.vga._q_xcount[5] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[6]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net275),
    .D(_0154_),
    .Q_N(_4508_),
    .Q(\main.demo.vga._q_xcount[6] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[7]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net276),
    .D(_0155_),
    .Q_N(_4507_),
    .Q(\main.demo.vga._q_xcount[7] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[8]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net277),
    .D(_0156_),
    .Q_N(_4506_),
    .Q(\main.demo.vga._q_xcount[8] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[9]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net278),
    .D(_0157_),
    .Q_N(_4505_),
    .Q(\main.demo.vga._q_xcount[9] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net279),
    .D(_0158_),
    .Q_N(_4504_),
    .Q(\main.demo.vga._q_ycount[0] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net280),
    .D(_0159_),
    .Q_N(_4503_),
    .Q(\main.demo.vga._q_ycount[1] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net281),
    .D(_0160_),
    .Q_N(_4502_),
    .Q(\main.demo.vga._q_ycount[2] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net282),
    .D(_0161_),
    .Q_N(_4501_),
    .Q(\main.demo.vga._q_ycount[3] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net283),
    .D(_0162_),
    .Q_N(_4500_),
    .Q(\main.demo.vga._q_ycount[4] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net284),
    .D(_0163_),
    .Q_N(_4499_),
    .Q(\main.demo.vga._q_ycount[5] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net285),
    .D(_0164_),
    .Q_N(_4498_),
    .Q(\main.demo.vga._q_ycount[6] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net286),
    .D(_0165_),
    .Q_N(_4497_),
    .Q(\main.demo.vga._q_ycount[7] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net287),
    .D(_0166_),
    .Q_N(_4496_),
    .Q(\main.demo.vga._q_ycount[8] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net288),
    .D(_0167_),
    .Q_N(_4495_),
    .Q(\main.demo.vga._d_vblank ));
 sg13g2_dfrbp_1 \main.demo.zic._q_clock_count[0]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net289),
    .D(_0168_),
    .Q_N(_0066_),
    .Q(\main.demo.zic._q_clock_count[0] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_clock_count[1]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net290),
    .D(_0169_),
    .Q_N(_4494_),
    .Q(\main.demo.zic._q_clock_count[1] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_clock_count[2]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net291),
    .D(_0170_),
    .Q_N(_4493_),
    .Q(\main.demo.zic._q_clock_count[2] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_clock_count[3]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net292),
    .D(_0171_),
    .Q_N(_4492_),
    .Q(\main.demo.zic._q_clock_count[3] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_clock_count[4]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net293),
    .D(_0172_),
    .Q_N(_4491_),
    .Q(\main.demo.zic._q_clock_count[4] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_clock_count[5]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net294),
    .D(_0173_),
    .Q_N(_4490_),
    .Q(\main.demo.zic._q_clock_count[5] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_clock_count[6]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net295),
    .D(_0174_),
    .Q_N(_0041_),
    .Q(\main.demo.zic._q_clock_count[6] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_clock_count[7]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net296),
    .D(_0175_),
    .Q_N(_4489_),
    .Q(\main.demo.zic._q_clock_count[7] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_clock_count[8]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net297),
    .D(_0176_),
    .Q_N(_4488_),
    .Q(\main.demo.zic._q_clock_count[8] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_drum_inc[0]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net298),
    .D(_0177_),
    .Q_N(_4487_),
    .Q(\main.demo.zic._q_drum_inc[0] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_drum_inc[1]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net299),
    .D(_0178_),
    .Q_N(_4486_),
    .Q(\main.demo.zic._q_drum_inc[1] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_drum_inc[2]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net300),
    .D(_0179_),
    .Q_N(_4485_),
    .Q(\main.demo.zic._q_drum_inc[2] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_drum_inc[3]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net301),
    .D(_0180_),
    .Q_N(_4484_),
    .Q(\main.demo.zic._q_drum_inc[3] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_idx[0]$_SDFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net302),
    .D(_0181_),
    .Q_N(_0045_),
    .Q(\main.demo.zic._q_idx[0] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_idx[1]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net303),
    .D(_0182_),
    .Q_N(_4483_),
    .Q(\main.demo.zic._q_idx[1] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_idx[2]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net304),
    .D(_0183_),
    .Q_N(_4482_),
    .Q(\main.demo.zic._q_idx[2] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_idx[3]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net305),
    .D(_0184_),
    .Q_N(_4481_),
    .Q(\main.demo.zic._q_idx[3] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_idx[4]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net306),
    .D(_0185_),
    .Q_N(_0055_),
    .Q(\main.demo.zic._q_idx[4] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_idx[5]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net307),
    .D(_0186_),
    .Q_N(_4480_),
    .Q(\main.demo.zic._q_idx[5] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_idx[6]$_SDFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net308),
    .D(_0187_),
    .Q_N(_0044_),
    .Q(\main.demo.zic._q_idx[6] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net309),
    .D(_0188_),
    .Q_N(_4479_),
    .Q(\main.demo.zic._q_qpos[0] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net310),
    .D(_0189_),
    .Q_N(_4478_),
    .Q(\main.demo.zic._q_qpos[10] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net311),
    .D(_0190_),
    .Q_N(_4477_),
    .Q(\main.demo.zic._q_qpos[11] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net312),
    .D(_0191_),
    .Q_N(_4476_),
    .Q(\main.demo.zic._q_qpos[12] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net313),
    .D(_0192_),
    .Q_N(_4475_),
    .Q(\main.demo.zic._q_qpos[1] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net314),
    .D(_0193_),
    .Q_N(_4474_),
    .Q(\main.demo.zic._q_qpos[2] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net315),
    .D(_0194_),
    .Q_N(_4473_),
    .Q(\main.demo.zic._q_qpos[3] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net316),
    .D(_0195_),
    .Q_N(_4472_),
    .Q(\main.demo.zic._q_qpos[4] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net317),
    .D(_0196_),
    .Q_N(_4471_),
    .Q(\main.demo.zic._q_qpos[5] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net318),
    .D(_0197_),
    .Q_N(_4470_),
    .Q(\main.demo.zic._q_qpos[6] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net319),
    .D(_0198_),
    .Q_N(_0043_),
    .Q(\main.demo.zic._q_qpos[7] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net320),
    .D(_0199_),
    .Q_N(_4469_),
    .Q(\main.demo.zic._q_qpos[8] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_qpos[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net321),
    .D(_0200_),
    .Q_N(_4468_),
    .Q(\main.demo.zic._q_qpos[9] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net322),
    .D(_0201_),
    .Q_N(_0068_),
    .Q(\main.demo.zic._q_rythm_count[0] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net323),
    .D(_0202_),
    .Q_N(_4467_),
    .Q(\main.demo.zic._q_rythm_count[10] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net324),
    .D(_0203_),
    .Q_N(_4466_),
    .Q(\main.demo.zic._q_rythm_count[11] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net325),
    .D(_0204_),
    .Q_N(_4465_),
    .Q(\main.demo.zic._q_rythm_count[12] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net326),
    .D(_0205_),
    .Q_N(_4464_),
    .Q(\main.demo.zic._q_rythm_count[1] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net327),
    .D(_0206_),
    .Q_N(_4463_),
    .Q(\main.demo.zic._q_rythm_count[2] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net328),
    .D(_0207_),
    .Q_N(_4462_),
    .Q(\main.demo.zic._q_rythm_count[3] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net329),
    .D(_0208_),
    .Q_N(_4461_),
    .Q(\main.demo.zic._q_rythm_count[4] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net330),
    .D(_0209_),
    .Q_N(_4460_),
    .Q(\main.demo.zic._q_rythm_count[5] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net331),
    .D(_0210_),
    .Q_N(_4459_),
    .Q(\main.demo.zic._q_rythm_count[6] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net332),
    .D(_0211_),
    .Q_N(_4458_),
    .Q(\main.demo.zic._q_rythm_count[7] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net333),
    .D(_0212_),
    .Q_N(_4457_),
    .Q(\main.demo.zic._q_rythm_count[8] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_rythm_count[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net334),
    .D(_0213_),
    .Q_N(_4456_),
    .Q(\main.demo.zic._q_rythm_count[9] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_squ_env[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net335),
    .D(_0214_),
    .Q_N(_4455_),
    .Q(\main.demo.zic._q_squ_env[0] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_squ_env[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net336),
    .D(_0215_),
    .Q_N(_4454_),
    .Q(\main.demo.zic._q_squ_env[1] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_squ_env[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net337),
    .D(_0216_),
    .Q_N(_4453_),
    .Q(\main.demo.zic._q_squ_env[2] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_squ_env[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net338),
    .D(_0217_),
    .Q_N(_0038_),
    .Q(\main.demo.zic._q_squ_env[3] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_squ_env[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net339),
    .D(_0218_),
    .Q_N(_0039_),
    .Q(\main.demo.zic._q_squ_env[4] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_squ_env[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net340),
    .D(_0219_),
    .Q_N(_0040_),
    .Q(\main.demo.zic._q_squ_env[5] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net341),
    .D(_0220_),
    .Q_N(_4452_),
    .Q(\main.demo.zic._q_tpos[0] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net342),
    .D(_0221_),
    .Q_N(_4451_),
    .Q(\main.demo.zic._q_tpos[10] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net343),
    .D(_0222_),
    .Q_N(_0042_),
    .Q(\main.demo.zic._q_tpos[11] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net344),
    .D(_0223_),
    .Q_N(_4450_),
    .Q(\main.demo.zic._q_tpos[1] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net345),
    .D(_0224_),
    .Q_N(_4449_),
    .Q(\main.demo.zic._q_tpos[2] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net346),
    .D(_0225_),
    .Q_N(_4448_),
    .Q(\main.demo.zic._q_tpos[3] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net347),
    .D(_0226_),
    .Q_N(_4447_),
    .Q(\main.demo.zic._q_tpos[4] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net348),
    .D(_0227_),
    .Q_N(_0056_),
    .Q(\main.demo.zic._q_tpos[5] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net349),
    .D(_0228_),
    .Q_N(_4446_),
    .Q(\main.demo.zic._q_tpos[6] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net350),
    .D(_0229_),
    .Q_N(_4445_),
    .Q(\main.demo.zic._q_tpos[7] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net351),
    .D(_0230_),
    .Q_N(_4444_),
    .Q(\main.demo.zic._q_tpos[8] ));
 sg13g2_dfrbp_1 \main.demo.zic._q_tpos[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net352),
    .D(_0231_),
    .Q_N(_4634_),
    .Q(\main.demo.zic._q_tpos[9] ));
 sg13g2_dfrbp_1 \rst_n_q$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net353),
    .D(net1),
    .Q_N(_0012_),
    .Q(rst_n_q));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uio_out[7]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout11 (.A(_3773_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_3160_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_1453_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_2059_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_1977_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_1913_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_1811_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_3945_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1810_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_3924_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_3920_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_3926_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_2374_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0416_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0413_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0288_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_4286_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_4282_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_2204_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0809_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_3598_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_4287_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_2313_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1011_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0436_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0408_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0387_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0308_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_4154_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0793_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0601_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_4411_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_3266_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_2208_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1734_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0798_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0797_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0615_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_4424_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2228_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2176_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1733_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1719_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1241_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0816_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0801_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0799_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0796_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_4423_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_2516_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1718_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1240_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1233_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0800_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0786_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0463_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0451_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_2525_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_2191_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2190_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0587_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0464_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0454_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_4132_),
    .X(net77));
 sg13g2_tielo _9098__78 (.L_LO(net78));
 sg13g2_tielo _9099__79 (.L_LO(net79));
 sg13g2_tielo _9100__80 (.L_LO(net80));
 sg13g2_tielo _9101__81 (.L_LO(net81));
 sg13g2_tielo _9102__82 (.L_LO(net82));
 sg13g2_tielo _9103__83 (.L_LO(net83));
 sg13g2_tielo _9104__84 (.L_LO(net84));
 sg13g2_tielo _9106__85 (.L_LO(net85));
 sg13g2_tielo _9107__86 (.L_LO(net86));
 sg13g2_tielo _9108__87 (.L_LO(net87));
 sg13g2_tielo _9109__88 (.L_LO(net88));
 sg13g2_tielo _9110__89 (.L_LO(net89));
 sg13g2_tielo _9111__90 (.L_LO(net90));
 sg13g2_tielo _9112__91 (.L_LO(net91));
 sg13g2_tiehi _9095__93 (.L_HI(net93));
 sg13g2_tiehi _9105__94 (.L_HI(net94));
 sg13g2_tiehi \main._q_uio_o[7]$_DFF_P__95  (.L_HI(net95));
 sg13g2_tiehi \main._q_uo[0]$_SDFF_PN0__96  (.L_HI(net96));
 sg13g2_tiehi \main._q_uo[1]$_SDFF_PN0__97  (.L_HI(net97));
 sg13g2_tiehi \main._q_uo[2]$_SDFF_PN0__98  (.L_HI(net98));
 sg13g2_tiehi \main._q_uo[3]$_DFF_P__99  (.L_HI(net99));
 sg13g2_tiehi \main._q_uo[4]$_SDFF_PN0__100  (.L_HI(net100));
 sg13g2_tiehi \main._q_uo[5]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_tiehi \main._q_uo[6]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \main._q_uo[7]$_DFF_P__103  (.L_HI(net103));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[0]$_DFF_P__104  (.L_HI(net104));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[10]$_DFF_P__105  (.L_HI(net105));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[1]$_DFF_P__106  (.L_HI(net106));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[2]$_DFF_P__107  (.L_HI(net107));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[3]$_DFF_P__108  (.L_HI(net108));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[4]$_DFF_P__109  (.L_HI(net109));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[5]$_DFF_P__110  (.L_HI(net110));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[6]$_DFF_P__111  (.L_HI(net111));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[7]$_DFF_P__112  (.L_HI(net112));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[8]$_DFF_P__113  (.L_HI(net113));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cx[9]$_DFF_P__114  (.L_HI(net114));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[0]$_DFF_P__115  (.L_HI(net115));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[10]$_DFF_P__116  (.L_HI(net116));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[1]$_DFF_P__117  (.L_HI(net117));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[2]$_DFF_P__118  (.L_HI(net118));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[3]$_DFF_P__119  (.L_HI(net119));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[4]$_DFF_P__120  (.L_HI(net120));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[5]$_DFF_P__121  (.L_HI(net121));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[6]$_DFF_P__122  (.L_HI(net122));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[7]$_DFF_P__123  (.L_HI(net123));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[8]$_DFF_P__124  (.L_HI(net124));
 sg13g2_tiehi \main.demo._q___pip_58_1_1___stage___block_3_cy[9]$_DFF_P__125  (.L_HI(net125));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_a[1]$_DFF_P__126  (.L_HI(net126));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_a[2]$_DFF_P__127  (.L_HI(net127));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_a[3]$_DFF_P__128  (.L_HI(net128));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_a[4]$_DFF_P__129  (.L_HI(net129));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_a[6]$_DFF_P__130  (.L_HI(net130));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_a[7]$_DFF_P__131  (.L_HI(net131));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[0]$_DFF_P__132  (.L_HI(net132));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[10]$_DFF_P__133  (.L_HI(net133));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[1]$_DFF_P__134  (.L_HI(net134));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[2]$_DFF_P__135  (.L_HI(net135));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[3]$_DFF_P__136  (.L_HI(net136));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[4]$_DFF_P__137  (.L_HI(net137));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[5]$_DFF_P__138  (.L_HI(net138));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[6]$_DFF_P__139  (.L_HI(net139));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[7]$_DFF_P__140  (.L_HI(net140));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[8]$_DFF_P__141  (.L_HI(net141));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cx[9]$_DFF_P__142  (.L_HI(net142));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[0]$_DFF_P__143  (.L_HI(net143));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[10]$_DFF_P__144  (.L_HI(net144));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[1]$_DFF_P__145  (.L_HI(net145));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[2]$_DFF_P__146  (.L_HI(net146));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[3]$_DFF_P__147  (.L_HI(net147));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[4]$_DFF_P__148  (.L_HI(net148));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[5]$_DFF_P__149  (.L_HI(net149));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[6]$_DFF_P__150  (.L_HI(net150));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[7]$_DFF_P__151  (.L_HI(net151));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[8]$_DFF_P__152  (.L_HI(net152));
 sg13g2_tiehi \main.demo._q___pip_58_1_2___stage___block_3_cy[9]$_DFF_P__153  (.L_HI(net153));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_a[1]$_DFF_P__154  (.L_HI(net154));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_a[2]$_DFF_P__155  (.L_HI(net155));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_a[3]$_DFF_P__156  (.L_HI(net156));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_a[4]$_DFF_P__157  (.L_HI(net157));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_a[5]$_DFF_P__158  (.L_HI(net158));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_a[6]$_DFF_P__159  (.L_HI(net159));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_a[7]$_DFF_P__160  (.L_HI(net160));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[0]$_DFF_P__161  (.L_HI(net161));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[10]$_DFF_P__162  (.L_HI(net162));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[1]$_DFF_P__163  (.L_HI(net163));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[2]$_DFF_P__164  (.L_HI(net164));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[3]$_DFF_P__165  (.L_HI(net165));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[4]$_DFF_P__166  (.L_HI(net166));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[5]$_DFF_P__167  (.L_HI(net167));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[6]$_DFF_P__168  (.L_HI(net168));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[7]$_DFF_P__169  (.L_HI(net169));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[8]$_DFF_P__170  (.L_HI(net170));
 sg13g2_tiehi \main.demo._q___pip_58_1_3___stage___block_3_cx[9]$_DFF_P__171  (.L_HI(net171));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_68_frag[0]$_DFF_P__172  (.L_HI(net172));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_68_frag[1]$_DFF_P__173  (.L_HI(net173));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_68_frag[2]$_DFF_P__174  (.L_HI(net174));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_68_frag[3]$_DFF_P__175  (.L_HI(net175));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_68_frag[4]$_DFF_P__176  (.L_HI(net176));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_68_frag[5]$_DFF_P__177  (.L_HI(net177));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_87_atten_h[0]$_DFF_P__178  (.L_HI(net178));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_87_atten_h[1]$_DFF_P__179  (.L_HI(net179));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_87_atten_h[2]$_DFF_P__180  (.L_HI(net180));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_87_atten_l[0]$_DFF_P__181  (.L_HI(net181));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___block_87_atten_l[1]$_DFF_P__182  (.L_HI(net182));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___stage___block_3_cx[1]$_DFF_P__183  (.L_HI(net183));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___stage___block_3_cx[2]$_DFF_P__184  (.L_HI(net184));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___stage___block_3_cx[3]$_DFF_P__185  (.L_HI(net185));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___stage___block_3_cx[4]$_DFF_P__186  (.L_HI(net186));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___stage___block_3_cx[5]$_DFF_P__187  (.L_HI(net187));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___stage___block_3_cx[6]$_DFF_P__188  (.L_HI(net188));
 sg13g2_tiehi \main.demo._q___pip_58_1_4___stage___block_3_cx[9]$_DFF_P__189  (.L_HI(net189));
 sg13g2_tiehi \main.demo._q_effect[0]$_SDFFE_PN0P__190  (.L_HI(net190));
 sg13g2_tiehi \main.demo._q_effect[1]$_SDFFE_PN1P__191  (.L_HI(net191));
 sg13g2_tiehi \main.demo._q_frame[0]$_SDFF_PN0__192  (.L_HI(net192));
 sg13g2_tiehi \main.demo._q_frame[10]$_SDFF_PN0__193  (.L_HI(net193));
 sg13g2_tiehi \main.demo._q_frame[11]$_SDFF_PN0__194  (.L_HI(net194));
 sg13g2_tiehi \main.demo._q_frame[12]$_SDFF_PN0__195  (.L_HI(net195));
 sg13g2_tiehi \main.demo._q_frame[13]$_SDFF_PN0__196  (.L_HI(net196));
 sg13g2_tiehi \main.demo._q_frame[14]$_SDFF_PN0__197  (.L_HI(net197));
 sg13g2_tiehi \main.demo._q_frame[1]$_SDFF_PN0__198  (.L_HI(net198));
 sg13g2_tiehi \main.demo._q_frame[2]$_SDFF_PN0__199  (.L_HI(net199));
 sg13g2_tiehi \main.demo._q_frame[3]$_SDFF_PN0__200  (.L_HI(net200));
 sg13g2_tiehi \main.demo._q_frame[4]$_SDFF_PN0__201  (.L_HI(net201));
 sg13g2_tiehi \main.demo._q_frame[5]$_SDFF_PN0__202  (.L_HI(net202));
 sg13g2_tiehi \main.demo._q_frame[6]$_SDFF_PN0__203  (.L_HI(net203));
 sg13g2_tiehi \main.demo._q_frame[7]$_SDFF_PN0__204  (.L_HI(net204));
 sg13g2_tiehi \main.demo._q_frame[8]$_SDFF_PN0__205  (.L_HI(net205));
 sg13g2_tiehi \main.demo._q_frame[9]$_SDFF_PN0__206  (.L_HI(net206));
 sg13g2_tiehi \main.demo._q_go$_SDFF_PN0__207  (.L_HI(net207));
 sg13g2_tiehi \main.demo._q_prev_b[0]$_DFF_P__208  (.L_HI(net208));
 sg13g2_tiehi \main.demo._q_prev_b[1]$_DFF_P__209  (.L_HI(net209));
 sg13g2_tiehi \main.demo._q_prev_b[2]$_DFF_P__210  (.L_HI(net210));
 sg13g2_tiehi \main.demo._q_prev_b[3]$_DFF_P__211  (.L_HI(net211));
 sg13g2_tiehi \main.demo._q_prev_b[4]$_DFF_P__212  (.L_HI(net212));
 sg13g2_tiehi \main.demo._q_prev_b[5]$_DFF_P__213  (.L_HI(net213));
 sg13g2_tiehi \main.demo._q_prev_b[6]$_DFF_P__214  (.L_HI(net214));
 sg13g2_tiehi \main.demo._q_prev_b[7]$_DFF_P__215  (.L_HI(net215));
 sg13g2_tiehi \main.demo._q_rot_en$_SDFFE_PN0P__216  (.L_HI(net216));
 sg13g2_tiehi \main.demo._q_speed[0]$_SDFFE_PP0P__217  (.L_HI(net217));
 sg13g2_tiehi \main.demo._q_speed[10]$_DFFE_PP__218  (.L_HI(net218));
 sg13g2_tiehi \main.demo._q_speed[11]$_DFFE_PP__219  (.L_HI(net219));
 sg13g2_tiehi \main.demo._q_speed[12]$_DFFE_PP__220  (.L_HI(net220));
 sg13g2_tiehi \main.demo._q_speed[13]$_DFFE_PP__221  (.L_HI(net221));
 sg13g2_tiehi \main.demo._q_speed[14]$_DFFE_PP__222  (.L_HI(net222));
 sg13g2_tiehi \main.demo._q_speed[15]$_DFFE_PP__223  (.L_HI(net223));
 sg13g2_tiehi \main.demo._q_speed[1]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \main.demo._q_speed[2]$_DFFE_PP__225  (.L_HI(net225));
 sg13g2_tiehi \main.demo._q_speed[3]$_DFFE_PP__226  (.L_HI(net226));
 sg13g2_tiehi \main.demo._q_speed[4]$_DFFE_PP__227  (.L_HI(net227));
 sg13g2_tiehi \main.demo._q_speed[5]$_DFFE_PP__228  (.L_HI(net228));
 sg13g2_tiehi \main.demo._q_speed[6]$_DFFE_PP__229  (.L_HI(net229));
 sg13g2_tiehi \main.demo._q_speed[7]$_DFFE_PP__230  (.L_HI(net230));
 sg13g2_tiehi \main.demo._q_speed[8]$_DFFE_PP__231  (.L_HI(net231));
 sg13g2_tiehi \main.demo._q_speed[9]$_DFFE_PP__232  (.L_HI(net232));
 sg13g2_tiehi \main.demo._q_th[0]$_SDFFE_PP0P__233  (.L_HI(net233));
 sg13g2_tiehi \main.demo._q_th[1]$_SDFFE_PP0P__234  (.L_HI(net234));
 sg13g2_tiehi \main.demo._q_th[2]$_SDFFE_PP0P__235  (.L_HI(net235));
 sg13g2_tiehi \main.demo._q_th[3]$_SDFFE_PP0P__236  (.L_HI(net236));
 sg13g2_tiehi \main.demo._q_th[4]$_SDFFE_PP0P__237  (.L_HI(net237));
 sg13g2_tiehi \main.demo._q_th[5]$_SDFFE_PP0P__238  (.L_HI(net238));
 sg13g2_tiehi \main.demo._q_th[6]$_SDFFE_PP0P__239  (.L_HI(net239));
 sg13g2_tiehi \main.demo._q_th[7]$_SDFFE_PP0P__240  (.L_HI(net240));
 sg13g2_tiehi \main.demo._q_th[8]$_SDFFE_PP0P__241  (.L_HI(net241));
 sg13g2_tiehi \main.demo.vga._q_active$_DFF_P__242  (.L_HI(net242));
 sg13g2_tiehi \main.demo.vga._q_active_h$_SDFF_PN0__243  (.L_HI(net243));
 sg13g2_tiehi \main.demo.vga._q_active_v$_SDFF_PN0__244  (.L_HI(net244));
 sg13g2_tiehi \main.demo.vga._q_vga_hs$_SDFFE_PP0N__245  (.L_HI(net245));
 sg13g2_tiehi \main.demo.vga._q_vga_vs$_SDFFE_PP0N__246  (.L_HI(net246));
 sg13g2_tiehi \main.demo.vga._q_vga_x[0]$_SDFF_PN0__247  (.L_HI(net247));
 sg13g2_tiehi \main.demo.vga._q_vga_x[10]$_SDFF_PN0__248  (.L_HI(net248));
 sg13g2_tiehi \main.demo.vga._q_vga_x[1]$_SDFF_PN0__249  (.L_HI(net249));
 sg13g2_tiehi \main.demo.vga._q_vga_x[2]$_SDFF_PN0__250  (.L_HI(net250));
 sg13g2_tiehi \main.demo.vga._q_vga_x[3]$_SDFF_PN0__251  (.L_HI(net251));
 sg13g2_tiehi \main.demo.vga._q_vga_x[4]$_SDFF_PN0__252  (.L_HI(net252));
 sg13g2_tiehi \main.demo.vga._q_vga_x[5]$_SDFF_PN0__253  (.L_HI(net253));
 sg13g2_tiehi \main.demo.vga._q_vga_x[6]$_SDFF_PN0__254  (.L_HI(net254));
 sg13g2_tiehi \main.demo.vga._q_vga_x[7]$_SDFF_PN0__255  (.L_HI(net255));
 sg13g2_tiehi \main.demo.vga._q_vga_x[8]$_SDFF_PN0__256  (.L_HI(net256));
 sg13g2_tiehi \main.demo.vga._q_vga_x[9]$_SDFF_PN0__257  (.L_HI(net257));
 sg13g2_tiehi \main.demo.vga._q_vga_y[0]$_SDFF_PP0__258  (.L_HI(net258));
 sg13g2_tiehi \main.demo.vga._q_vga_y[1]$_SDFF_PP0__259  (.L_HI(net259));
 sg13g2_tiehi \main.demo.vga._q_vga_y[2]$_SDFF_PP0__260  (.L_HI(net260));
 sg13g2_tiehi \main.demo.vga._q_vga_y[3]$_SDFF_PP0__261  (.L_HI(net261));
 sg13g2_tiehi \main.demo.vga._q_vga_y[4]$_SDFF_PP0__262  (.L_HI(net262));
 sg13g2_tiehi \main.demo.vga._q_vga_y[5]$_SDFF_PP0__263  (.L_HI(net263));
 sg13g2_tiehi \main.demo.vga._q_vga_y[6]$_SDFF_PP0__264  (.L_HI(net264));
 sg13g2_tiehi \main.demo.vga._q_vga_y[7]$_SDFF_PP0__265  (.L_HI(net265));
 sg13g2_tiehi \main.demo.vga._q_vga_y[8]$_SDFF_PP0__266  (.L_HI(net266));
 sg13g2_tiehi \main.demo.vga._q_vga_y[9]$_SDFF_PP0__267  (.L_HI(net267));
 sg13g2_tiehi \main.demo.vga._q_xcount[0]$_SDFF_PN0__268  (.L_HI(net268));
 sg13g2_tiehi \main.demo.vga._q_xcount[10]$_SDFF_PN0__269  (.L_HI(net269));
 sg13g2_tiehi \main.demo.vga._q_xcount[1]$_SDFF_PP0__270  (.L_HI(net270));
 sg13g2_tiehi \main.demo.vga._q_xcount[2]$_SDFF_PP0__271  (.L_HI(net271));
 sg13g2_tiehi \main.demo.vga._q_xcount[3]$_SDFF_PP0__272  (.L_HI(net272));
 sg13g2_tiehi \main.demo.vga._q_xcount[4]$_SDFF_PP0__273  (.L_HI(net273));
 sg13g2_tiehi \main.demo.vga._q_xcount[5]$_SDFF_PN0__274  (.L_HI(net274));
 sg13g2_tiehi \main.demo.vga._q_xcount[6]$_SDFF_PN0__275  (.L_HI(net275));
 sg13g2_tiehi \main.demo.vga._q_xcount[7]$_SDFF_PP0__276  (.L_HI(net276));
 sg13g2_tiehi \main.demo.vga._q_xcount[8]$_SDFF_PN0__277  (.L_HI(net277));
 sg13g2_tiehi \main.demo.vga._q_xcount[9]$_SDFF_PN0__278  (.L_HI(net278));
 sg13g2_tiehi \main.demo.vga._q_ycount[0]$_SDFFE_PN0P__279  (.L_HI(net279));
 sg13g2_tiehi \main.demo.vga._q_ycount[1]$_SDFFE_PN0P__280  (.L_HI(net280));
 sg13g2_tiehi \main.demo.vga._q_ycount[2]$_SDFFE_PN0P__281  (.L_HI(net281));
 sg13g2_tiehi \main.demo.vga._q_ycount[3]$_SDFFE_PN0P__282  (.L_HI(net282));
 sg13g2_tiehi \main.demo.vga._q_ycount[4]$_SDFFE_PN0P__283  (.L_HI(net283));
 sg13g2_tiehi \main.demo.vga._q_ycount[5]$_SDFFE_PN0P__284  (.L_HI(net284));
 sg13g2_tiehi \main.demo.vga._q_ycount[6]$_SDFFE_PN0P__285  (.L_HI(net285));
 sg13g2_tiehi \main.demo.vga._q_ycount[7]$_SDFFE_PN0P__286  (.L_HI(net286));
 sg13g2_tiehi \main.demo.vga._q_ycount[8]$_SDFFE_PN0P__287  (.L_HI(net287));
 sg13g2_tiehi \main.demo.vga._q_ycount[9]$_SDFFE_PN0P__288  (.L_HI(net288));
 sg13g2_tiehi \main.demo.zic._q_clock_count[0]$_SDFF_PN0__289  (.L_HI(net289));
 sg13g2_tiehi \main.demo.zic._q_clock_count[1]$_SDFF_PN0__290  (.L_HI(net290));
 sg13g2_tiehi \main.demo.zic._q_clock_count[2]$_SDFF_PN0__291  (.L_HI(net291));
 sg13g2_tiehi \main.demo.zic._q_clock_count[3]$_SDFF_PN0__292  (.L_HI(net292));
 sg13g2_tiehi \main.demo.zic._q_clock_count[4]$_SDFF_PN0__293  (.L_HI(net293));
 sg13g2_tiehi \main.demo.zic._q_clock_count[5]$_SDFF_PN0__294  (.L_HI(net294));
 sg13g2_tiehi \main.demo.zic._q_clock_count[6]$_SDFF_PN0__295  (.L_HI(net295));
 sg13g2_tiehi \main.demo.zic._q_clock_count[7]$_SDFF_PN0__296  (.L_HI(net296));
 sg13g2_tiehi \main.demo.zic._q_clock_count[8]$_SDFF_PN0__297  (.L_HI(net297));
 sg13g2_tiehi \main.demo.zic._q_drum_inc[0]$_DFFE_PP__298  (.L_HI(net298));
 sg13g2_tiehi \main.demo.zic._q_drum_inc[1]$_DFFE_PP__299  (.L_HI(net299));
 sg13g2_tiehi \main.demo.zic._q_drum_inc[2]$_DFFE_PP__300  (.L_HI(net300));
 sg13g2_tiehi \main.demo.zic._q_drum_inc[3]$_DFFE_PP__301  (.L_HI(net301));
 sg13g2_tiehi \main.demo.zic._q_idx[0]$_SDFF_PN0__302  (.L_HI(net302));
 sg13g2_tiehi \main.demo.zic._q_idx[1]$_SDFF_PN0__303  (.L_HI(net303));
 sg13g2_tiehi \main.demo.zic._q_idx[2]$_SDFF_PN0__304  (.L_HI(net304));
 sg13g2_tiehi \main.demo.zic._q_idx[3]$_SDFF_PN0__305  (.L_HI(net305));
 sg13g2_tiehi \main.demo.zic._q_idx[4]$_SDFF_PN0__306  (.L_HI(net306));
 sg13g2_tiehi \main.demo.zic._q_idx[5]$_SDFF_PN0__307  (.L_HI(net307));
 sg13g2_tiehi \main.demo.zic._q_idx[6]$_SDFF_PN0__308  (.L_HI(net308));
 sg13g2_tiehi \main.demo.zic._q_qpos[0]$_SDFFE_PN0P__309  (.L_HI(net309));
 sg13g2_tiehi \main.demo.zic._q_qpos[10]$_SDFFE_PN0P__310  (.L_HI(net310));
 sg13g2_tiehi \main.demo.zic._q_qpos[11]$_SDFFE_PN0P__311  (.L_HI(net311));
 sg13g2_tiehi \main.demo.zic._q_qpos[12]$_SDFFE_PN0P__312  (.L_HI(net312));
 sg13g2_tiehi \main.demo.zic._q_qpos[1]$_SDFFE_PN0P__313  (.L_HI(net313));
 sg13g2_tiehi \main.demo.zic._q_qpos[2]$_SDFFE_PN0P__314  (.L_HI(net314));
 sg13g2_tiehi \main.demo.zic._q_qpos[3]$_SDFFE_PN0P__315  (.L_HI(net315));
 sg13g2_tiehi \main.demo.zic._q_qpos[4]$_SDFFE_PN0P__316  (.L_HI(net316));
 sg13g2_tiehi \main.demo.zic._q_qpos[5]$_SDFFE_PN0P__317  (.L_HI(net317));
 sg13g2_tiehi \main.demo.zic._q_qpos[6]$_SDFFE_PN0P__318  (.L_HI(net318));
 sg13g2_tiehi \main.demo.zic._q_qpos[7]$_SDFFE_PN0P__319  (.L_HI(net319));
 sg13g2_tiehi \main.demo.zic._q_qpos[8]$_SDFFE_PN0P__320  (.L_HI(net320));
 sg13g2_tiehi \main.demo.zic._q_qpos[9]$_SDFFE_PN0P__321  (.L_HI(net321));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[0]$_SDFFE_PP0P__322  (.L_HI(net322));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[10]$_SDFFE_PP0P__323  (.L_HI(net323));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[11]$_SDFFE_PP0P__324  (.L_HI(net324));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[12]$_SDFFE_PP0P__325  (.L_HI(net325));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[1]$_SDFFE_PP0P__326  (.L_HI(net326));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[2]$_SDFFE_PP0P__327  (.L_HI(net327));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[3]$_SDFFE_PP0P__328  (.L_HI(net328));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[4]$_SDFFE_PP0P__329  (.L_HI(net329));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[5]$_SDFFE_PP0P__330  (.L_HI(net330));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[6]$_SDFFE_PP0P__331  (.L_HI(net331));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[7]$_SDFFE_PP0P__332  (.L_HI(net332));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[8]$_SDFFE_PP0P__333  (.L_HI(net333));
 sg13g2_tiehi \main.demo.zic._q_rythm_count[9]$_SDFFE_PP0P__334  (.L_HI(net334));
 sg13g2_tiehi \main.demo.zic._q_squ_env[0]$_SDFFE_PN0P__335  (.L_HI(net335));
 sg13g2_tiehi \main.demo.zic._q_squ_env[1]$_SDFFE_PN0P__336  (.L_HI(net336));
 sg13g2_tiehi \main.demo.zic._q_squ_env[2]$_SDFFE_PN0P__337  (.L_HI(net337));
 sg13g2_tiehi \main.demo.zic._q_squ_env[3]$_SDFFE_PN0P__338  (.L_HI(net338));
 sg13g2_tiehi \main.demo.zic._q_squ_env[4]$_SDFFE_PN0P__339  (.L_HI(net339));
 sg13g2_tiehi \main.demo.zic._q_squ_env[5]$_SDFFE_PN0P__340  (.L_HI(net340));
 sg13g2_tiehi \main.demo.zic._q_tpos[0]$_SDFFE_PN0P__341  (.L_HI(net341));
 sg13g2_tiehi \main.demo.zic._q_tpos[10]$_SDFFE_PN0P__342  (.L_HI(net342));
 sg13g2_tiehi \main.demo.zic._q_tpos[11]$_SDFFE_PN0P__343  (.L_HI(net343));
 sg13g2_tiehi \main.demo.zic._q_tpos[1]$_SDFFE_PN0P__344  (.L_HI(net344));
 sg13g2_tiehi \main.demo.zic._q_tpos[2]$_SDFFE_PN0P__345  (.L_HI(net345));
 sg13g2_tiehi \main.demo.zic._q_tpos[3]$_SDFFE_PN0P__346  (.L_HI(net346));
 sg13g2_tiehi \main.demo.zic._q_tpos[4]$_SDFFE_PN0P__347  (.L_HI(net347));
 sg13g2_tiehi \main.demo.zic._q_tpos[5]$_SDFFE_PN0P__348  (.L_HI(net348));
 sg13g2_tiehi \main.demo.zic._q_tpos[6]$_SDFFE_PN0P__349  (.L_HI(net349));
 sg13g2_tiehi \main.demo.zic._q_tpos[7]$_SDFFE_PN0P__350  (.L_HI(net350));
 sg13g2_tiehi \main.demo.zic._q_tpos[8]$_SDFFE_PN0P__351  (.L_HI(net351));
 sg13g2_tiehi \main.demo.zic._q_tpos[9]$_SDFFE_PN0P__352  (.L_HI(net352));
 sg13g2_tiehi \rst_n_q$_DFF_P__353  (.L_HI(net353));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_0_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_34_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_35_clk));
 sg13g2_buf_16 clkload7 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_26_clk));
 sg13g2_buf_16 clkload9 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_14_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_leaf_19_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0129_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(_0129_));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_antennanp ANTENNA_7 (.A(_0129_));
 sg13g2_antennanp ANTENNA_8 (.A(clk));
 sg13g2_antennanp ANTENNA_9 (.A(_0129_));
 sg13g2_antennanp ANTENNA_10 (.A(clk));
 sg13g2_antennanp ANTENNA_11 (.A(_0129_));
 sg13g2_antennanp ANTENNA_12 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_35 ();
 sg13g2_fill_2 FILLER_0_45 ();
 sg13g2_fill_1 FILLER_0_47 ();
 sg13g2_fill_1 FILLER_0_56 ();
 sg13g2_fill_1 FILLER_0_83 ();
 sg13g2_fill_1 FILLER_0_129 ();
 sg13g2_fill_1 FILLER_0_147 ();
 sg13g2_fill_2 FILLER_0_161 ();
 sg13g2_fill_2 FILLER_0_168 ();
 sg13g2_decap_4 FILLER_0_178 ();
 sg13g2_fill_2 FILLER_0_190 ();
 sg13g2_fill_1 FILLER_0_206 ();
 sg13g2_fill_2 FILLER_0_220 ();
 sg13g2_decap_4 FILLER_0_230 ();
 sg13g2_fill_1 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_243 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_fill_2 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_fill_2 FILLER_0_316 ();
 sg13g2_fill_1 FILLER_0_318 ();
 sg13g2_fill_1 FILLER_0_322 ();
 sg13g2_fill_1 FILLER_0_333 ();
 sg13g2_fill_2 FILLER_0_342 ();
 sg13g2_fill_1 FILLER_0_344 ();
 sg13g2_fill_1 FILLER_0_380 ();
 sg13g2_fill_1 FILLER_0_385 ();
 sg13g2_fill_2 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_decap_8 FILLER_0_422 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_4 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_46 ();
 sg13g2_decap_4 FILLER_1_55 ();
 sg13g2_fill_2 FILLER_1_115 ();
 sg13g2_fill_1 FILLER_1_128 ();
 sg13g2_fill_2 FILLER_1_142 ();
 sg13g2_fill_1 FILLER_1_144 ();
 sg13g2_decap_4 FILLER_1_154 ();
 sg13g2_fill_2 FILLER_1_179 ();
 sg13g2_fill_1 FILLER_1_181 ();
 sg13g2_fill_1 FILLER_1_234 ();
 sg13g2_fill_2 FILLER_1_238 ();
 sg13g2_fill_2 FILLER_1_244 ();
 sg13g2_fill_1 FILLER_1_254 ();
 sg13g2_decap_8 FILLER_1_260 ();
 sg13g2_decap_8 FILLER_1_267 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_decap_8 FILLER_1_288 ();
 sg13g2_fill_2 FILLER_1_299 ();
 sg13g2_fill_1 FILLER_1_301 ();
 sg13g2_fill_1 FILLER_1_329 ();
 sg13g2_fill_1 FILLER_1_334 ();
 sg13g2_fill_2 FILLER_1_342 ();
 sg13g2_fill_1 FILLER_1_348 ();
 sg13g2_fill_1 FILLER_1_382 ();
 sg13g2_fill_1 FILLER_1_388 ();
 sg13g2_fill_1 FILLER_1_401 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_417 ();
 sg13g2_decap_4 FILLER_1_424 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_4 FILLER_2_21 ();
 sg13g2_fill_2 FILLER_2_25 ();
 sg13g2_fill_2 FILLER_2_64 ();
 sg13g2_fill_1 FILLER_2_66 ();
 sg13g2_fill_2 FILLER_2_135 ();
 sg13g2_fill_1 FILLER_2_142 ();
 sg13g2_fill_1 FILLER_2_158 ();
 sg13g2_fill_2 FILLER_2_182 ();
 sg13g2_fill_1 FILLER_2_193 ();
 sg13g2_fill_1 FILLER_2_198 ();
 sg13g2_fill_2 FILLER_2_203 ();
 sg13g2_fill_1 FILLER_2_205 ();
 sg13g2_decap_8 FILLER_2_223 ();
 sg13g2_fill_1 FILLER_2_230 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_fill_2 FILLER_2_287 ();
 sg13g2_fill_1 FILLER_2_302 ();
 sg13g2_decap_4 FILLER_2_311 ();
 sg13g2_fill_1 FILLER_2_315 ();
 sg13g2_fill_2 FILLER_2_324 ();
 sg13g2_fill_1 FILLER_2_326 ();
 sg13g2_fill_1 FILLER_2_337 ();
 sg13g2_fill_2 FILLER_2_350 ();
 sg13g2_decap_4 FILLER_2_355 ();
 sg13g2_fill_1 FILLER_2_371 ();
 sg13g2_fill_1 FILLER_2_376 ();
 sg13g2_fill_1 FILLER_2_384 ();
 sg13g2_fill_2 FILLER_2_388 ();
 sg13g2_fill_1 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_419 ();
 sg13g2_decap_4 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_93 ();
 sg13g2_fill_1 FILLER_3_98 ();
 sg13g2_fill_2 FILLER_3_107 ();
 sg13g2_fill_1 FILLER_3_112 ();
 sg13g2_fill_1 FILLER_3_117 ();
 sg13g2_fill_1 FILLER_3_136 ();
 sg13g2_fill_2 FILLER_3_141 ();
 sg13g2_fill_1 FILLER_3_179 ();
 sg13g2_fill_1 FILLER_3_205 ();
 sg13g2_fill_2 FILLER_3_214 ();
 sg13g2_fill_1 FILLER_3_220 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_fill_1 FILLER_3_235 ();
 sg13g2_fill_2 FILLER_3_244 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_4 FILLER_3_266 ();
 sg13g2_fill_1 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_275 ();
 sg13g2_decap_8 FILLER_3_282 ();
 sg13g2_decap_4 FILLER_3_289 ();
 sg13g2_fill_2 FILLER_3_293 ();
 sg13g2_fill_1 FILLER_3_316 ();
 sg13g2_decap_4 FILLER_3_362 ();
 sg13g2_fill_2 FILLER_3_392 ();
 sg13g2_fill_2 FILLER_3_398 ();
 sg13g2_fill_2 FILLER_3_408 ();
 sg13g2_fill_2 FILLER_3_415 ();
 sg13g2_fill_1 FILLER_3_417 ();
 sg13g2_decap_8 FILLER_3_422 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_47 ();
 sg13g2_fill_1 FILLER_4_71 ();
 sg13g2_fill_2 FILLER_4_98 ();
 sg13g2_fill_1 FILLER_4_100 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_fill_2 FILLER_4_156 ();
 sg13g2_fill_2 FILLER_4_173 ();
 sg13g2_fill_1 FILLER_4_175 ();
 sg13g2_fill_1 FILLER_4_191 ();
 sg13g2_fill_1 FILLER_4_200 ();
 sg13g2_fill_1 FILLER_4_213 ();
 sg13g2_fill_2 FILLER_4_223 ();
 sg13g2_fill_1 FILLER_4_225 ();
 sg13g2_fill_2 FILLER_4_230 ();
 sg13g2_fill_1 FILLER_4_236 ();
 sg13g2_fill_2 FILLER_4_262 ();
 sg13g2_fill_2 FILLER_4_290 ();
 sg13g2_fill_1 FILLER_4_292 ();
 sg13g2_fill_2 FILLER_4_309 ();
 sg13g2_fill_1 FILLER_4_321 ();
 sg13g2_fill_1 FILLER_4_326 ();
 sg13g2_fill_1 FILLER_4_335 ();
 sg13g2_fill_1 FILLER_4_340 ();
 sg13g2_fill_1 FILLER_4_351 ();
 sg13g2_fill_1 FILLER_4_371 ();
 sg13g2_fill_1 FILLER_4_377 ();
 sg13g2_fill_1 FILLER_4_382 ();
 sg13g2_fill_1 FILLER_4_396 ();
 sg13g2_fill_1 FILLER_4_405 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_fill_2 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_26 ();
 sg13g2_fill_1 FILLER_5_32 ();
 sg13g2_fill_2 FILLER_5_53 ();
 sg13g2_fill_2 FILLER_5_59 ();
 sg13g2_fill_1 FILLER_5_69 ();
 sg13g2_fill_1 FILLER_5_74 ();
 sg13g2_fill_2 FILLER_5_116 ();
 sg13g2_fill_2 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_170 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_207 ();
 sg13g2_fill_1 FILLER_5_224 ();
 sg13g2_fill_1 FILLER_5_229 ();
 sg13g2_fill_1 FILLER_5_235 ();
 sg13g2_fill_1 FILLER_5_240 ();
 sg13g2_fill_1 FILLER_5_245 ();
 sg13g2_fill_1 FILLER_5_249 ();
 sg13g2_fill_1 FILLER_5_254 ();
 sg13g2_decap_4 FILLER_5_281 ();
 sg13g2_fill_2 FILLER_5_285 ();
 sg13g2_decap_4 FILLER_5_292 ();
 sg13g2_fill_1 FILLER_5_308 ();
 sg13g2_fill_1 FILLER_5_340 ();
 sg13g2_decap_4 FILLER_5_349 ();
 sg13g2_fill_2 FILLER_5_353 ();
 sg13g2_fill_2 FILLER_5_359 ();
 sg13g2_fill_1 FILLER_5_366 ();
 sg13g2_fill_1 FILLER_5_371 ();
 sg13g2_decap_4 FILLER_5_377 ();
 sg13g2_fill_1 FILLER_5_381 ();
 sg13g2_fill_1 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_2 FILLER_5_418 ();
 sg13g2_fill_1 FILLER_5_420 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_39 ();
 sg13g2_fill_1 FILLER_6_48 ();
 sg13g2_fill_1 FILLER_6_57 ();
 sg13g2_fill_1 FILLER_6_62 ();
 sg13g2_fill_1 FILLER_6_66 ();
 sg13g2_fill_2 FILLER_6_71 ();
 sg13g2_fill_1 FILLER_6_73 ();
 sg13g2_fill_1 FILLER_6_104 ();
 sg13g2_fill_2 FILLER_6_118 ();
 sg13g2_fill_2 FILLER_6_125 ();
 sg13g2_fill_2 FILLER_6_131 ();
 sg13g2_fill_1 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_144 ();
 sg13g2_fill_1 FILLER_6_150 ();
 sg13g2_fill_1 FILLER_6_156 ();
 sg13g2_fill_1 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_192 ();
 sg13g2_fill_2 FILLER_6_204 ();
 sg13g2_decap_4 FILLER_6_210 ();
 sg13g2_fill_2 FILLER_6_214 ();
 sg13g2_fill_1 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_227 ();
 sg13g2_fill_1 FILLER_6_236 ();
 sg13g2_fill_1 FILLER_6_245 ();
 sg13g2_fill_2 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_269 ();
 sg13g2_decap_4 FILLER_6_276 ();
 sg13g2_fill_2 FILLER_6_288 ();
 sg13g2_fill_1 FILLER_6_290 ();
 sg13g2_fill_1 FILLER_6_303 ();
 sg13g2_fill_1 FILLER_6_312 ();
 sg13g2_fill_1 FILLER_6_337 ();
 sg13g2_fill_1 FILLER_6_342 ();
 sg13g2_fill_1 FILLER_6_346 ();
 sg13g2_fill_2 FILLER_6_352 ();
 sg13g2_decap_4 FILLER_6_359 ();
 sg13g2_fill_2 FILLER_6_378 ();
 sg13g2_decap_4 FILLER_6_393 ();
 sg13g2_fill_1 FILLER_6_417 ();
 sg13g2_fill_2 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_4 FILLER_7_21 ();
 sg13g2_fill_1 FILLER_7_49 ();
 sg13g2_fill_2 FILLER_7_58 ();
 sg13g2_fill_2 FILLER_7_69 ();
 sg13g2_fill_1 FILLER_7_79 ();
 sg13g2_fill_1 FILLER_7_110 ();
 sg13g2_fill_1 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_131 ();
 sg13g2_fill_1 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_172 ();
 sg13g2_fill_1 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_184 ();
 sg13g2_fill_1 FILLER_7_217 ();
 sg13g2_fill_1 FILLER_7_226 ();
 sg13g2_fill_1 FILLER_7_235 ();
 sg13g2_fill_1 FILLER_7_241 ();
 sg13g2_fill_1 FILLER_7_247 ();
 sg13g2_decap_4 FILLER_7_285 ();
 sg13g2_fill_2 FILLER_7_289 ();
 sg13g2_fill_2 FILLER_7_325 ();
 sg13g2_fill_2 FILLER_7_347 ();
 sg13g2_fill_1 FILLER_7_374 ();
 sg13g2_fill_2 FILLER_7_389 ();
 sg13g2_fill_1 FILLER_7_400 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_1 FILLER_7_414 ();
 sg13g2_fill_1 FILLER_7_423 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_4 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_64 ();
 sg13g2_fill_1 FILLER_8_69 ();
 sg13g2_fill_1 FILLER_8_78 ();
 sg13g2_decap_8 FILLER_8_96 ();
 sg13g2_fill_1 FILLER_8_146 ();
 sg13g2_fill_1 FILLER_8_179 ();
 sg13g2_fill_1 FILLER_8_184 ();
 sg13g2_fill_2 FILLER_8_189 ();
 sg13g2_fill_1 FILLER_8_191 ();
 sg13g2_fill_1 FILLER_8_197 ();
 sg13g2_fill_2 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_210 ();
 sg13g2_fill_1 FILLER_8_228 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_fill_2 FILLER_8_285 ();
 sg13g2_fill_1 FILLER_8_287 ();
 sg13g2_fill_1 FILLER_8_295 ();
 sg13g2_fill_1 FILLER_8_322 ();
 sg13g2_fill_2 FILLER_8_349 ();
 sg13g2_fill_2 FILLER_8_355 ();
 sg13g2_fill_1 FILLER_8_357 ();
 sg13g2_fill_1 FILLER_8_367 ();
 sg13g2_fill_2 FILLER_8_372 ();
 sg13g2_fill_1 FILLER_8_374 ();
 sg13g2_fill_1 FILLER_8_379 ();
 sg13g2_fill_2 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_418 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_4 FILLER_9_21 ();
 sg13g2_fill_1 FILLER_9_25 ();
 sg13g2_fill_1 FILLER_9_40 ();
 sg13g2_fill_2 FILLER_9_53 ();
 sg13g2_decap_4 FILLER_9_59 ();
 sg13g2_fill_2 FILLER_9_117 ();
 sg13g2_fill_1 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_fill_2 FILLER_9_186 ();
 sg13g2_fill_1 FILLER_9_199 ();
 sg13g2_fill_2 FILLER_9_212 ();
 sg13g2_fill_2 FILLER_9_251 ();
 sg13g2_fill_1 FILLER_9_266 ();
 sg13g2_fill_1 FILLER_9_272 ();
 sg13g2_fill_1 FILLER_9_278 ();
 sg13g2_fill_1 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_287 ();
 sg13g2_fill_2 FILLER_9_293 ();
 sg13g2_fill_2 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_337 ();
 sg13g2_fill_2 FILLER_9_357 ();
 sg13g2_fill_1 FILLER_9_363 ();
 sg13g2_fill_2 FILLER_9_368 ();
 sg13g2_fill_1 FILLER_9_381 ();
 sg13g2_fill_1 FILLER_9_386 ();
 sg13g2_fill_2 FILLER_9_390 ();
 sg13g2_decap_4 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_38 ();
 sg13g2_fill_2 FILLER_10_62 ();
 sg13g2_fill_1 FILLER_10_72 ();
 sg13g2_fill_1 FILLER_10_86 ();
 sg13g2_fill_2 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_104 ();
 sg13g2_fill_2 FILLER_10_111 ();
 sg13g2_fill_1 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_129 ();
 sg13g2_fill_1 FILLER_10_160 ();
 sg13g2_fill_1 FILLER_10_164 ();
 sg13g2_fill_1 FILLER_10_170 ();
 sg13g2_fill_1 FILLER_10_179 ();
 sg13g2_fill_1 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_216 ();
 sg13g2_fill_2 FILLER_10_223 ();
 sg13g2_fill_2 FILLER_10_276 ();
 sg13g2_fill_1 FILLER_10_278 ();
 sg13g2_decap_4 FILLER_10_282 ();
 sg13g2_fill_2 FILLER_10_298 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_fill_1 FILLER_10_311 ();
 sg13g2_fill_1 FILLER_10_315 ();
 sg13g2_fill_1 FILLER_10_338 ();
 sg13g2_fill_2 FILLER_10_345 ();
 sg13g2_fill_2 FILLER_10_350 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_fill_2 FILLER_10_394 ();
 sg13g2_fill_1 FILLER_10_396 ();
 sg13g2_fill_2 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_10_418 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_13 ();
 sg13g2_fill_1 FILLER_11_19 ();
 sg13g2_fill_1 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_63 ();
 sg13g2_fill_1 FILLER_11_67 ();
 sg13g2_fill_1 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_171 ();
 sg13g2_fill_1 FILLER_11_173 ();
 sg13g2_fill_2 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_184 ();
 sg13g2_fill_2 FILLER_11_233 ();
 sg13g2_fill_2 FILLER_11_245 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_fill_2 FILLER_11_278 ();
 sg13g2_fill_2 FILLER_11_298 ();
 sg13g2_fill_1 FILLER_11_300 ();
 sg13g2_fill_2 FILLER_11_310 ();
 sg13g2_fill_2 FILLER_11_328 ();
 sg13g2_fill_1 FILLER_11_330 ();
 sg13g2_fill_1 FILLER_11_341 ();
 sg13g2_fill_2 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_381 ();
 sg13g2_fill_1 FILLER_11_383 ();
 sg13g2_fill_2 FILLER_11_390 ();
 sg13g2_fill_2 FILLER_11_396 ();
 sg13g2_fill_1 FILLER_11_418 ();
 sg13g2_fill_1 FILLER_11_423 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_5 ();
 sg13g2_fill_1 FILLER_12_10 ();
 sg13g2_fill_1 FILLER_12_16 ();
 sg13g2_fill_1 FILLER_12_22 ();
 sg13g2_decap_4 FILLER_12_27 ();
 sg13g2_fill_1 FILLER_12_31 ();
 sg13g2_fill_1 FILLER_12_35 ();
 sg13g2_fill_1 FILLER_12_57 ();
 sg13g2_fill_1 FILLER_12_61 ();
 sg13g2_fill_1 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_112 ();
 sg13g2_fill_1 FILLER_12_154 ();
 sg13g2_fill_2 FILLER_12_163 ();
 sg13g2_fill_1 FILLER_12_165 ();
 sg13g2_fill_1 FILLER_12_191 ();
 sg13g2_fill_1 FILLER_12_195 ();
 sg13g2_fill_2 FILLER_12_201 ();
 sg13g2_fill_1 FILLER_12_215 ();
 sg13g2_fill_2 FILLER_12_224 ();
 sg13g2_fill_1 FILLER_12_234 ();
 sg13g2_fill_2 FILLER_12_261 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_272 ();
 sg13g2_fill_1 FILLER_12_274 ();
 sg13g2_fill_1 FILLER_12_294 ();
 sg13g2_decap_4 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_fill_2 FILLER_12_373 ();
 sg13g2_decap_4 FILLER_12_381 ();
 sg13g2_fill_1 FILLER_12_385 ();
 sg13g2_fill_2 FILLER_12_391 ();
 sg13g2_fill_2 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_18 ();
 sg13g2_fill_1 FILLER_13_20 ();
 sg13g2_fill_1 FILLER_13_47 ();
 sg13g2_fill_1 FILLER_13_65 ();
 sg13g2_fill_1 FILLER_13_74 ();
 sg13g2_decap_4 FILLER_13_87 ();
 sg13g2_decap_4 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_decap_4 FILLER_13_148 ();
 sg13g2_fill_1 FILLER_13_152 ();
 sg13g2_fill_2 FILLER_13_187 ();
 sg13g2_fill_2 FILLER_13_211 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_232 ();
 sg13g2_decap_4 FILLER_13_239 ();
 sg13g2_fill_2 FILLER_13_251 ();
 sg13g2_fill_1 FILLER_13_253 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_265 ();
 sg13g2_fill_1 FILLER_13_282 ();
 sg13g2_fill_2 FILLER_13_291 ();
 sg13g2_fill_1 FILLER_13_301 ();
 sg13g2_fill_1 FILLER_13_348 ();
 sg13g2_fill_1 FILLER_13_362 ();
 sg13g2_fill_1 FILLER_13_379 ();
 sg13g2_fill_2 FILLER_13_383 ();
 sg13g2_fill_1 FILLER_13_385 ();
 sg13g2_fill_2 FILLER_13_390 ();
 sg13g2_fill_1 FILLER_13_392 ();
 sg13g2_fill_2 FILLER_13_408 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_24 ();
 sg13g2_fill_2 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_44 ();
 sg13g2_decap_4 FILLER_14_73 ();
 sg13g2_fill_2 FILLER_14_94 ();
 sg13g2_fill_1 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_108 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_162 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_fill_2 FILLER_14_210 ();
 sg13g2_fill_2 FILLER_14_217 ();
 sg13g2_fill_1 FILLER_14_219 ();
 sg13g2_fill_2 FILLER_14_259 ();
 sg13g2_fill_2 FILLER_14_274 ();
 sg13g2_fill_1 FILLER_14_276 ();
 sg13g2_fill_2 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_decap_4 FILLER_14_328 ();
 sg13g2_fill_1 FILLER_14_349 ();
 sg13g2_fill_1 FILLER_14_354 ();
 sg13g2_fill_1 FILLER_14_363 ();
 sg13g2_fill_2 FILLER_14_368 ();
 sg13g2_fill_1 FILLER_14_374 ();
 sg13g2_fill_1 FILLER_14_378 ();
 sg13g2_fill_2 FILLER_14_383 ();
 sg13g2_fill_2 FILLER_14_389 ();
 sg13g2_fill_2 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_424 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_15 ();
 sg13g2_fill_2 FILLER_15_33 ();
 sg13g2_fill_2 FILLER_15_45 ();
 sg13g2_fill_1 FILLER_15_47 ();
 sg13g2_fill_1 FILLER_15_86 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_99 ();
 sg13g2_fill_1 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_fill_1 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_226 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_decap_4 FILLER_15_278 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_fill_2 FILLER_15_302 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_fill_1 FILLER_15_317 ();
 sg13g2_fill_1 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_fill_2 FILLER_15_342 ();
 sg13g2_fill_1 FILLER_15_344 ();
 sg13g2_fill_2 FILLER_15_354 ();
 sg13g2_fill_2 FILLER_15_379 ();
 sg13g2_fill_1 FILLER_15_393 ();
 sg13g2_fill_2 FILLER_15_402 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_33 ();
 sg13g2_fill_1 FILLER_16_38 ();
 sg13g2_fill_1 FILLER_16_51 ();
 sg13g2_decap_4 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_fill_2 FILLER_16_161 ();
 sg13g2_fill_2 FILLER_16_171 ();
 sg13g2_fill_2 FILLER_16_202 ();
 sg13g2_fill_2 FILLER_16_220 ();
 sg13g2_fill_1 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_267 ();
 sg13g2_fill_1 FILLER_16_269 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_fill_2 FILLER_16_281 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_decap_4 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_decap_4 FILLER_16_343 ();
 sg13g2_fill_2 FILLER_16_347 ();
 sg13g2_fill_1 FILLER_16_378 ();
 sg13g2_fill_1 FILLER_16_383 ();
 sg13g2_fill_1 FILLER_16_411 ();
 sg13g2_fill_2 FILLER_16_416 ();
 sg13g2_fill_1 FILLER_16_423 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_1 FILLER_17_69 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_2 FILLER_17_128 ();
 sg13g2_decap_4 FILLER_17_156 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_265 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_decap_4 FILLER_17_277 ();
 sg13g2_fill_2 FILLER_17_281 ();
 sg13g2_decap_4 FILLER_17_287 ();
 sg13g2_fill_2 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_305 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_fill_2 FILLER_17_330 ();
 sg13g2_fill_2 FILLER_17_394 ();
 sg13g2_decap_4 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_405 ();
 sg13g2_decap_4 FILLER_17_415 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_11 ();
 sg13g2_fill_1 FILLER_18_16 ();
 sg13g2_fill_1 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_27 ();
 sg13g2_fill_2 FILLER_18_36 ();
 sg13g2_fill_1 FILLER_18_38 ();
 sg13g2_fill_1 FILLER_18_58 ();
 sg13g2_decap_4 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_67 ();
 sg13g2_fill_2 FILLER_18_81 ();
 sg13g2_fill_1 FILLER_18_83 ();
 sg13g2_decap_4 FILLER_18_87 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_decap_4 FILLER_18_96 ();
 sg13g2_fill_1 FILLER_18_100 ();
 sg13g2_fill_2 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_2 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_182 ();
 sg13g2_fill_2 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_225 ();
 sg13g2_fill_1 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_301 ();
 sg13g2_fill_2 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_332 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_fill_1 FILLER_18_364 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_399 ();
 sg13g2_fill_1 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_405 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_10 ();
 sg13g2_fill_1 FILLER_19_15 ();
 sg13g2_fill_1 FILLER_19_24 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_1 FILLER_19_41 ();
 sg13g2_fill_2 FILLER_19_45 ();
 sg13g2_fill_1 FILLER_19_47 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_fill_1 FILLER_19_117 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_decap_4 FILLER_19_196 ();
 sg13g2_fill_2 FILLER_19_200 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_320 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_fill_2 FILLER_19_340 ();
 sg13g2_decap_4 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_364 ();
 sg13g2_fill_1 FILLER_19_370 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_fill_1 FILLER_19_400 ();
 sg13g2_fill_1 FILLER_19_415 ();
 sg13g2_fill_1 FILLER_19_419 ();
 sg13g2_fill_2 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_13 ();
 sg13g2_fill_2 FILLER_20_40 ();
 sg13g2_fill_2 FILLER_20_45 ();
 sg13g2_fill_1 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_87 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_fill_1 FILLER_20_130 ();
 sg13g2_fill_1 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_4 FILLER_20_235 ();
 sg13g2_fill_2 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_254 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_296 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_338 ();
 sg13g2_fill_2 FILLER_20_377 ();
 sg13g2_fill_1 FILLER_20_383 ();
 sg13g2_fill_1 FILLER_20_400 ();
 sg13g2_decap_8 FILLER_20_405 ();
 sg13g2_decap_4 FILLER_20_412 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_72 ();
 sg13g2_fill_2 FILLER_21_81 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_241 ();
 sg13g2_decap_4 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_264 ();
 sg13g2_fill_1 FILLER_21_270 ();
 sg13g2_decap_4 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_284 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_2 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_326 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_fill_1 FILLER_21_336 ();
 sg13g2_fill_2 FILLER_21_353 ();
 sg13g2_decap_4 FILLER_21_392 ();
 sg13g2_fill_1 FILLER_21_405 ();
 sg13g2_decap_4 FILLER_21_415 ();
 sg13g2_decap_4 FILLER_21_423 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_22 ();
 sg13g2_fill_1 FILLER_22_24 ();
 sg13g2_fill_2 FILLER_22_30 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_fill_1 FILLER_22_52 ();
 sg13g2_fill_1 FILLER_22_57 ();
 sg13g2_fill_1 FILLER_22_88 ();
 sg13g2_fill_1 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_107 ();
 sg13g2_fill_2 FILLER_22_111 ();
 sg13g2_fill_1 FILLER_22_113 ();
 sg13g2_fill_2 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_4 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_144 ();
 sg13g2_decap_4 FILLER_22_149 ();
 sg13g2_decap_4 FILLER_22_157 ();
 sg13g2_fill_2 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_171 ();
 sg13g2_fill_2 FILLER_22_177 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_decap_4 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_decap_4 FILLER_22_231 ();
 sg13g2_fill_2 FILLER_22_235 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_fill_1 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_fill_2 FILLER_22_286 ();
 sg13g2_decap_4 FILLER_22_292 ();
 sg13g2_fill_1 FILLER_22_296 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_decap_4 FILLER_22_333 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_fill_1 FILLER_22_409 ();
 sg13g2_fill_1 FILLER_22_422 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_29 ();
 sg13g2_fill_1 FILLER_23_31 ();
 sg13g2_decap_8 FILLER_23_43 ();
 sg13g2_fill_2 FILLER_23_50 ();
 sg13g2_fill_1 FILLER_23_52 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_95 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_decap_8 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_244 ();
 sg13g2_fill_1 FILLER_23_246 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_fill_2 FILLER_23_334 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_386 ();
 sg13g2_fill_1 FILLER_23_391 ();
 sg13g2_fill_1 FILLER_23_396 ();
 sg13g2_fill_2 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_19 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_33 ();
 sg13g2_fill_2 FILLER_24_62 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_119 ();
 sg13g2_fill_1 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_245 ();
 sg13g2_decap_4 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_281 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_311 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_fill_2 FILLER_24_356 ();
 sg13g2_fill_1 FILLER_24_358 ();
 sg13g2_fill_2 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_379 ();
 sg13g2_fill_1 FILLER_24_392 ();
 sg13g2_fill_1 FILLER_24_397 ();
 sg13g2_fill_1 FILLER_24_402 ();
 sg13g2_fill_1 FILLER_24_413 ();
 sg13g2_fill_1 FILLER_25_8 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_fill_1 FILLER_25_25 ();
 sg13g2_decap_4 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_fill_1 FILLER_25_67 ();
 sg13g2_fill_1 FILLER_25_88 ();
 sg13g2_fill_1 FILLER_25_101 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_decap_4 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_fill_2 FILLER_25_260 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_fill_1 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_291 ();
 sg13g2_fill_2 FILLER_25_297 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_347 ();
 sg13g2_fill_1 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_decap_4 FILLER_25_367 ();
 sg13g2_fill_1 FILLER_25_371 ();
 sg13g2_decap_4 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_25_406 ();
 sg13g2_fill_2 FILLER_25_425 ();
 sg13g2_fill_2 FILLER_26_20 ();
 sg13g2_fill_2 FILLER_26_30 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_fill_1 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_86 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_fill_1 FILLER_26_122 ();
 sg13g2_fill_2 FILLER_26_153 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_decap_4 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_decap_4 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_fill_2 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_fill_2 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_350 ();
 sg13g2_fill_2 FILLER_26_355 ();
 sg13g2_decap_4 FILLER_26_365 ();
 sg13g2_fill_1 FILLER_26_369 ();
 sg13g2_fill_1 FILLER_26_379 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_27 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_fill_2 FILLER_27_61 ();
 sg13g2_fill_1 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_1 FILLER_27_128 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_fill_2 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_decap_4 FILLER_27_227 ();
 sg13g2_decap_4 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_fill_2 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_fill_2 FILLER_27_287 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_326 ();
 sg13g2_fill_2 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_352 ();
 sg13g2_decap_4 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_1 FILLER_27_409 ();
 sg13g2_fill_1 FILLER_27_414 ();
 sg13g2_fill_2 FILLER_27_424 ();
 sg13g2_fill_2 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_76 ();
 sg13g2_fill_2 FILLER_28_138 ();
 sg13g2_fill_1 FILLER_28_166 ();
 sg13g2_fill_2 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_fill_2 FILLER_28_321 ();
 sg13g2_decap_4 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_336 ();
 sg13g2_decap_4 FILLER_28_352 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_decap_4 FILLER_28_369 ();
 sg13g2_decap_4 FILLER_28_390 ();
 sg13g2_fill_1 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_1 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_410 ();
 sg13g2_fill_2 FILLER_28_415 ();
 sg13g2_fill_1 FILLER_28_417 ();
 sg13g2_decap_8 FILLER_28_422 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_51 ();
 sg13g2_fill_2 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_fill_1 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_157 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_decap_4 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_213 ();
 sg13g2_fill_2 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_226 ();
 sg13g2_decap_4 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_fill_2 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_323 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_fill_2 FILLER_29_347 ();
 sg13g2_fill_1 FILLER_29_372 ();
 sg13g2_fill_2 FILLER_29_377 ();
 sg13g2_fill_2 FILLER_29_392 ();
 sg13g2_decap_4 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_416 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_1 FILLER_30_18 ();
 sg13g2_fill_1 FILLER_30_51 ();
 sg13g2_fill_1 FILLER_30_64 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_171 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_decap_8 FILLER_30_241 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_4 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_decap_4 FILLER_30_319 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_fill_2 FILLER_30_344 ();
 sg13g2_fill_2 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_decap_4 FILLER_30_390 ();
 sg13g2_fill_2 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_406 ();
 sg13g2_fill_2 FILLER_30_420 ();
 sg13g2_fill_1 FILLER_30_422 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_111 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_fill_2 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_271 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_294 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_fill_2 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_358 ();
 sg13g2_decap_4 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_387 ();
 sg13g2_decap_4 FILLER_31_392 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_decap_4 FILLER_31_410 ();
 sg13g2_fill_1 FILLER_31_414 ();
 sg13g2_fill_2 FILLER_31_427 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_32 ();
 sg13g2_fill_1 FILLER_32_59 ();
 sg13g2_fill_1 FILLER_32_64 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_fill_2 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_decap_4 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_284 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_fill_1 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_319 ();
 sg13g2_fill_2 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_357 ();
 sg13g2_decap_4 FILLER_32_388 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_decap_4 FILLER_32_410 ();
 sg13g2_fill_1 FILLER_32_419 ();
 sg13g2_fill_1 FILLER_33_51 ();
 sg13g2_fill_2 FILLER_33_62 ();
 sg13g2_fill_1 FILLER_33_64 ();
 sg13g2_fill_2 FILLER_33_94 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_167 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_fill_2 FILLER_33_230 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_fill_1 FILLER_33_297 ();
 sg13g2_fill_2 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_333 ();
 sg13g2_fill_1 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_fill_1 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_1 FILLER_33_383 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_fill_1 FILLER_33_395 ();
 sg13g2_fill_2 FILLER_33_400 ();
 sg13g2_fill_1 FILLER_33_402 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_1 FILLER_33_409 ();
 sg13g2_fill_2 FILLER_33_414 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_fill_2 FILLER_34_104 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_176 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_decap_4 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_268 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_289 ();
 sg13g2_decap_8 FILLER_34_295 ();
 sg13g2_decap_4 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_311 ();
 sg13g2_fill_2 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_1 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_388 ();
 sg13g2_fill_2 FILLER_34_393 ();
 sg13g2_fill_1 FILLER_34_395 ();
 sg13g2_decap_4 FILLER_34_411 ();
 sg13g2_fill_2 FILLER_34_419 ();
 sg13g2_fill_1 FILLER_35_30 ();
 sg13g2_fill_1 FILLER_35_46 ();
 sg13g2_fill_2 FILLER_35_60 ();
 sg13g2_fill_2 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_179 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_fill_2 FILLER_35_189 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_decap_4 FILLER_35_265 ();
 sg13g2_fill_1 FILLER_35_269 ();
 sg13g2_decap_4 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_decap_4 FILLER_35_301 ();
 sg13g2_fill_1 FILLER_35_335 ();
 sg13g2_fill_2 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_381 ();
 sg13g2_fill_1 FILLER_35_390 ();
 sg13g2_decap_4 FILLER_35_399 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_fill_1 FILLER_35_415 ();
 sg13g2_decap_4 FILLER_35_425 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_22 ();
 sg13g2_fill_2 FILLER_36_39 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_fill_1 FILLER_36_108 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_143 ();
 sg13g2_fill_1 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_163 ();
 sg13g2_fill_2 FILLER_36_169 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_fill_2 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_229 ();
 sg13g2_fill_2 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_346 ();
 sg13g2_fill_1 FILLER_36_348 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_fill_2 FILLER_36_416 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_1 FILLER_37_26 ();
 sg13g2_fill_2 FILLER_37_37 ();
 sg13g2_fill_2 FILLER_37_46 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_2 FILLER_37_144 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_2 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_295 ();
 sg13g2_fill_1 FILLER_37_305 ();
 sg13g2_fill_1 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_374 ();
 sg13g2_fill_2 FILLER_37_380 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_decap_4 FILLER_37_392 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_1 FILLER_38_26 ();
 sg13g2_fill_1 FILLER_38_88 ();
 sg13g2_fill_2 FILLER_38_93 ();
 sg13g2_fill_2 FILLER_38_99 ();
 sg13g2_fill_2 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_114 ();
 sg13g2_fill_1 FILLER_38_129 ();
 sg13g2_fill_1 FILLER_38_168 ();
 sg13g2_fill_2 FILLER_38_173 ();
 sg13g2_fill_1 FILLER_38_182 ();
 sg13g2_fill_1 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_fill_1 FILLER_38_207 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_238 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_fill_2 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_283 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_fill_2 FILLER_38_353 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_363 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_fill_2 FILLER_38_383 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_2 ();
 sg13g2_fill_1 FILLER_39_15 ();
 sg13g2_fill_2 FILLER_39_60 ();
 sg13g2_decap_8 FILLER_39_73 ();
 sg13g2_decap_4 FILLER_39_80 ();
 sg13g2_fill_2 FILLER_39_84 ();
 sg13g2_fill_1 FILLER_39_117 ();
 sg13g2_fill_1 FILLER_39_157 ();
 sg13g2_fill_1 FILLER_39_166 ();
 sg13g2_fill_1 FILLER_39_183 ();
 sg13g2_fill_1 FILLER_39_191 ();
 sg13g2_fill_1 FILLER_39_200 ();
 sg13g2_fill_1 FILLER_39_209 ();
 sg13g2_fill_1 FILLER_39_236 ();
 sg13g2_fill_1 FILLER_39_242 ();
 sg13g2_fill_2 FILLER_39_316 ();
 sg13g2_fill_2 FILLER_39_325 ();
 sg13g2_fill_1 FILLER_39_327 ();
 sg13g2_fill_2 FILLER_39_354 ();
 sg13g2_fill_1 FILLER_39_356 ();
 sg13g2_fill_1 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_385 ();
 sg13g2_fill_1 FILLER_39_390 ();
 sg13g2_fill_1 FILLER_39_394 ();
 sg13g2_fill_1 FILLER_39_399 ();
 sg13g2_fill_1 FILLER_39_404 ();
 sg13g2_fill_2 FILLER_39_413 ();
 sg13g2_fill_1 FILLER_39_423 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_fill_1 FILLER_40_43 ();
 sg13g2_fill_2 FILLER_40_48 ();
 sg13g2_fill_1 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_81 ();
 sg13g2_fill_1 FILLER_40_117 ();
 sg13g2_fill_1 FILLER_40_131 ();
 sg13g2_fill_1 FILLER_40_151 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_2 FILLER_40_207 ();
 sg13g2_fill_1 FILLER_40_223 ();
 sg13g2_fill_1 FILLER_40_252 ();
 sg13g2_fill_2 FILLER_40_280 ();
 sg13g2_fill_1 FILLER_40_292 ();
 sg13g2_fill_1 FILLER_40_300 ();
 sg13g2_fill_2 FILLER_40_322 ();
 sg13g2_fill_1 FILLER_40_371 ();
 sg13g2_fill_2 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_fill_1 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_406 ();
 sg13g2_fill_2 FILLER_40_415 ();
 sg13g2_fill_1 FILLER_40_417 ();
 sg13g2_fill_2 FILLER_41_16 ();
 sg13g2_fill_2 FILLER_41_56 ();
 sg13g2_fill_2 FILLER_41_89 ();
 sg13g2_fill_1 FILLER_41_95 ();
 sg13g2_fill_2 FILLER_41_100 ();
 sg13g2_fill_1 FILLER_41_102 ();
 sg13g2_fill_1 FILLER_41_115 ();
 sg13g2_fill_1 FILLER_41_128 ();
 sg13g2_fill_1 FILLER_41_134 ();
 sg13g2_fill_2 FILLER_41_140 ();
 sg13g2_fill_1 FILLER_41_142 ();
 sg13g2_fill_1 FILLER_41_150 ();
 sg13g2_decap_8 FILLER_41_184 ();
 sg13g2_fill_2 FILLER_41_191 ();
 sg13g2_fill_1 FILLER_41_193 ();
 sg13g2_fill_1 FILLER_41_230 ();
 sg13g2_fill_1 FILLER_41_236 ();
 sg13g2_fill_2 FILLER_41_298 ();
 sg13g2_fill_2 FILLER_41_352 ();
 sg13g2_fill_2 FILLER_41_389 ();
 sg13g2_fill_2 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_fill_2 FILLER_42_18 ();
 sg13g2_fill_1 FILLER_42_25 ();
 sg13g2_fill_1 FILLER_42_34 ();
 sg13g2_fill_2 FILLER_42_42 ();
 sg13g2_fill_2 FILLER_42_74 ();
 sg13g2_fill_1 FILLER_42_110 ();
 sg13g2_fill_1 FILLER_42_137 ();
 sg13g2_fill_2 FILLER_42_142 ();
 sg13g2_fill_1 FILLER_42_154 ();
 sg13g2_decap_4 FILLER_42_176 ();
 sg13g2_fill_1 FILLER_42_180 ();
 sg13g2_fill_2 FILLER_42_202 ();
 sg13g2_fill_2 FILLER_42_253 ();
 sg13g2_fill_1 FILLER_42_255 ();
 sg13g2_fill_2 FILLER_42_260 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_fill_2 FILLER_42_273 ();
 sg13g2_fill_1 FILLER_42_341 ();
 sg13g2_fill_2 FILLER_42_375 ();
 sg13g2_fill_1 FILLER_42_386 ();
 sg13g2_fill_1 FILLER_42_395 ();
 sg13g2_fill_1 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_409 ();
 sg13g2_fill_1 FILLER_42_414 ();
 sg13g2_fill_1 FILLER_42_419 ();
 sg13g2_fill_1 FILLER_42_424 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_fill_1 FILLER_43_15 ();
 sg13g2_fill_1 FILLER_43_20 ();
 sg13g2_fill_1 FILLER_43_68 ();
 sg13g2_fill_1 FILLER_43_74 ();
 sg13g2_fill_1 FILLER_43_79 ();
 sg13g2_fill_1 FILLER_43_85 ();
 sg13g2_fill_1 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_96 ();
 sg13g2_fill_1 FILLER_43_160 ();
 sg13g2_fill_2 FILLER_43_182 ();
 sg13g2_fill_1 FILLER_43_184 ();
 sg13g2_decap_4 FILLER_43_197 ();
 sg13g2_fill_2 FILLER_43_201 ();
 sg13g2_fill_2 FILLER_43_211 ();
 sg13g2_fill_1 FILLER_43_218 ();
 sg13g2_fill_1 FILLER_43_224 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_fill_1 FILLER_43_235 ();
 sg13g2_decap_4 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_277 ();
 sg13g2_fill_1 FILLER_43_302 ();
 sg13g2_fill_1 FILLER_43_344 ();
 sg13g2_fill_2 FILLER_43_356 ();
 sg13g2_fill_2 FILLER_43_364 ();
 sg13g2_fill_1 FILLER_43_366 ();
 sg13g2_decap_4 FILLER_43_371 ();
 sg13g2_fill_1 FILLER_43_375 ();
 sg13g2_fill_1 FILLER_43_381 ();
 sg13g2_fill_2 FILLER_43_398 ();
 sg13g2_fill_1 FILLER_43_400 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_fill_2 FILLER_43_414 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_40 ();
 sg13g2_fill_2 FILLER_44_46 ();
 sg13g2_fill_1 FILLER_44_54 ();
 sg13g2_fill_2 FILLER_44_169 ();
 sg13g2_fill_2 FILLER_44_208 ();
 sg13g2_fill_1 FILLER_44_210 ();
 sg13g2_fill_1 FILLER_44_216 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_fill_2 FILLER_44_226 ();
 sg13g2_fill_1 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_250 ();
 sg13g2_fill_2 FILLER_44_294 ();
 sg13g2_decap_4 FILLER_44_329 ();
 sg13g2_decap_4 FILLER_44_371 ();
 sg13g2_fill_1 FILLER_44_375 ();
 sg13g2_fill_1 FILLER_44_381 ();
 sg13g2_fill_2 FILLER_44_409 ();
 sg13g2_fill_1 FILLER_44_424 ();
 sg13g2_fill_2 FILLER_45_15 ();
 sg13g2_fill_2 FILLER_45_21 ();
 sg13g2_fill_1 FILLER_45_23 ();
 sg13g2_fill_2 FILLER_45_44 ();
 sg13g2_fill_2 FILLER_45_67 ();
 sg13g2_fill_1 FILLER_45_90 ();
 sg13g2_fill_2 FILLER_45_138 ();
 sg13g2_fill_1 FILLER_45_166 ();
 sg13g2_fill_1 FILLER_45_197 ();
 sg13g2_fill_1 FILLER_45_205 ();
 sg13g2_fill_1 FILLER_45_246 ();
 sg13g2_decap_4 FILLER_45_303 ();
 sg13g2_fill_1 FILLER_45_321 ();
 sg13g2_fill_2 FILLER_45_327 ();
 sg13g2_decap_4 FILLER_45_342 ();
 sg13g2_fill_2 FILLER_45_346 ();
 sg13g2_fill_2 FILLER_45_356 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_fill_2 FILLER_45_381 ();
 sg13g2_fill_1 FILLER_45_383 ();
 sg13g2_fill_1 FILLER_45_410 ();
 sg13g2_decap_4 FILLER_45_426 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_8 ();
 sg13g2_fill_1 FILLER_46_19 ();
 sg13g2_fill_2 FILLER_46_69 ();
 sg13g2_fill_2 FILLER_46_117 ();
 sg13g2_fill_2 FILLER_46_169 ();
 sg13g2_fill_1 FILLER_46_175 ();
 sg13g2_fill_2 FILLER_46_180 ();
 sg13g2_fill_1 FILLER_46_182 ();
 sg13g2_fill_2 FILLER_46_217 ();
 sg13g2_fill_2 FILLER_46_232 ();
 sg13g2_fill_2 FILLER_46_238 ();
 sg13g2_fill_2 FILLER_46_248 ();
 sg13g2_fill_1 FILLER_46_290 ();
 sg13g2_fill_1 FILLER_46_300 ();
 sg13g2_fill_1 FILLER_46_309 ();
 sg13g2_fill_1 FILLER_46_369 ();
 sg13g2_fill_1 FILLER_46_375 ();
 sg13g2_fill_2 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_395 ();
 sg13g2_fill_1 FILLER_46_400 ();
 sg13g2_fill_2 FILLER_46_427 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_10 ();
 sg13g2_fill_2 FILLER_47_17 ();
 sg13g2_fill_1 FILLER_47_19 ();
 sg13g2_fill_1 FILLER_47_73 ();
 sg13g2_fill_1 FILLER_47_91 ();
 sg13g2_fill_1 FILLER_47_118 ();
 sg13g2_fill_2 FILLER_47_138 ();
 sg13g2_decap_4 FILLER_47_170 ();
 sg13g2_fill_1 FILLER_47_174 ();
 sg13g2_decap_4 FILLER_47_183 ();
 sg13g2_fill_2 FILLER_47_195 ();
 sg13g2_fill_1 FILLER_47_197 ();
 sg13g2_decap_4 FILLER_47_202 ();
 sg13g2_fill_1 FILLER_47_206 ();
 sg13g2_fill_1 FILLER_47_234 ();
 sg13g2_fill_1 FILLER_47_251 ();
 sg13g2_fill_2 FILLER_47_279 ();
 sg13g2_fill_2 FILLER_47_289 ();
 sg13g2_fill_1 FILLER_47_300 ();
 sg13g2_fill_2 FILLER_47_315 ();
 sg13g2_fill_1 FILLER_47_353 ();
 sg13g2_fill_1 FILLER_47_358 ();
 sg13g2_fill_1 FILLER_47_362 ();
 sg13g2_fill_1 FILLER_47_379 ();
 sg13g2_fill_2 FILLER_47_385 ();
 sg13g2_fill_2 FILLER_47_391 ();
 sg13g2_fill_1 FILLER_47_398 ();
 sg13g2_fill_1 FILLER_47_412 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_12 ();
 sg13g2_fill_1 FILLER_48_14 ();
 sg13g2_fill_2 FILLER_48_27 ();
 sg13g2_fill_1 FILLER_48_33 ();
 sg13g2_fill_1 FILLER_48_38 ();
 sg13g2_fill_1 FILLER_48_137 ();
 sg13g2_fill_2 FILLER_48_151 ();
 sg13g2_fill_1 FILLER_48_206 ();
 sg13g2_fill_1 FILLER_48_217 ();
 sg13g2_fill_1 FILLER_48_223 ();
 sg13g2_fill_1 FILLER_48_228 ();
 sg13g2_decap_4 FILLER_48_234 ();
 sg13g2_fill_2 FILLER_48_289 ();
 sg13g2_fill_1 FILLER_48_291 ();
 sg13g2_fill_1 FILLER_48_332 ();
 sg13g2_fill_2 FILLER_48_342 ();
 sg13g2_fill_1 FILLER_48_344 ();
 sg13g2_fill_2 FILLER_48_349 ();
 sg13g2_fill_1 FILLER_48_359 ();
 sg13g2_fill_1 FILLER_48_372 ();
 sg13g2_fill_1 FILLER_48_381 ();
 sg13g2_fill_2 FILLER_48_405 ();
 sg13g2_fill_1 FILLER_48_407 ();
 sg13g2_decap_4 FILLER_48_411 ();
 sg13g2_fill_1 FILLER_48_415 ();
 sg13g2_decap_4 FILLER_48_425 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_fill_1 FILLER_49_15 ();
 sg13g2_fill_1 FILLER_49_31 ();
 sg13g2_fill_2 FILLER_49_47 ();
 sg13g2_fill_1 FILLER_49_74 ();
 sg13g2_fill_1 FILLER_49_85 ();
 sg13g2_fill_2 FILLER_49_160 ();
 sg13g2_fill_1 FILLER_49_162 ();
 sg13g2_fill_1 FILLER_49_167 ();
 sg13g2_fill_1 FILLER_49_172 ();
 sg13g2_fill_1 FILLER_49_177 ();
 sg13g2_fill_2 FILLER_49_182 ();
 sg13g2_fill_1 FILLER_49_188 ();
 sg13g2_fill_1 FILLER_49_192 ();
 sg13g2_fill_1 FILLER_49_218 ();
 sg13g2_decap_4 FILLER_49_227 ();
 sg13g2_fill_1 FILLER_49_231 ();
 sg13g2_fill_2 FILLER_49_250 ();
 sg13g2_fill_1 FILLER_49_255 ();
 sg13g2_fill_2 FILLER_49_261 ();
 sg13g2_fill_2 FILLER_49_267 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_275 ();
 sg13g2_fill_1 FILLER_49_290 ();
 sg13g2_decap_4 FILLER_49_301 ();
 sg13g2_fill_1 FILLER_49_313 ();
 sg13g2_fill_2 FILLER_49_318 ();
 sg13g2_fill_1 FILLER_49_346 ();
 sg13g2_fill_2 FILLER_49_351 ();
 sg13g2_decap_4 FILLER_49_363 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_fill_1 FILLER_49_373 ();
 sg13g2_fill_1 FILLER_49_378 ();
 sg13g2_fill_2 FILLER_49_383 ();
 sg13g2_fill_1 FILLER_49_391 ();
 sg13g2_fill_2 FILLER_49_396 ();
 sg13g2_fill_2 FILLER_49_402 ();
 sg13g2_fill_2 FILLER_49_413 ();
 sg13g2_decap_4 FILLER_49_426 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_19 ();
 sg13g2_fill_1 FILLER_50_29 ();
 sg13g2_fill_1 FILLER_50_46 ();
 sg13g2_fill_1 FILLER_50_71 ();
 sg13g2_fill_1 FILLER_50_147 ();
 sg13g2_fill_2 FILLER_50_194 ();
 sg13g2_fill_2 FILLER_50_214 ();
 sg13g2_decap_4 FILLER_50_220 ();
 sg13g2_fill_1 FILLER_50_224 ();
 sg13g2_fill_1 FILLER_50_314 ();
 sg13g2_decap_4 FILLER_50_318 ();
 sg13g2_fill_1 FILLER_50_326 ();
 sg13g2_fill_2 FILLER_50_331 ();
 sg13g2_fill_2 FILLER_50_339 ();
 sg13g2_fill_2 FILLER_50_353 ();
 sg13g2_fill_1 FILLER_50_355 ();
 sg13g2_fill_2 FILLER_50_381 ();
 sg13g2_fill_1 FILLER_50_383 ();
 sg13g2_fill_1 FILLER_50_389 ();
 sg13g2_fill_1 FILLER_50_400 ();
 sg13g2_fill_1 FILLER_50_405 ();
 sg13g2_fill_1 FILLER_50_410 ();
 sg13g2_decap_8 FILLER_50_423 ();
 sg13g2_fill_2 FILLER_51_18 ();
 sg13g2_fill_1 FILLER_51_41 ();
 sg13g2_fill_1 FILLER_51_46 ();
 sg13g2_fill_1 FILLER_51_63 ();
 sg13g2_fill_1 FILLER_51_67 ();
 sg13g2_fill_1 FILLER_51_91 ();
 sg13g2_fill_2 FILLER_51_126 ();
 sg13g2_fill_2 FILLER_51_173 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_decap_4 FILLER_51_180 ();
 sg13g2_fill_2 FILLER_51_184 ();
 sg13g2_fill_1 FILLER_51_192 ();
 sg13g2_fill_1 FILLER_51_198 ();
 sg13g2_fill_2 FILLER_51_221 ();
 sg13g2_fill_2 FILLER_51_233 ();
 sg13g2_fill_2 FILLER_51_239 ();
 sg13g2_decap_8 FILLER_51_245 ();
 sg13g2_fill_2 FILLER_51_294 ();
 sg13g2_fill_1 FILLER_51_296 ();
 sg13g2_fill_2 FILLER_51_318 ();
 sg13g2_fill_2 FILLER_51_387 ();
 sg13g2_fill_1 FILLER_51_396 ();
 sg13g2_fill_1 FILLER_51_420 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_fill_1 FILLER_52_29 ();
 sg13g2_fill_1 FILLER_52_37 ();
 sg13g2_fill_1 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_60 ();
 sg13g2_fill_2 FILLER_52_81 ();
 sg13g2_fill_2 FILLER_52_109 ();
 sg13g2_fill_1 FILLER_52_120 ();
 sg13g2_fill_2 FILLER_52_156 ();
 sg13g2_fill_2 FILLER_52_163 ();
 sg13g2_fill_1 FILLER_52_165 ();
 sg13g2_fill_2 FILLER_52_194 ();
 sg13g2_fill_1 FILLER_52_202 ();
 sg13g2_fill_2 FILLER_52_207 ();
 sg13g2_fill_1 FILLER_52_257 ();
 sg13g2_decap_4 FILLER_52_266 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_fill_1 FILLER_52_280 ();
 sg13g2_fill_2 FILLER_52_297 ();
 sg13g2_fill_1 FILLER_52_299 ();
 sg13g2_fill_2 FILLER_52_313 ();
 sg13g2_fill_1 FILLER_52_315 ();
 sg13g2_fill_1 FILLER_52_342 ();
 sg13g2_decap_4 FILLER_52_374 ();
 sg13g2_fill_2 FILLER_52_394 ();
 sg13g2_decap_8 FILLER_52_421 ();
 sg13g2_fill_2 FILLER_52_428 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_21 ();
 sg13g2_fill_1 FILLER_53_42 ();
 sg13g2_fill_2 FILLER_53_57 ();
 sg13g2_fill_1 FILLER_53_88 ();
 sg13g2_fill_1 FILLER_53_182 ();
 sg13g2_fill_2 FILLER_53_228 ();
 sg13g2_fill_2 FILLER_53_270 ();
 sg13g2_fill_1 FILLER_53_272 ();
 sg13g2_fill_1 FILLER_53_286 ();
 sg13g2_fill_2 FILLER_53_333 ();
 sg13g2_fill_2 FILLER_53_342 ();
 sg13g2_fill_1 FILLER_53_344 ();
 sg13g2_fill_1 FILLER_53_375 ();
 sg13g2_fill_2 FILLER_53_384 ();
 sg13g2_fill_1 FILLER_53_389 ();
 sg13g2_decap_8 FILLER_53_394 ();
 sg13g2_fill_1 FILLER_53_401 ();
 sg13g2_fill_2 FILLER_53_410 ();
 sg13g2_fill_1 FILLER_53_412 ();
 sg13g2_decap_4 FILLER_53_418 ();
 sg13g2_fill_1 FILLER_54_41 ();
 sg13g2_fill_2 FILLER_54_61 ();
 sg13g2_decap_4 FILLER_54_71 ();
 sg13g2_fill_1 FILLER_54_96 ();
 sg13g2_fill_1 FILLER_54_110 ();
 sg13g2_fill_1 FILLER_54_116 ();
 sg13g2_fill_1 FILLER_54_129 ();
 sg13g2_fill_2 FILLER_54_134 ();
 sg13g2_fill_1 FILLER_54_178 ();
 sg13g2_fill_1 FILLER_54_193 ();
 sg13g2_fill_2 FILLER_54_204 ();
 sg13g2_fill_1 FILLER_54_206 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_1 FILLER_54_225 ();
 sg13g2_fill_1 FILLER_54_234 ();
 sg13g2_fill_2 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_246 ();
 sg13g2_fill_1 FILLER_54_269 ();
 sg13g2_fill_2 FILLER_54_306 ();
 sg13g2_fill_1 FILLER_54_317 ();
 sg13g2_fill_2 FILLER_54_343 ();
 sg13g2_fill_1 FILLER_54_345 ();
 sg13g2_fill_2 FILLER_54_358 ();
 sg13g2_fill_1 FILLER_54_360 ();
 sg13g2_fill_2 FILLER_54_364 ();
 sg13g2_fill_1 FILLER_54_366 ();
 sg13g2_fill_1 FILLER_54_375 ();
 sg13g2_fill_1 FILLER_54_380 ();
 sg13g2_fill_2 FILLER_54_385 ();
 sg13g2_fill_2 FILLER_54_390 ();
 sg13g2_fill_2 FILLER_54_409 ();
 sg13g2_fill_1 FILLER_54_415 ();
 sg13g2_fill_2 FILLER_54_427 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_fill_2 FILLER_55_25 ();
 sg13g2_fill_2 FILLER_55_148 ();
 sg13g2_fill_1 FILLER_55_150 ();
 sg13g2_fill_1 FILLER_55_216 ();
 sg13g2_fill_1 FILLER_55_243 ();
 sg13g2_decap_4 FILLER_55_274 ();
 sg13g2_fill_1 FILLER_55_325 ();
 sg13g2_fill_1 FILLER_55_343 ();
 sg13g2_fill_2 FILLER_55_352 ();
 sg13g2_fill_1 FILLER_55_359 ();
 sg13g2_fill_2 FILLER_55_368 ();
 sg13g2_fill_1 FILLER_55_388 ();
 sg13g2_fill_1 FILLER_56_47 ();
 sg13g2_fill_2 FILLER_56_52 ();
 sg13g2_fill_1 FILLER_56_63 ();
 sg13g2_fill_2 FILLER_56_71 ();
 sg13g2_fill_1 FILLER_56_81 ();
 sg13g2_fill_2 FILLER_56_86 ();
 sg13g2_fill_1 FILLER_56_96 ();
 sg13g2_fill_2 FILLER_56_106 ();
 sg13g2_fill_1 FILLER_56_116 ();
 sg13g2_fill_2 FILLER_56_133 ();
 sg13g2_fill_1 FILLER_56_135 ();
 sg13g2_fill_1 FILLER_56_141 ();
 sg13g2_fill_1 FILLER_56_172 ();
 sg13g2_fill_1 FILLER_56_204 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_fill_2 FILLER_56_228 ();
 sg13g2_fill_1 FILLER_56_235 ();
 sg13g2_fill_1 FILLER_56_270 ();
 sg13g2_decap_4 FILLER_56_292 ();
 sg13g2_fill_1 FILLER_56_302 ();
 sg13g2_fill_1 FILLER_56_308 ();
 sg13g2_fill_1 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_344 ();
 sg13g2_fill_1 FILLER_56_353 ();
 sg13g2_fill_2 FILLER_56_359 ();
 sg13g2_fill_1 FILLER_56_366 ();
 sg13g2_fill_1 FILLER_56_371 ();
 sg13g2_fill_1 FILLER_56_388 ();
 sg13g2_decap_4 FILLER_56_393 ();
 sg13g2_fill_1 FILLER_56_397 ();
 sg13g2_decap_8 FILLER_56_411 ();
 sg13g2_fill_1 FILLER_56_418 ();
 sg13g2_fill_2 FILLER_57_4 ();
 sg13g2_fill_1 FILLER_57_40 ();
 sg13g2_fill_1 FILLER_57_46 ();
 sg13g2_fill_1 FILLER_57_73 ();
 sg13g2_fill_2 FILLER_57_79 ();
 sg13g2_fill_1 FILLER_57_112 ();
 sg13g2_fill_1 FILLER_57_120 ();
 sg13g2_fill_2 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_216 ();
 sg13g2_fill_1 FILLER_57_245 ();
 sg13g2_fill_2 FILLER_57_250 ();
 sg13g2_fill_1 FILLER_57_252 ();
 sg13g2_fill_2 FILLER_57_256 ();
 sg13g2_fill_1 FILLER_57_258 ();
 sg13g2_fill_1 FILLER_57_264 ();
 sg13g2_fill_1 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_279 ();
 sg13g2_fill_2 FILLER_57_285 ();
 sg13g2_fill_2 FILLER_57_325 ();
 sg13g2_fill_1 FILLER_57_335 ();
 sg13g2_fill_2 FILLER_57_344 ();
 sg13g2_decap_4 FILLER_57_350 ();
 sg13g2_fill_2 FILLER_57_362 ();
 sg13g2_decap_4 FILLER_57_369 ();
 sg13g2_decap_8 FILLER_57_415 ();
 sg13g2_fill_2 FILLER_57_422 ();
 sg13g2_fill_2 FILLER_57_428 ();
 sg13g2_fill_1 FILLER_58_18 ();
 sg13g2_fill_1 FILLER_58_23 ();
 sg13g2_fill_1 FILLER_58_32 ();
 sg13g2_fill_1 FILLER_58_37 ();
 sg13g2_fill_1 FILLER_58_93 ();
 sg13g2_fill_2 FILLER_58_154 ();
 sg13g2_fill_1 FILLER_58_164 ();
 sg13g2_fill_1 FILLER_58_169 ();
 sg13g2_fill_2 FILLER_58_185 ();
 sg13g2_fill_1 FILLER_58_277 ();
 sg13g2_fill_1 FILLER_58_328 ();
 sg13g2_fill_1 FILLER_58_356 ();
 sg13g2_fill_1 FILLER_58_362 ();
 sg13g2_fill_1 FILLER_58_368 ();
 sg13g2_fill_1 FILLER_58_372 ();
 sg13g2_fill_1 FILLER_58_377 ();
 sg13g2_fill_1 FILLER_58_382 ();
 sg13g2_fill_2 FILLER_58_388 ();
 sg13g2_fill_1 FILLER_58_398 ();
 sg13g2_fill_2 FILLER_58_402 ();
 sg13g2_fill_2 FILLER_58_409 ();
 sg13g2_decap_4 FILLER_58_416 ();
 sg13g2_fill_1 FILLER_59_38 ();
 sg13g2_fill_1 FILLER_59_42 ();
 sg13g2_fill_1 FILLER_59_48 ();
 sg13g2_fill_2 FILLER_59_54 ();
 sg13g2_decap_4 FILLER_59_156 ();
 sg13g2_fill_2 FILLER_59_191 ();
 sg13g2_fill_2 FILLER_59_222 ();
 sg13g2_fill_2 FILLER_59_229 ();
 sg13g2_fill_1 FILLER_59_231 ();
 sg13g2_fill_1 FILLER_59_240 ();
 sg13g2_fill_1 FILLER_59_244 ();
 sg13g2_fill_1 FILLER_59_250 ();
 sg13g2_fill_2 FILLER_59_255 ();
 sg13g2_fill_1 FILLER_59_261 ();
 sg13g2_fill_2 FILLER_59_266 ();
 sg13g2_fill_2 FILLER_59_280 ();
 sg13g2_fill_1 FILLER_59_358 ();
 sg13g2_fill_1 FILLER_59_367 ();
 sg13g2_fill_1 FILLER_59_372 ();
 sg13g2_fill_2 FILLER_59_390 ();
 sg13g2_fill_2 FILLER_59_396 ();
 sg13g2_fill_1 FILLER_59_398 ();
 sg13g2_fill_2 FILLER_59_408 ();
 sg13g2_fill_1 FILLER_59_410 ();
 sg13g2_fill_1 FILLER_59_419 ();
 sg13g2_fill_1 FILLER_60_30 ();
 sg13g2_fill_1 FILLER_60_101 ();
 sg13g2_decap_4 FILLER_60_121 ();
 sg13g2_fill_1 FILLER_60_151 ();
 sg13g2_fill_2 FILLER_60_155 ();
 sg13g2_fill_1 FILLER_60_157 ();
 sg13g2_fill_2 FILLER_60_166 ();
 sg13g2_fill_1 FILLER_60_168 ();
 sg13g2_fill_1 FILLER_60_198 ();
 sg13g2_fill_1 FILLER_60_203 ();
 sg13g2_fill_2 FILLER_60_208 ();
 sg13g2_fill_2 FILLER_60_213 ();
 sg13g2_fill_1 FILLER_60_215 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_fill_2 FILLER_60_250 ();
 sg13g2_fill_2 FILLER_60_312 ();
 sg13g2_fill_1 FILLER_60_327 ();
 sg13g2_fill_1 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_337 ();
 sg13g2_fill_2 FILLER_60_342 ();
 sg13g2_fill_2 FILLER_60_349 ();
 sg13g2_fill_2 FILLER_60_373 ();
 sg13g2_fill_2 FILLER_60_379 ();
 sg13g2_fill_2 FILLER_60_386 ();
 sg13g2_fill_1 FILLER_60_388 ();
 sg13g2_decap_4 FILLER_60_414 ();
 sg13g2_fill_1 FILLER_60_418 ();
 sg13g2_fill_1 FILLER_60_424 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_39 ();
 sg13g2_fill_2 FILLER_61_144 ();
 sg13g2_fill_1 FILLER_61_146 ();
 sg13g2_fill_2 FILLER_61_167 ();
 sg13g2_fill_1 FILLER_61_169 ();
 sg13g2_fill_2 FILLER_61_174 ();
 sg13g2_fill_1 FILLER_61_176 ();
 sg13g2_fill_2 FILLER_61_229 ();
 sg13g2_fill_1 FILLER_61_279 ();
 sg13g2_fill_2 FILLER_61_311 ();
 sg13g2_fill_1 FILLER_61_374 ();
 sg13g2_fill_1 FILLER_61_387 ();
 sg13g2_fill_2 FILLER_61_392 ();
 sg13g2_fill_1 FILLER_61_417 ();
 sg13g2_decap_4 FILLER_61_426 ();
 sg13g2_fill_1 FILLER_62_22 ();
 sg13g2_fill_1 FILLER_62_34 ();
 sg13g2_fill_1 FILLER_62_53 ();
 sg13g2_fill_2 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_168 ();
 sg13g2_fill_1 FILLER_62_172 ();
 sg13g2_fill_1 FILLER_62_178 ();
 sg13g2_fill_2 FILLER_62_183 ();
 sg13g2_fill_2 FILLER_62_189 ();
 sg13g2_fill_2 FILLER_62_195 ();
 sg13g2_fill_1 FILLER_62_197 ();
 sg13g2_fill_1 FILLER_62_203 ();
 sg13g2_fill_1 FILLER_62_230 ();
 sg13g2_fill_1 FILLER_62_239 ();
 sg13g2_fill_1 FILLER_62_244 ();
 sg13g2_fill_2 FILLER_62_281 ();
 sg13g2_fill_1 FILLER_62_288 ();
 sg13g2_decap_4 FILLER_62_330 ();
 sg13g2_fill_1 FILLER_62_347 ();
 sg13g2_fill_1 FILLER_62_353 ();
 sg13g2_fill_1 FILLER_62_362 ();
 sg13g2_fill_1 FILLER_62_401 ();
 sg13g2_fill_2 FILLER_62_427 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_24 ();
 sg13g2_fill_1 FILLER_63_96 ();
 sg13g2_fill_1 FILLER_63_137 ();
 sg13g2_fill_1 FILLER_63_157 ();
 sg13g2_fill_2 FILLER_63_220 ();
 sg13g2_fill_1 FILLER_63_245 ();
 sg13g2_decap_4 FILLER_63_250 ();
 sg13g2_fill_2 FILLER_63_254 ();
 sg13g2_decap_4 FILLER_63_317 ();
 sg13g2_decap_8 FILLER_63_325 ();
 sg13g2_decap_8 FILLER_63_332 ();
 sg13g2_fill_1 FILLER_63_370 ();
 sg13g2_fill_2 FILLER_63_375 ();
 sg13g2_fill_1 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_63_397 ();
 sg13g2_fill_1 FILLER_63_413 ();
 sg13g2_fill_2 FILLER_63_428 ();
 sg13g2_fill_1 FILLER_64_51 ();
 sg13g2_fill_1 FILLER_64_56 ();
 sg13g2_fill_1 FILLER_64_62 ();
 sg13g2_fill_1 FILLER_64_77 ();
 sg13g2_fill_1 FILLER_64_92 ();
 sg13g2_fill_1 FILLER_64_101 ();
 sg13g2_fill_1 FILLER_64_107 ();
 sg13g2_fill_1 FILLER_64_113 ();
 sg13g2_fill_2 FILLER_64_118 ();
 sg13g2_fill_1 FILLER_64_165 ();
 sg13g2_fill_1 FILLER_64_170 ();
 sg13g2_fill_1 FILLER_64_180 ();
 sg13g2_fill_2 FILLER_64_192 ();
 sg13g2_fill_1 FILLER_64_272 ();
 sg13g2_fill_2 FILLER_64_291 ();
 sg13g2_decap_8 FILLER_64_328 ();
 sg13g2_fill_1 FILLER_64_335 ();
 sg13g2_fill_2 FILLER_64_340 ();
 sg13g2_fill_1 FILLER_64_342 ();
 sg13g2_fill_2 FILLER_64_350 ();
 sg13g2_fill_1 FILLER_64_352 ();
 sg13g2_fill_2 FILLER_64_357 ();
 sg13g2_fill_1 FILLER_64_359 ();
 sg13g2_fill_1 FILLER_64_364 ();
 sg13g2_fill_2 FILLER_64_386 ();
 sg13g2_fill_1 FILLER_64_388 ();
 sg13g2_fill_2 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_427 ();
 sg13g2_fill_1 FILLER_64_429 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_40 ();
 sg13g2_fill_1 FILLER_65_50 ();
 sg13g2_fill_2 FILLER_65_94 ();
 sg13g2_fill_1 FILLER_65_145 ();
 sg13g2_fill_1 FILLER_65_149 ();
 sg13g2_fill_1 FILLER_65_173 ();
 sg13g2_fill_2 FILLER_65_179 ();
 sg13g2_fill_1 FILLER_65_249 ();
 sg13g2_fill_1 FILLER_65_262 ();
 sg13g2_decap_4 FILLER_65_267 ();
 sg13g2_fill_2 FILLER_65_271 ();
 sg13g2_fill_2 FILLER_65_282 ();
 sg13g2_fill_1 FILLER_65_296 ();
 sg13g2_fill_1 FILLER_65_335 ();
 sg13g2_fill_2 FILLER_65_344 ();
 sg13g2_decap_4 FILLER_65_374 ();
 sg13g2_fill_2 FILLER_65_404 ();
 sg13g2_fill_2 FILLER_65_419 ();
 sg13g2_fill_1 FILLER_65_421 ();
 sg13g2_decap_4 FILLER_65_426 ();
 sg13g2_fill_1 FILLER_66_94 ();
 sg13g2_fill_1 FILLER_66_175 ();
 sg13g2_fill_2 FILLER_66_180 ();
 sg13g2_fill_1 FILLER_66_186 ();
 sg13g2_fill_1 FILLER_66_192 ();
 sg13g2_fill_1 FILLER_66_219 ();
 sg13g2_fill_2 FILLER_66_224 ();
 sg13g2_fill_1 FILLER_66_226 ();
 sg13g2_fill_2 FILLER_66_231 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_fill_2 FILLER_66_242 ();
 sg13g2_fill_1 FILLER_66_290 ();
 sg13g2_fill_1 FILLER_66_295 ();
 sg13g2_fill_1 FILLER_66_336 ();
 sg13g2_fill_2 FILLER_66_357 ();
 sg13g2_fill_1 FILLER_66_389 ();
 sg13g2_fill_1 FILLER_66_398 ();
 sg13g2_fill_1 FILLER_66_404 ();
 sg13g2_fill_2 FILLER_66_411 ();
 sg13g2_fill_2 FILLER_66_417 ();
 sg13g2_fill_1 FILLER_66_419 ();
 sg13g2_fill_2 FILLER_66_428 ();
 sg13g2_fill_1 FILLER_67_31 ();
 sg13g2_fill_1 FILLER_67_39 ();
 sg13g2_fill_1 FILLER_67_105 ();
 sg13g2_fill_1 FILLER_67_114 ();
 sg13g2_fill_1 FILLER_67_119 ();
 sg13g2_fill_1 FILLER_67_124 ();
 sg13g2_fill_1 FILLER_67_135 ();
 sg13g2_fill_1 FILLER_67_141 ();
 sg13g2_fill_1 FILLER_67_148 ();
 sg13g2_fill_1 FILLER_67_154 ();
 sg13g2_fill_1 FILLER_67_159 ();
 sg13g2_fill_1 FILLER_67_168 ();
 sg13g2_fill_2 FILLER_67_216 ();
 sg13g2_fill_1 FILLER_67_218 ();
 sg13g2_fill_2 FILLER_67_310 ();
 sg13g2_fill_2 FILLER_67_316 ();
 sg13g2_fill_2 FILLER_67_322 ();
 sg13g2_fill_1 FILLER_67_324 ();
 sg13g2_fill_1 FILLER_67_330 ();
 sg13g2_fill_2 FILLER_67_335 ();
 sg13g2_fill_1 FILLER_67_337 ();
 sg13g2_fill_2 FILLER_67_381 ();
 sg13g2_fill_2 FILLER_67_427 ();
 sg13g2_fill_1 FILLER_67_429 ();
 sg13g2_fill_1 FILLER_68_19 ();
 sg13g2_fill_2 FILLER_68_64 ();
 sg13g2_decap_8 FILLER_68_234 ();
 sg13g2_fill_1 FILLER_68_241 ();
 sg13g2_fill_2 FILLER_68_246 ();
 sg13g2_fill_1 FILLER_68_298 ();
 sg13g2_fill_1 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_336 ();
 sg13g2_fill_1 FILLER_68_348 ();
 sg13g2_fill_2 FILLER_68_355 ();
 sg13g2_fill_2 FILLER_68_366 ();
 sg13g2_fill_1 FILLER_68_368 ();
 sg13g2_fill_1 FILLER_68_376 ();
 sg13g2_fill_1 FILLER_68_380 ();
 sg13g2_fill_2 FILLER_68_412 ();
 sg13g2_fill_2 FILLER_68_427 ();
 sg13g2_fill_1 FILLER_68_429 ();
 sg13g2_fill_1 FILLER_69_34 ();
 sg13g2_fill_2 FILLER_69_90 ();
 sg13g2_fill_1 FILLER_69_109 ();
 sg13g2_fill_1 FILLER_69_115 ();
 sg13g2_fill_1 FILLER_69_120 ();
 sg13g2_fill_1 FILLER_69_126 ();
 sg13g2_fill_2 FILLER_69_136 ();
 sg13g2_fill_1 FILLER_69_159 ();
 sg13g2_fill_1 FILLER_69_218 ();
 sg13g2_decap_8 FILLER_69_223 ();
 sg13g2_decap_8 FILLER_69_230 ();
 sg13g2_fill_2 FILLER_69_245 ();
 sg13g2_fill_1 FILLER_69_247 ();
 sg13g2_fill_2 FILLER_69_253 ();
 sg13g2_fill_2 FILLER_69_297 ();
 sg13g2_fill_1 FILLER_69_320 ();
 sg13g2_fill_2 FILLER_69_344 ();
 sg13g2_fill_2 FILLER_69_350 ();
 sg13g2_fill_2 FILLER_69_356 ();
 sg13g2_decap_4 FILLER_69_366 ();
 sg13g2_fill_2 FILLER_69_370 ();
 sg13g2_decap_8 FILLER_69_380 ();
 sg13g2_fill_2 FILLER_69_387 ();
 sg13g2_fill_1 FILLER_69_403 ();
 sg13g2_fill_1 FILLER_69_412 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_fill_1 FILLER_70_68 ();
 sg13g2_fill_2 FILLER_70_87 ();
 sg13g2_fill_2 FILLER_70_97 ();
 sg13g2_fill_1 FILLER_70_126 ();
 sg13g2_fill_1 FILLER_70_170 ();
 sg13g2_fill_1 FILLER_70_175 ();
 sg13g2_fill_1 FILLER_70_207 ();
 sg13g2_fill_1 FILLER_70_248 ();
 sg13g2_fill_2 FILLER_70_263 ();
 sg13g2_fill_2 FILLER_70_274 ();
 sg13g2_fill_1 FILLER_70_321 ();
 sg13g2_fill_1 FILLER_70_326 ();
 sg13g2_fill_1 FILLER_70_332 ();
 sg13g2_fill_1 FILLER_70_337 ();
 sg13g2_fill_1 FILLER_70_346 ();
 sg13g2_fill_1 FILLER_70_357 ();
 sg13g2_fill_1 FILLER_70_365 ();
 sg13g2_fill_2 FILLER_70_370 ();
 sg13g2_decap_4 FILLER_70_384 ();
 sg13g2_fill_1 FILLER_70_388 ();
 sg13g2_fill_2 FILLER_70_394 ();
 sg13g2_fill_2 FILLER_70_404 ();
 sg13g2_fill_1 FILLER_70_406 ();
 sg13g2_fill_2 FILLER_70_415 ();
 sg13g2_fill_1 FILLER_70_417 ();
 sg13g2_fill_1 FILLER_71_40 ();
 sg13g2_fill_1 FILLER_71_49 ();
 sg13g2_fill_1 FILLER_71_55 ();
 sg13g2_fill_1 FILLER_71_85 ();
 sg13g2_fill_1 FILLER_71_97 ();
 sg13g2_fill_2 FILLER_71_143 ();
 sg13g2_fill_2 FILLER_71_179 ();
 sg13g2_fill_2 FILLER_71_236 ();
 sg13g2_fill_1 FILLER_71_238 ();
 sg13g2_fill_1 FILLER_71_247 ();
 sg13g2_fill_1 FILLER_71_261 ();
 sg13g2_fill_1 FILLER_71_271 ();
 sg13g2_fill_1 FILLER_71_305 ();
 sg13g2_fill_1 FILLER_71_311 ();
 sg13g2_fill_1 FILLER_71_362 ();
 sg13g2_fill_2 FILLER_71_374 ();
 sg13g2_fill_1 FILLER_71_376 ();
 sg13g2_fill_2 FILLER_71_390 ();
 sg13g2_fill_2 FILLER_71_419 ();
 sg13g2_decap_4 FILLER_71_426 ();
 sg13g2_fill_1 FILLER_72_5 ();
 sg13g2_fill_1 FILLER_72_19 ();
 sg13g2_fill_2 FILLER_72_126 ();
 sg13g2_fill_1 FILLER_72_195 ();
 sg13g2_fill_1 FILLER_72_207 ();
 sg13g2_fill_1 FILLER_72_218 ();
 sg13g2_fill_2 FILLER_72_223 ();
 sg13g2_fill_2 FILLER_72_230 ();
 sg13g2_fill_2 FILLER_72_237 ();
 sg13g2_fill_2 FILLER_72_259 ();
 sg13g2_fill_2 FILLER_72_329 ();
 sg13g2_fill_1 FILLER_72_331 ();
 sg13g2_fill_2 FILLER_72_337 ();
 sg13g2_fill_1 FILLER_72_339 ();
 sg13g2_fill_2 FILLER_72_349 ();
 sg13g2_fill_1 FILLER_72_355 ();
 sg13g2_fill_2 FILLER_72_361 ();
 sg13g2_fill_2 FILLER_72_366 ();
 sg13g2_decap_4 FILLER_72_381 ();
 sg13g2_fill_1 FILLER_72_388 ();
 sg13g2_fill_1 FILLER_72_394 ();
 sg13g2_fill_1 FILLER_72_399 ();
 sg13g2_fill_1 FILLER_72_412 ();
 sg13g2_fill_1 FILLER_72_425 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_85 ();
 sg13g2_fill_1 FILLER_73_96 ();
 sg13g2_fill_2 FILLER_73_175 ();
 sg13g2_fill_1 FILLER_73_181 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_fill_2 FILLER_73_302 ();
 sg13g2_fill_1 FILLER_73_304 ();
 sg13g2_decap_4 FILLER_73_309 ();
 sg13g2_fill_1 FILLER_73_313 ();
 sg13g2_fill_1 FILLER_73_330 ();
 sg13g2_decap_4 FILLER_73_418 ();
 sg13g2_fill_1 FILLER_73_422 ();
 sg13g2_fill_2 FILLER_73_427 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_fill_1 FILLER_74_31 ();
 sg13g2_fill_1 FILLER_74_118 ();
 sg13g2_fill_1 FILLER_74_133 ();
 sg13g2_fill_2 FILLER_74_189 ();
 sg13g2_fill_2 FILLER_74_195 ();
 sg13g2_fill_1 FILLER_74_219 ();
 sg13g2_fill_1 FILLER_74_230 ();
 sg13g2_fill_1 FILLER_74_235 ();
 sg13g2_fill_1 FILLER_74_265 ();
 sg13g2_fill_1 FILLER_74_276 ();
 sg13g2_fill_1 FILLER_74_285 ();
 sg13g2_fill_1 FILLER_74_317 ();
 sg13g2_fill_1 FILLER_74_331 ();
 sg13g2_fill_2 FILLER_74_337 ();
 sg13g2_fill_1 FILLER_74_343 ();
 sg13g2_fill_1 FILLER_74_348 ();
 sg13g2_fill_1 FILLER_74_353 ();
 sg13g2_fill_2 FILLER_74_359 ();
 sg13g2_fill_2 FILLER_74_386 ();
 sg13g2_decap_4 FILLER_74_397 ();
 sg13g2_fill_1 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_411 ();
 sg13g2_decap_4 FILLER_74_426 ();
 sg13g2_fill_1 FILLER_75_32 ();
 sg13g2_fill_1 FILLER_75_39 ();
 sg13g2_fill_1 FILLER_75_46 ();
 sg13g2_fill_2 FILLER_75_69 ();
 sg13g2_fill_2 FILLER_75_87 ();
 sg13g2_fill_2 FILLER_75_111 ();
 sg13g2_fill_2 FILLER_75_122 ();
 sg13g2_fill_1 FILLER_75_219 ();
 sg13g2_fill_1 FILLER_75_224 ();
 sg13g2_fill_2 FILLER_75_235 ();
 sg13g2_fill_2 FILLER_75_267 ();
 sg13g2_fill_1 FILLER_75_333 ();
 sg13g2_fill_1 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_358 ();
 sg13g2_decap_4 FILLER_75_375 ();
 sg13g2_fill_2 FILLER_75_379 ();
 sg13g2_fill_1 FILLER_75_398 ();
 sg13g2_fill_1 FILLER_75_404 ();
 sg13g2_decap_4 FILLER_75_409 ();
 sg13g2_decap_4 FILLER_75_416 ();
 sg13g2_fill_2 FILLER_75_420 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_27 ();
 sg13g2_fill_2 FILLER_76_54 ();
 sg13g2_fill_2 FILLER_76_70 ();
 sg13g2_fill_2 FILLER_76_173 ();
 sg13g2_fill_1 FILLER_76_201 ();
 sg13g2_fill_2 FILLER_76_212 ();
 sg13g2_fill_2 FILLER_76_272 ();
 sg13g2_fill_1 FILLER_76_303 ();
 sg13g2_fill_2 FILLER_76_308 ();
 sg13g2_fill_1 FILLER_76_323 ();
 sg13g2_fill_1 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_344 ();
 sg13g2_decap_4 FILLER_76_351 ();
 sg13g2_decap_4 FILLER_76_359 ();
 sg13g2_fill_2 FILLER_76_363 ();
 sg13g2_fill_1 FILLER_76_369 ();
 sg13g2_fill_1 FILLER_76_374 ();
 sg13g2_decap_8 FILLER_76_383 ();
 sg13g2_fill_1 FILLER_76_398 ();
 sg13g2_fill_1 FILLER_76_403 ();
 sg13g2_fill_1 FILLER_76_425 ();
 sg13g2_fill_2 FILLER_77_128 ();
 sg13g2_fill_1 FILLER_77_142 ();
 sg13g2_fill_1 FILLER_77_173 ();
 sg13g2_fill_1 FILLER_77_244 ();
 sg13g2_fill_1 FILLER_77_254 ();
 sg13g2_fill_1 FILLER_77_297 ();
 sg13g2_fill_1 FILLER_77_302 ();
 sg13g2_fill_1 FILLER_77_317 ();
 sg13g2_fill_1 FILLER_77_323 ();
 sg13g2_fill_2 FILLER_77_358 ();
 sg13g2_decap_4 FILLER_77_365 ();
 sg13g2_fill_2 FILLER_77_369 ();
 sg13g2_fill_1 FILLER_77_384 ();
 sg13g2_fill_2 FILLER_77_390 ();
 sg13g2_fill_2 FILLER_77_409 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_10 ();
 sg13g2_fill_1 FILLER_78_43 ();
 sg13g2_fill_1 FILLER_78_152 ();
 sg13g2_fill_1 FILLER_78_186 ();
 sg13g2_fill_1 FILLER_78_254 ();
 sg13g2_fill_1 FILLER_78_259 ();
 sg13g2_fill_1 FILLER_78_264 ();
 sg13g2_fill_1 FILLER_78_282 ();
 sg13g2_fill_2 FILLER_78_295 ();
 sg13g2_fill_2 FILLER_78_316 ();
 sg13g2_fill_2 FILLER_78_347 ();
 sg13g2_fill_1 FILLER_78_349 ();
 sg13g2_decap_8 FILLER_78_354 ();
 sg13g2_decap_4 FILLER_78_361 ();
 sg13g2_fill_2 FILLER_78_389 ();
 sg13g2_fill_1 FILLER_78_391 ();
 sg13g2_fill_2 FILLER_78_413 ();
 sg13g2_fill_1 FILLER_78_415 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_fill_1 FILLER_79_5 ();
 sg13g2_fill_1 FILLER_79_68 ();
 sg13g2_fill_1 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_145 ();
 sg13g2_fill_1 FILLER_79_158 ();
 sg13g2_fill_1 FILLER_79_167 ();
 sg13g2_fill_2 FILLER_79_279 ();
 sg13g2_fill_1 FILLER_79_289 ();
 sg13g2_fill_2 FILLER_79_316 ();
 sg13g2_fill_2 FILLER_79_323 ();
 sg13g2_fill_2 FILLER_79_330 ();
 sg13g2_fill_1 FILLER_79_332 ();
 sg13g2_fill_1 FILLER_79_337 ();
 sg13g2_fill_2 FILLER_79_343 ();
 sg13g2_fill_1 FILLER_79_345 ();
 sg13g2_fill_2 FILLER_79_380 ();
 sg13g2_fill_1 FILLER_79_392 ();
 sg13g2_fill_2 FILLER_79_409 ();
 sg13g2_fill_2 FILLER_79_417 ();
 sg13g2_fill_1 FILLER_79_419 ();
 sg13g2_decap_8 FILLER_79_423 ();
 sg13g2_fill_2 FILLER_80_82 ();
 sg13g2_fill_2 FILLER_80_184 ();
 sg13g2_fill_2 FILLER_80_318 ();
 sg13g2_decap_8 FILLER_80_324 ();
 sg13g2_decap_4 FILLER_80_331 ();
 sg13g2_decap_8 FILLER_80_352 ();
 sg13g2_decap_4 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_363 ();
 sg13g2_fill_2 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_decap_8 FILLER_80_406 ();
 sg13g2_decap_8 FILLER_80_413 ();
 sg13g2_decap_8 FILLER_80_420 ();
 sg13g2_fill_2 FILLER_80_427 ();
 sg13g2_fill_1 FILLER_80_429 ();
endmodule
