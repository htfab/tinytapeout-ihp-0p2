module tt_um_phansel_laplace_lut (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire clknet_0_clk;
 wire net221;
 wire \chars_remaining[0] ;
 wire \chars_remaining[1] ;
 wire \chars_remaining[2] ;
 wire \chars_remaining[3] ;
 wire \chars_remaining[4] ;
 wire \chars_remaining[5] ;
 wire \chars_remaining[6] ;
 wire \chars_remaining[7] ;
 wire \chars_remaining[8] ;
 wire \chars_remaining[9] ;
 wire clk_buffered;
 wire \clk_picker.clk_slow ;
 wire \clk_picker.counter[0] ;
 wire \clk_picker.counter[10] ;
 wire \clk_picker.counter[11] ;
 wire \clk_picker.counter[12] ;
 wire \clk_picker.counter[13] ;
 wire \clk_picker.counter[14] ;
 wire \clk_picker.counter[15] ;
 wire \clk_picker.counter[16] ;
 wire \clk_picker.counter[17] ;
 wire \clk_picker.counter[18] ;
 wire \clk_picker.counter[19] ;
 wire \clk_picker.counter[1] ;
 wire \clk_picker.counter[20] ;
 wire \clk_picker.counter[21] ;
 wire \clk_picker.counter[22] ;
 wire \clk_picker.counter[23] ;
 wire \clk_picker.counter[24] ;
 wire \clk_picker.counter[25] ;
 wire \clk_picker.counter[2] ;
 wire \clk_picker.counter[3] ;
 wire \clk_picker.counter[4] ;
 wire \clk_picker.counter[5] ;
 wire \clk_picker.counter[6] ;
 wire \clk_picker.counter[7] ;
 wire \clk_picker.counter[8] ;
 wire \clk_picker.counter[9] ;
 wire \line_mapper_1.pointer_addr[0] ;
 wire \line_mapper_1.pointer_addr[10] ;
 wire \line_mapper_1.pointer_addr[11] ;
 wire \line_mapper_1.pointer_addr[12] ;
 wire \line_mapper_1.pointer_addr[13] ;
 wire \line_mapper_1.pointer_addr[14] ;
 wire \line_mapper_1.pointer_addr[15] ;
 wire \line_mapper_1.pointer_addr[1] ;
 wire \line_mapper_1.pointer_addr[2] ;
 wire \line_mapper_1.pointer_addr[3] ;
 wire \line_mapper_1.pointer_addr[4] ;
 wire \line_mapper_1.pointer_addr[5] ;
 wire \line_mapper_1.pointer_addr[6] ;
 wire \line_mapper_1.pointer_addr[7] ;
 wire \line_mapper_1.pointer_addr[8] ;
 wire \line_mapper_1.pointer_addr[9] ;
 wire \mem_addr[0] ;
 wire \mem_addr[1] ;
 wire \mem_addr[2] ;
 wire \mem_addr[3] ;
 wire \mem_addr[4] ;
 wire \mem_addr[5] ;
 wire \mem_addr[6] ;
 wire \mem_addr[7] ;
 wire \mem_addr[8] ;
 wire \memory_1.mem_addr[9] ;
 wire \transformer_1.started ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_level_0_1_10_clk;
 wire clknet_level_1_1_11_clk;
 wire clknet_level_2_1_12_clk;
 wire clknet_level_0_1_23_clk;
 wire clknet_level_1_1_24_clk;
 wire clknet_level_2_1_25_clk;
 wire clknet_level_0_1_36_clk;
 wire clknet_level_1_1_37_clk;
 wire clknet_level_2_1_38_clk;
 wire clknet_level_0_1_49_clk;
 wire clknet_level_1_1_410_clk;
 wire clknet_level_2_1_411_clk;
 wire clknet_0_clk_buffered;
 wire clknet_3_0_0_clk_buffered;
 wire clknet_3_1_0_clk_buffered;
 wire clknet_3_2_0_clk_buffered;
 wire clknet_3_3_0_clk_buffered;
 wire clknet_3_4_0_clk_buffered;
 wire clknet_3_5_0_clk_buffered;
 wire clknet_3_6_0_clk_buffered;
 wire clknet_3_7_0_clk_buffered;

 sg13g2_buf_8 _3120_ (.A(\mem_addr[2] ),
    .X(_0725_));
 sg13g2_inv_2 _3121_ (.Y(_0736_),
    .A(_0725_));
 sg13g2_buf_8 _3122_ (.A(_0736_),
    .X(_0746_));
 sg13g2_buf_8 _3123_ (.A(net190),
    .X(_0757_));
 sg13g2_buf_8 _3124_ (.A(\mem_addr[1] ),
    .X(_0768_));
 sg13g2_inv_4 _3125_ (.A(_0768_),
    .Y(_0779_));
 sg13g2_buf_1 _3126_ (.A(_0779_),
    .X(_0790_));
 sg13g2_nand2_1 _3127_ (.Y(_0801_),
    .A(net158),
    .B(net189));
 sg13g2_buf_2 _3128_ (.A(\mem_addr[3] ),
    .X(_0812_));
 sg13g2_inv_2 _3129_ (.Y(_0823_),
    .A(_0812_));
 sg13g2_buf_8 _3130_ (.A(_0823_),
    .X(_0834_));
 sg13g2_buf_8 _3131_ (.A(net188),
    .X(_0845_));
 sg13g2_buf_8 _3132_ (.A(net157),
    .X(_0856_));
 sg13g2_buf_8 _3133_ (.A(_0725_),
    .X(_0867_));
 sg13g2_buf_8 _3134_ (.A(\mem_addr[0] ),
    .X(_0878_));
 sg13g2_buf_8 _3135_ (.A(_0878_),
    .X(_0889_));
 sg13g2_nand2_1 _3136_ (.Y(_0900_),
    .A(_0867_),
    .B(net207));
 sg13g2_buf_1 _3137_ (.A(_0900_),
    .X(_0910_));
 sg13g2_nand3_1 _3138_ (.B(net111),
    .C(net156),
    .A(_0801_),
    .Y(_0921_));
 sg13g2_buf_2 _3139_ (.A(_0037_),
    .X(_0932_));
 sg13g2_buf_2 _3140_ (.A(_0932_),
    .X(_0943_));
 sg13g2_nor2_1 _3141_ (.A(_0768_),
    .B(_0878_),
    .Y(_0954_));
 sg13g2_buf_2 _3142_ (.A(_0954_),
    .X(_0965_));
 sg13g2_buf_1 _3143_ (.A(_0965_),
    .X(_0976_));
 sg13g2_nor2_2 _3144_ (.A(net206),
    .B(net155),
    .Y(_0987_));
 sg13g2_buf_8 _3145_ (.A(_0812_),
    .X(_0998_));
 sg13g2_buf_8 _3146_ (.A(net205),
    .X(_1009_));
 sg13g2_buf_8 _3147_ (.A(net187),
    .X(_1020_));
 sg13g2_nand2_1 _3148_ (.Y(_1031_),
    .A(_0987_),
    .B(net154));
 sg13g2_buf_2 _3149_ (.A(\mem_addr[4] ),
    .X(_1042_));
 sg13g2_buf_8 _3150_ (.A(\mem_addr[5] ),
    .X(_1053_));
 sg13g2_inv_1 _3151_ (.Y(_1064_),
    .A(_1053_));
 sg13g2_nor2_1 _3152_ (.A(_1042_),
    .B(_1064_),
    .Y(_1074_));
 sg13g2_buf_2 _3153_ (.A(_1074_),
    .X(_1085_));
 sg13g2_inv_2 _3154_ (.Y(_1096_),
    .A(_1085_));
 sg13g2_buf_1 _3155_ (.A(_1096_),
    .X(_1107_));
 sg13g2_a21oi_1 _3156_ (.A1(_0921_),
    .A2(_1031_),
    .Y(_1118_),
    .B1(net64));
 sg13g2_inv_4 _3157_ (.A(_0878_),
    .Y(_1129_));
 sg13g2_nand2_1 _3158_ (.Y(_1140_),
    .A(_0746_),
    .B(_1129_));
 sg13g2_buf_2 _3159_ (.A(_1140_),
    .X(_1151_));
 sg13g2_buf_2 _3160_ (.A(_0032_),
    .X(_1162_));
 sg13g2_nand2_1 _3161_ (.Y(_1173_),
    .A(net208),
    .B(_1162_));
 sg13g2_buf_2 _3162_ (.A(_1173_),
    .X(_1184_));
 sg13g2_nand2_1 _3163_ (.Y(_1195_),
    .A(_1151_),
    .B(_1184_));
 sg13g2_buf_8 _3164_ (.A(_0768_),
    .X(_1205_));
 sg13g2_nor2_2 _3165_ (.A(net208),
    .B(net204),
    .Y(_1216_));
 sg13g2_nor2_2 _3166_ (.A(net205),
    .B(_1216_),
    .Y(_1227_));
 sg13g2_nand2_2 _3167_ (.Y(_1238_),
    .A(_1195_),
    .B(_1227_));
 sg13g2_buf_8 _3168_ (.A(_1205_),
    .X(_1249_));
 sg13g2_buf_8 _3169_ (.A(net207),
    .X(_1260_));
 sg13g2_a21oi_2 _3170_ (.B1(net206),
    .Y(_1271_),
    .A2(net185),
    .A1(net186));
 sg13g2_buf_1 _3171_ (.A(net205),
    .X(_1282_));
 sg13g2_nand2_2 _3172_ (.Y(_1293_),
    .A(_1271_),
    .B(net184));
 sg13g2_nand2_1 _3173_ (.Y(_1304_),
    .A(_1238_),
    .B(_1293_));
 sg13g2_nand2_1 _3174_ (.Y(_1315_),
    .A(_1042_),
    .B(net210));
 sg13g2_buf_2 _3175_ (.A(_1315_),
    .X(_1326_));
 sg13g2_inv_1 _3176_ (.Y(_1336_),
    .A(_1326_));
 sg13g2_buf_1 _3177_ (.A(_1336_),
    .X(_1347_));
 sg13g2_nand2_1 _3178_ (.Y(_1358_),
    .A(_1304_),
    .B(net110));
 sg13g2_buf_1 _3179_ (.A(\mem_addr[6] ),
    .X(_1369_));
 sg13g2_buf_1 _3180_ (.A(net209),
    .X(_1380_));
 sg13g2_nand2_1 _3181_ (.Y(_1391_),
    .A(_1358_),
    .B(net203));
 sg13g2_nor2_1 _3182_ (.A(_1118_),
    .B(_1391_),
    .Y(_1402_));
 sg13g2_xnor2_1 _3183_ (.Y(_1413_),
    .A(net204),
    .B(_0878_));
 sg13g2_buf_8 _3184_ (.A(net208),
    .X(_1424_));
 sg13g2_buf_8 _3185_ (.A(net183),
    .X(_1435_));
 sg13g2_nand2_1 _3186_ (.Y(_1446_),
    .A(_1413_),
    .B(net153));
 sg13g2_inv_1 _3187_ (.Y(_1457_),
    .A(_1162_));
 sg13g2_nor2_1 _3188_ (.A(net208),
    .B(_1457_),
    .Y(_1467_));
 sg13g2_buf_2 _3189_ (.A(_1467_),
    .X(_1478_));
 sg13g2_nor2_1 _3190_ (.A(net157),
    .B(_1478_),
    .Y(_1489_));
 sg13g2_nand2_1 _3191_ (.Y(_1500_),
    .A(_1446_),
    .B(_1489_));
 sg13g2_buf_8 _3192_ (.A(net188),
    .X(_1511_));
 sg13g2_buf_1 _3193_ (.A(net152),
    .X(_1522_));
 sg13g2_inv_2 _3194_ (.Y(_1533_),
    .A(_1042_));
 sg13g2_buf_8 _3195_ (.A(_1533_),
    .X(_1544_));
 sg13g2_buf_1 _3196_ (.A(net182),
    .X(_1555_));
 sg13g2_a21oi_1 _3197_ (.A1(_0987_),
    .A2(net109),
    .Y(_1566_),
    .B1(net151));
 sg13g2_nand2_1 _3198_ (.Y(_1577_),
    .A(_1500_),
    .B(_1566_));
 sg13g2_buf_8 _3199_ (.A(_1129_),
    .X(_1588_));
 sg13g2_nor2_1 _3200_ (.A(_0725_),
    .B(_0779_),
    .Y(_1599_));
 sg13g2_buf_2 _3201_ (.A(_1599_),
    .X(_1609_));
 sg13g2_nor2_1 _3202_ (.A(net181),
    .B(_1609_),
    .Y(_1620_));
 sg13g2_buf_1 _3203_ (.A(_1555_),
    .X(_1631_));
 sg13g2_nand2_1 _3204_ (.Y(_1642_),
    .A(_0812_),
    .B(_0725_));
 sg13g2_buf_2 _3205_ (.A(_1642_),
    .X(_1653_));
 sg13g2_nand3_1 _3206_ (.B(net108),
    .C(_1653_),
    .A(_1620_),
    .Y(_1664_));
 sg13g2_nand2_1 _3207_ (.Y(_1675_),
    .A(_1577_),
    .B(_1664_));
 sg13g2_buf_1 _3208_ (.A(_1064_),
    .X(_1685_));
 sg13g2_buf_1 _3209_ (.A(net180),
    .X(_1696_));
 sg13g2_buf_1 _3210_ (.A(net150),
    .X(_1707_));
 sg13g2_nand2_1 _3211_ (.Y(_1718_),
    .A(_1675_),
    .B(net107));
 sg13g2_nand2_1 _3212_ (.Y(_1729_),
    .A(_1402_),
    .B(_1718_));
 sg13g2_buf_1 _3213_ (.A(_1042_),
    .X(_1740_));
 sg13g2_buf_1 _3214_ (.A(net202),
    .X(_1751_));
 sg13g2_nand2_1 _3215_ (.Y(_1762_),
    .A(_0768_),
    .B(_0878_));
 sg13g2_buf_8 _3216_ (.A(_1762_),
    .X(_1773_));
 sg13g2_nand2_1 _3217_ (.Y(_1784_),
    .A(net178),
    .B(net190));
 sg13g2_buf_2 _3218_ (.A(_1784_),
    .X(_1795_));
 sg13g2_nor2_2 _3219_ (.A(net188),
    .B(_1795_),
    .Y(_1805_));
 sg13g2_nor2_1 _3220_ (.A(net179),
    .B(_1805_),
    .Y(_1816_));
 sg13g2_nand2_1 _3221_ (.Y(_1827_),
    .A(net188),
    .B(net204));
 sg13g2_buf_8 _3222_ (.A(_1827_),
    .X(_1838_));
 sg13g2_inv_4 _3223_ (.A(_0932_),
    .Y(_1848_));
 sg13g2_nand2_2 _3224_ (.Y(_1859_),
    .A(net201),
    .B(net185));
 sg13g2_nor2_2 _3225_ (.A(net106),
    .B(_1859_),
    .Y(_1869_));
 sg13g2_inv_1 _3226_ (.Y(_1880_),
    .A(_1869_));
 sg13g2_nand2_1 _3227_ (.Y(_1890_),
    .A(_1816_),
    .B(_1880_));
 sg13g2_nand2_1 _3228_ (.Y(_1901_),
    .A(_0725_),
    .B(_1205_));
 sg13g2_buf_2 _3229_ (.A(_1901_),
    .X(_1911_));
 sg13g2_nand2_1 _3230_ (.Y(_1921_),
    .A(_1911_),
    .B(net188));
 sg13g2_nor2_1 _3231_ (.A(net185),
    .B(_1921_),
    .Y(_1930_));
 sg13g2_nand2_1 _3232_ (.Y(_1938_),
    .A(_1216_),
    .B(net188));
 sg13g2_buf_2 _3233_ (.A(_1938_),
    .X(_1948_));
 sg13g2_nand2_1 _3234_ (.Y(_1958_),
    .A(_1948_),
    .B(_1740_));
 sg13g2_nor2_2 _3235_ (.A(_1930_),
    .B(_1958_),
    .Y(_1968_));
 sg13g2_inv_1 _3236_ (.Y(_1976_),
    .A(_1968_));
 sg13g2_nand2_1 _3237_ (.Y(_1987_),
    .A(_0998_),
    .B(_1042_));
 sg13g2_buf_4 _3238_ (.X(_1998_),
    .A(_1987_));
 sg13g2_nand3_1 _3239_ (.B(net186),
    .C(net207),
    .A(net183),
    .Y(_2009_));
 sg13g2_buf_2 _3240_ (.A(_2009_),
    .X(_2020_));
 sg13g2_nand2_1 _3241_ (.Y(_2031_),
    .A(_1795_),
    .B(_2020_));
 sg13g2_nor2_1 _3242_ (.A(net209),
    .B(net180),
    .Y(_2042_));
 sg13g2_buf_1 _3243_ (.A(_2042_),
    .X(_2053_));
 sg13g2_o21ai_1 _3244_ (.B1(net105),
    .Y(_2064_),
    .A1(_1998_),
    .A2(_2031_));
 sg13g2_a21oi_1 _3245_ (.A1(_1890_),
    .A2(_1976_),
    .Y(_2075_),
    .B1(_2064_));
 sg13g2_nand2_2 _3246_ (.Y(_2086_),
    .A(_1413_),
    .B(net158));
 sg13g2_nand2_2 _3247_ (.Y(_2097_),
    .A(net178),
    .B(net183));
 sg13g2_nand3_1 _3248_ (.B(net152),
    .C(_2097_),
    .A(_2086_),
    .Y(_2108_));
 sg13g2_buf_2 _3249_ (.A(_2108_),
    .X(_2119_));
 sg13g2_nor2_1 _3250_ (.A(net210),
    .B(_1369_),
    .Y(_2130_));
 sg13g2_buf_2 _3251_ (.A(_2130_),
    .X(_2141_));
 sg13g2_nand2_1 _3252_ (.Y(_2151_),
    .A(_2119_),
    .B(_2141_));
 sg13g2_buf_1 _3253_ (.A(net202),
    .X(_2162_));
 sg13g2_buf_1 _3254_ (.A(net177),
    .X(_2173_));
 sg13g2_nand2_1 _3255_ (.Y(_2183_),
    .A(_0812_),
    .B(_0878_));
 sg13g2_buf_1 _3256_ (.A(_2183_),
    .X(_2193_));
 sg13g2_nor2_2 _3257_ (.A(net153),
    .B(net176),
    .Y(_2203_));
 sg13g2_nand2_1 _3258_ (.Y(_2212_),
    .A(_1216_),
    .B(net205));
 sg13g2_buf_2 _3259_ (.A(_2212_),
    .X(_2221_));
 sg13g2_inv_1 _3260_ (.Y(_2230_),
    .A(_2221_));
 sg13g2_nor2_2 _3261_ (.A(_2203_),
    .B(_2230_),
    .Y(_2239_));
 sg13g2_nand2_1 _3262_ (.Y(_2248_),
    .A(_0779_),
    .B(_0812_));
 sg13g2_buf_1 _3263_ (.A(_2248_),
    .X(_2257_));
 sg13g2_xnor2_1 _3264_ (.Y(_2266_),
    .A(_1424_),
    .B(_0889_));
 sg13g2_buf_2 _3265_ (.A(_2266_),
    .X(_2273_));
 sg13g2_nor2_1 _3266_ (.A(net148),
    .B(_2273_),
    .Y(_2279_));
 sg13g2_nor2_1 _3267_ (.A(net177),
    .B(_2279_),
    .Y(_2289_));
 sg13g2_a21oi_1 _3268_ (.A1(net149),
    .A2(_2239_),
    .Y(_2299_),
    .B1(_2289_));
 sg13g2_nor2_1 _3269_ (.A(_2151_),
    .B(_2299_),
    .Y(_2308_));
 sg13g2_nor2_1 _3270_ (.A(_2075_),
    .B(_2308_),
    .Y(_2317_));
 sg13g2_nand2_1 _3271_ (.Y(_2325_),
    .A(_1729_),
    .B(_2317_));
 sg13g2_buf_1 _3272_ (.A(\mem_addr[7] ),
    .X(_2332_));
 sg13g2_inv_1 _3273_ (.Y(_2341_),
    .A(_2332_));
 sg13g2_buf_1 _3274_ (.A(_2341_),
    .X(_2351_));
 sg13g2_buf_1 _3275_ (.A(net175),
    .X(_2360_));
 sg13g2_nand2_1 _3276_ (.Y(_2369_),
    .A(_2325_),
    .B(net147));
 sg13g2_nor2_1 _3277_ (.A(net209),
    .B(_2341_),
    .Y(_2372_));
 sg13g2_buf_2 _3278_ (.A(_2372_),
    .X(_2373_));
 sg13g2_inv_1 _3279_ (.Y(_2374_),
    .A(_2373_));
 sg13g2_buf_1 _3280_ (.A(_2374_),
    .X(_2375_));
 sg13g2_buf_2 _3281_ (.A(_0036_),
    .X(_2376_));
 sg13g2_nand2_1 _3282_ (.Y(_2377_),
    .A(_0998_),
    .B(_2376_));
 sg13g2_inv_1 _3283_ (.Y(_2378_),
    .A(_2377_));
 sg13g2_nand2_2 _3284_ (.Y(_2379_),
    .A(net178),
    .B(_1848_));
 sg13g2_nor3_1 _3285_ (.A(_2378_),
    .B(net64),
    .C(_2379_),
    .Y(_2380_));
 sg13g2_nor2_1 _3286_ (.A(net210),
    .B(net182),
    .Y(_2381_));
 sg13g2_buf_1 _3287_ (.A(_2381_),
    .X(_2382_));
 sg13g2_inv_2 _3288_ (.Y(_2383_),
    .A(net104));
 sg13g2_buf_2 _3289_ (.A(net62),
    .X(_2384_));
 sg13g2_nand2_1 _3290_ (.Y(_2385_),
    .A(_0812_),
    .B(net204));
 sg13g2_buf_1 _3291_ (.A(_2385_),
    .X(_2386_));
 sg13g2_inv_2 _3292_ (.Y(_2387_),
    .A(net146));
 sg13g2_nor2_1 _3293_ (.A(_2387_),
    .B(_2203_),
    .Y(_2388_));
 sg13g2_nor2_1 _3294_ (.A(net31),
    .B(_2388_),
    .Y(_2389_));
 sg13g2_buf_1 _3295_ (.A(_1326_),
    .X(_2390_));
 sg13g2_nor2_1 _3296_ (.A(net207),
    .B(net190),
    .Y(_2391_));
 sg13g2_buf_2 _3297_ (.A(_2391_),
    .X(_2392_));
 sg13g2_nor2_1 _3298_ (.A(net146),
    .B(_2392_),
    .Y(_2393_));
 sg13g2_nor2_2 _3299_ (.A(_2203_),
    .B(_2393_),
    .Y(_2394_));
 sg13g2_nor2_1 _3300_ (.A(net145),
    .B(_2394_),
    .Y(_2395_));
 sg13g2_nor4_1 _3301_ (.A(_2375_),
    .B(_2380_),
    .C(_2389_),
    .D(_2395_),
    .Y(_2396_));
 sg13g2_inv_1 _3302_ (.Y(_2397_),
    .A(_0038_));
 sg13g2_nor2_1 _3303_ (.A(net208),
    .B(_2397_),
    .Y(_2398_));
 sg13g2_inv_2 _3304_ (.Y(_2399_),
    .A(_2398_));
 sg13g2_nand2_1 _3305_ (.Y(_2400_),
    .A(_2097_),
    .B(net144));
 sg13g2_buf_8 _3306_ (.A(net184),
    .X(_2401_));
 sg13g2_buf_1 _3307_ (.A(net143),
    .X(_2402_));
 sg13g2_nand2_1 _3308_ (.Y(_2403_),
    .A(_2400_),
    .B(net102));
 sg13g2_nor2_1 _3309_ (.A(_1042_),
    .B(net210),
    .Y(_2404_));
 sg13g2_buf_2 _3310_ (.A(_2404_),
    .X(_2405_));
 sg13g2_inv_1 _3311_ (.Y(_2406_),
    .A(_2405_));
 sg13g2_buf_1 _3312_ (.A(_2406_),
    .X(_2407_));
 sg13g2_buf_1 _3313_ (.A(net101),
    .X(_2408_));
 sg13g2_a21o_1 _3314_ (.A2(_1238_),
    .A1(_2403_),
    .B1(net61),
    .X(_2409_));
 sg13g2_nor2_1 _3315_ (.A(_0725_),
    .B(_0878_),
    .Y(_2410_));
 sg13g2_buf_2 _3316_ (.A(_2410_),
    .X(_2411_));
 sg13g2_nand2_1 _3317_ (.Y(_2412_),
    .A(_2411_),
    .B(net189));
 sg13g2_buf_1 _3318_ (.A(_2412_),
    .X(_2413_));
 sg13g2_nand2_1 _3319_ (.Y(_2414_),
    .A(net100),
    .B(_2020_));
 sg13g2_buf_2 _3320_ (.A(net111),
    .X(_2415_));
 sg13g2_buf_1 _3321_ (.A(net60),
    .X(_2416_));
 sg13g2_buf_1 _3322_ (.A(net202),
    .X(_2417_));
 sg13g2_buf_1 _3323_ (.A(net174),
    .X(_2418_));
 sg13g2_buf_1 _3324_ (.A(net142),
    .X(_2419_));
 sg13g2_nand3_1 _3325_ (.B(net30),
    .C(net99),
    .A(_2414_),
    .Y(_2420_));
 sg13g2_nand3_1 _3326_ (.B(_2409_),
    .C(_2420_),
    .A(_2396_),
    .Y(_2421_));
 sg13g2_nand2_1 _3327_ (.Y(_2422_),
    .A(_2369_),
    .B(_2421_));
 sg13g2_buf_2 _3328_ (.A(\mem_addr[8] ),
    .X(_2423_));
 sg13g2_buf_1 _3329_ (.A(_2423_),
    .X(_2424_));
 sg13g2_nand2_1 _3330_ (.Y(_2425_),
    .A(_2422_),
    .B(net200));
 sg13g2_buf_1 _3331_ (.A(net181),
    .X(_2426_));
 sg13g2_nand4_1 _3332_ (.B(_1911_),
    .C(_1511_),
    .A(_0801_),
    .Y(_2427_),
    .D(net141));
 sg13g2_buf_1 _3333_ (.A(_2427_),
    .X(_2428_));
 sg13g2_nor2_1 _3334_ (.A(net146),
    .B(_1859_),
    .Y(_2429_));
 sg13g2_inv_2 _3335_ (.Y(_2430_),
    .A(_2429_));
 sg13g2_a21oi_1 _3336_ (.A1(_2428_),
    .A2(_2430_),
    .Y(_2431_),
    .B1(net101));
 sg13g2_nand2_1 _3337_ (.Y(_2432_),
    .A(net190),
    .B(net204));
 sg13g2_buf_2 _3338_ (.A(_2432_),
    .X(_2433_));
 sg13g2_nand2_1 _3339_ (.Y(_2434_),
    .A(net189),
    .B(net183));
 sg13g2_buf_1 _3340_ (.A(_2434_),
    .X(_2435_));
 sg13g2_nand2_2 _3341_ (.Y(_2436_),
    .A(_2433_),
    .B(net98));
 sg13g2_buf_1 _3342_ (.A(_1282_),
    .X(_2437_));
 sg13g2_nand3_1 _3343_ (.B(net140),
    .C(net141),
    .A(_2436_),
    .Y(_2438_));
 sg13g2_nor2_1 _3344_ (.A(net208),
    .B(net181),
    .Y(_2439_));
 sg13g2_buf_2 _3345_ (.A(_2439_),
    .X(_2440_));
 sg13g2_nor2_2 _3346_ (.A(_0812_),
    .B(net204),
    .Y(_2441_));
 sg13g2_buf_1 _3347_ (.A(_2441_),
    .X(_2442_));
 sg13g2_nand2_1 _3348_ (.Y(_2443_),
    .A(_2440_),
    .B(net139));
 sg13g2_buf_2 _3349_ (.A(_2443_),
    .X(_2444_));
 sg13g2_buf_1 _3350_ (.A(_1326_),
    .X(_2445_));
 sg13g2_a21oi_1 _3351_ (.A1(_2438_),
    .A2(_2444_),
    .Y(_2446_),
    .B1(net138));
 sg13g2_nor2_1 _3352_ (.A(_2431_),
    .B(_2446_),
    .Y(_2447_));
 sg13g2_nand2_1 _3353_ (.Y(_2448_),
    .A(_1424_),
    .B(_0038_));
 sg13g2_buf_1 _3354_ (.A(_2448_),
    .X(_2449_));
 sg13g2_nor2_2 _3355_ (.A(net187),
    .B(net97),
    .Y(_2450_));
 sg13g2_nand2_1 _3356_ (.Y(_2451_),
    .A(_0834_),
    .B(net207));
 sg13g2_buf_1 _3357_ (.A(_2451_),
    .X(_2452_));
 sg13g2_nor2_2 _3358_ (.A(_2433_),
    .B(_2452_),
    .Y(_2453_));
 sg13g2_nor2_1 _3359_ (.A(_2450_),
    .B(_2453_),
    .Y(_2454_));
 sg13g2_inv_1 _3360_ (.Y(_2455_),
    .A(_2393_));
 sg13g2_a21oi_1 _3361_ (.A1(_2454_),
    .A2(_2455_),
    .Y(_2456_),
    .B1(net64));
 sg13g2_inv_2 _3362_ (.Y(_2457_),
    .A(_0965_));
 sg13g2_buf_1 _3363_ (.A(_2457_),
    .X(_2458_));
 sg13g2_nand3_1 _3364_ (.B(net95),
    .C(net104),
    .A(_1805_),
    .Y(_2459_));
 sg13g2_inv_2 _3365_ (.Y(_2460_),
    .A(net209));
 sg13g2_nand2_2 _3366_ (.Y(_2461_),
    .A(net104),
    .B(net157));
 sg13g2_nor2_2 _3367_ (.A(net100),
    .B(_2461_),
    .Y(_2462_));
 sg13g2_nor2_1 _3368_ (.A(_2460_),
    .B(_2462_),
    .Y(_2463_));
 sg13g2_nand2_1 _3369_ (.Y(_2464_),
    .A(_2459_),
    .B(_2463_));
 sg13g2_nor2_1 _3370_ (.A(_2456_),
    .B(_2464_),
    .Y(_2465_));
 sg13g2_nand2_1 _3371_ (.Y(_2466_),
    .A(_2447_),
    .B(_2465_));
 sg13g2_nor2_2 _3372_ (.A(net152),
    .B(net156),
    .Y(_2467_));
 sg13g2_xnor2_1 _3373_ (.Y(_2468_),
    .A(net208),
    .B(net186));
 sg13g2_buf_2 _3374_ (.A(_2468_),
    .X(_2469_));
 sg13g2_nor2_2 _3375_ (.A(net96),
    .B(_2469_),
    .Y(_2470_));
 sg13g2_nor2_1 _3376_ (.A(_2467_),
    .B(_2470_),
    .Y(_2471_));
 sg13g2_nor2_1 _3377_ (.A(net62),
    .B(_2471_),
    .Y(_2472_));
 sg13g2_nand2_1 _3378_ (.Y(_2473_),
    .A(net190),
    .B(net207));
 sg13g2_nand2_1 _3379_ (.Y(_2474_),
    .A(_2473_),
    .B(_0834_));
 sg13g2_buf_1 _3380_ (.A(_2474_),
    .X(_2475_));
 sg13g2_nand2_1 _3381_ (.Y(_2476_),
    .A(_1129_),
    .B(_0725_));
 sg13g2_buf_1 _3382_ (.A(_2476_),
    .X(_2477_));
 sg13g2_nand2_2 _3383_ (.Y(_2478_),
    .A(net137),
    .B(net187));
 sg13g2_nand3_1 _3384_ (.B(_2478_),
    .C(_1085_),
    .A(net59),
    .Y(_2479_));
 sg13g2_buf_1 _3385_ (.A(_2460_),
    .X(_2480_));
 sg13g2_nor2_1 _3386_ (.A(_1042_),
    .B(_2376_),
    .Y(_2481_));
 sg13g2_buf_2 _3387_ (.A(_2481_),
    .X(_2482_));
 sg13g2_nand3_1 _3388_ (.B(net150),
    .C(_2482_),
    .A(_0987_),
    .Y(_2483_));
 sg13g2_nand3_1 _3389_ (.B(net173),
    .C(_2483_),
    .A(_2479_),
    .Y(_2484_));
 sg13g2_nor2_1 _3390_ (.A(_2472_),
    .B(_2484_),
    .Y(_2485_));
 sg13g2_nand2_1 _3391_ (.Y(_2486_),
    .A(_0965_),
    .B(net183));
 sg13g2_buf_2 _3392_ (.A(_2486_),
    .X(_2487_));
 sg13g2_inv_1 _3393_ (.Y(_2488_),
    .A(_1478_));
 sg13g2_nand2_1 _3394_ (.Y(_2489_),
    .A(net94),
    .B(_2488_));
 sg13g2_buf_8 _3395_ (.A(net157),
    .X(_2490_));
 sg13g2_buf_8 _3396_ (.A(net93),
    .X(_2491_));
 sg13g2_nand2_1 _3397_ (.Y(_2492_),
    .A(_2489_),
    .B(_2491_));
 sg13g2_nor2_1 _3398_ (.A(net204),
    .B(_0736_),
    .Y(_2493_));
 sg13g2_buf_2 _3399_ (.A(_2493_),
    .X(_2494_));
 sg13g2_buf_1 _3400_ (.A(net187),
    .X(_2495_));
 sg13g2_nand2_2 _3401_ (.Y(_2496_),
    .A(_2494_),
    .B(net136));
 sg13g2_a21o_1 _3402_ (.A2(_2496_),
    .A1(_2492_),
    .B1(net138),
    .X(_2497_));
 sg13g2_nand2_1 _3403_ (.Y(_2498_),
    .A(_2485_),
    .B(_2497_));
 sg13g2_nand2_1 _3404_ (.Y(_2499_),
    .A(_2466_),
    .B(_2498_));
 sg13g2_nand2_1 _3405_ (.Y(_2500_),
    .A(_2499_),
    .B(net147));
 sg13g2_a21oi_2 _3406_ (.B1(net190),
    .Y(_2501_),
    .A2(net185),
    .A1(net186));
 sg13g2_nand2_1 _3407_ (.Y(_2502_),
    .A(_2501_),
    .B(_2457_));
 sg13g2_buf_1 _3408_ (.A(_2502_),
    .X(_2503_));
 sg13g2_nand2_1 _3409_ (.Y(_2504_),
    .A(net57),
    .B(net100));
 sg13g2_buf_1 _3410_ (.A(net154),
    .X(_2505_));
 sg13g2_buf_1 _3411_ (.A(net92),
    .X(_2506_));
 sg13g2_nand2_1 _3412_ (.Y(_2507_),
    .A(_2504_),
    .B(net56));
 sg13g2_buf_1 _3413_ (.A(net182),
    .X(_2508_));
 sg13g2_buf_1 _3414_ (.A(net135),
    .X(_2509_));
 sg13g2_buf_1 _3415_ (.A(net91),
    .X(_2510_));
 sg13g2_inv_1 _3416_ (.Y(_2511_),
    .A(_1838_));
 sg13g2_buf_1 _3417_ (.A(_2511_),
    .X(_2512_));
 sg13g2_buf_1 _3418_ (.A(_2473_),
    .X(_2513_));
 sg13g2_nand2_1 _3419_ (.Y(_2514_),
    .A(net29),
    .B(net90));
 sg13g2_nand3_1 _3420_ (.B(net55),
    .C(_2514_),
    .A(_2507_),
    .Y(_2515_));
 sg13g2_buf_1 _3421_ (.A(net210),
    .X(_2516_));
 sg13g2_buf_1 _3422_ (.A(net199),
    .X(_2517_));
 sg13g2_buf_1 _3423_ (.A(net135),
    .X(_2518_));
 sg13g2_nor2_2 _3424_ (.A(net187),
    .B(_1911_),
    .Y(_2519_));
 sg13g2_inv_1 _3425_ (.Y(_2520_),
    .A(_1031_));
 sg13g2_nor3_1 _3426_ (.A(net89),
    .B(_2519_),
    .C(_2520_),
    .Y(_2521_));
 sg13g2_nor2_1 _3427_ (.A(net172),
    .B(_2521_),
    .Y(_2522_));
 sg13g2_nand2_1 _3428_ (.Y(_2523_),
    .A(_2515_),
    .B(_2522_));
 sg13g2_nand2_2 _3429_ (.Y(_2524_),
    .A(_0779_),
    .B(_0878_));
 sg13g2_nand2_2 _3430_ (.Y(_2525_),
    .A(_2524_),
    .B(net201));
 sg13g2_nand2_2 _3431_ (.Y(_2526_),
    .A(_2411_),
    .B(net205));
 sg13g2_nand2_1 _3432_ (.Y(_2527_),
    .A(net110),
    .B(net146));
 sg13g2_a21oi_1 _3433_ (.A1(_2525_),
    .A2(_2526_),
    .Y(_2528_),
    .B1(_2527_));
 sg13g2_a21oi_2 _3434_ (.B1(net181),
    .Y(_2529_),
    .A2(net153),
    .A1(net206));
 sg13g2_nand2_2 _3435_ (.Y(_2530_),
    .A(_2529_),
    .B(net29));
 sg13g2_nand3_1 _3436_ (.B(_0867_),
    .C(_1249_),
    .A(_0812_),
    .Y(_2531_));
 sg13g2_buf_2 _3437_ (.A(_2531_),
    .X(_2532_));
 sg13g2_buf_1 _3438_ (.A(_1096_),
    .X(_2533_));
 sg13g2_a21oi_1 _3439_ (.A1(_2530_),
    .A2(_2532_),
    .Y(_2534_),
    .B1(net54));
 sg13g2_nor3_1 _3440_ (.A(net63),
    .B(_2528_),
    .C(_2534_),
    .Y(_2535_));
 sg13g2_inv_1 _3441_ (.Y(_2536_),
    .A(_1958_));
 sg13g2_nor2_1 _3442_ (.A(net157),
    .B(_2379_),
    .Y(_2537_));
 sg13g2_nand2_1 _3443_ (.Y(_2538_),
    .A(_2537_),
    .B(net95));
 sg13g2_nor2_1 _3444_ (.A(net202),
    .B(_2429_),
    .Y(_2539_));
 sg13g2_nor2_1 _3445_ (.A(net96),
    .B(_1609_),
    .Y(_2540_));
 sg13g2_inv_1 _3446_ (.Y(_2541_),
    .A(_2540_));
 sg13g2_nand2_1 _3447_ (.Y(_2542_),
    .A(_2539_),
    .B(_2541_));
 sg13g2_buf_1 _3448_ (.A(_1053_),
    .X(_2543_));
 sg13g2_buf_1 _3449_ (.A(net198),
    .X(_2544_));
 sg13g2_nand2_1 _3450_ (.Y(_2545_),
    .A(_2542_),
    .B(net171));
 sg13g2_a21oi_1 _3451_ (.A1(_2536_),
    .A2(_2538_),
    .Y(_2546_),
    .B1(_2545_));
 sg13g2_nand2_1 _3452_ (.Y(_2547_),
    .A(_2221_),
    .B(net176));
 sg13g2_inv_1 _3453_ (.Y(_2548_),
    .A(_2547_));
 sg13g2_a21oi_1 _3454_ (.A1(net183),
    .A2(net186),
    .Y(_2549_),
    .B1(net205));
 sg13g2_buf_2 _3455_ (.A(_2549_),
    .X(_2550_));
 sg13g2_nand2_1 _3456_ (.Y(_2551_),
    .A(_2550_),
    .B(net100));
 sg13g2_buf_1 _3457_ (.A(_2405_),
    .X(_2552_));
 sg13g2_nand3_1 _3458_ (.B(_2551_),
    .C(net134),
    .A(_2548_),
    .Y(_2553_));
 sg13g2_buf_1 _3459_ (.A(net178),
    .X(_2554_));
 sg13g2_a21oi_1 _3460_ (.A1(net133),
    .A2(net98),
    .Y(_2555_),
    .B1(_2461_));
 sg13g2_inv_1 _3461_ (.Y(_2556_),
    .A(_2555_));
 sg13g2_buf_1 _3462_ (.A(_2332_),
    .X(_2557_));
 sg13g2_nand2_1 _3463_ (.Y(_2558_),
    .A(net209),
    .B(net197));
 sg13g2_inv_2 _3464_ (.Y(_2559_),
    .A(_2558_));
 sg13g2_nand3_1 _3465_ (.B(_2556_),
    .C(_2559_),
    .A(_2553_),
    .Y(_2560_));
 sg13g2_nor2_1 _3466_ (.A(_2546_),
    .B(_2560_),
    .Y(_2561_));
 sg13g2_a21oi_1 _3467_ (.A1(_2523_),
    .A2(_2535_),
    .Y(_2562_),
    .B1(_2561_));
 sg13g2_nand2_1 _3468_ (.Y(_2563_),
    .A(_2500_),
    .B(_2562_));
 sg13g2_inv_2 _3469_ (.Y(_2564_),
    .A(_2423_));
 sg13g2_buf_1 _3470_ (.A(_2564_),
    .X(_2565_));
 sg13g2_buf_2 _3471_ (.A(net170),
    .X(_2566_));
 sg13g2_nand2_1 _3472_ (.Y(_2567_),
    .A(_2563_),
    .B(net132));
 sg13g2_buf_1 _3473_ (.A(_1085_),
    .X(_2568_));
 sg13g2_buf_1 _3474_ (.A(net88),
    .X(_2569_));
 sg13g2_nor2_1 _3475_ (.A(net188),
    .B(_2440_),
    .Y(_2570_));
 sg13g2_buf_2 _3476_ (.A(_2570_),
    .X(_2571_));
 sg13g2_inv_1 _3477_ (.Y(_2572_),
    .A(_2571_));
 sg13g2_nor2_1 _3478_ (.A(_0965_),
    .B(_2097_),
    .Y(_2573_));
 sg13g2_nor2_1 _3479_ (.A(_2572_),
    .B(_2573_),
    .Y(_2574_));
 sg13g2_inv_1 _3480_ (.Y(_2575_),
    .A(net97));
 sg13g2_nor2_1 _3481_ (.A(net208),
    .B(_0965_),
    .Y(_2576_));
 sg13g2_buf_2 _3482_ (.A(_2576_),
    .X(_2577_));
 sg13g2_o21ai_1 _3483_ (.B1(net60),
    .Y(_2578_),
    .A1(_2575_),
    .A2(_2577_));
 sg13g2_buf_1 _3484_ (.A(_2578_),
    .X(_2579_));
 sg13g2_nand2b_1 _3485_ (.Y(_2580_),
    .B(_2579_),
    .A_N(_2574_));
 sg13g2_nand2_1 _3486_ (.Y(_2581_),
    .A(net90),
    .B(net137));
 sg13g2_buf_2 _3487_ (.A(_2581_),
    .X(_2582_));
 sg13g2_buf_1 _3488_ (.A(_0801_),
    .X(_2583_));
 sg13g2_nor2_1 _3489_ (.A(net189),
    .B(_0900_),
    .Y(_2584_));
 sg13g2_nor2_2 _3490_ (.A(net93),
    .B(_2584_),
    .Y(_2585_));
 sg13g2_a22oi_1 _3491_ (.Y(_2586_),
    .B1(net52),
    .B2(_2585_),
    .A2(net139),
    .A1(_2582_));
 sg13g2_nor2_1 _3492_ (.A(net145),
    .B(_2586_),
    .Y(_2587_));
 sg13g2_a21oi_1 _3493_ (.A1(net53),
    .A2(_2580_),
    .Y(_2588_),
    .B1(_2587_));
 sg13g2_buf_1 _3494_ (.A(_0856_),
    .X(_2589_));
 sg13g2_nand2_1 _3495_ (.Y(_2590_),
    .A(_2273_),
    .B(net51));
 sg13g2_nand2_2 _3496_ (.Y(_2591_),
    .A(net103),
    .B(_2411_));
 sg13g2_nand2_1 _3497_ (.Y(_2592_),
    .A(_2590_),
    .B(_2591_));
 sg13g2_buf_1 _3498_ (.A(net104),
    .X(_2593_));
 sg13g2_nand2_1 _3499_ (.Y(_2594_),
    .A(_2592_),
    .B(net50));
 sg13g2_buf_2 _3500_ (.A(net203),
    .X(_2595_));
 sg13g2_buf_1 _3501_ (.A(net169),
    .X(_2596_));
 sg13g2_nand2_2 _3502_ (.Y(_2597_),
    .A(net197),
    .B(_2423_));
 sg13g2_inv_2 _3503_ (.Y(_2598_),
    .A(_2597_));
 sg13g2_nand3_1 _3504_ (.B(net131),
    .C(_2598_),
    .A(_2594_),
    .Y(_2599_));
 sg13g2_buf_1 _3505_ (.A(net198),
    .X(_2600_));
 sg13g2_buf_1 _3506_ (.A(net168),
    .X(_2601_));
 sg13g2_nor2_1 _3507_ (.A(net143),
    .B(net98),
    .Y(_2602_));
 sg13g2_buf_1 _3508_ (.A(_1911_),
    .X(_2603_));
 sg13g2_nand2_1 _3509_ (.Y(_2604_),
    .A(_1489_),
    .B(net87));
 sg13g2_nand2_2 _3510_ (.Y(_2605_),
    .A(_2411_),
    .B(net93));
 sg13g2_nand3_1 _3511_ (.B(net135),
    .C(_2605_),
    .A(_2604_),
    .Y(_2606_));
 sg13g2_nor3_1 _3512_ (.A(net130),
    .B(_2602_),
    .C(_2606_),
    .Y(_2607_));
 sg13g2_nor2_1 _3513_ (.A(_2599_),
    .B(_2607_),
    .Y(_2608_));
 sg13g2_buf_1 _3514_ (.A(\memory_1.mem_addr[9] ),
    .X(_2609_));
 sg13g2_buf_1 _3515_ (.A(_2609_),
    .X(_2610_));
 sg13g2_a21oi_1 _3516_ (.A1(_2588_),
    .A2(_2608_),
    .Y(_2611_),
    .B1(net196));
 sg13g2_nand3_1 _3517_ (.B(_2567_),
    .C(_2611_),
    .A(_2425_),
    .Y(_2612_));
 sg13g2_a21oi_2 _3518_ (.B1(_1609_),
    .Y(_2613_),
    .A2(net153),
    .A1(_0976_));
 sg13g2_nand2_1 _3519_ (.Y(_2614_),
    .A(_2613_),
    .B(_2571_));
 sg13g2_buf_1 _3520_ (.A(net104),
    .X(_2615_));
 sg13g2_nor2_2 _3521_ (.A(net187),
    .B(_2469_),
    .Y(_2616_));
 sg13g2_inv_1 _3522_ (.Y(_2617_),
    .A(_2616_));
 sg13g2_nand3_1 _3523_ (.B(net49),
    .C(_2617_),
    .A(_2614_),
    .Y(_2618_));
 sg13g2_buf_1 _3524_ (.A(net203),
    .X(_2619_));
 sg13g2_nand2_1 _3525_ (.Y(_2620_),
    .A(_2618_),
    .B(net167));
 sg13g2_nand2_1 _3526_ (.Y(_2621_),
    .A(_2577_),
    .B(net178));
 sg13g2_buf_2 _3527_ (.A(_2621_),
    .X(_2622_));
 sg13g2_nand2_1 _3528_ (.Y(_2623_),
    .A(net137),
    .B(net188));
 sg13g2_inv_1 _3529_ (.Y(_2624_),
    .A(_2623_));
 sg13g2_nand2_1 _3530_ (.Y(_2625_),
    .A(_2622_),
    .B(_2624_));
 sg13g2_buf_2 _3531_ (.A(_2405_),
    .X(_2626_));
 sg13g2_nand2_1 _3532_ (.Y(_2627_),
    .A(_1653_),
    .B(_2193_));
 sg13g2_buf_1 _3533_ (.A(_2627_),
    .X(_2628_));
 sg13g2_inv_1 _3534_ (.Y(_2629_),
    .A(_2628_));
 sg13g2_nand3_1 _3535_ (.B(net129),
    .C(_2629_),
    .A(_2625_),
    .Y(_2630_));
 sg13g2_nor2b_1 _3536_ (.A(_2620_),
    .B_N(_2630_),
    .Y(_2631_));
 sg13g2_nor2_1 _3537_ (.A(_0932_),
    .B(net207),
    .Y(_2632_));
 sg13g2_buf_2 _3538_ (.A(_2632_),
    .X(_2633_));
 sg13g2_inv_2 _3539_ (.Y(_2634_),
    .A(_2633_));
 sg13g2_nor2_2 _3540_ (.A(net148),
    .B(_2634_),
    .Y(_2635_));
 sg13g2_nor2_1 _3541_ (.A(_0932_),
    .B(_1588_),
    .Y(_2636_));
 sg13g2_nand2_2 _3542_ (.Y(_2637_),
    .A(_2636_),
    .B(_2441_));
 sg13g2_inv_1 _3543_ (.Y(_2638_),
    .A(_2637_));
 sg13g2_nor2_1 _3544_ (.A(_2635_),
    .B(_2638_),
    .Y(_2639_));
 sg13g2_inv_1 _3545_ (.Y(_2640_),
    .A(_2639_));
 sg13g2_nand2_2 _3546_ (.Y(_2641_),
    .A(net184),
    .B(net210));
 sg13g2_nand2_2 _3547_ (.Y(_2642_),
    .A(_2637_),
    .B(net202));
 sg13g2_nand2_1 _3548_ (.Y(_2643_),
    .A(_2642_),
    .B(net199));
 sg13g2_o21ai_1 _3549_ (.B1(_2643_),
    .Y(_2644_),
    .A1(_2641_),
    .A2(_2613_));
 sg13g2_o21ai_1 _3550_ (.B1(_2644_),
    .Y(_2645_),
    .A1(net99),
    .A2(_2640_));
 sg13g2_buf_1 _3551_ (.A(net197),
    .X(_2646_));
 sg13g2_a21oi_1 _3552_ (.A1(_2631_),
    .A2(_2645_),
    .Y(_2647_),
    .B1(net166));
 sg13g2_nor2_1 _3553_ (.A(net205),
    .B(_2411_),
    .Y(_2648_));
 sg13g2_buf_1 _3554_ (.A(_2648_),
    .X(_2649_));
 sg13g2_nand2_1 _3555_ (.Y(_2650_),
    .A(net85),
    .B(_2634_));
 sg13g2_nand2_1 _3556_ (.Y(_2651_),
    .A(net86),
    .B(_2433_));
 sg13g2_nand3_1 _3557_ (.B(_2651_),
    .C(net199),
    .A(_2650_),
    .Y(_2652_));
 sg13g2_buf_1 _3558_ (.A(net179),
    .X(_2653_));
 sg13g2_buf_2 _3559_ (.A(net128),
    .X(_2654_));
 sg13g2_nand2_1 _3560_ (.Y(_2655_),
    .A(_2652_),
    .B(net84));
 sg13g2_nand2_1 _3561_ (.Y(_2656_),
    .A(_2622_),
    .B(net143));
 sg13g2_inv_1 _3562_ (.Y(_2657_),
    .A(_2656_));
 sg13g2_nor3_1 _3563_ (.A(net168),
    .B(_2392_),
    .C(_2657_),
    .Y(_2658_));
 sg13g2_nand2_2 _3564_ (.Y(_2659_),
    .A(net155),
    .B(net201));
 sg13g2_inv_1 _3565_ (.Y(_2660_),
    .A(net96));
 sg13g2_nor2_1 _3566_ (.A(net179),
    .B(_2660_),
    .Y(_2661_));
 sg13g2_o21ai_1 _3567_ (.B1(_2661_),
    .Y(_2662_),
    .A1(_2641_),
    .A2(_2659_));
 sg13g2_o21ai_1 _3568_ (.B1(_2662_),
    .Y(_2663_),
    .A1(_2655_),
    .A2(_2658_));
 sg13g2_buf_1 _3569_ (.A(net173),
    .X(_2664_));
 sg13g2_buf_1 _3570_ (.A(net127),
    .X(_2665_));
 sg13g2_nand2_1 _3571_ (.Y(_2666_),
    .A(_2663_),
    .B(net83));
 sg13g2_nand2_1 _3572_ (.Y(_2667_),
    .A(_2647_),
    .B(_2666_));
 sg13g2_nand2_1 _3573_ (.Y(_2668_),
    .A(_1129_),
    .B(net204));
 sg13g2_buf_8 _3574_ (.A(_2668_),
    .X(_2669_));
 sg13g2_nand2_1 _3575_ (.Y(_2670_),
    .A(net126),
    .B(net190));
 sg13g2_buf_2 _3576_ (.A(_2670_),
    .X(_2671_));
 sg13g2_nand3_1 _3577_ (.B(net183),
    .C(_1249_),
    .A(_1588_),
    .Y(_2672_));
 sg13g2_buf_1 _3578_ (.A(_2672_),
    .X(_2673_));
 sg13g2_nand2_1 _3579_ (.Y(_2674_),
    .A(_2671_),
    .B(net82));
 sg13g2_nand2_1 _3580_ (.Y(_2675_),
    .A(net181),
    .B(_0038_));
 sg13g2_nand2_1 _3581_ (.Y(_2676_),
    .A(_0932_),
    .B(net185));
 sg13g2_nand2_1 _3582_ (.Y(_2677_),
    .A(_2675_),
    .B(_2676_));
 sg13g2_nor2_2 _3583_ (.A(net111),
    .B(_2677_),
    .Y(_2678_));
 sg13g2_nor2_1 _3584_ (.A(net99),
    .B(_2678_),
    .Y(_2679_));
 sg13g2_buf_1 _3585_ (.A(net109),
    .X(_2680_));
 sg13g2_nand2_1 _3586_ (.Y(_2681_),
    .A(net48),
    .B(net206));
 sg13g2_buf_1 _3587_ (.A(_2524_),
    .X(_2682_));
 sg13g2_nand2_1 _3588_ (.Y(_2683_),
    .A(net125),
    .B(net126));
 sg13g2_buf_1 _3589_ (.A(_2683_),
    .X(_2684_));
 sg13g2_nand2b_1 _3590_ (.Y(_2685_),
    .B(net47),
    .A_N(_2681_));
 sg13g2_nor2_2 _3591_ (.A(_2376_),
    .B(_1544_),
    .Y(_2686_));
 sg13g2_inv_1 _3592_ (.Y(_2687_),
    .A(_2686_));
 sg13g2_buf_1 _3593_ (.A(net180),
    .X(_2688_));
 sg13g2_buf_1 _3594_ (.A(net124),
    .X(_2689_));
 sg13g2_nand2_1 _3595_ (.Y(_2690_),
    .A(_2332_),
    .B(_0033_));
 sg13g2_inv_1 _3596_ (.Y(_2691_),
    .A(_2690_));
 sg13g2_nand3_1 _3597_ (.B(_2689_),
    .C(_2691_),
    .A(_2687_),
    .Y(_2692_));
 sg13g2_a221oi_1 _3598_ (.B2(_2685_),
    .C1(_2692_),
    .B1(_2679_),
    .A1(net99),
    .Y(_2693_),
    .A2(_2674_));
 sg13g2_nor2_1 _3599_ (.A(net170),
    .B(_2693_),
    .Y(_2694_));
 sg13g2_inv_1 _3600_ (.Y(_2695_),
    .A(_2609_));
 sg13g2_buf_1 _3601_ (.A(net195),
    .X(_2696_));
 sg13g2_a21oi_1 _3602_ (.A1(_2667_),
    .A2(_2694_),
    .Y(_2697_),
    .B1(net165));
 sg13g2_buf_1 _3603_ (.A(net173),
    .X(_2698_));
 sg13g2_buf_1 _3604_ (.A(net123),
    .X(_2699_));
 sg13g2_a21oi_1 _3605_ (.A1(_1238_),
    .A2(_2221_),
    .Y(_2700_),
    .B1(_2390_));
 sg13g2_inv_2 _3606_ (.Y(_2701_),
    .A(_2482_));
 sg13g2_nor2_1 _3607_ (.A(net87),
    .B(_2701_),
    .Y(_2702_));
 sg13g2_inv_1 _3608_ (.Y(_2703_),
    .A(_2702_));
 sg13g2_buf_1 _3609_ (.A(_1413_),
    .X(_2704_));
 sg13g2_nand2_1 _3610_ (.Y(_2705_),
    .A(net122),
    .B(net86));
 sg13g2_nand3_1 _3611_ (.B(net106),
    .C(_2626_),
    .A(_2705_),
    .Y(_2706_));
 sg13g2_o21ai_1 _3612_ (.B1(_2706_),
    .Y(_2707_),
    .A1(_2689_),
    .A2(_2703_));
 sg13g2_nor3_1 _3613_ (.A(net80),
    .B(_2700_),
    .C(_2707_),
    .Y(_2708_));
 sg13g2_nand2_2 _3614_ (.Y(_2709_),
    .A(_2440_),
    .B(net189));
 sg13g2_nand2_2 _3615_ (.Y(_2710_),
    .A(_2709_),
    .B(_2672_));
 sg13g2_buf_1 _3616_ (.A(net154),
    .X(_2711_));
 sg13g2_nand2_1 _3617_ (.Y(_2712_),
    .A(_2710_),
    .B(net79));
 sg13g2_nor2_1 _3618_ (.A(net187),
    .B(_0910_),
    .Y(_2713_));
 sg13g2_nor2_1 _3619_ (.A(net202),
    .B(_2713_),
    .Y(_2714_));
 sg13g2_buf_2 _3620_ (.A(_2714_),
    .X(_2715_));
 sg13g2_buf_1 _3621_ (.A(net124),
    .X(_2716_));
 sg13g2_a21oi_1 _3622_ (.A1(_2712_),
    .A2(_2715_),
    .Y(_2717_),
    .B1(net78));
 sg13g2_nand3_1 _3623_ (.B(net93),
    .C(net141),
    .A(_2469_),
    .Y(_2718_));
 sg13g2_buf_1 _3624_ (.A(_2718_),
    .X(_2719_));
 sg13g2_nand3_1 _3625_ (.B(net84),
    .C(_2705_),
    .A(_2719_),
    .Y(_2720_));
 sg13g2_nand2_1 _3626_ (.Y(_2721_),
    .A(_2717_),
    .B(_2720_));
 sg13g2_nand2_1 _3627_ (.Y(_2722_),
    .A(_2489_),
    .B(net102));
 sg13g2_nor2_2 _3628_ (.A(net106),
    .B(_2634_),
    .Y(_2723_));
 sg13g2_nor2_1 _3629_ (.A(net128),
    .B(_2723_),
    .Y(_2724_));
 sg13g2_nand2_1 _3630_ (.Y(_2725_),
    .A(_2722_),
    .B(_2724_));
 sg13g2_nor2_1 _3631_ (.A(net155),
    .B(_2379_),
    .Y(_2726_));
 sg13g2_nand2_2 _3632_ (.Y(_2727_),
    .A(_2726_),
    .B(_2415_));
 sg13g2_buf_1 _3633_ (.A(net136),
    .X(_2728_));
 sg13g2_buf_1 _3634_ (.A(net151),
    .X(_2729_));
 sg13g2_a21oi_1 _3635_ (.A1(_2494_),
    .A2(net77),
    .Y(_2730_),
    .B1(net76));
 sg13g2_nand2_1 _3636_ (.Y(_2731_),
    .A(_2727_),
    .B(_2730_));
 sg13g2_buf_1 _3637_ (.A(_1696_),
    .X(_2732_));
 sg13g2_buf_1 _3638_ (.A(_2732_),
    .X(_2733_));
 sg13g2_nand3_1 _3639_ (.B(_2731_),
    .C(net46),
    .A(_2725_),
    .Y(_2734_));
 sg13g2_nand3_1 _3640_ (.B(_2734_),
    .C(net80),
    .A(_2721_),
    .Y(_2735_));
 sg13g2_buf_1 _3641_ (.A(_2557_),
    .X(_2736_));
 sg13g2_nand3b_1 _3642_ (.B(_2735_),
    .C(net164),
    .Y(_2737_),
    .A_N(_2708_));
 sg13g2_buf_1 _3643_ (.A(_2564_),
    .X(_2738_));
 sg13g2_inv_1 _3644_ (.Y(_2739_),
    .A(_2526_));
 sg13g2_nor2_1 _3645_ (.A(net76),
    .B(_2739_),
    .Y(_2740_));
 sg13g2_a21oi_1 _3646_ (.A1(_2740_),
    .A2(_1238_),
    .Y(_2741_),
    .B1(net78));
 sg13g2_nand2_1 _3647_ (.Y(_2742_),
    .A(_2221_),
    .B(net135));
 sg13g2_inv_1 _3648_ (.Y(_2743_),
    .A(_2742_));
 sg13g2_nor2_1 _3649_ (.A(net205),
    .B(_2494_),
    .Y(_2744_));
 sg13g2_buf_2 _3650_ (.A(_2744_),
    .X(_2745_));
 sg13g2_nand2_1 _3651_ (.Y(_2746_),
    .A(_2745_),
    .B(net122));
 sg13g2_inv_1 _3652_ (.Y(_2747_),
    .A(_2203_));
 sg13g2_nand3_1 _3653_ (.B(_2746_),
    .C(_2747_),
    .A(_2743_),
    .Y(_2748_));
 sg13g2_buf_1 _3654_ (.A(net169),
    .X(_2749_));
 sg13g2_a21oi_1 _3655_ (.A1(_2741_),
    .A2(_2748_),
    .Y(_2750_),
    .B1(net121));
 sg13g2_inv_2 _3656_ (.Y(_2751_),
    .A(net176));
 sg13g2_nand2_1 _3657_ (.Y(_2752_),
    .A(net52),
    .B(_2751_));
 sg13g2_buf_1 _3658_ (.A(net76),
    .X(_2753_));
 sg13g2_nand2_1 _3659_ (.Y(_2754_),
    .A(_2752_),
    .B(net45));
 sg13g2_nand2_1 _3660_ (.Y(_2755_),
    .A(_2502_),
    .B(_2671_));
 sg13g2_nor2_1 _3661_ (.A(net79),
    .B(_2755_),
    .Y(_2756_));
 sg13g2_inv_1 _3662_ (.Y(_2757_),
    .A(_1805_));
 sg13g2_inv_1 _3663_ (.Y(_2758_),
    .A(net87));
 sg13g2_nor2_1 _3664_ (.A(net91),
    .B(_2758_),
    .Y(_2759_));
 sg13g2_buf_1 _3665_ (.A(net198),
    .X(_2760_));
 sg13g2_a21oi_1 _3666_ (.A1(_2757_),
    .A2(_2759_),
    .Y(_2761_),
    .B1(net162));
 sg13g2_o21ai_1 _3667_ (.B1(_2761_),
    .Y(_2762_),
    .A1(_2754_),
    .A2(_2756_));
 sg13g2_nand2_1 _3668_ (.Y(_2763_),
    .A(_2750_),
    .B(_2762_));
 sg13g2_a21oi_1 _3669_ (.A1(_2571_),
    .A2(net47),
    .Y(_2764_),
    .B1(net149));
 sg13g2_nand2_1 _3670_ (.Y(_2765_),
    .A(net94),
    .B(_2399_));
 sg13g2_nand2_1 _3671_ (.Y(_2766_),
    .A(_2765_),
    .B(net58));
 sg13g2_nand2_1 _3672_ (.Y(_2767_),
    .A(_2764_),
    .B(_2766_));
 sg13g2_nand2_1 _3673_ (.Y(_2768_),
    .A(_1609_),
    .B(net51));
 sg13g2_buf_1 _3674_ (.A(net174),
    .X(_2769_));
 sg13g2_a21oi_1 _3675_ (.A1(_2768_),
    .A2(net120),
    .Y(_2770_),
    .B1(net78));
 sg13g2_nand2_1 _3676_ (.Y(_2771_),
    .A(_2767_),
    .B(_2770_));
 sg13g2_nand2_1 _3677_ (.Y(_2772_),
    .A(_2629_),
    .B(net146));
 sg13g2_nand2_1 _3678_ (.Y(_2773_),
    .A(_2772_),
    .B(net97));
 sg13g2_buf_1 _3679_ (.A(net62),
    .X(_2774_));
 sg13g2_nor2_1 _3680_ (.A(_2711_),
    .B(_2636_),
    .Y(_2775_));
 sg13g2_nor3_1 _3681_ (.A(net139),
    .B(net28),
    .C(_2775_),
    .Y(_2776_));
 sg13g2_a21oi_1 _3682_ (.A1(_2773_),
    .A2(_2776_),
    .Y(_2777_),
    .B1(net127));
 sg13g2_buf_8 _3683_ (.A(_2469_),
    .X(_2778_));
 sg13g2_nand2_2 _3684_ (.Y(_2779_),
    .A(net44),
    .B(net154));
 sg13g2_inv_1 _3685_ (.Y(_2780_),
    .A(_2779_));
 sg13g2_a21oi_1 _3686_ (.A1(_2020_),
    .A2(net144),
    .Y(_2781_),
    .B1(net154));
 sg13g2_buf_1 _3687_ (.A(net134),
    .X(_2782_));
 sg13g2_o21ai_1 _3688_ (.B1(net74),
    .Y(_2783_),
    .A1(_2780_),
    .A2(_2781_));
 sg13g2_nand3_1 _3689_ (.B(_2777_),
    .C(_2783_),
    .A(_2771_),
    .Y(_2784_));
 sg13g2_buf_1 _3690_ (.A(net147),
    .X(_2785_));
 sg13g2_nand3_1 _3691_ (.B(_2784_),
    .C(net73),
    .A(_2763_),
    .Y(_2786_));
 sg13g2_nand3_1 _3692_ (.B(net163),
    .C(_2786_),
    .A(_2737_),
    .Y(_2787_));
 sg13g2_nand2_1 _3693_ (.Y(_2788_),
    .A(_2697_),
    .B(_2787_));
 sg13g2_nand2_1 _3694_ (.Y(_0021_),
    .A(_2612_),
    .B(_2788_));
 sg13g2_nand2_2 _3695_ (.Y(_2789_),
    .A(_2529_),
    .B(_2442_));
 sg13g2_inv_1 _3696_ (.Y(_2790_),
    .A(_2789_));
 sg13g2_nor2_1 _3697_ (.A(net89),
    .B(_2790_),
    .Y(_2791_));
 sg13g2_nand2_1 _3698_ (.Y(_2792_),
    .A(_1609_),
    .B(net181));
 sg13g2_buf_2 _3699_ (.A(_2792_),
    .X(_2793_));
 sg13g2_nand2_1 _3700_ (.Y(_2794_),
    .A(_2494_),
    .B(net207));
 sg13g2_buf_8 _3701_ (.A(_2794_),
    .X(_2795_));
 sg13g2_nand2_1 _3702_ (.Y(_2796_),
    .A(_2793_),
    .B(net43));
 sg13g2_nand2_2 _3703_ (.Y(_2797_),
    .A(_2796_),
    .B(net140));
 sg13g2_a21oi_1 _3704_ (.A1(_2791_),
    .A2(_2797_),
    .Y(_2798_),
    .B1(net81));
 sg13g2_nand2_1 _3705_ (.Y(_2799_),
    .A(_2524_),
    .B(net190));
 sg13g2_buf_2 _3706_ (.A(_2799_),
    .X(_2800_));
 sg13g2_inv_1 _3707_ (.Y(_2801_),
    .A(_2800_));
 sg13g2_nor2_1 _3708_ (.A(_2801_),
    .B(_2573_),
    .Y(_2802_));
 sg13g2_nand2_2 _3709_ (.Y(_2803_),
    .A(_2802_),
    .B(_2415_));
 sg13g2_nand2_1 _3710_ (.Y(_2804_),
    .A(_2803_),
    .B(_2764_));
 sg13g2_nand2_1 _3711_ (.Y(_2805_),
    .A(_2798_),
    .B(_2804_));
 sg13g2_nand2_1 _3712_ (.Y(_2806_),
    .A(net98),
    .B(net133));
 sg13g2_nand2_1 _3713_ (.Y(_2807_),
    .A(_2806_),
    .B(net79));
 sg13g2_buf_1 _3714_ (.A(net186),
    .X(_2808_));
 sg13g2_nand2_1 _3715_ (.Y(_2809_),
    .A(net156),
    .B(net119));
 sg13g2_nand2_1 _3716_ (.Y(_2810_),
    .A(net85),
    .B(_2809_));
 sg13g2_nand2_1 _3717_ (.Y(_2811_),
    .A(_2807_),
    .B(_2810_));
 sg13g2_inv_1 _3718_ (.Y(_2812_),
    .A(net85));
 sg13g2_nand2_1 _3719_ (.Y(_2813_),
    .A(_2751_),
    .B(_1609_));
 sg13g2_o21ai_1 _3720_ (.B1(_2813_),
    .Y(_2814_),
    .A1(net47),
    .A2(_2812_));
 sg13g2_a22oi_1 _3721_ (.Y(_2815_),
    .B1(net50),
    .B2(_2814_),
    .A2(net74),
    .A1(_2811_));
 sg13g2_buf_1 _3722_ (.A(_2558_),
    .X(_2816_));
 sg13g2_a21oi_1 _3723_ (.A1(_2805_),
    .A2(_2815_),
    .Y(_2817_),
    .B1(net118));
 sg13g2_nor2_1 _3724_ (.A(net198),
    .B(_2781_),
    .Y(_2818_));
 sg13g2_a21oi_1 _3725_ (.A1(_1151_),
    .A2(_1184_),
    .Y(_2819_),
    .B1(net152));
 sg13g2_nand2_1 _3726_ (.Y(_2820_),
    .A(_2819_),
    .B(net52));
 sg13g2_nand2_1 _3727_ (.Y(_2821_),
    .A(_2818_),
    .B(_2820_));
 sg13g2_a21oi_1 _3728_ (.A1(net44),
    .A2(_2660_),
    .Y(_2822_),
    .B1(net150));
 sg13g2_a22oi_1 _3729_ (.Y(_2823_),
    .B1(_2392_),
    .B2(net103),
    .A2(net143),
    .A1(_1478_));
 sg13g2_nand2_1 _3730_ (.Y(_2824_),
    .A(_2822_),
    .B(_2823_));
 sg13g2_nand2_1 _3731_ (.Y(_2825_),
    .A(_2821_),
    .B(_2824_));
 sg13g2_buf_2 _3732_ (.A(net149),
    .X(_2826_));
 sg13g2_nand2_1 _3733_ (.Y(_2827_),
    .A(_2825_),
    .B(net72));
 sg13g2_nand2_1 _3734_ (.Y(_2828_),
    .A(_2470_),
    .B(net198));
 sg13g2_nand2_1 _3735_ (.Y(_2829_),
    .A(net206),
    .B(net119));
 sg13g2_nand2_1 _3736_ (.Y(_2830_),
    .A(net125),
    .B(_2829_));
 sg13g2_a21oi_1 _3737_ (.A1(_2830_),
    .A2(net140),
    .Y(_2831_),
    .B1(net177));
 sg13g2_nand2_1 _3738_ (.Y(_2832_),
    .A(_2828_),
    .B(_2831_));
 sg13g2_nand2_1 _3739_ (.Y(_2833_),
    .A(net125),
    .B(net153));
 sg13g2_nand2_1 _3740_ (.Y(_2834_),
    .A(_2709_),
    .B(_2833_));
 sg13g2_nand2_1 _3741_ (.Y(_2835_),
    .A(_2834_),
    .B(net58));
 sg13g2_nor2_1 _3742_ (.A(net199),
    .B(_2835_),
    .Y(_2836_));
 sg13g2_nor2_1 _3743_ (.A(_2832_),
    .B(_2836_),
    .Y(_2837_));
 sg13g2_nor2_1 _3744_ (.A(_2374_),
    .B(_2837_),
    .Y(_2838_));
 sg13g2_nand2_1 _3745_ (.Y(_2839_),
    .A(_2827_),
    .B(_2838_));
 sg13g2_nand2_1 _3746_ (.Y(_2840_),
    .A(_2839_),
    .B(_2423_));
 sg13g2_nor2_1 _3747_ (.A(_2817_),
    .B(_2840_),
    .Y(_2841_));
 sg13g2_inv_2 _3748_ (.Y(_2842_),
    .A(_1998_));
 sg13g2_nand3_1 _3749_ (.B(net87),
    .C(_2842_),
    .A(net122),
    .Y(_2843_));
 sg13g2_buf_1 _3750_ (.A(net58),
    .X(_2844_));
 sg13g2_nand2_1 _3751_ (.Y(_2845_),
    .A(_2400_),
    .B(net27));
 sg13g2_nand2_1 _3752_ (.Y(_2846_),
    .A(_2843_),
    .B(_2845_));
 sg13g2_nor2_1 _3753_ (.A(net119),
    .B(net90),
    .Y(_2847_));
 sg13g2_buf_2 _3754_ (.A(_2847_),
    .X(_2848_));
 sg13g2_o21ai_1 _3755_ (.B1(net140),
    .Y(_2849_),
    .A1(_2575_),
    .A2(_2848_));
 sg13g2_buf_1 _3756_ (.A(_2849_),
    .X(_2850_));
 sg13g2_nor2_1 _3757_ (.A(net120),
    .B(_2850_),
    .Y(_2851_));
 sg13g2_o21ai_1 _3758_ (.B1(net46),
    .Y(_2852_),
    .A1(_2846_),
    .A2(_2851_));
 sg13g2_nand2_1 _3759_ (.Y(_2853_),
    .A(_1859_),
    .B(net152));
 sg13g2_inv_2 _3760_ (.Y(_2854_),
    .A(_2441_));
 sg13g2_nand3_1 _3761_ (.B(net76),
    .C(_2854_),
    .A(_2853_),
    .Y(_2855_));
 sg13g2_nand2_1 _3762_ (.Y(_2856_),
    .A(_2436_),
    .B(net140));
 sg13g2_nand2_1 _3763_ (.Y(_2857_),
    .A(_2856_),
    .B(net199));
 sg13g2_o21ai_1 _3764_ (.B1(net123),
    .Y(_2858_),
    .A1(_2855_),
    .A2(_2857_));
 sg13g2_nand3_1 _3765_ (.B(net186),
    .C(_0889_),
    .A(_0746_),
    .Y(_2859_));
 sg13g2_buf_1 _3766_ (.A(_2859_),
    .X(_2860_));
 sg13g2_nand2_2 _3767_ (.Y(_2861_),
    .A(net71),
    .B(net154));
 sg13g2_o21ai_1 _3768_ (.B1(_2861_),
    .Y(_2862_),
    .A1(net77),
    .A2(_2848_));
 sg13g2_a21oi_1 _3769_ (.A1(_2862_),
    .A2(net97),
    .Y(_2863_),
    .B1(net145));
 sg13g2_nor2_1 _3770_ (.A(_2858_),
    .B(_2863_),
    .Y(_2864_));
 sg13g2_nand2_1 _3771_ (.Y(_2865_),
    .A(_2852_),
    .B(_2864_));
 sg13g2_a21oi_1 _3772_ (.A1(_2634_),
    .A2(net125),
    .Y(_2866_),
    .B1(net154));
 sg13g2_nor2_1 _3773_ (.A(net62),
    .B(_2866_),
    .Y(_2867_));
 sg13g2_nand2_1 _3774_ (.Y(_2868_),
    .A(_2867_),
    .B(_2239_));
 sg13g2_nand2_1 _3775_ (.Y(_2869_),
    .A(net43),
    .B(_2800_));
 sg13g2_nand2_1 _3776_ (.Y(_2870_),
    .A(_2869_),
    .B(net51));
 sg13g2_nor2_2 _3777_ (.A(net157),
    .B(_2392_),
    .Y(_2871_));
 sg13g2_nor2_1 _3778_ (.A(_1326_),
    .B(_2871_),
    .Y(_2872_));
 sg13g2_nand2_1 _3779_ (.Y(_2873_),
    .A(_2870_),
    .B(_2872_));
 sg13g2_nand2_1 _3780_ (.Y(_2874_),
    .A(_2868_),
    .B(_2873_));
 sg13g2_a21oi_1 _3781_ (.A1(_2745_),
    .A2(_2793_),
    .Y(_2875_),
    .B1(_2467_));
 sg13g2_o21ai_1 _3782_ (.B1(net167),
    .Y(_2876_),
    .A1(net54),
    .A2(_2875_));
 sg13g2_nor2_1 _3783_ (.A(_2874_),
    .B(_2876_),
    .Y(_2877_));
 sg13g2_nand2_1 _3784_ (.Y(_2878_),
    .A(_1805_),
    .B(_2457_));
 sg13g2_buf_4 _3785_ (.X(_2879_),
    .A(_2878_));
 sg13g2_inv_4 _3786_ (.A(_2879_),
    .Y(_2880_));
 sg13g2_nor2_1 _3787_ (.A(net56),
    .B(_2504_),
    .Y(_2881_));
 sg13g2_buf_1 _3788_ (.A(net129),
    .X(_2882_));
 sg13g2_o21ai_1 _3789_ (.B1(net70),
    .Y(_2883_),
    .A1(_2880_),
    .A2(_2881_));
 sg13g2_nand2_1 _3790_ (.Y(_2884_),
    .A(_2877_),
    .B(_2883_));
 sg13g2_nand3_1 _3791_ (.B(_2884_),
    .C(net73),
    .A(_2865_),
    .Y(_2885_));
 sg13g2_a21oi_1 _3792_ (.A1(_2841_),
    .A2(_2885_),
    .Y(_2886_),
    .B1(net196));
 sg13g2_nor2_2 _3793_ (.A(net186),
    .B(net181),
    .Y(_2887_));
 sg13g2_nor2_1 _3794_ (.A(_2887_),
    .B(_2671_),
    .Y(_2888_));
 sg13g2_nor2_1 _3795_ (.A(net157),
    .B(_2888_),
    .Y(_2889_));
 sg13g2_nand2_1 _3796_ (.Y(_2890_),
    .A(_2889_),
    .B(net57));
 sg13g2_nor2_1 _3797_ (.A(_1009_),
    .B(_2584_),
    .Y(_2891_));
 sg13g2_buf_2 _3798_ (.A(_2891_),
    .X(_2892_));
 sg13g2_nand2_1 _3799_ (.Y(_2893_),
    .A(_2892_),
    .B(net95));
 sg13g2_nand2_1 _3800_ (.Y(_2894_),
    .A(_2890_),
    .B(_2893_));
 sg13g2_buf_2 _3801_ (.A(net110),
    .X(_2895_));
 sg13g2_nand2_1 _3802_ (.Y(_2896_),
    .A(_2894_),
    .B(net42));
 sg13g2_nand2_1 _3803_ (.Y(_2897_),
    .A(_1271_),
    .B(_2458_));
 sg13g2_a21oi_1 _3804_ (.A1(_2897_),
    .A2(net51),
    .Y(_2898_),
    .B1(_2406_));
 sg13g2_nor2_1 _3805_ (.A(net157),
    .B(_2494_),
    .Y(_2899_));
 sg13g2_buf_2 _3806_ (.A(_2899_),
    .X(_2900_));
 sg13g2_nand2_1 _3807_ (.Y(_2901_),
    .A(_2900_),
    .B(net90));
 sg13g2_nand2_1 _3808_ (.Y(_2902_),
    .A(_2898_),
    .B(_2901_));
 sg13g2_nand2_1 _3809_ (.Y(_2903_),
    .A(_2896_),
    .B(_2902_));
 sg13g2_nand2_1 _3810_ (.Y(_2904_),
    .A(_0845_),
    .B(net202));
 sg13g2_buf_1 _3811_ (.A(_2904_),
    .X(_2905_));
 sg13g2_nor2_1 _3812_ (.A(_2398_),
    .B(_2573_),
    .Y(_2906_));
 sg13g2_o21ai_1 _3813_ (.B1(_2842_),
    .Y(_2907_),
    .A1(_2575_),
    .A2(_2577_));
 sg13g2_o21ai_1 _3814_ (.B1(_2907_),
    .Y(_2908_),
    .A1(net41),
    .A2(_2906_));
 sg13g2_nand2_1 _3815_ (.Y(_2909_),
    .A(_2908_),
    .B(net107));
 sg13g2_nand3_1 _3816_ (.B(net82),
    .C(net111),
    .A(_2671_),
    .Y(_2910_));
 sg13g2_nand2_1 _3817_ (.Y(_2911_),
    .A(_2897_),
    .B(net143));
 sg13g2_nand3_1 _3818_ (.B(_2911_),
    .C(net88),
    .A(_2910_),
    .Y(_2912_));
 sg13g2_nand2_1 _3819_ (.Y(_2913_),
    .A(_2909_),
    .B(_2912_));
 sg13g2_nor2_1 _3820_ (.A(_2903_),
    .B(_2913_),
    .Y(_2914_));
 sg13g2_nor2_1 _3821_ (.A(net63),
    .B(_2914_),
    .Y(_2915_));
 sg13g2_nor2_1 _3822_ (.A(net146),
    .B(_2273_),
    .Y(_2916_));
 sg13g2_nor2_1 _3823_ (.A(net174),
    .B(_2916_),
    .Y(_2917_));
 sg13g2_nand2_1 _3824_ (.Y(_2918_),
    .A(_2803_),
    .B(_2917_));
 sg13g2_a21oi_1 _3825_ (.A1(_2726_),
    .A2(_1020_),
    .Y(_2919_),
    .B1(net151));
 sg13g2_nand2_2 _3826_ (.Y(_2920_),
    .A(_2273_),
    .B(net139));
 sg13g2_nand2_1 _3827_ (.Y(_2921_),
    .A(_2919_),
    .B(_2920_));
 sg13g2_nand3_1 _3828_ (.B(_2921_),
    .C(net168),
    .A(_2918_),
    .Y(_2922_));
 sg13g2_nand2_1 _3829_ (.Y(_2923_),
    .A(_2854_),
    .B(_2508_));
 sg13g2_nor2_1 _3830_ (.A(_2923_),
    .B(_2869_),
    .Y(_2924_));
 sg13g2_a22oi_1 _3831_ (.Y(_2925_),
    .B1(net49),
    .B2(_2756_),
    .A2(_2924_),
    .A1(net107));
 sg13g2_nand2_1 _3832_ (.Y(_2926_),
    .A(_2922_),
    .B(_2925_));
 sg13g2_nand2_1 _3833_ (.Y(_2927_),
    .A(_2926_),
    .B(_2559_));
 sg13g2_nand2_1 _3834_ (.Y(_2928_),
    .A(_2927_),
    .B(net170));
 sg13g2_nor2_1 _3835_ (.A(_2915_),
    .B(_2928_),
    .Y(_2929_));
 sg13g2_o21ai_1 _3836_ (.B1(_2524_),
    .Y(_2930_),
    .A1(net201),
    .A2(net158));
 sg13g2_nor2_1 _3837_ (.A(net93),
    .B(_2930_),
    .Y(_2931_));
 sg13g2_nand2_1 _3838_ (.Y(_2932_),
    .A(_2931_),
    .B(net126));
 sg13g2_nand2_1 _3839_ (.Y(_2933_),
    .A(net85),
    .B(net87));
 sg13g2_a21oi_1 _3840_ (.A1(_2932_),
    .A2(_2933_),
    .Y(_2934_),
    .B1(net145));
 sg13g2_buf_1 _3841_ (.A(_1085_),
    .X(_2935_));
 sg13g2_nor2_1 _3842_ (.A(_1380_),
    .B(net69),
    .Y(_2936_));
 sg13g2_nand2_1 _3843_ (.Y(_2937_),
    .A(_2795_),
    .B(net144));
 sg13g2_nand2_1 _3844_ (.Y(_2938_),
    .A(_2937_),
    .B(_2711_));
 sg13g2_nand3_1 _3845_ (.B(_2428_),
    .C(_2480_),
    .A(_2938_),
    .Y(_2939_));
 sg13g2_nand2b_1 _3846_ (.Y(_2940_),
    .B(_2939_),
    .A_N(_2936_));
 sg13g2_nor2b_1 _3847_ (.A(_2934_),
    .B_N(_2940_),
    .Y(_2941_));
 sg13g2_nand2_1 _3848_ (.Y(_2942_),
    .A(net57),
    .B(_2800_));
 sg13g2_nand2_1 _3849_ (.Y(_2943_),
    .A(_2942_),
    .B(net30));
 sg13g2_nand2_1 _3850_ (.Y(_2944_),
    .A(_2919_),
    .B(_2943_));
 sg13g2_nor2_1 _3851_ (.A(net174),
    .B(_2638_),
    .Y(_2945_));
 sg13g2_nand2_1 _3852_ (.Y(_2946_),
    .A(net126),
    .B(_1848_));
 sg13g2_buf_2 _3853_ (.A(_2946_),
    .X(_2947_));
 sg13g2_nor2_1 _3854_ (.A(net58),
    .B(_2947_),
    .Y(_2948_));
 sg13g2_inv_1 _3855_ (.Y(_2949_),
    .A(_2948_));
 sg13g2_a21oi_1 _3856_ (.A1(_2945_),
    .A2(_2949_),
    .Y(_2950_),
    .B1(net172));
 sg13g2_nand2_1 _3857_ (.Y(_2951_),
    .A(_2944_),
    .B(_2950_));
 sg13g2_a21oi_1 _3858_ (.A1(_2941_),
    .A2(_2951_),
    .Y(_2952_),
    .B1(net164));
 sg13g2_nand2_1 _3859_ (.Y(_2953_),
    .A(net71),
    .B(net94));
 sg13g2_nor2_1 _3860_ (.A(_2416_),
    .B(_2953_),
    .Y(_2954_));
 sg13g2_a21oi_1 _3861_ (.A1(_2503_),
    .A2(_2433_),
    .Y(_2955_),
    .B1(net56));
 sg13g2_o21ai_1 _3862_ (.B1(_2569_),
    .Y(_2956_),
    .A1(_2954_),
    .A2(_2955_));
 sg13g2_buf_1 _3863_ (.A(net167),
    .X(_2957_));
 sg13g2_nor2_1 _3864_ (.A(net184),
    .B(_1795_),
    .Y(_2958_));
 sg13g2_nand2_1 _3865_ (.Y(_2959_),
    .A(_2958_),
    .B(net95));
 sg13g2_nor2_1 _3866_ (.A(net185),
    .B(_1653_),
    .Y(_2960_));
 sg13g2_nor2_1 _3867_ (.A(net103),
    .B(_2960_),
    .Y(_2961_));
 sg13g2_a21o_1 _3868_ (.A2(_2961_),
    .A1(_2959_),
    .B1(net145),
    .X(_2962_));
 sg13g2_buf_1 _3869_ (.A(net101),
    .X(_2963_));
 sg13g2_nand2_1 _3870_ (.Y(_2964_),
    .A(_1911_),
    .B(_1009_));
 sg13g2_inv_1 _3871_ (.Y(_2965_),
    .A(_2964_));
 sg13g2_nor2_1 _3872_ (.A(_2963_),
    .B(_2965_),
    .Y(_2966_));
 sg13g2_nand2_2 _3873_ (.Y(_2967_),
    .A(_2273_),
    .B(_0790_));
 sg13g2_buf_1 _3874_ (.A(net49),
    .X(_2968_));
 sg13g2_nor2_2 _3875_ (.A(_1838_),
    .B(_2392_),
    .Y(_2969_));
 sg13g2_inv_1 _3876_ (.Y(_2970_),
    .A(_2969_));
 sg13g2_nand2_1 _3877_ (.Y(_2971_),
    .A(_2970_),
    .B(net148));
 sg13g2_a22oi_1 _3878_ (.Y(_2972_),
    .B1(net26),
    .B2(_2971_),
    .A2(_2967_),
    .A1(_2966_));
 sg13g2_nand4_1 _3879_ (.B(net117),
    .C(_2962_),
    .A(_2956_),
    .Y(_2973_),
    .D(_2972_));
 sg13g2_nand2_1 _3880_ (.Y(_2974_),
    .A(_2952_),
    .B(_2973_));
 sg13g2_nand2_1 _3881_ (.Y(_2975_),
    .A(_2929_),
    .B(_2974_));
 sg13g2_nand2_1 _3882_ (.Y(_2976_),
    .A(_2886_),
    .B(_2975_));
 sg13g2_a21oi_2 _3883_ (.B1(_2450_),
    .Y(_2977_),
    .A2(net95),
    .A1(_2958_));
 sg13g2_nand2_1 _3884_ (.Y(_2978_),
    .A(_2020_),
    .B(net144));
 sg13g2_nand2_1 _3885_ (.Y(_2979_),
    .A(_2978_),
    .B(net102));
 sg13g2_nand3_1 _3886_ (.B(net84),
    .C(_2979_),
    .A(_2977_),
    .Y(_2980_));
 sg13g2_nor2_1 _3887_ (.A(net176),
    .B(net44),
    .Y(_2981_));
 sg13g2_inv_1 _3888_ (.Y(_2982_),
    .A(_2981_));
 sg13g2_nor2_1 _3889_ (.A(net179),
    .B(_2519_),
    .Y(_2983_));
 sg13g2_a21oi_1 _3890_ (.A1(_2982_),
    .A2(_2983_),
    .Y(_2984_),
    .B1(net162));
 sg13g2_nand2_1 _3891_ (.Y(_2985_),
    .A(_2980_),
    .B(_2984_));
 sg13g2_a21oi_2 _3892_ (.B1(net154),
    .Y(_2986_),
    .A2(net201),
    .A1(net155));
 sg13g2_nor2_1 _3893_ (.A(net54),
    .B(_2986_),
    .Y(_2987_));
 sg13g2_nand2_1 _3894_ (.Y(_2988_),
    .A(net94),
    .B(net90));
 sg13g2_nand2_1 _3895_ (.Y(_2989_),
    .A(_2988_),
    .B(net56));
 sg13g2_buf_2 _3896_ (.A(net110),
    .X(_2990_));
 sg13g2_buf_1 _3897_ (.A(net39),
    .X(_2991_));
 sg13g2_nor2_2 _3898_ (.A(net187),
    .B(_2887_),
    .Y(_2992_));
 sg13g2_nand2_1 _3899_ (.Y(_2993_),
    .A(_2992_),
    .B(net158));
 sg13g2_nand2_1 _3900_ (.Y(_2994_),
    .A(_2993_),
    .B(_2455_));
 sg13g2_a22oi_1 _3901_ (.Y(_2995_),
    .B1(net25),
    .B2(_2994_),
    .A2(_2989_),
    .A1(_2987_));
 sg13g2_a21oi_1 _3902_ (.A1(_2985_),
    .A2(_2995_),
    .Y(_2996_),
    .B1(net63));
 sg13g2_buf_8 _3903_ (.A(_1151_),
    .X(_2997_));
 sg13g2_nor2_2 _3904_ (.A(net106),
    .B(net38),
    .Y(_2998_));
 sg13g2_nor2_1 _3905_ (.A(_2998_),
    .B(_2723_),
    .Y(_2999_));
 sg13g2_nand2_1 _3906_ (.Y(_3000_),
    .A(_2999_),
    .B(_2221_));
 sg13g2_nand2_1 _3907_ (.Y(_3001_),
    .A(_2579_),
    .B(_2979_));
 sg13g2_a22oi_1 _3908_ (.Y(_3002_),
    .B1(net53),
    .B2(_3001_),
    .A2(_3000_),
    .A1(net50));
 sg13g2_nand2_2 _3909_ (.Y(_3003_),
    .A(_1609_),
    .B(net136));
 sg13g2_nand2_1 _3910_ (.Y(_3004_),
    .A(_2530_),
    .B(_3003_));
 sg13g2_nand2_2 _3911_ (.Y(_3005_),
    .A(_1948_),
    .B(net96));
 sg13g2_nor2_1 _3912_ (.A(net40),
    .B(_3005_),
    .Y(_3006_));
 sg13g2_nand2_1 _3913_ (.Y(_3007_),
    .A(_2622_),
    .B(net137));
 sg13g2_nand2_1 _3914_ (.Y(_3008_),
    .A(_3007_),
    .B(net92));
 sg13g2_a22oi_1 _3915_ (.Y(_3009_),
    .B1(_3006_),
    .B2(_3008_),
    .A2(_3004_),
    .A1(net42));
 sg13g2_a21oi_1 _3916_ (.A1(_3002_),
    .A2(_3009_),
    .Y(_3010_),
    .B1(net118));
 sg13g2_nor3_1 _3917_ (.A(net200),
    .B(_2996_),
    .C(_3010_),
    .Y(_3011_));
 sg13g2_nand2_1 _3918_ (.Y(_3012_),
    .A(_2582_),
    .B(net139));
 sg13g2_nor2_2 _3919_ (.A(_0845_),
    .B(_2633_),
    .Y(_3013_));
 sg13g2_nand2_1 _3920_ (.Y(_3014_),
    .A(_2397_),
    .B(net185));
 sg13g2_nand2_1 _3921_ (.Y(_3015_),
    .A(_3013_),
    .B(_3014_));
 sg13g2_a21oi_1 _3922_ (.A1(_3012_),
    .A2(_3015_),
    .Y(_3016_),
    .B1(net61));
 sg13g2_nand3_1 _3923_ (.B(net100),
    .C(net60),
    .A(net82),
    .Y(_3017_));
 sg13g2_nor2_1 _3924_ (.A(net111),
    .B(_1620_),
    .Y(_3018_));
 sg13g2_inv_1 _3925_ (.Y(_3019_),
    .A(_3018_));
 sg13g2_and3_1 _3926_ (.X(_3020_),
    .A(_3017_),
    .B(net50),
    .C(_3019_));
 sg13g2_nor3_1 _3927_ (.A(net121),
    .B(_3016_),
    .C(_3020_),
    .Y(_3021_));
 sg13g2_buf_1 _3928_ (.A(net108),
    .X(_3022_));
 sg13g2_buf_1 _3929_ (.A(net37),
    .X(_3023_));
 sg13g2_nand2_1 _3930_ (.Y(_3024_),
    .A(_2796_),
    .B(net109));
 sg13g2_buf_2 _3931_ (.A(_3024_),
    .X(_3025_));
 sg13g2_nand2_1 _3932_ (.Y(_3026_),
    .A(_2751_),
    .B(net98));
 sg13g2_nand2_1 _3933_ (.Y(_3027_),
    .A(_3025_),
    .B(_3026_));
 sg13g2_nor2_1 _3934_ (.A(net184),
    .B(_2379_),
    .Y(_3028_));
 sg13g2_nor2_2 _3935_ (.A(net148),
    .B(_1151_),
    .Y(_3029_));
 sg13g2_nor2_2 _3936_ (.A(_1740_),
    .B(_3029_),
    .Y(_3030_));
 sg13g2_nand2b_1 _3937_ (.Y(_3031_),
    .B(_3030_),
    .A_N(_2635_));
 sg13g2_nor2_1 _3938_ (.A(_3028_),
    .B(_3031_),
    .Y(_3032_));
 sg13g2_nor2_1 _3939_ (.A(net81),
    .B(_3032_),
    .Y(_3033_));
 sg13g2_o21ai_1 _3940_ (.B1(_3033_),
    .Y(_3034_),
    .A1(net24),
    .A2(_3027_));
 sg13g2_nand2_1 _3941_ (.Y(_3035_),
    .A(_3021_),
    .B(_3034_));
 sg13g2_inv_1 _3942_ (.Y(_3036_),
    .A(_1930_));
 sg13g2_nand3_1 _3943_ (.B(net55),
    .C(_3036_),
    .A(_2850_),
    .Y(_3037_));
 sg13g2_a21oi_1 _3944_ (.A1(_2530_),
    .A2(net120),
    .Y(_3038_),
    .B1(net78));
 sg13g2_buf_1 _3945_ (.A(_2460_),
    .X(_3039_));
 sg13g2_buf_1 _3946_ (.A(net161),
    .X(_3040_));
 sg13g2_a21oi_1 _3947_ (.A1(_3037_),
    .A2(_3038_),
    .Y(_3041_),
    .B1(net116));
 sg13g2_nand2_1 _3948_ (.Y(_3042_),
    .A(_2086_),
    .B(_2745_));
 sg13g2_buf_8 _3949_ (.A(_3042_),
    .X(_3043_));
 sg13g2_nand2_1 _3950_ (.Y(_3044_),
    .A(net44),
    .B(_2751_));
 sg13g2_nand2_1 _3951_ (.Y(_3045_),
    .A(_3043_),
    .B(_3044_));
 sg13g2_a21oi_2 _3952_ (.B1(_2519_),
    .Y(_3046_),
    .A2(_1478_),
    .A1(net111));
 sg13g2_nor2_1 _3953_ (.A(net152),
    .B(_2809_),
    .Y(_3047_));
 sg13g2_inv_1 _3954_ (.Y(_3048_),
    .A(_3047_));
 sg13g2_nand3_1 _3955_ (.B(_3048_),
    .C(_2496_),
    .A(_3046_),
    .Y(_3049_));
 sg13g2_a22oi_1 _3956_ (.Y(_0088_),
    .B1(net70),
    .B2(_3049_),
    .A2(net26),
    .A1(_3045_));
 sg13g2_nand2_1 _3957_ (.Y(_0089_),
    .A(_3041_),
    .B(_0088_));
 sg13g2_buf_2 _3958_ (.A(net147),
    .X(_0090_));
 sg13g2_nand3_1 _3959_ (.B(_0089_),
    .C(net68),
    .A(_3035_),
    .Y(_0091_));
 sg13g2_nand2_1 _3960_ (.Y(_0092_),
    .A(_3011_),
    .B(_0091_));
 sg13g2_nand2_2 _3961_ (.Y(_0093_),
    .A(_2965_),
    .B(net122));
 sg13g2_a21oi_1 _3962_ (.A1(_3012_),
    .A2(_0093_),
    .Y(_0094_),
    .B1(net31));
 sg13g2_nor3_1 _3963_ (.A(_1096_),
    .B(_2577_),
    .C(_2478_),
    .Y(_0095_));
 sg13g2_nand2_1 _3964_ (.Y(_0096_),
    .A(_2745_),
    .B(_2683_));
 sg13g2_nor2_1 _3965_ (.A(net174),
    .B(_0096_),
    .Y(_0097_));
 sg13g2_nor2_1 _3966_ (.A(_0095_),
    .B(_0097_),
    .Y(_0098_));
 sg13g2_nand2_1 _3967_ (.Y(_0099_),
    .A(_2675_),
    .B(_0910_));
 sg13g2_nand2_2 _3968_ (.Y(_0100_),
    .A(_0099_),
    .B(net136));
 sg13g2_nor2_1 _3969_ (.A(_2406_),
    .B(_0100_),
    .Y(_0101_));
 sg13g2_nor2_1 _3970_ (.A(net203),
    .B(_0101_),
    .Y(_0102_));
 sg13g2_nand2_1 _3971_ (.Y(_0103_),
    .A(_0098_),
    .B(_0102_));
 sg13g2_a21oi_1 _3972_ (.A1(_2850_),
    .A2(_3025_),
    .Y(_0104_),
    .B1(net145));
 sg13g2_nor3_1 _3973_ (.A(_0094_),
    .B(_0103_),
    .C(_0104_),
    .Y(_0105_));
 sg13g2_nor2_1 _3974_ (.A(net166),
    .B(_0105_),
    .Y(_0106_));
 sg13g2_nand2_1 _3975_ (.Y(_0107_),
    .A(net82),
    .B(_0801_));
 sg13g2_nand2_1 _3976_ (.Y(_0108_),
    .A(net43),
    .B(net86));
 sg13g2_o21ai_1 _3977_ (.B1(_0108_),
    .Y(_0109_),
    .A1(net77),
    .A2(_0107_));
 sg13g2_buf_1 _3978_ (.A(net108),
    .X(_0110_));
 sg13g2_nand2_1 _3979_ (.Y(_0111_),
    .A(_0109_),
    .B(net36));
 sg13g2_nor2_1 _3980_ (.A(net183),
    .B(net178),
    .Y(_0112_));
 sg13g2_nor3_1 _3981_ (.A(net155),
    .B(_1998_),
    .C(_0112_),
    .Y(_0113_));
 sg13g2_nor2_1 _3982_ (.A(net41),
    .B(_2897_),
    .Y(_0114_));
 sg13g2_nor3_1 _3983_ (.A(net173),
    .B(_0113_),
    .C(_0114_),
    .Y(_0115_));
 sg13g2_nand2_1 _3984_ (.Y(_0116_),
    .A(_0111_),
    .B(_0115_));
 sg13g2_nand2_1 _3985_ (.Y(_0117_),
    .A(net180),
    .B(\mem_addr[6] ));
 sg13g2_buf_2 _3986_ (.A(_0117_),
    .X(_0118_));
 sg13g2_nand2_1 _3987_ (.Y(_0119_),
    .A(_0116_),
    .B(_0118_));
 sg13g2_nand3_1 _3988_ (.B(net38),
    .C(_1653_),
    .A(net57),
    .Y(_0120_));
 sg13g2_a22oi_1 _3989_ (.Y(_0121_),
    .B1(_2882_),
    .B2(_3027_),
    .A2(net50),
    .A1(_0120_));
 sg13g2_nand2_1 _3990_ (.Y(_0122_),
    .A(_0119_),
    .B(_0121_));
 sg13g2_nand2_1 _3991_ (.Y(_0123_),
    .A(_0106_),
    .B(_0122_));
 sg13g2_nand2_1 _3992_ (.Y(_0124_),
    .A(_2793_),
    .B(net156));
 sg13g2_nand2_1 _3993_ (.Y(_0125_),
    .A(_0124_),
    .B(net56));
 sg13g2_nand2_1 _3994_ (.Y(_0126_),
    .A(_0125_),
    .B(_2854_));
 sg13g2_buf_1 _3995_ (.A(_0035_),
    .X(_0127_));
 sg13g2_inv_2 _3996_ (.Y(_0128_),
    .A(_0127_));
 sg13g2_nor3_1 _3997_ (.A(_2601_),
    .B(_0128_),
    .C(_2690_),
    .Y(_0129_));
 sg13g2_a21oi_1 _3998_ (.A1(_0126_),
    .A2(_0129_),
    .Y(_0130_),
    .B1(net170));
 sg13g2_a21oi_1 _3999_ (.A1(_0123_),
    .A2(_0130_),
    .Y(_0131_),
    .B1(net165));
 sg13g2_nand2_1 _4000_ (.Y(_0132_),
    .A(_0092_),
    .B(_0131_));
 sg13g2_nand2_1 _4001_ (.Y(_0022_),
    .A(_2976_),
    .B(_0132_));
 sg13g2_nand2_1 _4002_ (.Y(_0133_),
    .A(net71),
    .B(net82));
 sg13g2_nor2_1 _4003_ (.A(net111),
    .B(_0133_),
    .Y(_0134_));
 sg13g2_nand2_1 _4004_ (.Y(_0135_),
    .A(_2683_),
    .B(_2550_));
 sg13g2_nand2_1 _4005_ (.Y(_0136_),
    .A(_0135_),
    .B(_2405_));
 sg13g2_nor2_1 _4006_ (.A(_0134_),
    .B(_0136_),
    .Y(_0137_));
 sg13g2_nand2_1 _4007_ (.Y(_0138_),
    .A(_2397_),
    .B(net181));
 sg13g2_nand2_1 _4008_ (.Y(_0139_),
    .A(_0138_),
    .B(_1859_));
 sg13g2_nand2_1 _4009_ (.Y(_0140_),
    .A(_0139_),
    .B(net93));
 sg13g2_nand2_1 _4010_ (.Y(_0141_),
    .A(_0140_),
    .B(_1336_));
 sg13g2_inv_2 _4011_ (.Y(_0142_),
    .A(net148));
 sg13g2_nor2_2 _4012_ (.A(_0142_),
    .B(net86),
    .Y(_0143_));
 sg13g2_nor2_1 _4013_ (.A(net158),
    .B(_2683_),
    .Y(_0144_));
 sg13g2_nor2_1 _4014_ (.A(_0143_),
    .B(_0144_),
    .Y(_0145_));
 sg13g2_nor2_1 _4015_ (.A(_0141_),
    .B(_0145_),
    .Y(_0146_));
 sg13g2_nor2_1 _4016_ (.A(_0137_),
    .B(_0146_),
    .Y(_0147_));
 sg13g2_nor2_2 _4017_ (.A(net136),
    .B(net90),
    .Y(_0148_));
 sg13g2_nand2_2 _4018_ (.Y(_0149_),
    .A(_2469_),
    .B(net185));
 sg13g2_nand2_2 _4019_ (.Y(_0150_),
    .A(_0149_),
    .B(_2547_));
 sg13g2_nand2b_1 _4020_ (.Y(_0151_),
    .B(_0150_),
    .A_N(_0148_));
 sg13g2_nand2_1 _4021_ (.Y(_0152_),
    .A(_0151_),
    .B(net88));
 sg13g2_inv_1 _4022_ (.Y(_0153_),
    .A(net126));
 sg13g2_nor3_1 _4023_ (.A(net109),
    .B(_0153_),
    .C(_2848_),
    .Y(_0154_));
 sg13g2_nor2_1 _4024_ (.A(net62),
    .B(_0154_),
    .Y(_0155_));
 sg13g2_nand2_1 _4025_ (.Y(_0156_),
    .A(_3007_),
    .B(_2550_));
 sg13g2_nand2_1 _4026_ (.Y(_0157_),
    .A(_0155_),
    .B(_0156_));
 sg13g2_nand3_1 _4027_ (.B(_0152_),
    .C(_0157_),
    .A(_0147_),
    .Y(_0158_));
 sg13g2_nand2_1 _4028_ (.Y(_0159_),
    .A(_0158_),
    .B(net131));
 sg13g2_nand2_2 _4029_ (.Y(_0160_),
    .A(_2710_),
    .B(net109));
 sg13g2_buf_2 _4030_ (.A(net149),
    .X(_0161_));
 sg13g2_nand3_1 _4031_ (.B(net67),
    .C(net176),
    .A(_0160_),
    .Y(_0162_));
 sg13g2_inv_2 _4032_ (.Y(_0163_),
    .A(_2053_));
 sg13g2_a21oi_1 _4033_ (.A1(_0108_),
    .A2(_2715_),
    .Y(_0164_),
    .B1(net35));
 sg13g2_buf_1 _4034_ (.A(_2141_),
    .X(_0165_));
 sg13g2_nor2_1 _4035_ (.A(net182),
    .B(_3029_),
    .Y(_0166_));
 sg13g2_buf_2 _4036_ (.A(_0166_),
    .X(_0167_));
 sg13g2_a21oi_2 _4037_ (.B1(net155),
    .Y(_0168_),
    .A2(net153),
    .A1(net206));
 sg13g2_nand3_1 _4038_ (.B(net51),
    .C(net133),
    .A(_0168_),
    .Y(_0169_));
 sg13g2_o21ai_1 _4039_ (.B1(_0169_),
    .Y(_0170_),
    .A1(_0167_),
    .A2(_1816_));
 sg13g2_a22oi_1 _4040_ (.Y(_0171_),
    .B1(net115),
    .B2(_0170_),
    .A2(_0164_),
    .A1(_0162_));
 sg13g2_nand2_1 _4041_ (.Y(_0172_),
    .A(_0159_),
    .B(_0171_));
 sg13g2_nand2_1 _4042_ (.Y(_0173_),
    .A(_0172_),
    .B(net68));
 sg13g2_nand2_2 _4043_ (.Y(_0174_),
    .A(_2871_),
    .B(_2436_));
 sg13g2_nand2_1 _4044_ (.Y(_0175_),
    .A(_2525_),
    .B(net93));
 sg13g2_nand2_1 _4045_ (.Y(_0176_),
    .A(_0174_),
    .B(_0175_));
 sg13g2_nand2_1 _4046_ (.Y(_0177_),
    .A(_0176_),
    .B(net91));
 sg13g2_nand2_1 _4047_ (.Y(_0178_),
    .A(net122),
    .B(net137));
 sg13g2_nand2_1 _4048_ (.Y(_0179_),
    .A(_0178_),
    .B(_2842_));
 sg13g2_a21oi_1 _4049_ (.A1(_0177_),
    .A2(_0179_),
    .Y(_0180_),
    .B1(net81));
 sg13g2_buf_8 _4050_ (.A(_2086_),
    .X(_0181_));
 sg13g2_nand3_1 _4051_ (.B(net79),
    .C(net43),
    .A(net34),
    .Y(_0182_));
 sg13g2_nand3_1 _4052_ (.B(net129),
    .C(_0140_),
    .A(_0182_),
    .Y(_0183_));
 sg13g2_nand2_1 _4053_ (.Y(_0184_),
    .A(_2819_),
    .B(net150));
 sg13g2_nand2_1 _4054_ (.Y(_0185_),
    .A(_2273_),
    .B(_1227_));
 sg13g2_nand2_1 _4055_ (.Y(_0186_),
    .A(_0184_),
    .B(_0185_));
 sg13g2_nand2_1 _4056_ (.Y(_0187_),
    .A(_0186_),
    .B(net142));
 sg13g2_nand2_1 _4057_ (.Y(_0188_),
    .A(_0183_),
    .B(_0187_));
 sg13g2_nor2_1 _4058_ (.A(_0180_),
    .B(_0188_),
    .Y(_0189_));
 sg13g2_nor2_1 _4059_ (.A(net63),
    .B(_0189_),
    .Y(_0190_));
 sg13g2_a21oi_1 _4060_ (.A1(net43),
    .A2(net85),
    .Y(_0191_),
    .B1(net150));
 sg13g2_nand2_1 _4061_ (.Y(_0192_),
    .A(_3008_),
    .B(_0191_));
 sg13g2_nor2_1 _4062_ (.A(net198),
    .B(_3005_),
    .Y(_0193_));
 sg13g2_o21ai_1 _4063_ (.B1(_0193_),
    .Y(_0194_),
    .A1(net48),
    .A2(_2674_));
 sg13g2_nand2_1 _4064_ (.Y(_0195_),
    .A(_0192_),
    .B(_0194_));
 sg13g2_nand2_1 _4065_ (.Y(_0196_),
    .A(_0195_),
    .B(net24));
 sg13g2_nand2_1 _4066_ (.Y(_0197_),
    .A(net137),
    .B(net189));
 sg13g2_inv_1 _4067_ (.Y(_0198_),
    .A(_0197_));
 sg13g2_nor2_1 _4068_ (.A(net59),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_nor3_1 _4069_ (.A(net28),
    .B(_0199_),
    .C(_2574_),
    .Y(_0200_));
 sg13g2_a21oi_1 _4070_ (.A1(_2571_),
    .A2(net82),
    .Y(_0201_),
    .B1(net150));
 sg13g2_nand2_1 _4071_ (.Y(_0202_),
    .A(_0201_),
    .B(_1968_));
 sg13g2_nand2_1 _4072_ (.Y(_0203_),
    .A(_0202_),
    .B(_2559_));
 sg13g2_nor2_1 _4073_ (.A(_0200_),
    .B(_0203_),
    .Y(_0204_));
 sg13g2_nand2_1 _4074_ (.Y(_0205_),
    .A(_0196_),
    .B(_0204_));
 sg13g2_nand2_1 _4075_ (.Y(_0206_),
    .A(_0205_),
    .B(_2423_));
 sg13g2_nor2_1 _4076_ (.A(_0190_),
    .B(_0206_),
    .Y(_0207_));
 sg13g2_nand2_1 _4077_ (.Y(_0208_),
    .A(_0173_),
    .B(_0207_));
 sg13g2_inv_1 _4078_ (.Y(_0209_),
    .A(_0143_));
 sg13g2_nand2_1 _4079_ (.Y(_0210_),
    .A(_0209_),
    .B(_1446_));
 sg13g2_nand2_1 _4080_ (.Y(_0211_),
    .A(_2967_),
    .B(net60));
 sg13g2_nand2_1 _4081_ (.Y(_0212_),
    .A(_0210_),
    .B(_0211_));
 sg13g2_nand2_1 _4082_ (.Y(_0213_),
    .A(_0212_),
    .B(net129));
 sg13g2_nor2_1 _4083_ (.A(net152),
    .B(net155),
    .Y(_0214_));
 sg13g2_nand2_1 _4084_ (.Y(_0215_),
    .A(_0149_),
    .B(_0214_));
 sg13g2_nand2_1 _4085_ (.Y(_0216_),
    .A(_2835_),
    .B(_0215_));
 sg13g2_nand2_1 _4086_ (.Y(_0217_),
    .A(_0216_),
    .B(net49));
 sg13g2_nand2_1 _4087_ (.Y(_0218_),
    .A(_0213_),
    .B(_0217_));
 sg13g2_nand2_2 _4088_ (.Y(_0219_),
    .A(_2812_),
    .B(net106));
 sg13g2_buf_1 _4089_ (.A(net177),
    .X(_0220_));
 sg13g2_a21oi_1 _4090_ (.A1(_0219_),
    .A2(net156),
    .Y(_0221_),
    .B1(net114));
 sg13g2_nand2_1 _4091_ (.Y(_0222_),
    .A(net34),
    .B(net87));
 sg13g2_nand2_1 _4092_ (.Y(_0223_),
    .A(_0222_),
    .B(net102));
 sg13g2_nor2_1 _4093_ (.A(net60),
    .B(net44),
    .Y(_0224_));
 sg13g2_nor2_1 _4094_ (.A(net182),
    .B(_2511_),
    .Y(_0225_));
 sg13g2_inv_1 _4095_ (.Y(_0226_),
    .A(_2467_));
 sg13g2_nand2_1 _4096_ (.Y(_0227_),
    .A(_0225_),
    .B(_0226_));
 sg13g2_o21ai_1 _4097_ (.B1(net171),
    .Y(_0228_),
    .A1(_0224_),
    .A2(_0227_));
 sg13g2_a21oi_1 _4098_ (.A1(_0221_),
    .A2(_0223_),
    .Y(_0229_),
    .B1(_0228_));
 sg13g2_nor2_1 _4099_ (.A(_0218_),
    .B(_0229_),
    .Y(_0230_));
 sg13g2_nor2_1 _4100_ (.A(net63),
    .B(_0230_),
    .Y(_0231_));
 sg13g2_nor2_1 _4101_ (.A(net101),
    .B(_2678_),
    .Y(_0232_));
 sg13g2_nand2_1 _4102_ (.Y(_0233_),
    .A(_2624_),
    .B(_2709_));
 sg13g2_buf_2 _4103_ (.A(_0233_),
    .X(_0234_));
 sg13g2_a21oi_1 _4104_ (.A1(_2752_),
    .A2(_2605_),
    .Y(_0235_),
    .B1(_1326_));
 sg13g2_a21oi_1 _4105_ (.A1(_0232_),
    .A2(_0234_),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_nand2_1 _4106_ (.Y(_0237_),
    .A(_2428_),
    .B(_2430_));
 sg13g2_nand2_1 _4107_ (.Y(_0238_),
    .A(_0237_),
    .B(net49));
 sg13g2_nand3_1 _4108_ (.B(net136),
    .C(_2426_),
    .A(_2778_),
    .Y(_0239_));
 sg13g2_nand2_1 _4109_ (.Y(_0240_),
    .A(net43),
    .B(_2649_));
 sg13g2_nand2_1 _4110_ (.Y(_0241_),
    .A(_0239_),
    .B(_0240_));
 sg13g2_nand2_1 _4111_ (.Y(_0242_),
    .A(_0241_),
    .B(net88));
 sg13g2_nand3_1 _4112_ (.B(_0238_),
    .C(_0242_),
    .A(_0236_),
    .Y(_0243_));
 sg13g2_nand2_1 _4113_ (.Y(_0244_),
    .A(_0243_),
    .B(_2559_));
 sg13g2_nand2_1 _4114_ (.Y(_0245_),
    .A(_0244_),
    .B(net170));
 sg13g2_nor2_1 _4115_ (.A(_0231_),
    .B(_0245_),
    .Y(_0246_));
 sg13g2_a21oi_1 _4116_ (.A1(_0099_),
    .A2(_2401_),
    .Y(_0247_),
    .B1(net135));
 sg13g2_nand2_1 _4117_ (.Y(_0248_),
    .A(_0247_),
    .B(_2910_));
 sg13g2_a21oi_1 _4118_ (.A1(_2529_),
    .A2(_0142_),
    .Y(_0249_),
    .B1(net177));
 sg13g2_nand2_1 _4119_ (.Y(_0250_),
    .A(_2582_),
    .B(_1227_));
 sg13g2_nand2_1 _4120_ (.Y(_0251_),
    .A(_0249_),
    .B(_0250_));
 sg13g2_nand3_1 _4121_ (.B(_0251_),
    .C(_2600_),
    .A(_0248_),
    .Y(_0252_));
 sg13g2_nand2_1 _4122_ (.Y(_0253_),
    .A(_2965_),
    .B(_0197_));
 sg13g2_nand3_1 _4123_ (.B(_0149_),
    .C(net104),
    .A(_0253_),
    .Y(_0254_));
 sg13g2_and2_1 _4124_ (.A(_0254_),
    .B(_2483_),
    .X(_0255_));
 sg13g2_nand2_1 _4125_ (.Y(_0256_),
    .A(_0252_),
    .B(_0255_));
 sg13g2_nand2_1 _4126_ (.Y(_0257_),
    .A(_0256_),
    .B(net80));
 sg13g2_inv_1 _4127_ (.Y(_0258_),
    .A(_2031_));
 sg13g2_a21oi_1 _4128_ (.A1(_0258_),
    .A2(net48),
    .Y(_0259_),
    .B1(net114));
 sg13g2_nand2_1 _4129_ (.Y(_0260_),
    .A(_2526_),
    .B(net146));
 sg13g2_nor2_1 _4130_ (.A(net75),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_o21ai_1 _4131_ (.B1(_0261_),
    .Y(_0262_),
    .A1(_1968_),
    .A2(_0259_));
 sg13g2_o21ai_1 _4132_ (.B1(net124),
    .Y(_0263_),
    .A1(net41),
    .A2(net34));
 sg13g2_nor2_1 _4133_ (.A(_2426_),
    .B(_2494_),
    .Y(_0264_));
 sg13g2_o21ai_1 _4134_ (.B1(net135),
    .Y(_0265_),
    .A1(net29),
    .A2(_0264_));
 sg13g2_nor2_2 _4135_ (.A(_2964_),
    .B(net122),
    .Y(_0266_));
 sg13g2_nand2_1 _4136_ (.Y(_0267_),
    .A(_0266_),
    .B(net177));
 sg13g2_nand2_1 _4137_ (.Y(_0268_),
    .A(_0265_),
    .B(_0267_));
 sg13g2_nor2_1 _4138_ (.A(_0263_),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_nor2_1 _4139_ (.A(net123),
    .B(_0269_),
    .Y(_0270_));
 sg13g2_nand2_1 _4140_ (.Y(_0271_),
    .A(_0262_),
    .B(_0270_));
 sg13g2_nand2_1 _4141_ (.Y(_0272_),
    .A(_0257_),
    .B(_0271_));
 sg13g2_nand2_1 _4142_ (.Y(_0273_),
    .A(_0272_),
    .B(net68));
 sg13g2_nand2_1 _4143_ (.Y(_0274_),
    .A(_0246_),
    .B(_0273_));
 sg13g2_nand3_1 _4144_ (.B(_0274_),
    .C(net165),
    .A(_0208_),
    .Y(_0275_));
 sg13g2_nand2_1 _4145_ (.Y(_0276_),
    .A(_2532_),
    .B(net176));
 sg13g2_nand2_1 _4146_ (.Y(_0277_),
    .A(_0149_),
    .B(_0276_));
 sg13g2_nand2_1 _4147_ (.Y(_0278_),
    .A(_2930_),
    .B(_1511_));
 sg13g2_nand3_1 _4148_ (.B(_0278_),
    .C(net114),
    .A(_0277_),
    .Y(_0279_));
 sg13g2_nand2_1 _4149_ (.Y(_0280_),
    .A(_0279_),
    .B(_0177_));
 sg13g2_nand2_1 _4150_ (.Y(_0281_),
    .A(_0280_),
    .B(net46));
 sg13g2_inv_1 _4151_ (.Y(_0282_),
    .A(_0260_));
 sg13g2_nand2_1 _4152_ (.Y(_0283_),
    .A(_2660_),
    .B(net52));
 sg13g2_a21oi_1 _4153_ (.A1(_0282_),
    .A2(_0283_),
    .Y(_0284_),
    .B1(net138));
 sg13g2_nand2_1 _4154_ (.Y(_0285_),
    .A(_2900_),
    .B(net38));
 sg13g2_a21oi_1 _4155_ (.A1(_2617_),
    .A2(_0285_),
    .Y(_0286_),
    .B1(net54));
 sg13g2_nor3_1 _4156_ (.A(net127),
    .B(_0284_),
    .C(_0286_),
    .Y(_0287_));
 sg13g2_a21oi_1 _4157_ (.A1(_0281_),
    .A2(_0287_),
    .Y(_0288_),
    .B1(net166));
 sg13g2_nand2_1 _4158_ (.Y(_0289_),
    .A(_0900_),
    .B(_1911_));
 sg13g2_o21ai_1 _4159_ (.B1(net56),
    .Y(_0290_),
    .A1(_1478_),
    .A2(_0289_));
 sg13g2_nand2_1 _4160_ (.Y(_0291_),
    .A(_2119_),
    .B(_0290_));
 sg13g2_nand2_1 _4161_ (.Y(_0292_),
    .A(_2890_),
    .B(_3012_));
 sg13g2_a22oi_1 _4162_ (.Y(_0293_),
    .B1(net26),
    .B2(_0292_),
    .A2(net70),
    .A1(_0291_));
 sg13g2_buf_1 _4163_ (.A(net64),
    .X(_0294_));
 sg13g2_a21oi_1 _4164_ (.A1(_2119_),
    .A2(_2572_),
    .Y(_0295_),
    .B1(net23));
 sg13g2_nand2_1 _4165_ (.Y(_0296_),
    .A(_2830_),
    .B(net51));
 sg13g2_nand2_1 _4166_ (.Y(_0297_),
    .A(_0174_),
    .B(_0296_));
 sg13g2_a21oi_1 _4167_ (.A1(_0297_),
    .A2(net42),
    .Y(_0298_),
    .B1(net169));
 sg13g2_nor2b_1 _4168_ (.A(_0295_),
    .B_N(_0298_),
    .Y(_0299_));
 sg13g2_nand2_1 _4169_ (.Y(_0300_),
    .A(_0293_),
    .B(_0299_));
 sg13g2_nand2_1 _4170_ (.Y(_0301_),
    .A(_0288_),
    .B(_0300_));
 sg13g2_a21oi_1 _4171_ (.A1(_2387_),
    .A2(_2633_),
    .Y(_0302_),
    .B1(_2173_));
 sg13g2_nand2_2 _4172_ (.Y(_0303_),
    .A(_2691_),
    .B(_0034_));
 sg13g2_a221oi_1 _4173_ (.B2(_0302_),
    .C1(_0303_),
    .B1(_0169_),
    .A1(_0167_),
    .Y(_0304_),
    .A2(_1880_));
 sg13g2_nor2_1 _4174_ (.A(net170),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_a21oi_1 _4175_ (.A1(_0301_),
    .A2(_0305_),
    .Y(_0306_),
    .B1(net165));
 sg13g2_a21oi_1 _4176_ (.A1(_2803_),
    .A2(_0285_),
    .Y(_0307_),
    .B1(net23));
 sg13g2_a21oi_1 _4177_ (.A1(_2746_),
    .A2(_2747_),
    .Y(_0308_),
    .B1(net28));
 sg13g2_inv_1 _4178_ (.Y(_0309_),
    .A(_2960_));
 sg13g2_nand3b_1 _4179_ (.B(net134),
    .C(_0309_),
    .Y(_0310_),
    .A_N(_2470_));
 sg13g2_nand2_1 _4180_ (.Y(_0311_),
    .A(_2440_),
    .B(net177));
 sg13g2_o21ai_1 _4181_ (.B1(_0311_),
    .Y(_0312_),
    .A1(_1998_),
    .A2(net47));
 sg13g2_nand2_1 _4182_ (.Y(_0313_),
    .A(_0312_),
    .B(net171));
 sg13g2_nand3b_1 _4183_ (.B(_0310_),
    .C(_0313_),
    .Y(_0314_),
    .A_N(_0308_));
 sg13g2_nor2_1 _4184_ (.A(_0307_),
    .B(_0314_),
    .Y(_0315_));
 sg13g2_nor2_1 _4185_ (.A(net118),
    .B(_0315_),
    .Y(_0316_));
 sg13g2_nor2_1 _4186_ (.A(net200),
    .B(_0316_),
    .Y(_0317_));
 sg13g2_nand2_1 _4187_ (.Y(_0318_),
    .A(_2086_),
    .B(net140));
 sg13g2_nand2_1 _4188_ (.Y(_0319_),
    .A(net122),
    .B(_2550_));
 sg13g2_nand2_1 _4189_ (.Y(_0320_),
    .A(_0318_),
    .B(_0319_));
 sg13g2_nor2_2 _4190_ (.A(_2512_),
    .B(_2713_),
    .Y(_0321_));
 sg13g2_o21ai_1 _4191_ (.B1(_0321_),
    .Y(_0322_),
    .A1(_2494_),
    .A2(_0143_));
 sg13g2_a22oi_1 _4192_ (.Y(_0323_),
    .B1(net25),
    .B2(_0322_),
    .A2(net53),
    .A1(_0320_));
 sg13g2_a21oi_2 _4193_ (.B1(net51),
    .Y(_0324_),
    .A2(net94),
    .A1(_2622_));
 sg13g2_o21ai_1 _4194_ (.B1(net26),
    .Y(_0325_),
    .A1(_2955_),
    .A2(_0324_));
 sg13g2_buf_1 _4195_ (.A(net79),
    .X(_0326_));
 sg13g2_nor2_1 _4196_ (.A(net33),
    .B(_2525_),
    .Y(_0327_));
 sg13g2_o21ai_1 _4197_ (.B1(net70),
    .Y(_0328_),
    .A1(_0327_),
    .A2(_2948_));
 sg13g2_nand3_1 _4198_ (.B(_0325_),
    .C(_0328_),
    .A(_0323_),
    .Y(_0329_));
 sg13g2_nand2_1 _4199_ (.Y(_0330_),
    .A(_0329_),
    .B(_2373_));
 sg13g2_nand3_1 _4200_ (.B(net42),
    .C(_0174_),
    .A(_2870_),
    .Y(_0331_));
 sg13g2_nand2_2 _4201_ (.Y(_0332_),
    .A(net87),
    .B(net141));
 sg13g2_nand2_1 _4202_ (.Y(_0333_),
    .A(_2892_),
    .B(_0332_));
 sg13g2_buf_2 _4203_ (.A(net69),
    .X(_0334_));
 sg13g2_nand3_1 _4204_ (.B(_0333_),
    .C(net32),
    .A(_0150_),
    .Y(_0335_));
 sg13g2_a21oi_1 _4205_ (.A1(_0331_),
    .A2(_0335_),
    .Y(_0336_),
    .B1(net131));
 sg13g2_inv_1 _4206_ (.Y(_0337_),
    .A(_2141_));
 sg13g2_buf_1 _4207_ (.A(_0337_),
    .X(_0338_));
 sg13g2_nand2_1 _4208_ (.Y(_0339_),
    .A(_2671_),
    .B(_2947_));
 sg13g2_nor2_1 _4209_ (.A(net48),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_nand2_1 _4210_ (.Y(_0341_),
    .A(_0234_),
    .B(net114));
 sg13g2_nor2_1 _4211_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_nor2_1 _4212_ (.A(net66),
    .B(_0342_),
    .Y(_0343_));
 sg13g2_nand2_1 _4213_ (.Y(_0344_),
    .A(_2436_),
    .B(net141));
 sg13g2_nand2_1 _4214_ (.Y(_0345_),
    .A(_3018_),
    .B(_0344_));
 sg13g2_nor2_2 _4215_ (.A(_1216_),
    .B(net59),
    .Y(_0346_));
 sg13g2_nand2_1 _4216_ (.Y(_0347_),
    .A(_0346_),
    .B(_2947_));
 sg13g2_nand3_1 _4217_ (.B(_0347_),
    .C(net24),
    .A(_0345_),
    .Y(_0348_));
 sg13g2_a21oi_1 _4218_ (.A1(_0343_),
    .A2(_0348_),
    .Y(_0349_),
    .B1(_2646_));
 sg13g2_nand2_2 _4219_ (.Y(_0350_),
    .A(_2800_),
    .B(_2525_));
 sg13g2_nand2_1 _4220_ (.Y(_0351_),
    .A(_0350_),
    .B(_2844_));
 sg13g2_nor2_1 _4221_ (.A(net179),
    .B(_2751_),
    .Y(_0352_));
 sg13g2_nand2_1 _4222_ (.Y(_0353_),
    .A(_0351_),
    .B(_0352_));
 sg13g2_nand2_1 _4223_ (.Y(_0354_),
    .A(_2616_),
    .B(net95));
 sg13g2_nand2_1 _4224_ (.Y(_0355_),
    .A(_0354_),
    .B(_0167_));
 sg13g2_nand3_1 _4225_ (.B(_0355_),
    .C(net130),
    .A(_0353_),
    .Y(_0356_));
 sg13g2_nor2_1 _4226_ (.A(net101),
    .B(_0266_),
    .Y(_0357_));
 sg13g2_a21oi_1 _4227_ (.A1(_2969_),
    .A2(net104),
    .Y(_0358_),
    .B1(net173));
 sg13g2_nand2_1 _4228_ (.Y(_0359_),
    .A(_1795_),
    .B(_1184_));
 sg13g2_nor2_2 _4229_ (.A(_2543_),
    .B(_1998_),
    .Y(_0360_));
 sg13g2_nand2_1 _4230_ (.Y(_0361_),
    .A(_0359_),
    .B(_0360_));
 sg13g2_nand2_1 _4231_ (.Y(_0362_),
    .A(_0358_),
    .B(_0361_));
 sg13g2_a21oi_1 _4232_ (.A1(_0160_),
    .A2(_0357_),
    .Y(_0363_),
    .B1(_0362_));
 sg13g2_nand2_1 _4233_ (.Y(_0364_),
    .A(_0356_),
    .B(_0363_));
 sg13g2_nand3b_1 _4234_ (.B(_0349_),
    .C(_0364_),
    .Y(_0365_),
    .A_N(_0336_));
 sg13g2_nand3_1 _4235_ (.B(_0330_),
    .C(_0365_),
    .A(_0317_),
    .Y(_0366_));
 sg13g2_nand2_1 _4236_ (.Y(_0367_),
    .A(_0306_),
    .B(_0366_));
 sg13g2_nand2_1 _4237_ (.Y(_0023_),
    .A(_0275_),
    .B(_0367_));
 sg13g2_nor2_1 _4238_ (.A(net128),
    .B(_2602_),
    .Y(_0368_));
 sg13g2_a21oi_1 _4239_ (.A1(_0150_),
    .A2(_0368_),
    .Y(_0369_),
    .B1(net162));
 sg13g2_nand2_1 _4240_ (.Y(_0370_),
    .A(_2086_),
    .B(net97));
 sg13g2_nand2_1 _4241_ (.Y(_0371_),
    .A(_0370_),
    .B(net27));
 sg13g2_inv_1 _4242_ (.Y(_0372_),
    .A(_2813_));
 sg13g2_nor2_1 _4243_ (.A(net37),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_nand2_1 _4244_ (.Y(_0374_),
    .A(_0371_),
    .B(_0373_));
 sg13g2_nand2_1 _4245_ (.Y(_0375_),
    .A(_0369_),
    .B(_0374_));
 sg13g2_nand2_1 _4246_ (.Y(_0376_),
    .A(net126),
    .B(net153));
 sg13g2_nand2_1 _4247_ (.Y(_0377_),
    .A(_0376_),
    .B(_2488_));
 sg13g2_nand2_1 _4248_ (.Y(_0378_),
    .A(_0377_),
    .B(net27));
 sg13g2_nand3_1 _4249_ (.B(_2614_),
    .C(net45),
    .A(_0378_),
    .Y(_0379_));
 sg13g2_nand3_1 _4250_ (.B(net198),
    .C(_2020_),
    .A(_0276_),
    .Y(_0380_));
 sg13g2_nand2_1 _4251_ (.Y(_0381_),
    .A(_0380_),
    .B(_2643_));
 sg13g2_nand2_1 _4252_ (.Y(_0382_),
    .A(_0379_),
    .B(_0381_));
 sg13g2_a21oi_1 _4253_ (.A1(_0375_),
    .A2(_0382_),
    .Y(_0383_),
    .B1(net118));
 sg13g2_nor2_1 _4254_ (.A(_1326_),
    .B(_0260_),
    .Y(_0384_));
 sg13g2_nand2_1 _4255_ (.Y(_0385_),
    .A(_0160_),
    .B(_0384_));
 sg13g2_nand2_1 _4256_ (.Y(_0386_),
    .A(_0385_),
    .B(_2373_));
 sg13g2_nand2_2 _4257_ (.Y(_0387_),
    .A(_2582_),
    .B(net29));
 sg13g2_nand2_1 _4258_ (.Y(_0388_),
    .A(_2582_),
    .B(_0214_));
 sg13g2_nand3_1 _4259_ (.B(_0388_),
    .C(net69),
    .A(_0387_),
    .Y(_0389_));
 sg13g2_nor2b_1 _4260_ (.A(_0386_),
    .B_N(_0389_),
    .Y(_0390_));
 sg13g2_a21oi_1 _4261_ (.A1(_0214_),
    .A2(_1859_),
    .Y(_0391_),
    .B1(net174));
 sg13g2_nand2_1 _4262_ (.Y(_0392_),
    .A(_3043_),
    .B(_0391_));
 sg13g2_nand2_1 _4263_ (.Y(_0393_),
    .A(net144),
    .B(net137));
 sg13g2_nand2_1 _4264_ (.Y(_0394_),
    .A(_0393_),
    .B(_2745_));
 sg13g2_nor2_1 _4265_ (.A(net151),
    .B(net103),
    .Y(_0395_));
 sg13g2_nand2_1 _4266_ (.Y(_0396_),
    .A(_0394_),
    .B(_0395_));
 sg13g2_nand2_1 _4267_ (.Y(_0397_),
    .A(_0392_),
    .B(_0396_));
 sg13g2_nand2_1 _4268_ (.Y(_0398_),
    .A(_0397_),
    .B(net46));
 sg13g2_nand2_1 _4269_ (.Y(_0399_),
    .A(_0390_),
    .B(_0398_));
 sg13g2_nand2_1 _4270_ (.Y(_0400_),
    .A(_0399_),
    .B(_2423_));
 sg13g2_nor2_1 _4271_ (.A(_0383_),
    .B(_0400_),
    .Y(_0401_));
 sg13g2_nand2_1 _4272_ (.Y(_0402_),
    .A(_2833_),
    .B(net144));
 sg13g2_nand2_1 _4273_ (.Y(_0403_),
    .A(_0402_),
    .B(net27));
 sg13g2_inv_1 _4274_ (.Y(_0404_),
    .A(_2525_));
 sg13g2_nand2_1 _4275_ (.Y(_0405_),
    .A(_0404_),
    .B(net79));
 sg13g2_a21oi_1 _4276_ (.A1(_0403_),
    .A2(_0405_),
    .Y(_0406_),
    .B1(net23));
 sg13g2_a21oi_1 _4277_ (.A1(_3043_),
    .A2(_0277_),
    .Y(_0407_),
    .B1(net145));
 sg13g2_nor2_1 _4278_ (.A(_0406_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_nand2_1 _4279_ (.Y(_0409_),
    .A(_2889_),
    .B(_2097_));
 sg13g2_nand2_1 _4280_ (.Y(_0410_),
    .A(_0409_),
    .B(_2977_));
 sg13g2_nand2_1 _4281_ (.Y(_0411_),
    .A(_0410_),
    .B(net70));
 sg13g2_nand3_1 _4282_ (.B(net30),
    .C(net100),
    .A(net57),
    .Y(_0412_));
 sg13g2_nand2_1 _4283_ (.Y(_0413_),
    .A(_0412_),
    .B(_0100_));
 sg13g2_nand2_1 _4284_ (.Y(_0414_),
    .A(_0413_),
    .B(net26));
 sg13g2_nand3_1 _4285_ (.B(_0411_),
    .C(_0414_),
    .A(_0408_),
    .Y(_0415_));
 sg13g2_nor2_1 _4286_ (.A(net166),
    .B(net83),
    .Y(_0416_));
 sg13g2_nand2_1 _4287_ (.Y(_0417_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_inv_1 _4288_ (.Y(_0418_),
    .A(_2900_));
 sg13g2_nand3_1 _4289_ (.B(net37),
    .C(_0418_),
    .A(net34),
    .Y(_0419_));
 sg13g2_nand2_1 _4290_ (.Y(_0420_),
    .A(_2988_),
    .B(_2842_));
 sg13g2_nor2_1 _4291_ (.A(_1282_),
    .B(_1544_),
    .Y(_0421_));
 sg13g2_buf_2 _4292_ (.A(_0421_),
    .X(_0422_));
 sg13g2_nand2_1 _4293_ (.Y(_0423_),
    .A(_0178_),
    .B(_0422_));
 sg13g2_nand3_1 _4294_ (.B(_0420_),
    .C(_0423_),
    .A(_0419_),
    .Y(_0424_));
 sg13g2_nand2_1 _4295_ (.Y(_0425_),
    .A(_0424_),
    .B(net115));
 sg13g2_a21oi_1 _4296_ (.A1(_1609_),
    .A2(net141),
    .Y(_0426_),
    .B1(_2575_));
 sg13g2_nor2_1 _4297_ (.A(net33),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_nand2_1 _4298_ (.Y(_0428_),
    .A(net103),
    .B(_1162_));
 sg13g2_nand2_1 _4299_ (.Y(_0429_),
    .A(_2730_),
    .B(_0428_));
 sg13g2_nand2_1 _4300_ (.Y(_0430_),
    .A(_2871_),
    .B(net71));
 sg13g2_a21oi_1 _4301_ (.A1(_2724_),
    .A2(_0430_),
    .Y(_0431_),
    .B1(net35));
 sg13g2_o21ai_1 _4302_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0427_),
    .A2(_0429_));
 sg13g2_nand2_1 _4303_ (.Y(_0433_),
    .A(_0425_),
    .B(_0432_));
 sg13g2_nand2_1 _4304_ (.Y(_0434_),
    .A(_0433_),
    .B(net73));
 sg13g2_nand3_1 _4305_ (.B(_0417_),
    .C(_0434_),
    .A(_0401_),
    .Y(_0435_));
 sg13g2_nand2_1 _4306_ (.Y(_0436_),
    .A(_0370_),
    .B(_2842_));
 sg13g2_a21oi_1 _4307_ (.A1(_2983_),
    .A2(_3003_),
    .Y(_0437_),
    .B1(net35));
 sg13g2_nor2_2 _4308_ (.A(_0932_),
    .B(_1773_),
    .Y(_0438_));
 sg13g2_inv_1 _4309_ (.Y(_0439_),
    .A(_0438_));
 sg13g2_nand3_1 _4310_ (.B(net114),
    .C(_0439_),
    .A(_2986_),
    .Y(_0440_));
 sg13g2_nand3_1 _4311_ (.B(_0437_),
    .C(_0440_),
    .A(_0436_),
    .Y(_0441_));
 sg13g2_nand2_1 _4312_ (.Y(_0442_),
    .A(_0441_),
    .B(net175));
 sg13g2_nand3_1 _4313_ (.B(net111),
    .C(net158),
    .A(net126),
    .Y(_0443_));
 sg13g2_nand2_1 _4314_ (.Y(_0444_),
    .A(_0443_),
    .B(_2430_));
 sg13g2_a21oi_1 _4315_ (.A1(_0444_),
    .A2(net134),
    .Y(_0445_),
    .B1(net173));
 sg13g2_nand3_1 _4316_ (.B(net77),
    .C(net97),
    .A(_2622_),
    .Y(_0446_));
 sg13g2_nand2_1 _4317_ (.Y(_0447_),
    .A(_0446_),
    .B(_2867_));
 sg13g2_nand2_1 _4318_ (.Y(_0448_),
    .A(_0445_),
    .B(_0447_));
 sg13g2_nor2b_1 _4319_ (.A(_0107_),
    .B_N(_2992_),
    .Y(_0449_));
 sg13g2_nor2_1 _4320_ (.A(net114),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_nand2_1 _4321_ (.Y(_0451_),
    .A(_2942_),
    .B(net56));
 sg13g2_nor2_1 _4322_ (.A(_2641_),
    .B(_2513_),
    .Y(_0452_));
 sg13g2_nor2_2 _4323_ (.A(net182),
    .B(_2453_),
    .Y(_0453_));
 sg13g2_nor2_1 _4324_ (.A(net150),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_nor2_1 _4325_ (.A(_0452_),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_a21oi_1 _4326_ (.A1(_0450_),
    .A2(_0451_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_nor2_1 _4327_ (.A(_0448_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_nor2_1 _4328_ (.A(_0442_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_nand3_1 _4329_ (.B(net72),
    .C(_0405_),
    .A(_2119_),
    .Y(_0459_));
 sg13g2_nor2_1 _4330_ (.A(net149),
    .B(_2537_),
    .Y(_0460_));
 sg13g2_nand2_1 _4331_ (.Y(_0461_),
    .A(_0460_),
    .B(_2920_));
 sg13g2_nand2_1 _4332_ (.Y(_0462_),
    .A(_0459_),
    .B(_0461_));
 sg13g2_nand2_1 _4333_ (.Y(_0463_),
    .A(_0462_),
    .B(net115));
 sg13g2_nand2_1 _4334_ (.Y(_0464_),
    .A(_0458_),
    .B(_0463_));
 sg13g2_nand2_1 _4335_ (.Y(_0465_),
    .A(_3043_),
    .B(_2879_));
 sg13g2_a21oi_1 _4336_ (.A1(_1948_),
    .A2(_2532_),
    .Y(_0466_),
    .B1(net23));
 sg13g2_a21oi_1 _4337_ (.A1(_0465_),
    .A2(net25),
    .Y(_0467_),
    .B1(_0466_));
 sg13g2_nand2_1 _4338_ (.Y(_0468_),
    .A(_0987_),
    .B(_0856_));
 sg13g2_a21o_1 _4339_ (.A2(_0468_),
    .A1(_0215_),
    .B1(net61),
    .X(_0469_));
 sg13g2_nand3_1 _4340_ (.B(net136),
    .C(_1773_),
    .A(_0168_),
    .Y(_0470_));
 sg13g2_nand2_1 _4341_ (.Y(_0471_),
    .A(_2778_),
    .B(net109));
 sg13g2_nand2_1 _4342_ (.Y(_0472_),
    .A(_0470_),
    .B(_0471_));
 sg13g2_nand2_1 _4343_ (.Y(_0473_),
    .A(_0472_),
    .B(_2968_));
 sg13g2_nand3_1 _4344_ (.B(_0469_),
    .C(_0473_),
    .A(_0467_),
    .Y(_0474_));
 sg13g2_nand2_1 _4345_ (.Y(_0475_),
    .A(_0474_),
    .B(_2373_));
 sg13g2_nor2_1 _4346_ (.A(_1151_),
    .B(_2854_),
    .Y(_0476_));
 sg13g2_buf_2 _4347_ (.A(_0476_),
    .X(_0477_));
 sg13g2_nand2_2 _4348_ (.Y(_0478_),
    .A(_0477_),
    .B(net182));
 sg13g2_o21ai_1 _4349_ (.B1(_0478_),
    .Y(_0479_),
    .A1(_1998_),
    .A2(_2634_));
 sg13g2_nor2_1 _4350_ (.A(_2450_),
    .B(_2916_),
    .Y(_0480_));
 sg13g2_nor2_1 _4351_ (.A(net120),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_nand2_1 _4352_ (.Y(_0482_),
    .A(net210),
    .B(_1369_));
 sg13g2_buf_1 _4353_ (.A(_0482_),
    .X(_0483_));
 sg13g2_nor2_1 _4354_ (.A(net175),
    .B(net160),
    .Y(_0484_));
 sg13g2_o21ai_1 _4355_ (.B1(_0484_),
    .Y(_0485_),
    .A1(_0479_),
    .A2(_0481_));
 sg13g2_nand2_1 _4356_ (.Y(_0486_),
    .A(_0485_),
    .B(_2564_));
 sg13g2_nand2_1 _4357_ (.Y(_0487_),
    .A(net34),
    .B(_2900_));
 sg13g2_nand2_1 _4358_ (.Y(_0488_),
    .A(_0487_),
    .B(_2715_));
 sg13g2_a21oi_1 _4359_ (.A1(_0185_),
    .A2(net120),
    .Y(_0489_),
    .B1(net162));
 sg13g2_a22oi_1 _4360_ (.Y(_0490_),
    .B1(_0488_),
    .B2(_0489_),
    .A2(_2790_),
    .A1(net25));
 sg13g2_nor2_1 _4361_ (.A(net118),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_nor2_1 _4362_ (.A(_0486_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_nand3_1 _4363_ (.B(_0475_),
    .C(_0492_),
    .A(_0464_),
    .Y(_0493_));
 sg13g2_nand3_1 _4364_ (.B(_0493_),
    .C(net165),
    .A(_0435_),
    .Y(_0494_));
 sg13g2_nand2_1 _4365_ (.Y(_0495_),
    .A(net100),
    .B(_1184_));
 sg13g2_nand2_1 _4366_ (.Y(_0496_),
    .A(_0495_),
    .B(net60));
 sg13g2_a21oi_1 _4367_ (.A1(_2289_),
    .A2(_0496_),
    .Y(_0497_),
    .B1(net75));
 sg13g2_nand2_1 _4368_ (.Y(_0498_),
    .A(_2538_),
    .B(_2993_));
 sg13g2_nand2_1 _4369_ (.Y(_0499_),
    .A(_0498_),
    .B(net114));
 sg13g2_nand2_1 _4370_ (.Y(_0500_),
    .A(_0497_),
    .B(_0499_));
 sg13g2_nor2_1 _4371_ (.A(_2577_),
    .B(_2623_),
    .Y(_0501_));
 sg13g2_nor2_1 _4372_ (.A(_0266_),
    .B(_0501_),
    .Y(_0502_));
 sg13g2_nor2_1 _4373_ (.A(net28),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_nand2_1 _4374_ (.Y(_0504_),
    .A(_2801_),
    .B(net143));
 sg13g2_a21oi_1 _4375_ (.A1(_2959_),
    .A2(_0504_),
    .Y(_0505_),
    .B1(net101));
 sg13g2_nor2_1 _4376_ (.A(_0503_),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_nand2_1 _4377_ (.Y(_0507_),
    .A(_0500_),
    .B(_0506_));
 sg13g2_nand2_1 _4378_ (.Y(_0508_),
    .A(_0507_),
    .B(net80));
 sg13g2_nor2_1 _4379_ (.A(net142),
    .B(_2960_),
    .Y(_0509_));
 sg13g2_nor2_1 _4380_ (.A(net47),
    .B(_2812_),
    .Y(_0510_));
 sg13g2_inv_1 _4381_ (.Y(_0511_),
    .A(net160));
 sg13g2_o21ai_1 _4382_ (.B1(net113),
    .Y(_0512_),
    .A1(net37),
    .A2(_0510_));
 sg13g2_a21oi_1 _4383_ (.A1(_2977_),
    .A2(_0509_),
    .Y(_0513_),
    .B1(_0512_));
 sg13g2_nand2_2 _4384_ (.Y(_0514_),
    .A(_2414_),
    .B(net136));
 sg13g2_nand2_1 _4385_ (.Y(_0515_),
    .A(_0514_),
    .B(net128));
 sg13g2_inv_2 _4386_ (.Y(_0516_),
    .A(_2119_));
 sg13g2_nor2_1 _4387_ (.A(_0515_),
    .B(_0516_),
    .Y(_0517_));
 sg13g2_nand2_1 _4388_ (.Y(_0518_),
    .A(_0282_),
    .B(net108));
 sg13g2_nor2_1 _4389_ (.A(net77),
    .B(_0258_),
    .Y(_0519_));
 sg13g2_inv_1 _4390_ (.Y(_0520_),
    .A(_0118_));
 sg13g2_buf_1 _4391_ (.A(_0520_),
    .X(_0521_));
 sg13g2_o21ai_1 _4392_ (.B1(net22),
    .Y(_0522_),
    .A1(_0518_),
    .A2(_0519_));
 sg13g2_nor2_1 _4393_ (.A(_0517_),
    .B(_0522_),
    .Y(_0523_));
 sg13g2_nor2_1 _4394_ (.A(_0513_),
    .B(_0523_),
    .Y(_0524_));
 sg13g2_nand2_1 _4395_ (.Y(_0525_),
    .A(_0508_),
    .B(_0524_));
 sg13g2_nand2_1 _4396_ (.Y(_0526_),
    .A(_0525_),
    .B(net68));
 sg13g2_nor2_2 _4397_ (.A(net184),
    .B(net158),
    .Y(_0527_));
 sg13g2_inv_1 _4398_ (.Y(_0528_),
    .A(_0527_));
 sg13g2_a21oi_1 _4399_ (.A1(_2478_),
    .A2(_0528_),
    .Y(_0529_),
    .B1(net64));
 sg13g2_buf_1 _4400_ (.A(_2376_),
    .X(_0530_));
 sg13g2_nor2_1 _4401_ (.A(net194),
    .B(_1326_),
    .Y(_0531_));
 sg13g2_buf_1 _4402_ (.A(_0531_),
    .X(_0532_));
 sg13g2_inv_1 _4403_ (.Y(_0533_),
    .A(net65));
 sg13g2_nor2_1 _4404_ (.A(_0533_),
    .B(_2755_),
    .Y(_0534_));
 sg13g2_nor3_1 _4405_ (.A(net167),
    .B(_0529_),
    .C(_0534_),
    .Y(_0535_));
 sg13g2_inv_1 _4406_ (.Y(_0536_),
    .A(_2585_));
 sg13g2_a21oi_1 _4407_ (.A1(_0536_),
    .A2(_2715_),
    .Y(_0537_),
    .B1(net162));
 sg13g2_nor2_1 _4408_ (.A(net89),
    .B(_2547_),
    .Y(_0538_));
 sg13g2_nand2_1 _4409_ (.Y(_0539_),
    .A(_0169_),
    .B(_0538_));
 sg13g2_nand2_1 _4410_ (.Y(_0540_),
    .A(_0537_),
    .B(_0539_));
 sg13g2_a21oi_1 _4411_ (.A1(_0535_),
    .A2(_0540_),
    .Y(_0541_),
    .B1(net147));
 sg13g2_nand2_1 _4412_ (.Y(_0542_),
    .A(_0402_),
    .B(net77));
 sg13g2_nand2_1 _4413_ (.Y(_0543_),
    .A(_0542_),
    .B(net36));
 sg13g2_a21oi_1 _4414_ (.A1(net34),
    .A2(net57),
    .Y(_0544_),
    .B1(net33));
 sg13g2_a21oi_1 _4415_ (.A1(_2999_),
    .A2(_0167_),
    .Y(_0545_),
    .B1(net162));
 sg13g2_o21ai_1 _4416_ (.B1(_0545_),
    .Y(_0546_),
    .A1(_0543_),
    .A2(_0544_));
 sg13g2_nand2_1 _4417_ (.Y(_0547_),
    .A(_1435_),
    .B(_2376_));
 sg13g2_inv_1 _4418_ (.Y(_0548_),
    .A(_0547_));
 sg13g2_o21ai_1 _4419_ (.B1(net110),
    .Y(_0549_),
    .A1(_0548_),
    .A2(_2801_));
 sg13g2_nand2_1 _4420_ (.Y(_0550_),
    .A(_0549_),
    .B(net169));
 sg13g2_a21oi_1 _4421_ (.A1(_0514_),
    .A2(_2789_),
    .Y(_0551_),
    .B1(net23));
 sg13g2_nor2_1 _4422_ (.A(_0550_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_nand2_1 _4423_ (.Y(_0553_),
    .A(_0546_),
    .B(_0552_));
 sg13g2_a21oi_1 _4424_ (.A1(_0541_),
    .A2(_0553_),
    .Y(_0554_),
    .B1(net200));
 sg13g2_nand2_1 _4425_ (.Y(_0555_),
    .A(_0526_),
    .B(_0554_));
 sg13g2_nand2_1 _4426_ (.Y(_0556_),
    .A(_0376_),
    .B(net144));
 sg13g2_nand3_1 _4427_ (.B(net92),
    .C(net150),
    .A(_0556_),
    .Y(_0557_));
 sg13g2_nand2_1 _4428_ (.Y(_0558_),
    .A(net59),
    .B(net106));
 sg13g2_a21oi_1 _4429_ (.A1(net52),
    .A2(net156),
    .Y(_0559_),
    .B1(_2641_));
 sg13g2_nor2_1 _4430_ (.A(_0558_),
    .B(_0559_),
    .Y(_0560_));
 sg13g2_nand2_1 _4431_ (.Y(_0561_),
    .A(_0557_),
    .B(_0560_));
 sg13g2_nand2_1 _4432_ (.Y(_0562_),
    .A(_0561_),
    .B(net36));
 sg13g2_nand2_1 _4433_ (.Y(_0563_),
    .A(_1795_),
    .B(_2449_));
 sg13g2_nand2_1 _4434_ (.Y(_0564_),
    .A(_0563_),
    .B(_2495_));
 sg13g2_nand2_1 _4435_ (.Y(_0565_),
    .A(net95),
    .B(_0757_));
 sg13g2_nand2_1 _4436_ (.Y(_0566_),
    .A(_0565_),
    .B(net58));
 sg13g2_nand2_1 _4437_ (.Y(_0567_),
    .A(_0564_),
    .B(_0566_));
 sg13g2_inv_1 _4438_ (.Y(_0568_),
    .A(_1948_));
 sg13g2_nor3_1 _4439_ (.A(_0568_),
    .B(net62),
    .C(_2678_),
    .Y(_0569_));
 sg13g2_a21oi_1 _4440_ (.A1(_0567_),
    .A2(net39),
    .Y(_0570_),
    .B1(_0569_));
 sg13g2_nand2_1 _4441_ (.Y(_0571_),
    .A(_0562_),
    .B(_0570_));
 sg13g2_nand2_1 _4442_ (.Y(_0572_),
    .A(_0571_),
    .B(net80));
 sg13g2_nand2_1 _4443_ (.Y(_0573_),
    .A(_2502_),
    .B(_2433_));
 sg13g2_nand2_1 _4444_ (.Y(_0574_),
    .A(_0573_),
    .B(_2842_));
 sg13g2_o21ai_1 _4445_ (.B1(_2518_),
    .Y(_0575_),
    .A1(_0112_),
    .A2(_1869_));
 sg13g2_nor2_1 _4446_ (.A(_2477_),
    .B(_2905_),
    .Y(_0576_));
 sg13g2_inv_1 _4447_ (.Y(_0577_),
    .A(_0576_));
 sg13g2_nand3_1 _4448_ (.B(_0575_),
    .C(_0577_),
    .A(_0574_),
    .Y(_0578_));
 sg13g2_nand2_1 _4449_ (.Y(_0579_),
    .A(net98),
    .B(net152));
 sg13g2_nor2_1 _4450_ (.A(_0112_),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_nand2_1 _4451_ (.Y(_0581_),
    .A(_0395_),
    .B(_0226_));
 sg13g2_o21ai_1 _4452_ (.B1(net22),
    .Y(_0582_),
    .A1(_0580_),
    .A2(_0581_));
 sg13g2_nor2_1 _4453_ (.A(_2162_),
    .B(_0527_),
    .Y(_0583_));
 sg13g2_nand2_1 _4454_ (.Y(_0584_),
    .A(_2911_),
    .B(_0583_));
 sg13g2_nor2b_1 _4455_ (.A(_0582_),
    .B_N(_0584_),
    .Y(_0585_));
 sg13g2_a21oi_1 _4456_ (.A1(_0578_),
    .A2(net113),
    .Y(_0586_),
    .B1(_0585_));
 sg13g2_nand2_1 _4457_ (.Y(_0587_),
    .A(_0572_),
    .B(_0586_));
 sg13g2_nand2_1 _4458_ (.Y(_0588_),
    .A(_0587_),
    .B(net68));
 sg13g2_nand3_1 _4459_ (.B(net52),
    .C(_0422_),
    .A(net82),
    .Y(_0589_));
 sg13g2_o21ai_1 _4460_ (.B1(_0589_),
    .Y(_0590_),
    .A1(net99),
    .A2(_2977_));
 sg13g2_inv_1 _4461_ (.Y(_0591_),
    .A(_0303_));
 sg13g2_a21oi_1 _4462_ (.A1(_0590_),
    .A2(_0591_),
    .Y(_0592_),
    .B1(net163));
 sg13g2_nand2_1 _4463_ (.Y(_0593_),
    .A(_0588_),
    .B(_0592_));
 sg13g2_nand3_1 _4464_ (.B(_0593_),
    .C(net196),
    .A(_0555_),
    .Y(_0594_));
 sg13g2_nand2_1 _4465_ (.Y(_0024_),
    .A(_0494_),
    .B(_0594_));
 sg13g2_a21oi_1 _4466_ (.A1(net178),
    .A2(_0757_),
    .Y(_0595_),
    .B1(net184));
 sg13g2_inv_1 _4467_ (.Y(_0596_),
    .A(_0289_));
 sg13g2_nand2_2 _4468_ (.Y(_0597_),
    .A(_0595_),
    .B(_0596_));
 sg13g2_nor2_2 _4469_ (.A(_1653_),
    .B(net178),
    .Y(_0598_));
 sg13g2_inv_1 _4470_ (.Y(_0599_),
    .A(_0598_));
 sg13g2_nor2_2 _4471_ (.A(_2460_),
    .B(_2406_),
    .Y(_0600_));
 sg13g2_nand3_1 _4472_ (.B(_0599_),
    .C(_0600_),
    .A(_0597_),
    .Y(_0601_));
 sg13g2_inv_1 _4473_ (.Y(_0602_),
    .A(_2376_));
 sg13g2_nand2_1 _4474_ (.Y(_0603_),
    .A(_2848_),
    .B(net193));
 sg13g2_nor2_1 _4475_ (.A(_1555_),
    .B(_0118_),
    .Y(_0604_));
 sg13g2_a21oi_1 _4476_ (.A1(_0603_),
    .A2(_0604_),
    .Y(_0605_),
    .B1(_2423_));
 sg13g2_nand2_1 _4477_ (.Y(_0606_),
    .A(_0601_),
    .B(_0605_));
 sg13g2_nor2_2 _4478_ (.A(_0943_),
    .B(_2682_),
    .Y(_0607_));
 sg13g2_nand2_1 _4479_ (.Y(_0608_),
    .A(_0607_),
    .B(net193));
 sg13g2_nand2_2 _4480_ (.Y(_0609_),
    .A(_2633_),
    .B(_2808_));
 sg13g2_nor2_1 _4481_ (.A(net194),
    .B(_0609_),
    .Y(_0610_));
 sg13g2_nor2_1 _4482_ (.A(_1631_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_a21oi_1 _4483_ (.A1(_3022_),
    .A2(_0608_),
    .Y(_0612_),
    .B1(_0611_));
 sg13g2_nor2_1 _4484_ (.A(net66),
    .B(_0612_),
    .Y(_0613_));
 sg13g2_nor2_1 _4485_ (.A(_0606_),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_nor2_1 _4486_ (.A(_2445_),
    .B(_2640_),
    .Y(_0615_));
 sg13g2_nand2_2 _4487_ (.Y(_0616_),
    .A(_2887_),
    .B(net201));
 sg13g2_nand2_1 _4488_ (.Y(_0617_),
    .A(_0616_),
    .B(_2495_));
 sg13g2_nand2_2 _4489_ (.Y(_0618_),
    .A(_2659_),
    .B(_2589_));
 sg13g2_a21oi_1 _4490_ (.A1(_0617_),
    .A2(_0618_),
    .Y(_0619_),
    .B1(net54));
 sg13g2_o21ai_1 _4491_ (.B1(net116),
    .Y(_0620_),
    .A1(_0615_),
    .A2(_0619_));
 sg13g2_nor2_1 _4492_ (.A(net184),
    .B(_0112_),
    .Y(_0621_));
 sg13g2_inv_2 _4493_ (.Y(_0622_),
    .A(_0621_));
 sg13g2_nand3_1 _4494_ (.B(_2753_),
    .C(_0143_),
    .A(_0622_),
    .Y(_0623_));
 sg13g2_nand2_1 _4495_ (.Y(_0624_),
    .A(_2953_),
    .B(_2686_));
 sg13g2_nand3_1 _4496_ (.B(net113),
    .C(_0624_),
    .A(_0623_),
    .Y(_0625_));
 sg13g2_nand3_1 _4497_ (.B(_0620_),
    .C(_0625_),
    .A(_0614_),
    .Y(_0626_));
 sg13g2_nand2_1 _4498_ (.Y(_0627_),
    .A(_1795_),
    .B(_2490_));
 sg13g2_nor2_2 _4499_ (.A(_1271_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nand2_1 _4500_ (.Y(_0629_),
    .A(_2442_),
    .B(_2633_));
 sg13g2_a21oi_1 _4501_ (.A1(_1631_),
    .A2(_0128_),
    .Y(_0630_),
    .B1(net124));
 sg13g2_nand2_1 _4502_ (.Y(_0631_),
    .A(_2848_),
    .B(_0530_));
 sg13g2_a22oi_1 _4503_ (.Y(_0632_),
    .B1(_0630_),
    .B2(_0631_),
    .A2(_0629_),
    .A1(net134));
 sg13g2_o21ai_1 _4504_ (.B1(_0632_),
    .Y(_0633_),
    .A1(_2384_),
    .A2(_0628_));
 sg13g2_nand2_1 _4505_ (.Y(_0634_),
    .A(_0633_),
    .B(_2749_));
 sg13g2_a22oi_1 _4506_ (.Y(_0635_),
    .B1(_2701_),
    .B2(_0608_),
    .A2(net89),
    .A1(_0149_));
 sg13g2_nor2_1 _4507_ (.A(net35),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_nand2_1 _4508_ (.Y(_0637_),
    .A(_2710_),
    .B(net194));
 sg13g2_a21oi_1 _4509_ (.A1(_2729_),
    .A2(_0128_),
    .Y(_0638_),
    .B1(_0337_));
 sg13g2_a21oi_1 _4510_ (.A1(_0637_),
    .A2(_0638_),
    .Y(_0639_),
    .B1(_2564_));
 sg13g2_nor2b_1 _4511_ (.A(_0636_),
    .B_N(_0639_),
    .Y(_0640_));
 sg13g2_nand2_1 _4512_ (.Y(_0641_),
    .A(_0634_),
    .B(_0640_));
 sg13g2_nand2_1 _4513_ (.Y(_0642_),
    .A(_0626_),
    .B(_0641_));
 sg13g2_nand2_1 _4514_ (.Y(_0643_),
    .A(_0642_),
    .B(net68));
 sg13g2_nor3_2 _4515_ (.A(net177),
    .B(_0142_),
    .C(_3013_),
    .Y(_0644_));
 sg13g2_a21o_1 _4516_ (.A2(_0618_),
    .A1(_0644_),
    .B1(net160),
    .X(_0645_));
 sg13g2_nor2_1 _4517_ (.A(_0943_),
    .B(_2669_),
    .Y(_0646_));
 sg13g2_o21ai_1 _4518_ (.B1(_0646_),
    .Y(_0647_),
    .A1(_0422_),
    .A2(_2482_));
 sg13g2_nand2_1 _4519_ (.Y(_0648_),
    .A(_0609_),
    .B(_2490_));
 sg13g2_nand2_1 _4520_ (.Y(_0649_),
    .A(_0617_),
    .B(_0648_));
 sg13g2_nand2_1 _4521_ (.Y(_0650_),
    .A(net180),
    .B(_0128_));
 sg13g2_buf_2 _4522_ (.A(_0650_),
    .X(_0651_));
 sg13g2_a21oi_1 _4523_ (.A1(_2407_),
    .A2(_0651_),
    .Y(_0652_),
    .B1(_2595_));
 sg13g2_a22oi_1 _4524_ (.Y(_0653_),
    .B1(_0649_),
    .B2(_0652_),
    .A2(net105),
    .A1(_0647_));
 sg13g2_nand2_1 _4525_ (.Y(_0654_),
    .A(_0603_),
    .B(_2509_));
 sg13g2_inv_1 _4526_ (.Y(_0655_),
    .A(_2998_));
 sg13g2_nand2_1 _4527_ (.Y(_0656_),
    .A(_0655_),
    .B(_2173_));
 sg13g2_nand2_1 _4528_ (.Y(_0657_),
    .A(_0654_),
    .B(_0656_));
 sg13g2_nand2_1 _4529_ (.Y(_0658_),
    .A(_0657_),
    .B(net22));
 sg13g2_nand3_1 _4530_ (.B(_0653_),
    .C(_0658_),
    .A(_0645_),
    .Y(_0659_));
 sg13g2_nand2_1 _4531_ (.Y(_0660_),
    .A(_0659_),
    .B(_2565_));
 sg13g2_nand2_1 _4532_ (.Y(_0661_),
    .A(_0339_),
    .B(net128));
 sg13g2_nand2_1 _4533_ (.Y(_0662_),
    .A(_2417_),
    .B(net194));
 sg13g2_nand2_1 _4534_ (.Y(_0663_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_nand2_1 _4535_ (.Y(_0664_),
    .A(net71),
    .B(_2377_));
 sg13g2_o21ai_1 _4536_ (.B1(net161),
    .Y(_0665_),
    .A1(_1107_),
    .A2(_0664_));
 sg13g2_nor2_1 _4537_ (.A(_0663_),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_nand2_1 _4538_ (.Y(_0667_),
    .A(_2862_),
    .B(net74));
 sg13g2_a21oi_1 _4539_ (.A1(_0666_),
    .A2(_0667_),
    .Y(_0668_),
    .B1(_2564_));
 sg13g2_nand2_2 _4540_ (.Y(_0669_),
    .A(_0609_),
    .B(_2401_));
 sg13g2_o21ai_1 _4541_ (.B1(_0669_),
    .Y(_0670_),
    .A1(_0438_),
    .A2(_0618_));
 sg13g2_nand2_1 _4542_ (.Y(_0671_),
    .A(_0670_),
    .B(_0334_));
 sg13g2_nor3_1 _4543_ (.A(_2407_),
    .B(_2378_),
    .C(_0607_),
    .Y(_0672_));
 sg13g2_nand2_2 _4544_ (.Y(_0673_),
    .A(_0629_),
    .B(net179));
 sg13g2_nor2_1 _4545_ (.A(net171),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_nor2_1 _4546_ (.A(_0672_),
    .B(_0674_),
    .Y(_0675_));
 sg13g2_a21oi_1 _4547_ (.A1(_0608_),
    .A2(net42),
    .Y(_0676_),
    .B1(_2664_));
 sg13g2_nand3_1 _4548_ (.B(_0675_),
    .C(_0676_),
    .A(_0671_),
    .Y(_0677_));
 sg13g2_nand2_1 _4549_ (.Y(_0678_),
    .A(_0668_),
    .B(_0677_));
 sg13g2_nand3_1 _4550_ (.B(_0678_),
    .C(_2736_),
    .A(_0660_),
    .Y(_0679_));
 sg13g2_a21oi_1 _4551_ (.A1(_0643_),
    .A2(_0679_),
    .Y(_0680_),
    .B1(_2610_));
 sg13g2_nor2_1 _4552_ (.A(net133),
    .B(_0547_),
    .Y(_0681_));
 sg13g2_nand2_1 _4553_ (.Y(_0682_),
    .A(_0565_),
    .B(_2097_));
 sg13g2_nand2_1 _4554_ (.Y(_0683_),
    .A(_0682_),
    .B(net27));
 sg13g2_a22oi_1 _4555_ (.Y(_0684_),
    .B1(_0644_),
    .B2(_0683_),
    .A2(_0681_),
    .A1(_2654_));
 sg13g2_nand2_1 _4556_ (.Y(_0685_),
    .A(_0597_),
    .B(net37));
 sg13g2_nand2_1 _4557_ (.Y(_0686_),
    .A(_2768_),
    .B(net114));
 sg13g2_a21oi_1 _4558_ (.A1(_0685_),
    .A2(_0686_),
    .Y(_0687_),
    .B1(net160));
 sg13g2_a21oi_1 _4559_ (.A1(_0684_),
    .A2(net22),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_nor2_1 _4560_ (.A(_1107_),
    .B(_2723_),
    .Y(_0689_));
 sg13g2_nand3_1 _4561_ (.B(_2444_),
    .C(_2405_),
    .A(_2591_),
    .Y(_0690_));
 sg13g2_nor2b_1 _4562_ (.A(_0689_),
    .B_N(_0690_),
    .Y(_0691_));
 sg13g2_o21ai_1 _4563_ (.B1(_2861_),
    .Y(_0692_),
    .A1(_2505_),
    .A2(_0607_));
 sg13g2_nand2_1 _4564_ (.Y(_0693_),
    .A(_0692_),
    .B(net39));
 sg13g2_o21ai_1 _4565_ (.B1(net49),
    .Y(_0694_),
    .A1(net194),
    .A2(_0350_));
 sg13g2_nand3_1 _4566_ (.B(_0693_),
    .C(_0694_),
    .A(_0691_),
    .Y(_0695_));
 sg13g2_nand2_1 _4567_ (.Y(_0696_),
    .A(_0695_),
    .B(net116));
 sg13g2_nand2_1 _4568_ (.Y(_0697_),
    .A(_0688_),
    .B(_0696_));
 sg13g2_nand2_1 _4569_ (.Y(_0698_),
    .A(_0697_),
    .B(_0090_));
 sg13g2_nor2_1 _4570_ (.A(_2408_),
    .B(_2892_),
    .Y(_0699_));
 sg13g2_nand2_1 _4571_ (.Y(_0700_),
    .A(_2413_),
    .B(net193));
 sg13g2_nand3_1 _4572_ (.B(net55),
    .C(_2532_),
    .A(_2444_),
    .Y(_0701_));
 sg13g2_a221oi_1 _4573_ (.B2(_0701_),
    .C1(net118),
    .B1(_0454_),
    .A1(_0699_),
    .Y(_0702_),
    .A2(_0700_));
 sg13g2_nand2_1 _4574_ (.Y(_0703_),
    .A(_2273_),
    .B(net119));
 sg13g2_nand2_1 _4575_ (.Y(_0704_),
    .A(_0703_),
    .B(net92));
 sg13g2_a21oi_1 _4576_ (.A1(_0704_),
    .A2(_0618_),
    .Y(_0705_),
    .B1(net54));
 sg13g2_nand2_1 _4577_ (.Y(_0706_),
    .A(_0599_),
    .B(net128));
 sg13g2_nor3_1 _4578_ (.A(net107),
    .B(_0477_),
    .C(_0706_),
    .Y(_0707_));
 sg13g2_nor2_1 _4579_ (.A(_2383_),
    .B(_2638_),
    .Y(_0708_));
 sg13g2_nor2_1 _4580_ (.A(_0530_),
    .B(_0607_),
    .Y(_0709_));
 sg13g2_o21ai_1 _4581_ (.B1(_2552_),
    .Y(_0710_),
    .A1(_2892_),
    .A2(_0709_));
 sg13g2_nand2b_1 _4582_ (.Y(_0711_),
    .B(_0710_),
    .A_N(_0708_));
 sg13g2_nor3_1 _4583_ (.A(_0705_),
    .B(_0707_),
    .C(_0711_),
    .Y(_0712_));
 sg13g2_nor2_1 _4584_ (.A(_2375_),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_nor2_1 _4585_ (.A(_0702_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_nand2_1 _4586_ (.Y(_0715_),
    .A(_0698_),
    .B(_0714_));
 sg13g2_nor2_2 _4587_ (.A(net179),
    .B(_2998_),
    .Y(_0716_));
 sg13g2_a22oi_1 _4588_ (.Y(_0717_),
    .B1(_0716_),
    .B2(_0514_),
    .A2(_2637_),
    .A1(net42));
 sg13g2_nand3b_1 _4589_ (.B(_0717_),
    .C(_2699_),
    .Y(_0718_),
    .A_N(_0674_));
 sg13g2_nand2_1 _4590_ (.Y(_0719_),
    .A(_0692_),
    .B(net24));
 sg13g2_nor2_1 _4591_ (.A(_2386_),
    .B(_1151_),
    .Y(_0720_));
 sg13g2_nor2_2 _4592_ (.A(net151),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_nand2_1 _4593_ (.Y(_0722_),
    .A(_2719_),
    .B(_0721_));
 sg13g2_nand3_1 _4594_ (.B(_0722_),
    .C(net22),
    .A(_0719_),
    .Y(_0723_));
 sg13g2_nand2_1 _4595_ (.Y(_0724_),
    .A(_0664_),
    .B(_0334_));
 sg13g2_o21ai_1 _4596_ (.B1(_0724_),
    .Y(_0726_),
    .A1(_2793_),
    .A2(_0533_));
 sg13g2_nor2_1 _4597_ (.A(net197),
    .B(_2564_),
    .Y(_0727_));
 sg13g2_buf_1 _4598_ (.A(_0727_),
    .X(_0728_));
 sg13g2_inv_1 _4599_ (.Y(_0729_),
    .A(net112));
 sg13g2_a21oi_1 _4600_ (.A1(_0726_),
    .A2(net131),
    .Y(_0730_),
    .B1(_0729_));
 sg13g2_nand3_1 _4601_ (.B(_0723_),
    .C(_0730_),
    .A(_0718_),
    .Y(_0731_));
 sg13g2_nand2_1 _4602_ (.Y(_0732_),
    .A(net115),
    .B(_0127_));
 sg13g2_o21ai_1 _4603_ (.B1(_2598_),
    .Y(_0733_),
    .A1(_0732_),
    .A2(_0631_));
 sg13g2_nand3_1 _4604_ (.B(_2610_),
    .C(_0733_),
    .A(_0731_),
    .Y(_0734_));
 sg13g2_a21oi_1 _4605_ (.A1(_0715_),
    .A2(_2566_),
    .Y(_0735_),
    .B1(_0734_));
 sg13g2_nor2_1 _4606_ (.A(_0680_),
    .B(_0735_),
    .Y(_0025_));
 sg13g2_nor2_1 _4607_ (.A(net108),
    .B(_0580_),
    .Y(_0737_));
 sg13g2_o21ai_1 _4608_ (.B1(_0737_),
    .Y(_0738_),
    .A1(_2392_),
    .A2(_2656_));
 sg13g2_nor3_1 _4609_ (.A(net179),
    .B(net103),
    .C(_3013_),
    .Y(_0739_));
 sg13g2_a21oi_1 _4610_ (.A1(_0739_),
    .A2(_3046_),
    .Y(_0740_),
    .B1(net173));
 sg13g2_nand2_1 _4611_ (.Y(_0741_),
    .A(_0738_),
    .B(_0740_));
 sg13g2_nand2_1 _4612_ (.Y(_0742_),
    .A(_0596_),
    .B(_2399_));
 sg13g2_nand2_1 _4613_ (.Y(_0743_),
    .A(_0742_),
    .B(net143));
 sg13g2_inv_1 _4614_ (.Y(_0744_),
    .A(_0477_));
 sg13g2_nand2_1 _4615_ (.Y(_0745_),
    .A(_0743_),
    .B(_0744_));
 sg13g2_nand3_1 _4616_ (.B(net142),
    .C(net161),
    .A(_0745_),
    .Y(_0747_));
 sg13g2_nor2_2 _4617_ (.A(_2417_),
    .B(net209),
    .Y(_0748_));
 sg13g2_nand3_1 _4618_ (.B(_2719_),
    .C(_0748_),
    .A(_2712_),
    .Y(_0749_));
 sg13g2_nand3_1 _4619_ (.B(_0747_),
    .C(_0749_),
    .A(_0741_),
    .Y(_0750_));
 sg13g2_nand2_1 _4620_ (.Y(_0751_),
    .A(_0750_),
    .B(net46));
 sg13g2_a21oi_1 _4621_ (.A1(_2489_),
    .A2(_2402_),
    .Y(_0752_),
    .B1(net142));
 sg13g2_nand2_1 _4622_ (.Y(_0753_),
    .A(_2616_),
    .B(net125));
 sg13g2_o21ai_1 _4623_ (.B1(net113),
    .Y(_0754_),
    .A1(net89),
    .A2(net29));
 sg13g2_a21oi_1 _4624_ (.A1(_0752_),
    .A2(_0753_),
    .Y(_0755_),
    .B1(_0754_));
 sg13g2_nand2_1 _4625_ (.Y(_0756_),
    .A(_0468_),
    .B(_0669_));
 sg13g2_nor2_1 _4626_ (.A(net64),
    .B(_2678_),
    .Y(_0758_));
 sg13g2_a22oi_1 _4627_ (.Y(_0759_),
    .B1(_0758_),
    .B2(_3025_),
    .A2(_1347_),
    .A1(_0756_));
 sg13g2_nor2_1 _4628_ (.A(_2619_),
    .B(_0759_),
    .Y(_0760_));
 sg13g2_nor3_1 _4629_ (.A(net197),
    .B(_0755_),
    .C(_0760_),
    .Y(_0761_));
 sg13g2_nand2_1 _4630_ (.Y(_0762_),
    .A(_0751_),
    .B(_0761_));
 sg13g2_a21oi_1 _4631_ (.A1(_0096_),
    .A2(_2526_),
    .Y(_0763_),
    .B1(net31));
 sg13g2_nor2_1 _4632_ (.A(_2844_),
    .B(_2031_),
    .Y(_0764_));
 sg13g2_nor3_1 _4633_ (.A(net40),
    .B(_2616_),
    .C(_0764_),
    .Y(_0765_));
 sg13g2_nor3_1 _4634_ (.A(_2816_),
    .B(_0763_),
    .C(_0765_),
    .Y(_0766_));
 sg13g2_nand3_1 _4635_ (.B(net55),
    .C(_2901_),
    .A(_0683_),
    .Y(_0767_));
 sg13g2_a21oi_1 _4636_ (.A1(net77),
    .A2(net206),
    .Y(_0769_),
    .B1(net76));
 sg13g2_a21oi_1 _4637_ (.A1(_0627_),
    .A2(_0769_),
    .Y(_0770_),
    .B1(net81));
 sg13g2_nand2_1 _4638_ (.Y(_0771_),
    .A(_0767_),
    .B(_0770_));
 sg13g2_nand3_1 _4639_ (.B(net72),
    .C(_2853_),
    .A(_0125_),
    .Y(_0772_));
 sg13g2_a21oi_1 _4640_ (.A1(_0669_),
    .A2(_0583_),
    .Y(_0773_),
    .B1(net46));
 sg13g2_nand2_1 _4641_ (.Y(_0774_),
    .A(_0772_),
    .B(_0773_));
 sg13g2_o21ai_1 _4642_ (.B1(_2779_),
    .Y(_0775_),
    .A1(net33),
    .A2(_2888_));
 sg13g2_o21ai_1 _4643_ (.B1(_2373_),
    .Y(_0776_),
    .A1(net172),
    .A2(_2855_));
 sg13g2_a21oi_1 _4644_ (.A1(_2968_),
    .A2(_0775_),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_a22oi_1 _4645_ (.Y(_0778_),
    .B1(_0774_),
    .B2(_0777_),
    .A2(_0771_),
    .A1(_0766_));
 sg13g2_nand2_1 _4646_ (.Y(_0780_),
    .A(_0762_),
    .B(_0778_));
 sg13g2_nand2_1 _4647_ (.Y(_0781_),
    .A(_0780_),
    .B(net132));
 sg13g2_nand3_1 _4648_ (.B(_2433_),
    .C(_1522_),
    .A(net95),
    .Y(_0782_));
 sg13g2_a21oi_1 _4649_ (.A1(_0644_),
    .A2(_0782_),
    .Y(_0783_),
    .B1(_0118_));
 sg13g2_inv_1 _4650_ (.Y(_0784_),
    .A(net59));
 sg13g2_nand2_1 _4651_ (.Y(_0785_),
    .A(_0784_),
    .B(net94));
 sg13g2_nand3_1 _4652_ (.B(_2769_),
    .C(_0785_),
    .A(_0487_),
    .Y(_0786_));
 sg13g2_nor4_1 _4653_ (.A(net36),
    .B(_0337_),
    .C(_2453_),
    .D(_2520_),
    .Y(_0787_));
 sg13g2_a21oi_1 _4654_ (.A1(_0783_),
    .A2(_0786_),
    .Y(_0788_),
    .B1(_0787_));
 sg13g2_nand3_1 _4655_ (.B(_0514_),
    .C(net110),
    .A(_3017_),
    .Y(_0789_));
 sg13g2_inv_1 _4656_ (.Y(_0791_),
    .A(_1653_));
 sg13g2_o21ai_1 _4657_ (.B1(net69),
    .Y(_0792_),
    .A1(_0791_),
    .A2(_2806_));
 sg13g2_nand2_1 _4658_ (.Y(_0793_),
    .A(_0789_),
    .B(_0792_));
 sg13g2_nand2_1 _4659_ (.Y(_0794_),
    .A(_0793_),
    .B(net121));
 sg13g2_nand2_1 _4660_ (.Y(_0795_),
    .A(_1948_),
    .B(net182));
 sg13g2_nor2_1 _4661_ (.A(_0795_),
    .B(_2916_),
    .Y(_0796_));
 sg13g2_inv_1 _4662_ (.Y(_0797_),
    .A(_2532_));
 sg13g2_nor3_1 _4663_ (.A(_2732_),
    .B(_0797_),
    .C(_0673_),
    .Y(_0798_));
 sg13g2_o21ai_1 _4664_ (.B1(_3040_),
    .Y(_0799_),
    .A1(_0796_),
    .A2(_0798_));
 sg13g2_nand3_1 _4665_ (.B(_0794_),
    .C(_0799_),
    .A(_0788_),
    .Y(_0800_));
 sg13g2_nand2_1 _4666_ (.Y(_0802_),
    .A(_0800_),
    .B(net73));
 sg13g2_nor2_1 _4667_ (.A(_2467_),
    .B(_2880_),
    .Y(_0803_));
 sg13g2_nand2_1 _4668_ (.Y(_0804_),
    .A(_0803_),
    .B(_1921_));
 sg13g2_a21oi_1 _4669_ (.A1(_0804_),
    .A2(_0129_),
    .Y(_0805_),
    .B1(_2565_));
 sg13g2_a21oi_1 _4670_ (.A1(_0802_),
    .A2(_0805_),
    .Y(_0806_),
    .B1(net165));
 sg13g2_nand2_1 _4671_ (.Y(_0807_),
    .A(_0781_),
    .B(_0806_));
 sg13g2_nand2_2 _4672_ (.Y(_0808_),
    .A(_2020_),
    .B(net109));
 sg13g2_nand2_1 _4673_ (.Y(_0809_),
    .A(_0743_),
    .B(_0808_));
 sg13g2_nand3_1 _4674_ (.B(_3039_),
    .C(net88),
    .A(_0809_),
    .Y(_0810_));
 sg13g2_nor2_1 _4675_ (.A(net35),
    .B(_0673_),
    .Y(_0811_));
 sg13g2_nand2_1 _4676_ (.Y(_0813_),
    .A(_0409_),
    .B(_0811_));
 sg13g2_nand2_1 _4677_ (.Y(_0814_),
    .A(_0810_),
    .B(_0813_));
 sg13g2_a21oi_1 _4678_ (.A1(_2945_),
    .A2(_1653_),
    .Y(_0815_),
    .B1(_0337_));
 sg13g2_nor2_1 _4679_ (.A(net151),
    .B(_0797_),
    .Y(_0816_));
 sg13g2_nand2_1 _4680_ (.Y(_0817_),
    .A(_3025_),
    .B(_0816_));
 sg13g2_nand2_1 _4681_ (.Y(_0818_),
    .A(_0815_),
    .B(_0817_));
 sg13g2_nor2b_1 _4682_ (.A(_0814_),
    .B_N(_0818_),
    .Y(_0819_));
 sg13g2_nand2b_1 _4683_ (.Y(_0820_),
    .B(_0816_),
    .A_N(_3028_));
 sg13g2_nand2_1 _4684_ (.Y(_0821_),
    .A(_2606_),
    .B(_0820_));
 sg13g2_nand2_1 _4685_ (.Y(_0822_),
    .A(_0821_),
    .B(net107));
 sg13g2_nor2_1 _4686_ (.A(_1096_),
    .B(_0598_),
    .Y(_0824_));
 sg13g2_nand2_1 _4687_ (.Y(_0825_),
    .A(_1795_),
    .B(_1020_));
 sg13g2_nand2_1 _4688_ (.Y(_0826_),
    .A(_0825_),
    .B(_2444_));
 sg13g2_a22oi_1 _4689_ (.Y(_0827_),
    .B1(net39),
    .B2(_0826_),
    .A2(_0824_),
    .A1(_0471_));
 sg13g2_nand2_1 _4690_ (.Y(_0828_),
    .A(_0822_),
    .B(_0827_));
 sg13g2_nand2_1 _4691_ (.Y(_0829_),
    .A(_0828_),
    .B(net131));
 sg13g2_nand2_1 _4692_ (.Y(_0830_),
    .A(_0819_),
    .B(_0829_));
 sg13g2_nand2_1 _4693_ (.Y(_0831_),
    .A(_0830_),
    .B(_0090_));
 sg13g2_nand2_1 _4694_ (.Y(_0832_),
    .A(_0563_),
    .B(_2589_));
 sg13g2_nand2_1 _4695_ (.Y(_0833_),
    .A(net103),
    .B(_2633_));
 sg13g2_and3_1 _4696_ (.X(_0835_),
    .A(_0832_),
    .B(net72),
    .C(_0833_));
 sg13g2_o21ai_1 _4697_ (.B1(net130),
    .Y(_0836_),
    .A1(_0346_),
    .A2(_0518_));
 sg13g2_o21ai_1 _4698_ (.B1(net169),
    .Y(_0837_),
    .A1(net168),
    .A2(_0589_));
 sg13g2_nand2_1 _4699_ (.Y(_0838_),
    .A(_2967_),
    .B(net92));
 sg13g2_nand2_1 _4700_ (.Y(_0839_),
    .A(_2414_),
    .B(net27));
 sg13g2_a21oi_1 _4701_ (.A1(_0838_),
    .A2(_0839_),
    .Y(_0840_),
    .B1(_2408_));
 sg13g2_nor2_1 _4702_ (.A(_0837_),
    .B(_0840_),
    .Y(_0841_));
 sg13g2_o21ai_1 _4703_ (.B1(_0841_),
    .Y(_0842_),
    .A1(_0835_),
    .A2(_0836_));
 sg13g2_a21o_1 _4704_ (.A2(_0785_),
    .A1(_2656_),
    .B1(net61),
    .X(_0843_));
 sg13g2_a22oi_1 _4705_ (.Y(_0844_),
    .B1(net201),
    .B2(_0142_),
    .A2(_1457_),
    .A1(net103));
 sg13g2_nor2_1 _4706_ (.A(net138),
    .B(_2453_),
    .Y(_0846_));
 sg13g2_nand2_1 _4707_ (.Y(_0847_),
    .A(_2854_),
    .B(net158));
 sg13g2_nand2_1 _4708_ (.Y(_0848_),
    .A(_2392_),
    .B(net58));
 sg13g2_nand3_1 _4709_ (.B(_0848_),
    .C(net69),
    .A(_0847_),
    .Y(_0849_));
 sg13g2_nand2_1 _4710_ (.Y(_0850_),
    .A(_0849_),
    .B(net123));
 sg13g2_a21oi_1 _4711_ (.A1(_0844_),
    .A2(_0846_),
    .Y(_0851_),
    .B1(_0850_));
 sg13g2_nand2_1 _4712_ (.Y(_0852_),
    .A(_0742_),
    .B(_2416_));
 sg13g2_nand2_1 _4713_ (.Y(_0853_),
    .A(_0852_),
    .B(_2861_));
 sg13g2_nand2_1 _4714_ (.Y(_0854_),
    .A(_0853_),
    .B(net26));
 sg13g2_nand3_1 _4715_ (.B(_0851_),
    .C(_0854_),
    .A(_0843_),
    .Y(_0855_));
 sg13g2_nand3_1 _4716_ (.B(_0855_),
    .C(net164),
    .A(_0842_),
    .Y(_0857_));
 sg13g2_nand3_1 _4717_ (.B(_0857_),
    .C(_2738_),
    .A(_0831_),
    .Y(_0858_));
 sg13g2_inv_1 _4718_ (.Y(_0859_),
    .A(_0470_));
 sg13g2_o21ai_1 _4719_ (.B1(net99),
    .Y(_0860_),
    .A1(_0568_),
    .A2(_0859_));
 sg13g2_nand3_1 _4720_ (.B(net24),
    .C(_2920_),
    .A(_0514_),
    .Y(_0861_));
 sg13g2_a21oi_1 _4721_ (.A1(_0860_),
    .A2(_0861_),
    .Y(_0862_),
    .B1(net66));
 sg13g2_inv_1 _4722_ (.Y(_0863_),
    .A(_0716_));
 sg13g2_o21ai_1 _4723_ (.B1(_0220_),
    .Y(_0864_),
    .A1(_0548_),
    .A2(_2801_));
 sg13g2_o21ai_1 _4724_ (.B1(_0864_),
    .Y(_0865_),
    .A1(_2279_),
    .A2(_0863_));
 sg13g2_nor2_1 _4725_ (.A(net202),
    .B(_0482_),
    .Y(_0866_));
 sg13g2_inv_1 _4726_ (.Y(_0868_),
    .A(_0866_));
 sg13g2_nor2b_1 _4727_ (.A(_0510_),
    .B_N(_2861_),
    .Y(_0869_));
 sg13g2_o21ai_1 _4728_ (.B1(_2598_),
    .Y(_0870_),
    .A1(_0868_),
    .A2(_0869_));
 sg13g2_a21oi_1 _4729_ (.A1(_0865_),
    .A2(_0521_),
    .Y(_0871_),
    .B1(_0870_));
 sg13g2_nand2_1 _4730_ (.Y(_0872_),
    .A(_0259_),
    .B(_0704_));
 sg13g2_a21oi_1 _4731_ (.A1(_0487_),
    .A2(_2536_),
    .Y(_0873_),
    .B1(net35));
 sg13g2_nand2_1 _4732_ (.Y(_0874_),
    .A(_0872_),
    .B(_0873_));
 sg13g2_a21o_1 _4733_ (.A2(_2496_),
    .A1(_0832_),
    .B1(net37),
    .X(_0875_));
 sg13g2_nand2b_1 _4734_ (.Y(_0876_),
    .B(net113),
    .A_N(_0875_));
 sg13g2_nand3_1 _4735_ (.B(_0874_),
    .C(_0876_),
    .A(_0871_),
    .Y(_0877_));
 sg13g2_nor2_1 _4736_ (.A(_0862_),
    .B(_0877_),
    .Y(_0879_));
 sg13g2_nand3_1 _4737_ (.B(_0669_),
    .C(_2990_),
    .A(_2967_),
    .Y(_0880_));
 sg13g2_o21ai_1 _4738_ (.B1(net88),
    .Y(_0881_),
    .A1(_0438_),
    .A2(_2775_));
 sg13g2_a21oi_1 _4739_ (.A1(_0880_),
    .A2(_0881_),
    .Y(_0882_),
    .B1(net127));
 sg13g2_nand2_1 _4740_ (.Y(_0883_),
    .A(_2970_),
    .B(net149));
 sg13g2_nor2_1 _4741_ (.A(net174),
    .B(_0548_),
    .Y(_0884_));
 sg13g2_a21oi_1 _4742_ (.A1(_2622_),
    .A2(_0884_),
    .Y(_0885_),
    .B1(_0118_));
 sg13g2_o21ai_1 _4743_ (.B1(_0885_),
    .Y(_0886_),
    .A1(_0134_),
    .A2(_0883_));
 sg13g2_nand2_1 _4744_ (.Y(_0887_),
    .A(_0886_),
    .B(net112));
 sg13g2_nor2_1 _4745_ (.A(_0882_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_a21oi_1 _4746_ (.A1(_2978_),
    .A2(_2482_),
    .Y(_0890_),
    .B1(net107));
 sg13g2_nand2_1 _4747_ (.Y(_0891_),
    .A(_0875_),
    .B(_0890_));
 sg13g2_nand2_1 _4748_ (.Y(_0892_),
    .A(net124),
    .B(net193));
 sg13g2_a21oi_1 _4749_ (.A1(_2677_),
    .A2(net142),
    .Y(_0893_),
    .B1(_0892_));
 sg13g2_nand2_1 _4750_ (.Y(_0894_),
    .A(_0563_),
    .B(net36));
 sg13g2_a21oi_1 _4751_ (.A1(_0893_),
    .A2(_0894_),
    .Y(_0895_),
    .B1(net167));
 sg13g2_nand2_1 _4752_ (.Y(_0896_),
    .A(_0891_),
    .B(_0895_));
 sg13g2_a21oi_1 _4753_ (.A1(_0888_),
    .A2(_0896_),
    .Y(_0897_),
    .B1(_2609_));
 sg13g2_nor2b_1 _4754_ (.A(_0879_),
    .B_N(_0897_),
    .Y(_0898_));
 sg13g2_nand2_1 _4755_ (.Y(_0899_),
    .A(_0858_),
    .B(_0898_));
 sg13g2_nand2_1 _4756_ (.Y(_0026_),
    .A(_0807_),
    .B(_0899_));
 sg13g2_nand2_1 _4757_ (.Y(_0901_),
    .A(_0573_),
    .B(_2491_));
 sg13g2_nand2_1 _4758_ (.Y(_0902_),
    .A(_0901_),
    .B(_0470_));
 sg13g2_nand2_1 _4759_ (.Y(_0903_),
    .A(_0902_),
    .B(net42));
 sg13g2_a21oi_1 _4760_ (.A1(_3036_),
    .A2(_1948_),
    .Y(_0904_),
    .B1(net101));
 sg13g2_nor2_1 _4761_ (.A(_1685_),
    .B(_2378_),
    .Y(_0905_));
 sg13g2_nand3_1 _4762_ (.B(net135),
    .C(_0905_),
    .A(_0563_),
    .Y(_0906_));
 sg13g2_nand2_1 _4763_ (.Y(_0907_),
    .A(_2603_),
    .B(net146));
 sg13g2_nand2_1 _4764_ (.Y(_0908_),
    .A(_0907_),
    .B(net104));
 sg13g2_nand2_1 _4765_ (.Y(_0909_),
    .A(_0906_),
    .B(_0908_));
 sg13g2_nor2_1 _4766_ (.A(_0904_),
    .B(_0909_),
    .Y(_0911_));
 sg13g2_nand2_1 _4767_ (.Y(_0912_),
    .A(_0903_),
    .B(_0911_));
 sg13g2_nand2_1 _4768_ (.Y(_0913_),
    .A(_0912_),
    .B(net121));
 sg13g2_o21ai_1 _4769_ (.B1(_0564_),
    .Y(_0914_),
    .A1(_0976_),
    .A2(_0622_));
 sg13g2_nor2_2 _4770_ (.A(_0127_),
    .B(net180),
    .Y(_0915_));
 sg13g2_nand2_1 _4771_ (.Y(_0916_),
    .A(_0915_),
    .B(_2460_));
 sg13g2_inv_1 _4772_ (.Y(_0917_),
    .A(_0916_));
 sg13g2_nor2_1 _4773_ (.A(net140),
    .B(_2947_),
    .Y(_0918_));
 sg13g2_nor2_1 _4774_ (.A(_3047_),
    .B(_0918_),
    .Y(_0919_));
 sg13g2_a21oi_1 _4775_ (.A1(_0919_),
    .A2(net84),
    .Y(_0920_),
    .B1(_0716_));
 sg13g2_a22oi_1 _4776_ (.Y(_0922_),
    .B1(net115),
    .B2(_0920_),
    .A2(_0917_),
    .A1(_0914_));
 sg13g2_nand2_1 _4777_ (.Y(_0923_),
    .A(_0913_),
    .B(_0922_));
 sg13g2_nand2_1 _4778_ (.Y(_0924_),
    .A(_0923_),
    .B(_2785_));
 sg13g2_nor2_1 _4779_ (.A(_1707_),
    .B(_0673_),
    .Y(_0925_));
 sg13g2_inv_1 _4780_ (.Y(_0926_),
    .A(_0648_));
 sg13g2_nor2_1 _4781_ (.A(_0598_),
    .B(_0926_),
    .Y(_0927_));
 sg13g2_a22oi_1 _4782_ (.Y(_0928_),
    .B1(net50),
    .B2(_0927_),
    .A2(_0825_),
    .A1(_0925_));
 sg13g2_o21ai_1 _4783_ (.B1(net32),
    .Y(_0929_),
    .A1(net85),
    .A2(_2429_));
 sg13g2_a21oi_1 _4784_ (.A1(_0928_),
    .A2(_0929_),
    .Y(_0930_),
    .B1(_2816_));
 sg13g2_nand2_1 _4785_ (.Y(_0931_),
    .A(_0803_),
    .B(_0250_));
 sg13g2_nand2_1 _4786_ (.Y(_0933_),
    .A(_0931_),
    .B(net53));
 sg13g2_nor2_1 _4787_ (.A(_2537_),
    .B(_1805_),
    .Y(_0934_));
 sg13g2_nand2_1 _4788_ (.Y(_0935_),
    .A(_0934_),
    .B(_2810_));
 sg13g2_a21oi_1 _4789_ (.A1(_0935_),
    .A2(net74),
    .Y(_0936_),
    .B1(_2462_));
 sg13g2_a21oi_1 _4790_ (.A1(_0933_),
    .A2(_0936_),
    .Y(_0937_),
    .B1(net63));
 sg13g2_nor2_1 _4791_ (.A(_0930_),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_nand2_1 _4792_ (.Y(_0939_),
    .A(_0924_),
    .B(_0938_));
 sg13g2_nor2_1 _4793_ (.A(net128),
    .B(_0372_),
    .Y(_0940_));
 sg13g2_o21ai_1 _4794_ (.B1(_0940_),
    .Y(_0941_),
    .A1(net33),
    .A2(_2031_));
 sg13g2_nand2_1 _4795_ (.Y(_0942_),
    .A(net193),
    .B(_2543_));
 sg13g2_o21ai_1 _4796_ (.B1(_2533_),
    .Y(_0944_),
    .A1(_0942_),
    .A2(_0607_));
 sg13g2_a21oi_1 _4797_ (.A1(_0351_),
    .A2(_2856_),
    .Y(_0945_),
    .B1(_2963_));
 sg13g2_a21oi_1 _4798_ (.A1(_0941_),
    .A2(_0944_),
    .Y(_0946_),
    .B1(_0945_));
 sg13g2_nor3_1 _4799_ (.A(net180),
    .B(net193),
    .C(_0128_),
    .Y(_0947_));
 sg13g2_inv_1 _4800_ (.Y(_0948_),
    .A(_0947_));
 sg13g2_nor2_1 _4801_ (.A(net203),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_nand4_1 _4802_ (.B(_1948_),
    .C(_2605_),
    .A(_2430_),
    .Y(_0950_),
    .D(net120));
 sg13g2_nand2_1 _4803_ (.Y(_0951_),
    .A(_2854_),
    .B(net96));
 sg13g2_nand2_1 _4804_ (.Y(_0952_),
    .A(_0951_),
    .B(_2795_));
 sg13g2_a21oi_1 _4805_ (.A1(_0739_),
    .A2(_0952_),
    .Y(_0953_),
    .B1(net66));
 sg13g2_a22oi_1 _4806_ (.Y(_0955_),
    .B1(_0950_),
    .B2(_0953_),
    .A2(_0949_),
    .A1(_0339_));
 sg13g2_o21ai_1 _4807_ (.B1(_0955_),
    .Y(_0956_),
    .A1(net83),
    .A2(_0946_));
 sg13g2_nand2_1 _4808_ (.Y(_0957_),
    .A(_0956_),
    .B(net112));
 sg13g2_a21oi_1 _4809_ (.A1(net44),
    .A2(net86),
    .Y(_0958_),
    .B1(net174));
 sg13g2_nor2_1 _4810_ (.A(_2564_),
    .B(_0303_),
    .Y(_0959_));
 sg13g2_inv_1 _4811_ (.Y(_0960_),
    .A(_0959_));
 sg13g2_a221oi_1 _4812_ (.B2(_2959_),
    .C1(_0960_),
    .B1(_0958_),
    .A1(_2740_),
    .Y(_0961_),
    .A2(_0321_));
 sg13g2_nor2_1 _4813_ (.A(net195),
    .B(_0961_),
    .Y(_0962_));
 sg13g2_nand2_1 _4814_ (.Y(_0963_),
    .A(_0957_),
    .B(_0962_));
 sg13g2_a21oi_1 _4815_ (.A1(_0939_),
    .A2(net132),
    .Y(_0964_),
    .B1(_0963_));
 sg13g2_a21oi_1 _4816_ (.A1(_1968_),
    .A2(_2807_),
    .Y(_0966_),
    .B1(net81));
 sg13g2_nand2_1 _4817_ (.Y(_0967_),
    .A(_0371_),
    .B(_0460_));
 sg13g2_nand2_1 _4818_ (.Y(_0968_),
    .A(_0966_),
    .B(_0967_));
 sg13g2_nand3_1 _4819_ (.B(net94),
    .C(net27),
    .A(net71),
    .Y(_0969_));
 sg13g2_a21oi_1 _4820_ (.A1(_0969_),
    .A2(_1293_),
    .Y(_0970_),
    .B1(net40));
 sg13g2_nor2_1 _4821_ (.A(net198),
    .B(_2687_),
    .Y(_0971_));
 sg13g2_inv_1 _4822_ (.Y(_0972_),
    .A(_2947_));
 sg13g2_a21oi_1 _4823_ (.A1(_0971_),
    .A2(_0972_),
    .Y(_0973_),
    .B1(net203));
 sg13g2_nor2b_1 _4824_ (.A(_0970_),
    .B_N(_0973_),
    .Y(_0974_));
 sg13g2_nand2_1 _4825_ (.Y(_0975_),
    .A(_0968_),
    .B(_0974_));
 sg13g2_nand2_1 _4826_ (.Y(_0977_),
    .A(_0142_),
    .B(_2411_));
 sg13g2_a21oi_1 _4827_ (.A1(_0321_),
    .A2(_0977_),
    .Y(_0978_),
    .B1(net54));
 sg13g2_nand2_1 _4828_ (.Y(_0979_),
    .A(_0703_),
    .B(net65));
 sg13g2_nand2_1 _4829_ (.Y(_0980_),
    .A(_0979_),
    .B(net169));
 sg13g2_nor2_1 _4830_ (.A(_0978_),
    .B(_0980_),
    .Y(_0981_));
 sg13g2_nand2_1 _4831_ (.Y(_0982_),
    .A(_2800_),
    .B(net97));
 sg13g2_nand2_1 _4832_ (.Y(_0983_),
    .A(_0982_),
    .B(_2842_));
 sg13g2_nand2_1 _4833_ (.Y(_0984_),
    .A(_0983_),
    .B(_2703_));
 sg13g2_nand2_1 _4834_ (.Y(_0985_),
    .A(_0984_),
    .B(net46));
 sg13g2_nand2_1 _4835_ (.Y(_0986_),
    .A(_2881_),
    .B(net50));
 sg13g2_nand3_1 _4836_ (.B(_0985_),
    .C(_0986_),
    .A(_0981_),
    .Y(_0988_));
 sg13g2_nand3_1 _4837_ (.B(_0988_),
    .C(net147),
    .A(_0975_),
    .Y(_0989_));
 sg13g2_nand2_1 _4838_ (.Y(_0990_),
    .A(_1446_),
    .B(net144));
 sg13g2_nand2_1 _4839_ (.Y(_0991_),
    .A(_0990_),
    .B(net56));
 sg13g2_nand3_1 _4840_ (.B(net67),
    .C(_0354_),
    .A(_0991_),
    .Y(_0992_));
 sg13g2_a21oi_1 _4841_ (.A1(_0919_),
    .A2(net45),
    .Y(_0993_),
    .B1(net172));
 sg13g2_nand2_1 _4842_ (.Y(_0994_),
    .A(_0992_),
    .B(_0993_));
 sg13g2_a21oi_2 _4843_ (.B1(_2450_),
    .Y(_0995_),
    .A2(net139),
    .A1(_2440_));
 sg13g2_nand3_1 _4844_ (.B(_0161_),
    .C(_0995_),
    .A(_2932_),
    .Y(_0996_));
 sg13g2_a22oi_1 _4845_ (.Y(_0997_),
    .B1(net86),
    .B2(net44),
    .A2(_1478_),
    .A1(net27));
 sg13g2_a21oi_1 _4846_ (.A1(net47),
    .A2(_0527_),
    .Y(_0999_),
    .B1(net128));
 sg13g2_a21oi_1 _4847_ (.A1(_0997_),
    .A2(_0999_),
    .Y(_1000_),
    .B1(_2716_));
 sg13g2_nand2_1 _4848_ (.Y(_1001_),
    .A(_0996_),
    .B(_1000_));
 sg13g2_nand2_1 _4849_ (.Y(_1002_),
    .A(_0994_),
    .B(_1001_));
 sg13g2_nand2_1 _4850_ (.Y(_1003_),
    .A(_1002_),
    .B(_2559_));
 sg13g2_nand2_1 _4851_ (.Y(_1004_),
    .A(_2948_),
    .B(net125));
 sg13g2_nor3_1 _4852_ (.A(net36),
    .B(net168),
    .C(_2745_),
    .Y(_1005_));
 sg13g2_nand3_1 _4853_ (.B(net82),
    .C(net48),
    .A(_2860_),
    .Y(_1006_));
 sg13g2_nand2_1 _4854_ (.Y(_1007_),
    .A(_1006_),
    .B(_0167_));
 sg13g2_inv_1 _4855_ (.Y(_1008_),
    .A(_0795_));
 sg13g2_a21oi_1 _4856_ (.A1(_1008_),
    .A2(_2705_),
    .Y(_1010_),
    .B1(net78));
 sg13g2_a22oi_1 _4857_ (.Y(_1011_),
    .B1(_1007_),
    .B2(_1010_),
    .A2(_1005_),
    .A1(_1004_));
 sg13g2_nor2_1 _4858_ (.A(net210),
    .B(_0478_),
    .Y(_1012_));
 sg13g2_inv_2 _4859_ (.Y(_1013_),
    .A(_1012_));
 sg13g2_nand2_1 _4860_ (.Y(_1014_),
    .A(_1011_),
    .B(_1013_));
 sg13g2_nand2_1 _4861_ (.Y(_1015_),
    .A(_1014_),
    .B(_2373_));
 sg13g2_nand3_1 _4862_ (.B(_1003_),
    .C(_1015_),
    .A(_0989_),
    .Y(_1016_));
 sg13g2_nand3_1 _4863_ (.B(_2727_),
    .C(net84),
    .A(_2850_),
    .Y(_1017_));
 sg13g2_nand2_1 _4864_ (.Y(_1018_),
    .A(_0350_),
    .B(_0951_));
 sg13g2_nand3_1 _4865_ (.B(net45),
    .C(_2591_),
    .A(_1018_),
    .Y(_1019_));
 sg13g2_nand3_1 _4866_ (.B(_1019_),
    .C(net46),
    .A(_1017_),
    .Y(_1021_));
 sg13g2_a21oi_1 _4867_ (.A1(_0150_),
    .A2(_2727_),
    .Y(_1022_),
    .B1(net145));
 sg13g2_nand2_1 _4868_ (.Y(_1023_),
    .A(_0240_),
    .B(_2935_));
 sg13g2_o21ai_1 _4869_ (.B1(_2698_),
    .Y(_1024_),
    .A1(_1023_),
    .A2(_2657_));
 sg13g2_nor2_1 _4870_ (.A(_1022_),
    .B(_1024_),
    .Y(_1025_));
 sg13g2_nand2_1 _4871_ (.Y(_1026_),
    .A(_1021_),
    .B(_1025_));
 sg13g2_nand2_1 _4872_ (.Y(_1027_),
    .A(_0438_),
    .B(_0602_));
 sg13g2_nand3_1 _4873_ (.B(net65),
    .C(_2435_),
    .A(_2793_),
    .Y(_1028_));
 sg13g2_o21ai_1 _4874_ (.B1(_1028_),
    .Y(_1029_),
    .A1(net28),
    .A2(_1027_));
 sg13g2_nand2_1 _4875_ (.Y(_1030_),
    .A(_1013_),
    .B(net169));
 sg13g2_nor2_1 _4876_ (.A(_1029_),
    .B(_1030_),
    .Y(_1032_));
 sg13g2_nand2_1 _4877_ (.Y(_1033_),
    .A(_2592_),
    .B(net53));
 sg13g2_a21oi_1 _4878_ (.A1(_1032_),
    .A2(_1033_),
    .Y(_1034_),
    .B1(_2597_));
 sg13g2_a21oi_1 _4879_ (.A1(_1026_),
    .A2(_1034_),
    .Y(_1035_),
    .B1(_2609_));
 sg13g2_nor2_1 _4880_ (.A(_2704_),
    .B(net59),
    .Y(_1036_));
 sg13g2_nor3_1 _4881_ (.A(net91),
    .B(_2279_),
    .C(_1036_),
    .Y(_1037_));
 sg13g2_nand2_1 _4882_ (.Y(_1038_),
    .A(_2571_),
    .B(net44));
 sg13g2_nand2_1 _4883_ (.Y(_1039_),
    .A(_1038_),
    .B(net108));
 sg13g2_a21oi_1 _4884_ (.A1(_0350_),
    .A2(_0951_),
    .Y(_1040_),
    .B1(_1039_));
 sg13g2_nor3_1 _4885_ (.A(net162),
    .B(_1037_),
    .C(_1040_),
    .Y(_1041_));
 sg13g2_a21oi_1 _4886_ (.A1(_2797_),
    .A2(_0135_),
    .Y(_1043_),
    .B1(_2445_));
 sg13g2_nand2_1 _4887_ (.Y(_1044_),
    .A(net71),
    .B(_1184_));
 sg13g2_nor2_2 _4888_ (.A(_1685_),
    .B(_2701_),
    .Y(_1045_));
 sg13g2_a21oi_1 _4889_ (.A1(_1044_),
    .A2(_1045_),
    .Y(_1046_),
    .B1(net161));
 sg13g2_nand2b_1 _4890_ (.Y(_1047_),
    .B(_1046_),
    .A_N(_1043_));
 sg13g2_nor2_1 _4891_ (.A(_1041_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_nor2_1 _4892_ (.A(_0729_),
    .B(_1048_),
    .Y(_1049_));
 sg13g2_nor2_1 _4893_ (.A(net140),
    .B(_2458_),
    .Y(_1050_));
 sg13g2_nor2_1 _4894_ (.A(_0264_),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_a21oi_1 _4895_ (.A1(_1051_),
    .A2(net36),
    .Y(_1052_),
    .B1(_2595_));
 sg13g2_nand3_1 _4896_ (.B(net133),
    .C(_0422_),
    .A(_2577_),
    .Y(_1054_));
 sg13g2_a21oi_1 _4897_ (.A1(_1052_),
    .A2(_1054_),
    .Y(_1055_),
    .B1(_2141_));
 sg13g2_nand3_1 _4898_ (.B(_1522_),
    .C(net133),
    .A(net94),
    .Y(_1056_));
 sg13g2_nor2_1 _4899_ (.A(net90),
    .B(_2257_),
    .Y(_1057_));
 sg13g2_nor2_1 _4900_ (.A(_1751_),
    .B(_1057_),
    .Y(_1058_));
 sg13g2_a21oi_1 _4901_ (.A1(_1056_),
    .A2(_1058_),
    .Y(_1059_),
    .B1(net172));
 sg13g2_nand3_1 _4902_ (.B(net67),
    .C(_0418_),
    .A(_2579_),
    .Y(_1060_));
 sg13g2_a22oi_1 _4903_ (.Y(_1061_),
    .B1(_1059_),
    .B2(_1060_),
    .A2(_0324_),
    .A1(net25));
 sg13g2_nand2b_1 _4904_ (.Y(_1062_),
    .B(_1061_),
    .A_N(_1055_));
 sg13g2_nand2_1 _4905_ (.Y(_1063_),
    .A(_1049_),
    .B(_1062_));
 sg13g2_nand2_1 _4906_ (.Y(_1065_),
    .A(_1035_),
    .B(_1063_));
 sg13g2_a21oi_1 _4907_ (.A1(_1016_),
    .A2(net132),
    .Y(_1066_),
    .B1(_1065_));
 sg13g2_nor2_1 _4908_ (.A(_0964_),
    .B(_1066_),
    .Y(_0027_));
 sg13g2_nand3_1 _4909_ (.B(_2727_),
    .C(_2654_),
    .A(_0838_),
    .Y(_1067_));
 sg13g2_a21oi_1 _4910_ (.A1(_2743_),
    .A2(_0808_),
    .Y(_1068_),
    .B1(_2760_));
 sg13g2_nand2_1 _4911_ (.Y(_1069_),
    .A(_1067_),
    .B(_1068_));
 sg13g2_o21ai_1 _4912_ (.B1(_2991_),
    .Y(_1070_),
    .A1(_2723_),
    .A2(_0145_));
 sg13g2_nor2_1 _4913_ (.A(net180),
    .B(_0795_),
    .Y(_1071_));
 sg13g2_nand2b_1 _4914_ (.Y(_1072_),
    .B(_1071_),
    .A_N(_2772_));
 sg13g2_nand4_1 _4915_ (.B(_1070_),
    .C(net80),
    .A(_1069_),
    .Y(_1073_),
    .D(_1072_));
 sg13g2_a21oi_1 _4916_ (.A1(_0234_),
    .A2(_0977_),
    .Y(_1075_),
    .B1(_0294_));
 sg13g2_nand3_1 _4917_ (.B(net38),
    .C(net65),
    .A(_2503_),
    .Y(_1076_));
 sg13g2_nor2_1 _4918_ (.A(_0651_),
    .B(_1027_),
    .Y(_1077_));
 sg13g2_nor2_1 _4919_ (.A(_2480_),
    .B(_1077_),
    .Y(_1078_));
 sg13g2_nand3b_1 _4920_ (.B(_1076_),
    .C(_1078_),
    .Y(_1079_),
    .A_N(_1075_));
 sg13g2_a21oi_1 _4921_ (.A1(_1073_),
    .A2(_1079_),
    .Y(_1080_),
    .B1(_2597_));
 sg13g2_nand2_1 _4922_ (.Y(_1081_),
    .A(_2477_),
    .B(net133));
 sg13g2_a22oi_1 _4923_ (.Y(_1082_),
    .B1(net134),
    .B2(_2892_),
    .A2(_1081_),
    .A1(_1045_));
 sg13g2_inv_1 _4924_ (.Y(_1083_),
    .A(_2642_));
 sg13g2_nand3_1 _4925_ (.B(_2779_),
    .C(_2516_),
    .A(_1083_),
    .Y(_1084_));
 sg13g2_a21oi_1 _4926_ (.A1(_1082_),
    .A2(_1084_),
    .Y(_1086_),
    .B1(net123));
 sg13g2_a221oi_1 _4927_ (.B2(_0627_),
    .C1(_0338_),
    .B1(_3030_),
    .A1(_2789_),
    .Y(_1087_),
    .A2(_2769_));
 sg13g2_nand2_1 _4928_ (.Y(_1088_),
    .A(_0438_),
    .B(_2482_));
 sg13g2_inv_1 _4929_ (.Y(_1089_),
    .A(_1088_));
 sg13g2_a21oi_1 _4930_ (.A1(_2728_),
    .A2(_2800_),
    .Y(_1090_),
    .B1(_1958_));
 sg13g2_o21ai_1 _4931_ (.B1(net22),
    .Y(_1091_),
    .A1(_1089_),
    .A2(_1090_));
 sg13g2_nand2_1 _4932_ (.Y(_1092_),
    .A(_1091_),
    .B(net112));
 sg13g2_nor3_1 _4933_ (.A(_1086_),
    .B(_1087_),
    .C(_1092_),
    .Y(_1093_));
 sg13g2_o21ai_1 _4934_ (.B1(_0394_),
    .Y(_1094_),
    .A1(net48),
    .A2(_2848_));
 sg13g2_a22oi_1 _4935_ (.Y(_1095_),
    .B1(_2568_),
    .B2(_1094_),
    .A2(_0360_),
    .A1(_0565_));
 sg13g2_nand2_1 _4936_ (.Y(_1097_),
    .A(_0428_),
    .B(_2496_));
 sg13g2_o21ai_1 _4937_ (.B1(_2895_),
    .Y(_1098_),
    .A1(_0477_),
    .A2(_1097_));
 sg13g2_nand2_1 _4938_ (.Y(_1099_),
    .A(_1095_),
    .B(_1098_));
 sg13g2_nand2_1 _4939_ (.Y(_1100_),
    .A(_1099_),
    .B(_2699_));
 sg13g2_nand2_1 _4940_ (.Y(_1101_),
    .A(_1093_),
    .B(_1100_));
 sg13g2_nand2_1 _4941_ (.Y(_1102_),
    .A(_1101_),
    .B(net195));
 sg13g2_nor2_1 _4942_ (.A(_1080_),
    .B(_1102_),
    .Y(_1103_));
 sg13g2_nor2_2 _4943_ (.A(_1751_),
    .B(_0477_),
    .Y(_1104_));
 sg13g2_nor2_1 _4944_ (.A(_2577_),
    .B(_2478_),
    .Y(_1105_));
 sg13g2_nor2_1 _4945_ (.A(_2642_),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_nor2_1 _4946_ (.A(_1104_),
    .B(_1106_),
    .Y(_1108_));
 sg13g2_nand2_1 _4947_ (.Y(_1109_),
    .A(_2487_),
    .B(_2554_));
 sg13g2_a21o_1 _4948_ (.A2(_2482_),
    .A1(_1109_),
    .B1(_0576_),
    .X(_1110_));
 sg13g2_a22oi_1 _4949_ (.Y(_1111_),
    .B1(net105),
    .B2(_1110_),
    .A2(_2141_),
    .A1(_1108_));
 sg13g2_nor3_1 _4950_ (.A(net89),
    .B(net29),
    .C(_0148_),
    .Y(_1112_));
 sg13g2_nand2_1 _4951_ (.Y(_1113_),
    .A(_1112_),
    .B(_1004_));
 sg13g2_nand2_1 _4952_ (.Y(_1114_),
    .A(_2992_),
    .B(_2673_));
 sg13g2_nand3_1 _4953_ (.B(_1114_),
    .C(net45),
    .A(_1038_),
    .Y(_1115_));
 sg13g2_nand3_1 _4954_ (.B(_1115_),
    .C(net113),
    .A(_1113_),
    .Y(_1116_));
 sg13g2_a22oi_1 _4955_ (.Y(_1117_),
    .B1(_0321_),
    .B2(_0769_),
    .A2(_2964_),
    .A1(_2715_));
 sg13g2_nand2_1 _4956_ (.Y(_1119_),
    .A(_1117_),
    .B(net22));
 sg13g2_nand3_1 _4957_ (.B(_1116_),
    .C(_1119_),
    .A(_1111_),
    .Y(_1120_));
 sg13g2_nand2_1 _4958_ (.Y(_1121_),
    .A(_1120_),
    .B(net164));
 sg13g2_a21oi_1 _4959_ (.A1(_0743_),
    .A2(_3043_),
    .Y(_1122_),
    .B1(net61));
 sg13g2_nor2_1 _4960_ (.A(net28),
    .B(_0226_),
    .Y(_1123_));
 sg13g2_inv_1 _4961_ (.Y(_1124_),
    .A(_2462_));
 sg13g2_nand2_1 _4962_ (.Y(_1125_),
    .A(_1124_),
    .B(net173));
 sg13g2_a21oi_1 _4963_ (.A1(_1293_),
    .A2(_2681_),
    .Y(_1126_),
    .B1(net138));
 sg13g2_nor3_1 _4964_ (.A(_1123_),
    .B(_1125_),
    .C(_1126_),
    .Y(_1127_));
 sg13g2_nor3_1 _4965_ (.A(_2506_),
    .B(_2411_),
    .C(_0289_),
    .Y(_1128_));
 sg13g2_o21ai_1 _4966_ (.B1(net53),
    .Y(_1130_),
    .A1(_2520_),
    .A2(_1128_));
 sg13g2_nand3b_1 _4967_ (.B(_1127_),
    .C(_1130_),
    .Y(_1131_),
    .A_N(_1122_));
 sg13g2_nand2_1 _4968_ (.Y(_1132_),
    .A(_2901_),
    .B(_2444_));
 sg13g2_a22oi_1 _4969_ (.Y(_1133_),
    .B1(net50),
    .B2(_1132_),
    .A2(net65),
    .A1(_0264_));
 sg13g2_o21ai_1 _4970_ (.B1(net32),
    .Y(_1134_),
    .A1(_2470_),
    .A2(_2880_));
 sg13g2_a21oi_2 _4971_ (.B1(_2460_),
    .Y(_1135_),
    .A2(net124),
    .A1(_1089_));
 sg13g2_nand3_1 _4972_ (.B(_1134_),
    .C(_1135_),
    .A(_1133_),
    .Y(_1136_));
 sg13g2_nand3_1 _4973_ (.B(net73),
    .C(_1136_),
    .A(_1131_),
    .Y(_1137_));
 sg13g2_nand3_1 _4974_ (.B(_1137_),
    .C(_2738_),
    .A(_1121_),
    .Y(_1138_));
 sg13g2_nand2_1 _4975_ (.Y(_1139_),
    .A(_1103_),
    .B(_1138_));
 sg13g2_a21oi_1 _4976_ (.A1(net52),
    .A2(_1260_),
    .Y(_1141_),
    .B1(net108));
 sg13g2_nand3_1 _4977_ (.B(_2856_),
    .C(net176),
    .A(_1141_),
    .Y(_1142_));
 sg13g2_nand3_1 _4978_ (.B(_2518_),
    .C(_0848_),
    .A(_2239_),
    .Y(_1143_));
 sg13g2_nand3_1 _4979_ (.B(_1143_),
    .C(_2760_),
    .A(_1142_),
    .Y(_1144_));
 sg13g2_nor2_1 _4980_ (.A(net151),
    .B(_1869_),
    .Y(_1145_));
 sg13g2_o21ai_1 _4981_ (.B1(_1145_),
    .Y(_1146_),
    .A1(_0198_),
    .A2(_2572_));
 sg13g2_a21oi_1 _4982_ (.A1(_0443_),
    .A2(net89),
    .Y(_1147_),
    .B1(net171));
 sg13g2_nand2_1 _4983_ (.Y(_1148_),
    .A(_1146_),
    .B(_1147_));
 sg13g2_a21oi_1 _4984_ (.A1(_1144_),
    .A2(_1148_),
    .Y(_1149_),
    .B1(net116));
 sg13g2_nor3_1 _4985_ (.A(net66),
    .B(net41),
    .C(_2947_),
    .Y(_1150_));
 sg13g2_a21oi_1 _4986_ (.A1(_2843_),
    .A2(_0478_),
    .Y(_1152_),
    .B1(net66));
 sg13g2_a21oi_1 _4987_ (.A1(_0333_),
    .A2(_0309_),
    .Y(_1153_),
    .B1(_0916_));
 sg13g2_nor4_1 _4988_ (.A(net197),
    .B(_1150_),
    .C(_1152_),
    .D(_1153_),
    .Y(_1154_));
 sg13g2_nand2b_1 _4989_ (.Y(_1155_),
    .B(_1154_),
    .A_N(_1149_));
 sg13g2_nand2_1 _4990_ (.Y(_1156_),
    .A(_0556_),
    .B(net30));
 sg13g2_nand3_1 _4991_ (.B(net67),
    .C(_2221_),
    .A(_1156_),
    .Y(_1157_));
 sg13g2_inv_1 _4992_ (.Y(_1158_),
    .A(net156));
 sg13g2_nor2_1 _4993_ (.A(net106),
    .B(_1158_),
    .Y(_1159_));
 sg13g2_inv_1 _4994_ (.Y(_1160_),
    .A(_1159_));
 sg13g2_a21oi_1 _4995_ (.A1(_1160_),
    .A2(net45),
    .Y(_1161_),
    .B1(net160));
 sg13g2_a21oi_1 _4996_ (.A1(_1157_),
    .A2(_1161_),
    .Y(_1163_),
    .B1(net175));
 sg13g2_nand2_1 _4997_ (.Y(_1164_),
    .A(net34),
    .B(net57));
 sg13g2_nand2_1 _4998_ (.Y(_1165_),
    .A(_1164_),
    .B(net102));
 sg13g2_nand2_1 _4999_ (.Y(_1166_),
    .A(_1165_),
    .B(_1880_));
 sg13g2_inv_2 _5000_ (.Y(_1167_),
    .A(_0651_));
 sg13g2_nand3_1 _5001_ (.B(net121),
    .C(_1167_),
    .A(_1166_),
    .Y(_1168_));
 sg13g2_inv_1 _5002_ (.Y(_1169_),
    .A(_0175_));
 sg13g2_o21ai_1 _5003_ (.B1(net172),
    .Y(_1170_),
    .A1(_0266_),
    .A2(_1169_));
 sg13g2_nand2_1 _5004_ (.Y(_1171_),
    .A(_0099_),
    .B(net58));
 sg13g2_nand3_1 _5005_ (.B(_0825_),
    .C(net78),
    .A(_1171_),
    .Y(_1172_));
 sg13g2_nand3_1 _5006_ (.B(_0748_),
    .C(_1172_),
    .A(_1170_),
    .Y(_1174_));
 sg13g2_nand3_1 _5007_ (.B(_1168_),
    .C(_1174_),
    .A(_1163_),
    .Y(_1175_));
 sg13g2_nand2_1 _5008_ (.Y(_1176_),
    .A(_1155_),
    .B(_1175_));
 sg13g2_nand2_1 _5009_ (.Y(_1177_),
    .A(_1176_),
    .B(net132));
 sg13g2_inv_1 _5010_ (.Y(_1178_),
    .A(_2678_));
 sg13g2_a221oi_1 _5011_ (.B2(_2740_),
    .C1(_0303_),
    .B1(_0901_),
    .A1(_1178_),
    .Y(_1179_),
    .A2(_1104_));
 sg13g2_nor2_1 _5012_ (.A(net163),
    .B(_1179_),
    .Y(_1180_));
 sg13g2_a21oi_1 _5013_ (.A1(_0495_),
    .A2(_0326_),
    .Y(_1181_),
    .B1(_2642_));
 sg13g2_nand2_1 _5014_ (.Y(_1182_),
    .A(_0368_),
    .B(_2747_));
 sg13g2_nand3b_1 _5015_ (.B(net130),
    .C(_1182_),
    .Y(_1183_),
    .A_N(_1181_));
 sg13g2_nand3_1 _5016_ (.B(net74),
    .C(_2651_),
    .A(_2625_),
    .Y(_1185_));
 sg13g2_nand3_1 _5017_ (.B(net117),
    .C(_1185_),
    .A(_1183_),
    .Y(_1186_));
 sg13g2_nor3_1 _5018_ (.A(net171),
    .B(net41),
    .C(_2583_),
    .Y(_1187_));
 sg13g2_nor3_1 _5019_ (.A(net75),
    .B(_0128_),
    .C(_0808_),
    .Y(_1188_));
 sg13g2_a21oi_1 _5020_ (.A1(_0100_),
    .A2(net96),
    .Y(_1189_),
    .B1(net40));
 sg13g2_nor3_1 _5021_ (.A(_1187_),
    .B(_1188_),
    .C(_1189_),
    .Y(_1190_));
 sg13g2_a21oi_1 _5022_ (.A1(_1190_),
    .A2(net80),
    .Y(_1191_),
    .B1(_2646_));
 sg13g2_nand2_1 _5023_ (.Y(_1192_),
    .A(_1186_),
    .B(_1191_));
 sg13g2_a21oi_1 _5024_ (.A1(_1180_),
    .A2(_1192_),
    .Y(_1193_),
    .B1(_2696_));
 sg13g2_nand2_1 _5025_ (.Y(_1194_),
    .A(_1177_),
    .B(_1193_));
 sg13g2_nand2_1 _5026_ (.Y(_0028_),
    .A(_1139_),
    .B(_1194_));
 sg13g2_nand3_1 _5027_ (.B(net93),
    .C(net201),
    .A(_1413_),
    .Y(_1196_));
 sg13g2_buf_2 _5028_ (.A(_1196_),
    .X(_1197_));
 sg13g2_nand2_1 _5029_ (.Y(_1198_),
    .A(_1197_),
    .B(_0388_));
 sg13g2_a21oi_1 _5030_ (.A1(_1198_),
    .A2(net32),
    .Y(_1199_),
    .B1(_1125_));
 sg13g2_nand2_1 _5031_ (.Y(_1200_),
    .A(_0345_),
    .B(_2789_));
 sg13g2_nand2_1 _5032_ (.Y(_1201_),
    .A(_1200_),
    .B(net74));
 sg13g2_a21oi_1 _5033_ (.A1(_1199_),
    .A2(_1201_),
    .Y(_1202_),
    .B1(net147));
 sg13g2_o21ai_1 _5034_ (.B1(net55),
    .Y(_1203_),
    .A1(net33),
    .A2(_1164_));
 sg13g2_nand2_1 _5035_ (.Y(_1204_),
    .A(_2671_),
    .B(_1184_));
 sg13g2_nand2_1 _5036_ (.Y(_1206_),
    .A(_0558_),
    .B(_1204_));
 sg13g2_a21oi_1 _5037_ (.A1(_1206_),
    .A2(_2740_),
    .Y(_1207_),
    .B1(net78));
 sg13g2_nand2_1 _5038_ (.Y(_1208_),
    .A(_1203_),
    .B(_1207_));
 sg13g2_nor3_1 _5039_ (.A(net51),
    .B(_2575_),
    .C(_2848_),
    .Y(_1209_));
 sg13g2_nor3_1 _5040_ (.A(_2550_),
    .B(_0651_),
    .C(_1209_),
    .Y(_1210_));
 sg13g2_nor2_1 _5041_ (.A(net116),
    .B(_1210_),
    .Y(_1211_));
 sg13g2_nand2_1 _5042_ (.Y(_1212_),
    .A(_1208_),
    .B(_1211_));
 sg13g2_a21oi_1 _5043_ (.A1(_1202_),
    .A2(_1212_),
    .Y(_1213_),
    .B1(net195));
 sg13g2_nand2_1 _5044_ (.Y(_1214_),
    .A(_2900_),
    .B(net122));
 sg13g2_nand2_1 _5045_ (.Y(_1215_),
    .A(_0597_),
    .B(_1214_));
 sg13g2_nor2_1 _5046_ (.A(_2751_),
    .B(_1096_),
    .Y(_1217_));
 sg13g2_nand2_1 _5047_ (.Y(_1218_),
    .A(_2779_),
    .B(_1217_));
 sg13g2_nor2_1 _5048_ (.A(_2866_),
    .B(_1218_),
    .Y(_1219_));
 sg13g2_a21oi_1 _5049_ (.A1(_1215_),
    .A2(net39),
    .Y(_1220_),
    .B1(_1219_));
 sg13g2_nand2_1 _5050_ (.Y(_1221_),
    .A(_2529_),
    .B(_0142_));
 sg13g2_a21oi_1 _5051_ (.A1(_1145_),
    .A2(_1221_),
    .Y(_1222_),
    .B1(net199));
 sg13g2_nand2_1 _5052_ (.Y(_1223_),
    .A(_2428_),
    .B(net91));
 sg13g2_nand2_1 _5053_ (.Y(_1224_),
    .A(_1222_),
    .B(_1223_));
 sg13g2_nand2_1 _5054_ (.Y(_1225_),
    .A(_1220_),
    .B(_1224_));
 sg13g2_nand2_1 _5055_ (.Y(_1226_),
    .A(_1225_),
    .B(net121));
 sg13g2_nand2_1 _5056_ (.Y(_1228_),
    .A(_0564_),
    .B(_1083_));
 sg13g2_nor2_1 _5057_ (.A(_0337_),
    .B(_1008_),
    .Y(_1229_));
 sg13g2_o21ai_1 _5058_ (.B1(_2394_),
    .Y(_1230_),
    .A1(_2684_),
    .A2(_2475_));
 sg13g2_a22oi_1 _5059_ (.Y(_1231_),
    .B1(_0917_),
    .B2(_1230_),
    .A2(_1229_),
    .A1(_1228_));
 sg13g2_nand2_1 _5060_ (.Y(_1232_),
    .A(_1226_),
    .B(_1231_));
 sg13g2_nand2_1 _5061_ (.Y(_1233_),
    .A(_1232_),
    .B(net73));
 sg13g2_a21oi_1 _5062_ (.A1(_1213_),
    .A2(_1233_),
    .Y(_1234_),
    .B1(net200));
 sg13g2_a21oi_1 _5063_ (.A1(_2879_),
    .A2(_0387_),
    .Y(_1235_),
    .B1(_0294_));
 sg13g2_nand2_1 _5064_ (.Y(_1236_),
    .A(_2802_),
    .B(net65));
 sg13g2_nand2_1 _5065_ (.Y(_1237_),
    .A(_1135_),
    .B(_1236_));
 sg13g2_a21oi_1 _5066_ (.A1(_0345_),
    .A2(_0655_),
    .Y(_1239_),
    .B1(net31));
 sg13g2_nor3_1 _5067_ (.A(_1235_),
    .B(_1237_),
    .C(_1239_),
    .Y(_1240_));
 sg13g2_nor2_1 _5068_ (.A(net166),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_nand2_1 _5069_ (.Y(_1242_),
    .A(_2428_),
    .B(_0309_));
 sg13g2_nand2_1 _5070_ (.Y(_1243_),
    .A(_3025_),
    .B(_0226_));
 sg13g2_a22oi_1 _5071_ (.Y(_1244_),
    .B1(net53),
    .B2(_1243_),
    .A2(_2991_),
    .A1(_1242_));
 sg13g2_nor2_1 _5072_ (.A(_2162_),
    .B(_1105_),
    .Y(_1245_));
 sg13g2_a21oi_1 _5073_ (.A1(_1245_),
    .A2(_0160_),
    .Y(_1246_),
    .B1(net199));
 sg13g2_nand2_1 _5074_ (.Y(_1247_),
    .A(_2919_),
    .B(_0744_));
 sg13g2_nand2_1 _5075_ (.Y(_1248_),
    .A(_1246_),
    .B(_1247_));
 sg13g2_nand3_1 _5076_ (.B(_1248_),
    .C(net83),
    .A(_1244_),
    .Y(_1250_));
 sg13g2_nand2_1 _5077_ (.Y(_1251_),
    .A(_1241_),
    .B(_1250_));
 sg13g2_a21oi_1 _5078_ (.A1(_2712_),
    .A2(_2637_),
    .Y(_1252_),
    .B1(_0651_));
 sg13g2_inv_1 _5079_ (.Y(_1253_),
    .A(_2659_));
 sg13g2_nor2_1 _5080_ (.A(_2390_),
    .B(_2920_),
    .Y(_1254_));
 sg13g2_a21oi_1 _5081_ (.A1(_1253_),
    .A2(_1045_),
    .Y(_1255_),
    .B1(_1254_));
 sg13g2_nand3b_1 _5082_ (.B(net83),
    .C(_1255_),
    .Y(_1256_),
    .A_N(_1252_));
 sg13g2_a21oi_1 _5083_ (.A1(_2879_),
    .A2(_0387_),
    .Y(_1257_),
    .B1(net31));
 sg13g2_nor2_1 _5084_ (.A(net91),
    .B(_2635_),
    .Y(_1258_));
 sg13g2_a21oi_1 _5085_ (.A1(_1258_),
    .A2(_1238_),
    .Y(_1259_),
    .B1(net78));
 sg13g2_nand2_1 _5086_ (.Y(_1261_),
    .A(_2625_),
    .B(_2539_));
 sg13g2_nand2_1 _5087_ (.Y(_1262_),
    .A(_1259_),
    .B(_1261_));
 sg13g2_nand2_1 _5088_ (.Y(_1263_),
    .A(_0093_),
    .B(_2637_));
 sg13g2_a21oi_1 _5089_ (.A1(_1263_),
    .A2(net74),
    .Y(_1264_),
    .B1(net127));
 sg13g2_nand3b_1 _5090_ (.B(_1262_),
    .C(_1264_),
    .Y(_1265_),
    .A_N(_1257_));
 sg13g2_nand3_1 _5091_ (.B(_1265_),
    .C(net164),
    .A(_1256_),
    .Y(_1266_));
 sg13g2_nand3_1 _5092_ (.B(_1266_),
    .C(_2696_),
    .A(_1251_),
    .Y(_1267_));
 sg13g2_nand2_1 _5093_ (.Y(_1268_),
    .A(_1234_),
    .B(_1267_));
 sg13g2_nand2_1 _5094_ (.Y(_1269_),
    .A(_2997_),
    .B(_2808_));
 sg13g2_o21ai_1 _5095_ (.B1(_2719_),
    .Y(_1270_),
    .A1(net48),
    .A2(_1269_));
 sg13g2_nand2_1 _5096_ (.Y(_1272_),
    .A(_1270_),
    .B(net32));
 sg13g2_nand2_1 _5097_ (.Y(_1273_),
    .A(_2796_),
    .B(_0532_));
 sg13g2_nand2_1 _5098_ (.Y(_1274_),
    .A(_1272_),
    .B(_1273_));
 sg13g2_nand2_1 _5099_ (.Y(_1275_),
    .A(_1274_),
    .B(net80));
 sg13g2_nand2_1 _5100_ (.Y(_1276_),
    .A(_0995_),
    .B(_2539_));
 sg13g2_nand2_1 _5101_ (.Y(_1277_),
    .A(net29),
    .B(net38));
 sg13g2_nand2_1 _5102_ (.Y(_1278_),
    .A(_0721_),
    .B(_1277_));
 sg13g2_nand3_1 _5103_ (.B(_1278_),
    .C(_0520_),
    .A(_1276_),
    .Y(_1279_));
 sg13g2_nand2_1 _5104_ (.Y(_1280_),
    .A(_1279_),
    .B(net175));
 sg13g2_o21ai_1 _5105_ (.B1(_1347_),
    .Y(_1281_),
    .A1(_1159_),
    .A2(_2981_));
 sg13g2_inv_1 _5106_ (.Y(_1283_),
    .A(_1045_));
 sg13g2_nor2_1 _5107_ (.A(_2947_),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_nand2_1 _5108_ (.Y(_1285_),
    .A(_1284_),
    .B(_2682_));
 sg13g2_a21oi_1 _5109_ (.A1(_1281_),
    .A2(_1285_),
    .Y(_1286_),
    .B1(net127));
 sg13g2_nor2_1 _5110_ (.A(_1280_),
    .B(_1286_),
    .Y(_1287_));
 sg13g2_nand2_1 _5111_ (.Y(_1288_),
    .A(_2802_),
    .B(net102));
 sg13g2_nand3_1 _5112_ (.B(net72),
    .C(_3025_),
    .A(_1288_),
    .Y(_1289_));
 sg13g2_o21ai_1 _5113_ (.B1(_2983_),
    .Y(_1290_),
    .A1(_0326_),
    .A2(_0181_));
 sg13g2_nand3_1 _5114_ (.B(_1290_),
    .C(net115),
    .A(_1289_),
    .Y(_1291_));
 sg13g2_nand3_1 _5115_ (.B(_1287_),
    .C(_1291_),
    .A(_1275_),
    .Y(_1292_));
 sg13g2_and3_1 _5116_ (.X(_1294_),
    .A(_2997_),
    .B(_2686_),
    .C(_3014_));
 sg13g2_a21oi_1 _5117_ (.A1(_1206_),
    .A2(_2221_),
    .Y(_1295_),
    .B1(net67));
 sg13g2_nor2_1 _5118_ (.A(_0034_),
    .B(net161),
    .Y(_1296_));
 sg13g2_o21ai_1 _5119_ (.B1(_1296_),
    .Y(_1297_),
    .A1(_1294_),
    .A2(_1295_));
 sg13g2_nor2_1 _5120_ (.A(net76),
    .B(_0926_),
    .Y(_1298_));
 sg13g2_nand2_1 _5121_ (.Y(_1299_),
    .A(_1298_),
    .B(_0150_));
 sg13g2_o21ai_1 _5122_ (.B1(_1299_),
    .Y(_1300_),
    .A1(net67),
    .A2(_2530_));
 sg13g2_nand2_1 _5123_ (.Y(_1301_),
    .A(_1300_),
    .B(net105));
 sg13g2_a22oi_1 _5124_ (.Y(_1302_),
    .B1(_3030_),
    .B2(_0995_),
    .A2(_0609_),
    .A1(_0721_));
 sg13g2_a21oi_1 _5125_ (.A1(_1302_),
    .A2(_2141_),
    .Y(_1303_),
    .B1(net175));
 sg13g2_nand3_1 _5126_ (.B(_1301_),
    .C(_1303_),
    .A(_1297_),
    .Y(_1305_));
 sg13g2_nand2_1 _5127_ (.Y(_1306_),
    .A(_1292_),
    .B(_1305_));
 sg13g2_nand2_1 _5128_ (.Y(_1307_),
    .A(_1306_),
    .B(net165));
 sg13g2_inv_1 _5129_ (.Y(_1308_),
    .A(_2450_));
 sg13g2_nand3_1 _5130_ (.B(_1308_),
    .C(_0453_),
    .A(_1288_),
    .Y(_1309_));
 sg13g2_a21oi_1 _5131_ (.A1(_1197_),
    .A2(_2743_),
    .Y(_1310_),
    .B1(net81));
 sg13g2_nand2_1 _5132_ (.Y(_1311_),
    .A(_1309_),
    .B(_1310_));
 sg13g2_inv_1 _5133_ (.Y(_1312_),
    .A(_0199_));
 sg13g2_nand3b_1 _5134_ (.B(net74),
    .C(_1312_),
    .Y(_1313_),
    .A_N(_1209_));
 sg13g2_nand3_1 _5135_ (.B(net117),
    .C(_1313_),
    .A(_1311_),
    .Y(_1314_));
 sg13g2_nor3_1 _5136_ (.A(net107),
    .B(_0128_),
    .C(_2590_),
    .Y(_1316_));
 sg13g2_o21ai_1 _5137_ (.B1(net161),
    .Y(_1317_),
    .A1(net38),
    .A2(_2461_));
 sg13g2_nand2_2 _5138_ (.Y(_1318_),
    .A(_2582_),
    .B(net143));
 sg13g2_a21oi_1 _5139_ (.A1(_0096_),
    .A2(_1318_),
    .Y(_1319_),
    .B1(net40));
 sg13g2_nor3_1 _5140_ (.A(_1316_),
    .B(_1317_),
    .C(_1319_),
    .Y(_1320_));
 sg13g2_nor2_1 _5141_ (.A(net166),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_nand2_1 _5142_ (.Y(_1322_),
    .A(_1314_),
    .B(_1321_));
 sg13g2_nor2_1 _5143_ (.A(_2739_),
    .B(_0656_),
    .Y(_1323_));
 sg13g2_a21oi_1 _5144_ (.A1(_0124_),
    .A2(net193),
    .Y(_1324_),
    .B1(_2419_));
 sg13g2_nor3_1 _5145_ (.A(_0303_),
    .B(_1323_),
    .C(_1324_),
    .Y(_1325_));
 sg13g2_nor2_1 _5146_ (.A(net195),
    .B(_1325_),
    .Y(_1327_));
 sg13g2_a21oi_1 _5147_ (.A1(_1322_),
    .A2(_1327_),
    .Y(_1328_),
    .B1(net132));
 sg13g2_nand2_1 _5148_ (.Y(_1329_),
    .A(_1307_),
    .B(_1328_));
 sg13g2_nand2_1 _5149_ (.Y(_0029_),
    .A(_1268_),
    .B(_1329_));
 sg13g2_nor2_1 _5150_ (.A(net135),
    .B(_2960_),
    .Y(_1330_));
 sg13g2_a21oi_1 _5151_ (.A1(_2492_),
    .A2(_1330_),
    .Y(_1331_),
    .B1(net124));
 sg13g2_nand2_1 _5152_ (.Y(_1332_),
    .A(_2471_),
    .B(_2509_));
 sg13g2_nand2_1 _5153_ (.Y(_1333_),
    .A(_1331_),
    .B(_1332_));
 sg13g2_nand3_1 _5154_ (.B(net127),
    .C(_1333_),
    .A(_1248_),
    .Y(_1334_));
 sg13g2_o21ai_1 _5155_ (.B1(_2593_),
    .Y(_1335_),
    .A1(_1930_),
    .A2(_0145_));
 sg13g2_nand2_1 _5156_ (.Y(_1337_),
    .A(_0825_),
    .B(_1085_));
 sg13g2_nor2_1 _5157_ (.A(net79),
    .B(_1044_),
    .Y(_1338_));
 sg13g2_nor2_1 _5158_ (.A(_1337_),
    .B(_1338_),
    .Y(_1339_));
 sg13g2_nand3_1 _5159_ (.B(net43),
    .C(_0531_),
    .A(_0181_),
    .Y(_1340_));
 sg13g2_nor2b_1 _5160_ (.A(_1339_),
    .B_N(_1340_),
    .Y(_1341_));
 sg13g2_nand3_1 _5161_ (.B(_1341_),
    .C(_1135_),
    .A(_1335_),
    .Y(_1342_));
 sg13g2_nand2_1 _5162_ (.Y(_1343_),
    .A(_1334_),
    .B(_1342_));
 sg13g2_nand2_1 _5163_ (.Y(_1344_),
    .A(_1343_),
    .B(net147));
 sg13g2_nor2_1 _5164_ (.A(_2437_),
    .B(_1162_),
    .Y(_1345_));
 sg13g2_nor3_1 _5165_ (.A(net76),
    .B(net160),
    .C(_1345_),
    .Y(_1346_));
 sg13g2_a21o_1 _5166_ (.A2(_1346_),
    .A1(_2394_),
    .B1(net175),
    .X(_1348_));
 sg13g2_o21ai_1 _5167_ (.B1(_0250_),
    .Y(_1349_),
    .A1(_2680_),
    .A2(_0332_));
 sg13g2_and2_1 _5168_ (.A(_1349_),
    .B(_0604_),
    .X(_1350_));
 sg13g2_nand2_1 _5169_ (.Y(_1351_),
    .A(_2897_),
    .B(_2680_));
 sg13g2_nand2_1 _5170_ (.Y(_1352_),
    .A(_1489_),
    .B(net137));
 sg13g2_nand3_1 _5171_ (.B(_0600_),
    .C(_1352_),
    .A(_1351_),
    .Y(_1353_));
 sg13g2_inv_1 _5172_ (.Y(_1354_),
    .A(_3005_));
 sg13g2_nand2_1 _5173_ (.Y(_1355_),
    .A(_1354_),
    .B(_3044_));
 sg13g2_nand2_1 _5174_ (.Y(_1356_),
    .A(_1355_),
    .B(_0866_));
 sg13g2_nand2_1 _5175_ (.Y(_1357_),
    .A(_1353_),
    .B(_1356_));
 sg13g2_nor3_1 _5176_ (.A(_1348_),
    .B(_1350_),
    .C(_1357_),
    .Y(_1359_));
 sg13g2_nand2_1 _5177_ (.Y(_1360_),
    .A(_0234_),
    .B(_0167_));
 sg13g2_nand2_1 _5178_ (.Y(_1361_),
    .A(_1008_),
    .B(_1293_));
 sg13g2_nand3_1 _5179_ (.B(_1361_),
    .C(_2544_),
    .A(_1360_),
    .Y(_1362_));
 sg13g2_nand2_1 _5180_ (.Y(_1363_),
    .A(_1318_),
    .B(_0468_));
 sg13g2_a21oi_1 _5181_ (.A1(_1363_),
    .A2(net49),
    .Y(_1364_),
    .B1(_1012_));
 sg13g2_nand2_1 _5182_ (.Y(_1365_),
    .A(_1362_),
    .B(_1364_));
 sg13g2_nand2_1 _5183_ (.Y(_1366_),
    .A(_1365_),
    .B(net116));
 sg13g2_a21oi_1 _5184_ (.A1(_1359_),
    .A2(_1366_),
    .Y(_1367_),
    .B1(_2424_));
 sg13g2_nand2_1 _5185_ (.Y(_1368_),
    .A(_1344_),
    .B(_1367_));
 sg13g2_inv_1 _5186_ (.Y(_1370_),
    .A(_2519_));
 sg13g2_nand3_1 _5187_ (.B(_1370_),
    .C(_0184_),
    .A(_0380_),
    .Y(_1371_));
 sg13g2_nor2_1 _5188_ (.A(net209),
    .B(_2729_),
    .Y(_1372_));
 sg13g2_nor2_1 _5189_ (.A(net75),
    .B(_3005_),
    .Y(_1373_));
 sg13g2_nand2_1 _5190_ (.Y(_1374_),
    .A(net96),
    .B(_1696_));
 sg13g2_o21ai_1 _5191_ (.B1(_0748_),
    .Y(_1375_),
    .A1(_1374_),
    .A2(_2739_));
 sg13g2_a21oi_1 _5192_ (.A1(_2879_),
    .A2(_1373_),
    .Y(_1376_),
    .B1(_1375_));
 sg13g2_a21oi_1 _5193_ (.A1(_1371_),
    .A2(_1372_),
    .Y(_1377_),
    .B1(_1376_));
 sg13g2_o21ai_1 _5194_ (.B1(net69),
    .Y(_1378_),
    .A1(_2739_),
    .A2(_3005_));
 sg13g2_nand3_1 _5195_ (.B(_1013_),
    .C(_1340_),
    .A(_1378_),
    .Y(_1379_));
 sg13g2_nand2_1 _5196_ (.Y(_1381_),
    .A(_1379_),
    .B(_2749_));
 sg13g2_a21oi_1 _5197_ (.A1(_1377_),
    .A2(_1381_),
    .Y(_1382_),
    .B1(_2597_));
 sg13g2_a21oi_1 _5198_ (.A1(_2871_),
    .A2(_2583_),
    .Y(_1383_),
    .B1(net108));
 sg13g2_nand2_1 _5199_ (.Y(_1384_),
    .A(_1383_),
    .B(_2959_));
 sg13g2_nand2_1 _5200_ (.Y(_1385_),
    .A(_3046_),
    .B(_0352_));
 sg13g2_nand3_1 _5201_ (.B(net168),
    .C(_1385_),
    .A(_1384_),
    .Y(_1386_));
 sg13g2_nor2_1 _5202_ (.A(_2508_),
    .B(_0784_),
    .Y(_1387_));
 sg13g2_nand2_1 _5203_ (.Y(_1388_),
    .A(_1387_),
    .B(_1318_));
 sg13g2_nand2_1 _5204_ (.Y(_1389_),
    .A(_0234_),
    .B(_1058_));
 sg13g2_nand3_1 _5205_ (.B(_1389_),
    .C(net75),
    .A(_1388_),
    .Y(_1390_));
 sg13g2_nand3_1 _5206_ (.B(_2664_),
    .C(_1390_),
    .A(_1386_),
    .Y(_1392_));
 sg13g2_nand2_1 _5207_ (.Y(_1393_),
    .A(_1354_),
    .B(_2653_));
 sg13g2_a21oi_1 _5208_ (.A1(_0514_),
    .A2(_2661_),
    .Y(_1394_),
    .B1(net199));
 sg13g2_o21ai_1 _5209_ (.B1(_1394_),
    .Y(_1395_),
    .A1(_0324_),
    .A2(_1393_));
 sg13g2_nand2_1 _5210_ (.Y(_1396_),
    .A(net52),
    .B(_2437_));
 sg13g2_nand2_1 _5211_ (.Y(_1397_),
    .A(_0332_),
    .B(_1336_));
 sg13g2_a21oi_1 _5212_ (.A1(_0808_),
    .A2(_1396_),
    .Y(_1398_),
    .B1(_1397_));
 sg13g2_nor3_1 _5213_ (.A(_3039_),
    .B(_1284_),
    .C(_1398_),
    .Y(_1399_));
 sg13g2_nand2_1 _5214_ (.Y(_1400_),
    .A(_1395_),
    .B(_1399_));
 sg13g2_nand2_1 _5215_ (.Y(_1401_),
    .A(_1392_),
    .B(_1400_));
 sg13g2_nor2_1 _5216_ (.A(_0729_),
    .B(_1401_),
    .Y(_1403_));
 sg13g2_nor2_1 _5217_ (.A(_1382_),
    .B(_1403_),
    .Y(_1404_));
 sg13g2_nand2_1 _5218_ (.Y(_1405_),
    .A(_1368_),
    .B(_1404_));
 sg13g2_nand2_1 _5219_ (.Y(_1406_),
    .A(_1405_),
    .B(net165));
 sg13g2_nand2_1 _5220_ (.Y(_1407_),
    .A(net47),
    .B(net85));
 sg13g2_a21oi_1 _5221_ (.A1(_3019_),
    .A2(_1407_),
    .Y(_1408_),
    .B1(net61));
 sg13g2_o21ai_1 _5222_ (.B1(net88),
    .Y(_1409_),
    .A1(_0276_),
    .A2(_0918_));
 sg13g2_nand2_1 _5223_ (.Y(_1410_),
    .A(_1409_),
    .B(_1124_));
 sg13g2_o21ai_1 _5224_ (.B1(_2373_),
    .Y(_1411_),
    .A1(_1408_),
    .A2(_1410_));
 sg13g2_nand2_1 _5225_ (.Y(_1412_),
    .A(_1411_),
    .B(net170));
 sg13g2_nor2b_1 _5226_ (.A(_0449_),
    .B_N(_0833_),
    .Y(_1414_));
 sg13g2_nand2_1 _5227_ (.Y(_1415_),
    .A(_0791_),
    .B(net133));
 sg13g2_nor2_1 _5228_ (.A(net138),
    .B(_2440_),
    .Y(_1416_));
 sg13g2_nand2_1 _5229_ (.Y(_1417_),
    .A(_1880_),
    .B(net148));
 sg13g2_a22oi_1 _5230_ (.Y(_1418_),
    .B1(_1167_),
    .B2(_1417_),
    .A2(_1416_),
    .A1(_1415_));
 sg13g2_o21ai_1 _5231_ (.B1(_1418_),
    .Y(_1419_),
    .A1(net23),
    .A2(_1414_));
 sg13g2_nand2_1 _5232_ (.Y(_1420_),
    .A(_1419_),
    .B(_2559_));
 sg13g2_nor2b_1 _5233_ (.A(_1412_),
    .B_N(_1420_),
    .Y(_1421_));
 sg13g2_nand3b_1 _5234_ (.B(_2747_),
    .C(_3003_),
    .Y(_1422_),
    .A_N(_0501_));
 sg13g2_a21oi_1 _5235_ (.A1(_1422_),
    .A2(_0915_),
    .Y(_1423_),
    .B1(net121));
 sg13g2_nor2b_1 _5236_ (.A(_2819_),
    .B_N(_3003_),
    .Y(_1425_));
 sg13g2_nand3_1 _5237_ (.B(net67),
    .C(_2727_),
    .A(_1425_),
    .Y(_1426_));
 sg13g2_a21oi_1 _5238_ (.A1(_2605_),
    .A2(net45),
    .Y(_1427_),
    .B1(net162));
 sg13g2_nand2_1 _5239_ (.Y(_1428_),
    .A(_1426_),
    .B(_1427_));
 sg13g2_nand4_1 _5240_ (.B(net67),
    .C(net176),
    .A(_0597_),
    .Y(_1429_),
    .D(net113));
 sg13g2_nand2_1 _5241_ (.Y(_1430_),
    .A(_1429_),
    .B(net175));
 sg13g2_a21oi_1 _5242_ (.A1(_1423_),
    .A2(_1428_),
    .Y(_1431_),
    .B1(_1430_));
 sg13g2_nand2_1 _5243_ (.Y(_1432_),
    .A(_0393_),
    .B(_2900_));
 sg13g2_a22oi_1 _5244_ (.Y(_1433_),
    .B1(_1145_),
    .B2(_1432_),
    .A2(net45),
    .A1(_3036_));
 sg13g2_nand2_1 _5245_ (.Y(_1434_),
    .A(_2571_),
    .B(net87));
 sg13g2_nand3_1 _5246_ (.B(_2993_),
    .C(net32),
    .A(_1434_),
    .Y(_1436_));
 sg13g2_o21ai_1 _5247_ (.B1(_1436_),
    .Y(_1437_),
    .A1(net130),
    .A2(_1433_));
 sg13g2_nand2_1 _5248_ (.Y(_1438_),
    .A(_1437_),
    .B(net117));
 sg13g2_nand2_1 _5249_ (.Y(_1439_),
    .A(_1431_),
    .B(_1438_));
 sg13g2_nand2_1 _5250_ (.Y(_1440_),
    .A(_1421_),
    .B(_1439_));
 sg13g2_o21ai_1 _5251_ (.B1(_2579_),
    .Y(_1441_),
    .A1(net30),
    .A2(_0426_));
 sg13g2_nand2_1 _5252_ (.Y(_1442_),
    .A(_1441_),
    .B(net70));
 sg13g2_nand2_1 _5253_ (.Y(_1443_),
    .A(_1312_),
    .B(_2743_));
 sg13g2_nand2_1 _5254_ (.Y(_1444_),
    .A(net38),
    .B(net126));
 sg13g2_nor2_1 _5255_ (.A(net91),
    .B(_0527_),
    .Y(_1445_));
 sg13g2_o21ai_1 _5256_ (.B1(_1445_),
    .Y(_1447_),
    .A1(net139),
    .A2(_1444_));
 sg13g2_nand3_1 _5257_ (.B(net130),
    .C(_1447_),
    .A(_1443_),
    .Y(_1448_));
 sg13g2_nand3_1 _5258_ (.B(_1448_),
    .C(net131),
    .A(_1442_),
    .Y(_1449_));
 sg13g2_o21ai_1 _5259_ (.B1(_2882_),
    .Y(_1450_),
    .A1(_2889_),
    .A2(_0516_));
 sg13g2_a21oi_1 _5260_ (.A1(net156),
    .A2(_2800_),
    .Y(_1451_),
    .B1(_0948_));
 sg13g2_nor2_1 _5261_ (.A(_1451_),
    .B(_1317_),
    .Y(_1452_));
 sg13g2_nand2_1 _5262_ (.Y(_1453_),
    .A(_1450_),
    .B(_1452_));
 sg13g2_nand3_1 _5263_ (.B(_1453_),
    .C(net73),
    .A(_1449_),
    .Y(_1454_));
 sg13g2_a221oi_1 _5264_ (.B2(_2685_),
    .C1(_2692_),
    .B1(_0302_),
    .A1(net99),
    .Y(_1455_),
    .A2(_0616_));
 sg13g2_nor2_1 _5265_ (.A(net163),
    .B(_1455_),
    .Y(_1456_));
 sg13g2_nand2_1 _5266_ (.Y(_1458_),
    .A(_1454_),
    .B(_1456_));
 sg13g2_nand3_1 _5267_ (.B(_1458_),
    .C(net196),
    .A(_1440_),
    .Y(_1459_));
 sg13g2_nand2_1 _5268_ (.Y(_0017_),
    .A(_1406_),
    .B(_1459_));
 sg13g2_nand3_1 _5269_ (.B(net60),
    .C(_2405_),
    .A(_2765_),
    .Y(_1460_));
 sg13g2_nand3_1 _5270_ (.B(_2413_),
    .C(_2382_),
    .A(_0648_),
    .Y(_1461_));
 sg13g2_nand2_1 _5271_ (.Y(_1462_),
    .A(_1460_),
    .B(_1461_));
 sg13g2_inv_1 _5272_ (.Y(_1463_),
    .A(_2765_));
 sg13g2_nand2_1 _5273_ (.Y(_1464_),
    .A(_1463_),
    .B(_2505_));
 sg13g2_nand2_1 _5274_ (.Y(_1465_),
    .A(_1464_),
    .B(_1071_));
 sg13g2_nor2b_1 _5275_ (.A(_1462_),
    .B_N(_1465_),
    .Y(_1466_));
 sg13g2_nand2b_1 _5276_ (.Y(_1468_),
    .B(_2911_),
    .A_N(_0346_));
 sg13g2_nand2_1 _5277_ (.Y(_1469_),
    .A(_1468_),
    .B(_2895_));
 sg13g2_nand2_1 _5278_ (.Y(_1470_),
    .A(_1466_),
    .B(_1469_));
 sg13g2_nand2_1 _5279_ (.Y(_1471_),
    .A(_1470_),
    .B(net131));
 sg13g2_nand2_1 _5280_ (.Y(_1472_),
    .A(_0808_),
    .B(_2629_));
 sg13g2_nand3_1 _5281_ (.B(net72),
    .C(net148),
    .A(_1197_),
    .Y(_1473_));
 sg13g2_a22oi_1 _5282_ (.Y(_1474_),
    .B1(_1229_),
    .B2(_1473_),
    .A2(_1472_),
    .A1(_0917_));
 sg13g2_nand2_1 _5283_ (.Y(_1475_),
    .A(_1471_),
    .B(_1474_));
 sg13g2_nand2_1 _5284_ (.Y(_1476_),
    .A(_1475_),
    .B(net68));
 sg13g2_a21oi_1 _5285_ (.A1(_0439_),
    .A2(net106),
    .Y(_1477_),
    .B1(net54));
 sg13g2_a21oi_1 _5286_ (.A1(_2879_),
    .A2(_0995_),
    .Y(_1479_),
    .B1(net138));
 sg13g2_nand2_1 _5287_ (.Y(_1480_),
    .A(_3018_),
    .B(_2793_));
 sg13g2_a21oi_1 _5288_ (.A1(_1480_),
    .A2(_1880_),
    .Y(_1481_),
    .B1(_0651_));
 sg13g2_nor3_1 _5289_ (.A(_1477_),
    .B(_1479_),
    .C(_1481_),
    .Y(_1482_));
 sg13g2_nor2_1 _5290_ (.A(net118),
    .B(_1482_),
    .Y(_1483_));
 sg13g2_nand2_1 _5291_ (.Y(_1484_),
    .A(_1480_),
    .B(_1277_));
 sg13g2_a21oi_1 _5292_ (.A1(_1484_),
    .A2(net32),
    .Y(_1485_),
    .B1(_2462_));
 sg13g2_nand2_1 _5293_ (.Y(_1486_),
    .A(_0990_),
    .B(net30));
 sg13g2_nand2_1 _5294_ (.Y(_1487_),
    .A(_1486_),
    .B(_2807_));
 sg13g2_nand2_1 _5295_ (.Y(_1488_),
    .A(_1487_),
    .B(net70));
 sg13g2_a21oi_1 _5296_ (.A1(_1485_),
    .A2(_1488_),
    .Y(_1490_),
    .B1(net63));
 sg13g2_nor2_1 _5297_ (.A(_1483_),
    .B(_1490_),
    .Y(_1491_));
 sg13g2_nand2_1 _5298_ (.Y(_1492_),
    .A(_1476_),
    .B(_1491_));
 sg13g2_nand2_1 _5299_ (.Y(_1493_),
    .A(_1492_),
    .B(net132));
 sg13g2_o21ai_1 _5300_ (.B1(_2552_),
    .Y(_1494_),
    .A1(_2965_),
    .A2(_0621_));
 sg13g2_nand2_1 _5301_ (.Y(_1495_),
    .A(_0239_),
    .B(_0453_));
 sg13g2_nand2_1 _5302_ (.Y(_1496_),
    .A(_0940_),
    .B(_0283_));
 sg13g2_nand3_1 _5303_ (.B(_1496_),
    .C(net172),
    .A(_1495_),
    .Y(_1497_));
 sg13g2_o21ai_1 _5304_ (.B1(_1497_),
    .Y(_1498_),
    .A1(_1050_),
    .A2(_1494_));
 sg13g2_nand2_1 _5305_ (.Y(_1499_),
    .A(_1498_),
    .B(_2957_));
 sg13g2_nor2_1 _5306_ (.A(net37),
    .B(_2430_),
    .Y(_1501_));
 sg13g2_nand3_1 _5307_ (.B(net55),
    .C(_2386_),
    .A(_2444_),
    .Y(_1502_));
 sg13g2_nand3b_1 _5308_ (.B(_1502_),
    .C(_1054_),
    .Y(_1503_),
    .A_N(_1501_));
 sg13g2_a22oi_1 _5309_ (.Y(_1504_),
    .B1(net115),
    .B2(_1503_),
    .A2(_0949_),
    .A1(_2967_));
 sg13g2_nand2_1 _5310_ (.Y(_1505_),
    .A(_1499_),
    .B(_1504_));
 sg13g2_a21oi_1 _5311_ (.A1(_2879_),
    .A2(_2970_),
    .Y(_1506_),
    .B1(net31));
 sg13g2_nand3_1 _5312_ (.B(net200),
    .C(_2691_),
    .A(_1506_),
    .Y(_1507_));
 sg13g2_nand2_1 _5313_ (.Y(_1508_),
    .A(_1507_),
    .B(net196));
 sg13g2_a21oi_1 _5314_ (.A1(_1505_),
    .A2(net112),
    .Y(_1509_),
    .B1(_1508_));
 sg13g2_a21oi_1 _5315_ (.A1(_0542_),
    .A2(_2590_),
    .Y(_1510_),
    .B1(net61));
 sg13g2_nor2_1 _5316_ (.A(net149),
    .B(_2550_),
    .Y(_1512_));
 sg13g2_a21oi_1 _5317_ (.A1(_0405_),
    .A2(_1512_),
    .Y(_1513_),
    .B1(net107));
 sg13g2_nor2_1 _5318_ (.A(net92),
    .B(_0139_),
    .Y(_1514_));
 sg13g2_nor2_1 _5319_ (.A(net89),
    .B(_1514_),
    .Y(_1515_));
 sg13g2_nand2_1 _5320_ (.Y(_1516_),
    .A(_1515_),
    .B(_0277_));
 sg13g2_nand2_1 _5321_ (.Y(_1517_),
    .A(_1513_),
    .B(_1516_));
 sg13g2_a21oi_1 _5322_ (.A1(_0971_),
    .A2(_0404_),
    .Y(_1518_),
    .B1(net167));
 sg13g2_nand3b_1 _5323_ (.B(_1517_),
    .C(_1518_),
    .Y(_1519_),
    .A_N(_1510_));
 sg13g2_nor3_1 _5324_ (.A(net96),
    .B(net28),
    .C(_2436_),
    .Y(_1520_));
 sg13g2_nand2_1 _5325_ (.Y(_1521_),
    .A(_0610_),
    .B(_2405_));
 sg13g2_nand3_1 _5326_ (.B(_0532_),
    .C(net98),
    .A(_2704_),
    .Y(_1523_));
 sg13g2_nand2_1 _5327_ (.Y(_1524_),
    .A(_1521_),
    .B(_1523_));
 sg13g2_nor2_1 _5328_ (.A(_0790_),
    .B(_2440_),
    .Y(_1525_));
 sg13g2_a21o_1 _5329_ (.A2(_0360_),
    .A1(_1525_),
    .B1(net161),
    .X(_1526_));
 sg13g2_nor3_1 _5330_ (.A(_1520_),
    .B(_1524_),
    .C(_1526_),
    .Y(_1527_));
 sg13g2_nand2b_1 _5331_ (.Y(_1528_),
    .B(_3025_),
    .A_N(_1057_));
 sg13g2_nand2_1 _5332_ (.Y(_1529_),
    .A(_1528_),
    .B(_2569_));
 sg13g2_nand2_1 _5333_ (.Y(_1530_),
    .A(_1527_),
    .B(_1529_));
 sg13g2_a21oi_1 _5334_ (.A1(_1519_),
    .A2(_1530_),
    .Y(_1531_),
    .B1(net164));
 sg13g2_nand3_1 _5335_ (.B(_2673_),
    .C(net109),
    .A(_0197_),
    .Y(_1532_));
 sg13g2_a21oi_1 _5336_ (.A1(_1532_),
    .A2(_0239_),
    .Y(_1534_),
    .B1(_0868_));
 sg13g2_nor3_1 _5337_ (.A(net209),
    .B(_0651_),
    .C(_2986_),
    .Y(_1535_));
 sg13g2_nand2_1 _5338_ (.Y(_1536_),
    .A(_0439_),
    .B(net71));
 sg13g2_nor2_1 _5339_ (.A(_1998_),
    .B(_0482_),
    .Y(_1537_));
 sg13g2_nand2_1 _5340_ (.Y(_1538_),
    .A(_1536_),
    .B(_1537_));
 sg13g2_nand2_1 _5341_ (.Y(_1539_),
    .A(_1538_),
    .B(net197));
 sg13g2_a21oi_1 _5342_ (.A1(_1535_),
    .A2(_0838_),
    .Y(_1540_),
    .B1(_1539_));
 sg13g2_nand2b_1 _5343_ (.Y(_1541_),
    .B(_1540_),
    .A_N(_1534_));
 sg13g2_nand2_1 _5344_ (.Y(_1542_),
    .A(_1536_),
    .B(_2482_));
 sg13g2_o21ai_1 _5345_ (.B1(_1542_),
    .Y(_1543_),
    .A1(net41),
    .A2(_2659_));
 sg13g2_nand2_1 _5346_ (.Y(_1545_),
    .A(_1543_),
    .B(net105));
 sg13g2_nor2b_1 _5347_ (.A(_1541_),
    .B_N(_1545_),
    .Y(_1546_));
 sg13g2_a21o_1 _5348_ (.A2(_0140_),
    .A1(_2394_),
    .B1(net28),
    .X(_1547_));
 sg13g2_nand2_1 _5349_ (.Y(_1548_),
    .A(_2671_),
    .B(net97));
 sg13g2_nand2_1 _5350_ (.Y(_1549_),
    .A(_1548_),
    .B(net92));
 sg13g2_nand2_1 _5351_ (.Y(_1550_),
    .A(_1549_),
    .B(_1197_));
 sg13g2_nand2_1 _5352_ (.Y(_1551_),
    .A(_1550_),
    .B(net129));
 sg13g2_o21ai_1 _5353_ (.B1(net110),
    .Y(_1552_),
    .A1(net29),
    .A2(_0148_));
 sg13g2_nand3_1 _5354_ (.B(_1551_),
    .C(_1552_),
    .A(_1547_),
    .Y(_1553_));
 sg13g2_nand2_1 _5355_ (.Y(_1554_),
    .A(_1553_),
    .B(net121));
 sg13g2_nand2_1 _5356_ (.Y(_1556_),
    .A(_1546_),
    .B(_1554_));
 sg13g2_nand2_1 _5357_ (.Y(_1557_),
    .A(_1556_),
    .B(net163));
 sg13g2_nor2_1 _5358_ (.A(_1531_),
    .B(_1557_),
    .Y(_1558_));
 sg13g2_nand2_1 _5359_ (.Y(_1559_),
    .A(_0197_),
    .B(net58));
 sg13g2_nand2_1 _5360_ (.Y(_1560_),
    .A(_0504_),
    .B(_1559_));
 sg13g2_nor2_1 _5361_ (.A(_1269_),
    .B(_1283_),
    .Y(_1561_));
 sg13g2_a21oi_1 _5362_ (.A1(_1560_),
    .A2(_2615_),
    .Y(_1562_),
    .B1(_1561_));
 sg13g2_inv_1 _5363_ (.Y(_1563_),
    .A(_0278_));
 sg13g2_nor2_1 _5364_ (.A(net91),
    .B(_1563_),
    .Y(_1564_));
 sg13g2_a21oi_1 _5365_ (.A1(_2613_),
    .A2(_2728_),
    .Y(_1565_),
    .B1(_2688_));
 sg13g2_nand2_1 _5366_ (.Y(_1567_),
    .A(_1564_),
    .B(_1565_));
 sg13g2_nand2_1 _5367_ (.Y(_1568_),
    .A(_1562_),
    .B(_1567_));
 sg13g2_nand2_1 _5368_ (.Y(_1569_),
    .A(_1568_),
    .B(net131));
 sg13g2_inv_1 _5369_ (.Y(_1570_),
    .A(_2931_));
 sg13g2_nand2_1 _5370_ (.Y(_1571_),
    .A(_2937_),
    .B(net60));
 sg13g2_nand2_1 _5371_ (.Y(_1572_),
    .A(_1570_),
    .B(_1571_));
 sg13g2_nand2_1 _5372_ (.Y(_1573_),
    .A(_1572_),
    .B(_2568_));
 sg13g2_a21oi_1 _5373_ (.A1(net86),
    .A2(_3014_),
    .Y(_1574_),
    .B1(_0477_));
 sg13g2_nand2b_1 _5374_ (.Y(_1575_),
    .B(_2990_),
    .A_N(_1574_));
 sg13g2_nand2_1 _5375_ (.Y(_1576_),
    .A(_1573_),
    .B(_1575_));
 sg13g2_nand2_1 _5376_ (.Y(_1578_),
    .A(_1576_),
    .B(net116));
 sg13g2_nor4_1 _5377_ (.A(net142),
    .B(_0118_),
    .C(_0142_),
    .D(_3013_),
    .Y(_1579_));
 sg13g2_inv_1 _5378_ (.Y(_1580_),
    .A(_0628_));
 sg13g2_nand2_1 _5379_ (.Y(_1581_),
    .A(_0247_),
    .B(_2444_));
 sg13g2_nand2_1 _5380_ (.Y(_1582_),
    .A(net85),
    .B(net125));
 sg13g2_a21oi_1 _5381_ (.A1(_3030_),
    .A2(_1582_),
    .Y(_1583_),
    .B1(net66));
 sg13g2_a22oi_1 _5382_ (.Y(_1584_),
    .B1(_1581_),
    .B2(_1583_),
    .A2(_1580_),
    .A1(_1579_));
 sg13g2_nand3_1 _5383_ (.B(_1578_),
    .C(_1584_),
    .A(_1569_),
    .Y(_1585_));
 sg13g2_nand2_1 _5384_ (.Y(_1586_),
    .A(_1585_),
    .B(net112));
 sg13g2_nand2_1 _5385_ (.Y(_1587_),
    .A(_0225_),
    .B(_2853_));
 sg13g2_inv_1 _5386_ (.Y(_1589_),
    .A(_1587_));
 sg13g2_a21oi_1 _5387_ (.A1(_1589_),
    .A2(_2982_),
    .Y(_1590_),
    .B1(net75));
 sg13g2_nand2_1 _5388_ (.Y(_1591_),
    .A(_1532_),
    .B(_0977_));
 sg13g2_nand2_1 _5389_ (.Y(_1592_),
    .A(_1591_),
    .B(net36));
 sg13g2_nand2_1 _5390_ (.Y(_1593_),
    .A(_1590_),
    .B(_1592_));
 sg13g2_nor2_1 _5391_ (.A(net171),
    .B(_3028_),
    .Y(_1594_));
 sg13g2_nor2_1 _5392_ (.A(_2958_),
    .B(_2742_),
    .Y(_1595_));
 sg13g2_a22oi_1 _5393_ (.Y(_1596_),
    .B1(_1594_),
    .B2(_1595_),
    .A2(_2388_),
    .A1(_0708_));
 sg13g2_nand2_1 _5394_ (.Y(_1597_),
    .A(_1593_),
    .B(_1596_));
 sg13g2_nand2_1 _5395_ (.Y(_1598_),
    .A(_1597_),
    .B(net83));
 sg13g2_nand2_1 _5396_ (.Y(_1600_),
    .A(_0921_),
    .B(_2221_));
 sg13g2_nand2_1 _5397_ (.Y(_1601_),
    .A(_1600_),
    .B(net69));
 sg13g2_nand2_1 _5398_ (.Y(_1602_),
    .A(_1601_),
    .B(_1078_));
 sg13g2_a21oi_1 _5399_ (.A1(_0370_),
    .A2(net65),
    .Y(_1603_),
    .B1(_1602_));
 sg13g2_nor2_1 _5400_ (.A(_2597_),
    .B(_1603_),
    .Y(_1604_));
 sg13g2_a21oi_1 _5401_ (.A1(_1598_),
    .A2(_1604_),
    .Y(_1605_),
    .B1(_2609_));
 sg13g2_nand2_1 _5402_ (.Y(_1606_),
    .A(_1586_),
    .B(_1605_));
 sg13g2_nor2_1 _5403_ (.A(_1558_),
    .B(_1606_),
    .Y(_1607_));
 sg13g2_a21oi_1 _5404_ (.A1(_1493_),
    .A2(_1509_),
    .Y(_0018_),
    .B1(_1607_));
 sg13g2_nand3_1 _5405_ (.B(net120),
    .C(_0618_),
    .A(_0934_),
    .Y(_1608_));
 sg13g2_nand2_1 _5406_ (.Y(_1610_),
    .A(_2453_),
    .B(_2753_));
 sg13g2_nand3_1 _5407_ (.B(_2601_),
    .C(_1610_),
    .A(_1608_),
    .Y(_1611_));
 sg13g2_o21ai_1 _5408_ (.B1(_2733_),
    .Y(_1612_),
    .A1(_0127_),
    .A2(_0603_));
 sg13g2_nand2_1 _5409_ (.Y(_1613_),
    .A(_1611_),
    .B(_1612_));
 sg13g2_nor2_1 _5410_ (.A(net48),
    .B(_0168_),
    .Y(_1614_));
 sg13g2_nand2_1 _5411_ (.Y(_1615_),
    .A(_1614_),
    .B(_0161_));
 sg13g2_nand3_1 _5412_ (.B(_2141_),
    .C(_0478_),
    .A(_1615_),
    .Y(_1616_));
 sg13g2_nand2_1 _5413_ (.Y(_1617_),
    .A(_2861_),
    .B(_0128_));
 sg13g2_o21ai_1 _5414_ (.B1(net105),
    .Y(_1618_),
    .A1(_0219_),
    .A2(_1617_));
 sg13g2_nand3_1 _5415_ (.B(_1618_),
    .C(_2360_),
    .A(_1616_),
    .Y(_1619_));
 sg13g2_a21oi_1 _5416_ (.A1(_1613_),
    .A2(net117),
    .Y(_1621_),
    .B1(_1619_));
 sg13g2_nand3_1 _5417_ (.B(_0673_),
    .C(net168),
    .A(_0863_),
    .Y(_1622_));
 sg13g2_a21oi_1 _5418_ (.A1(_0681_),
    .A2(_1167_),
    .Y(_1623_),
    .B1(_2698_));
 sg13g2_nand2_1 _5419_ (.Y(_1624_),
    .A(_1622_),
    .B(_1623_));
 sg13g2_o21ai_1 _5420_ (.B1(net105),
    .Y(_1625_),
    .A1(_2892_),
    .A2(_0134_));
 sg13g2_o21ai_1 _5421_ (.B1(_2936_),
    .Y(_1626_),
    .A1(_2701_),
    .A2(_2860_));
 sg13g2_nand3_1 _5422_ (.B(_1625_),
    .C(_1626_),
    .A(_1624_),
    .Y(_1627_));
 sg13g2_o21ai_1 _5423_ (.B1(net163),
    .Y(_1628_),
    .A1(_2785_),
    .A2(_1627_));
 sg13g2_nor2_1 _5424_ (.A(_1621_),
    .B(_1628_),
    .Y(_1629_));
 sg13g2_o21ai_1 _5425_ (.B1(_0454_),
    .Y(_1630_),
    .A1(net72),
    .A2(_0681_));
 sg13g2_a21oi_1 _5426_ (.A1(_1563_),
    .A2(_2782_),
    .Y(_1632_),
    .B1(net127));
 sg13g2_a221oi_1 _5427_ (.B2(_2635_),
    .C1(_2619_),
    .B1(_2782_),
    .A1(_2998_),
    .Y(_1633_),
    .A2(net55));
 sg13g2_a21oi_1 _5428_ (.A1(_1630_),
    .A2(_1632_),
    .Y(_1634_),
    .B1(_1633_));
 sg13g2_nand2b_1 _5429_ (.Y(_1635_),
    .B(net112),
    .A_N(_1634_));
 sg13g2_nor2_1 _5430_ (.A(_2701_),
    .B(_1204_),
    .Y(_1636_));
 sg13g2_a21oi_1 _5431_ (.A1(_2727_),
    .A2(_2757_),
    .Y(_1637_),
    .B1(_0110_));
 sg13g2_o21ai_1 _5432_ (.B1(net115),
    .Y(_1638_),
    .A1(_1636_),
    .A2(_1637_));
 sg13g2_nand2_1 _5433_ (.Y(_1639_),
    .A(_1638_),
    .B(_2598_));
 sg13g2_nand3_1 _5434_ (.B(net196),
    .C(_1639_),
    .A(_1635_),
    .Y(_1640_));
 sg13g2_nor2_1 _5435_ (.A(_1629_),
    .B(_1640_),
    .Y(_1641_));
 sg13g2_a21oi_1 _5436_ (.A1(_1006_),
    .A2(_2861_),
    .Y(_1643_),
    .B1(_2510_));
 sg13g2_a21oi_1 _5437_ (.A1(net24),
    .A2(_0599_),
    .Y(_1644_),
    .B1(_1643_));
 sg13g2_nor2_1 _5438_ (.A(_0220_),
    .B(_0219_),
    .Y(_1645_));
 sg13g2_o21ai_1 _5439_ (.B1(net171),
    .Y(_1646_),
    .A1(_2687_),
    .A2(_0616_));
 sg13g2_a21oi_1 _5440_ (.A1(_1645_),
    .A2(_0934_),
    .Y(_1647_),
    .B1(_1646_));
 sg13g2_nand2_1 _5441_ (.Y(_1648_),
    .A(_1253_),
    .B(net193));
 sg13g2_a21oi_1 _5442_ (.A1(_1648_),
    .A2(_2615_),
    .Y(_1649_),
    .B1(_1380_));
 sg13g2_o21ai_1 _5443_ (.B1(_1649_),
    .Y(_1650_),
    .A1(net40),
    .A2(_0628_));
 sg13g2_nor2_1 _5444_ (.A(_1647_),
    .B(_1650_),
    .Y(_1651_));
 sg13g2_a21oi_1 _5445_ (.A1(_1644_),
    .A2(_0511_),
    .Y(_1652_),
    .B1(_1651_));
 sg13g2_a21oi_1 _5446_ (.A1(_0278_),
    .A2(net24),
    .Y(_1654_),
    .B1(_0118_));
 sg13g2_nand2_1 _5447_ (.Y(_1655_),
    .A(_1580_),
    .B(_0721_));
 sg13g2_a21oi_1 _5448_ (.A1(_1654_),
    .A2(_1655_),
    .Y(_1656_),
    .B1(_0729_));
 sg13g2_a21oi_1 _5449_ (.A1(_1652_),
    .A2(_1656_),
    .Y(_1657_),
    .B1(_2609_));
 sg13g2_nand3_1 _5450_ (.B(_0706_),
    .C(_2517_),
    .A(_0654_),
    .Y(_1658_));
 sg13g2_a21oi_1 _5451_ (.A1(_0610_),
    .A2(_1167_),
    .Y(_1659_),
    .B1(net123));
 sg13g2_o21ai_1 _5452_ (.B1(_2626_),
    .Y(_1660_),
    .A1(net194),
    .A2(_0682_));
 sg13g2_nor2_1 _5453_ (.A(_0824_),
    .B(_0611_),
    .Y(_1661_));
 sg13g2_nand2_1 _5454_ (.Y(_1662_),
    .A(_1660_),
    .B(_1661_));
 sg13g2_a22oi_1 _5455_ (.Y(_1663_),
    .B1(_3040_),
    .B2(_1662_),
    .A2(_1659_),
    .A1(_1658_));
 sg13g2_nand2_1 _5456_ (.Y(_1665_),
    .A(_1663_),
    .B(_2360_));
 sg13g2_nor3_1 _5457_ (.A(_2774_),
    .B(_0720_),
    .C(_2723_),
    .Y(_1666_));
 sg13g2_nor2_1 _5458_ (.A(net40),
    .B(_1614_),
    .Y(_1667_));
 sg13g2_nor4_1 _5459_ (.A(_2351_),
    .B(_0033_),
    .C(_1666_),
    .D(_1667_),
    .Y(_1668_));
 sg13g2_a21oi_1 _5460_ (.A1(_0628_),
    .A2(_3022_),
    .Y(_1669_),
    .B1(_1707_));
 sg13g2_o21ai_1 _5461_ (.B1(_1669_),
    .Y(_1670_),
    .A1(_3023_),
    .A2(_0347_));
 sg13g2_a21oi_1 _5462_ (.A1(_1668_),
    .A2(_1670_),
    .Y(_1671_),
    .B1(_2423_));
 sg13g2_nand2_1 _5463_ (.Y(_1672_),
    .A(_1665_),
    .B(_1671_));
 sg13g2_nand2_1 _5464_ (.Y(_1673_),
    .A(_1657_),
    .B(_1672_));
 sg13g2_nor2_1 _5465_ (.A(_2418_),
    .B(_2772_),
    .Y(_1674_));
 sg13g2_a22oi_1 _5466_ (.Y(_1676_),
    .B1(_0622_),
    .B2(_1674_),
    .A2(_2686_),
    .A1(_1253_));
 sg13g2_nor2b_1 _5467_ (.A(_1676_),
    .B_N(_1296_),
    .Y(_1677_));
 sg13g2_nand2_1 _5468_ (.Y(_1678_),
    .A(_2710_),
    .B(_2686_));
 sg13g2_a21oi_1 _5469_ (.A1(_1669_),
    .A2(_1678_),
    .Y(_1679_),
    .B1(_2596_));
 sg13g2_nor3_1 _5470_ (.A(_2826_),
    .B(_3029_),
    .C(_1563_),
    .Y(_1680_));
 sg13g2_o21ai_1 _5471_ (.B1(_0165_),
    .Y(_1681_),
    .A1(_0663_),
    .A2(_1680_));
 sg13g2_o21ai_1 _5472_ (.B1(_1681_),
    .Y(_1682_),
    .A1(_1677_),
    .A2(_1679_));
 sg13g2_nand2_1 _5473_ (.Y(_1683_),
    .A(_1682_),
    .B(_2598_));
 sg13g2_nor2b_1 _5474_ (.A(_1673_),
    .B_N(_1683_),
    .Y(_1684_));
 sg13g2_nor2_1 _5475_ (.A(_1641_),
    .B(_1684_),
    .Y(_0019_));
 sg13g2_inv_1 _5476_ (.Y(_1686_),
    .A(_2715_));
 sg13g2_nor2_1 _5477_ (.A(_1686_),
    .B(_2880_),
    .Y(_1687_));
 sg13g2_nand3b_1 _5478_ (.B(net172),
    .C(_0662_),
    .Y(_1688_),
    .A_N(_1141_));
 sg13g2_nand3_1 _5479_ (.B(net59),
    .C(_1167_),
    .A(_2548_),
    .Y(_1689_));
 sg13g2_o21ai_1 _5480_ (.B1(_1689_),
    .Y(_1690_),
    .A1(_1687_),
    .A2(_1688_));
 sg13g2_nand2_1 _5481_ (.Y(_1691_),
    .A(_1690_),
    .B(net117));
 sg13g2_a21oi_1 _5482_ (.A1(_2513_),
    .A2(_2969_),
    .Y(_1692_),
    .B1(_1039_));
 sg13g2_a21oi_1 _5483_ (.A1(_0816_),
    .A2(_0744_),
    .Y(_1693_),
    .B1(_0338_));
 sg13g2_nor2b_1 _5484_ (.A(_1692_),
    .B_N(_1693_),
    .Y(_1694_));
 sg13g2_nor3_1 _5485_ (.A(net72),
    .B(_2550_),
    .C(_0797_),
    .Y(_1695_));
 sg13g2_nand2_1 _5486_ (.Y(_1697_),
    .A(_0744_),
    .B(_0629_));
 sg13g2_nor3_1 _5487_ (.A(net55),
    .B(_2520_),
    .C(_1697_),
    .Y(_1698_));
 sg13g2_nor3_1 _5488_ (.A(_0163_),
    .B(_1695_),
    .C(_1698_),
    .Y(_1699_));
 sg13g2_nor2_1 _5489_ (.A(_1694_),
    .B(_1699_),
    .Y(_1700_));
 sg13g2_nand3_1 _5490_ (.B(_1700_),
    .C(net68),
    .A(_1691_),
    .Y(_1701_));
 sg13g2_nor2b_1 _5491_ (.A(_2848_),
    .B_N(_1184_),
    .Y(_1702_));
 sg13g2_o21ai_1 _5492_ (.B1(_1542_),
    .Y(_1703_),
    .A1(net41),
    .A2(_1702_));
 sg13g2_nand2_1 _5493_ (.Y(_1704_),
    .A(_1703_),
    .B(net130));
 sg13g2_a21oi_1 _5494_ (.A1(_2273_),
    .A2(_0360_),
    .Y(_1705_),
    .B1(_1012_));
 sg13g2_nand2_1 _5495_ (.Y(_1706_),
    .A(_1704_),
    .B(_1705_));
 sg13g2_nand2_1 _5496_ (.Y(_1708_),
    .A(_1706_),
    .B(_2665_));
 sg13g2_nor2_1 _5497_ (.A(_2826_),
    .B(_1869_),
    .Y(_1709_));
 sg13g2_nor2_1 _5498_ (.A(_2510_),
    .B(_1036_),
    .Y(_1710_));
 sg13g2_a22oi_1 _5499_ (.Y(_1711_),
    .B1(_2879_),
    .B2(_1710_),
    .A2(_1709_),
    .A1(_0093_));
 sg13g2_nor3_1 _5500_ (.A(_2418_),
    .B(net189),
    .C(_3013_),
    .Y(_1712_));
 sg13g2_nor2_1 _5501_ (.A(_1501_),
    .B(_1712_),
    .Y(_1713_));
 sg13g2_nand3_1 _5502_ (.B(_2554_),
    .C(_0422_),
    .A(_0168_),
    .Y(_1714_));
 sg13g2_a21oi_1 _5503_ (.A1(_1713_),
    .A2(_1714_),
    .Y(_1715_),
    .B1(net160));
 sg13g2_a21oi_1 _5504_ (.A1(_1711_),
    .A2(_0521_),
    .Y(_1716_),
    .B1(_1715_));
 sg13g2_nand3_1 _5505_ (.B(_1716_),
    .C(_2736_),
    .A(_1708_),
    .Y(_1717_));
 sg13g2_nand3_1 _5506_ (.B(_1717_),
    .C(_2566_),
    .A(_1701_),
    .Y(_1719_));
 sg13g2_nor2_1 _5507_ (.A(_2774_),
    .B(_2793_),
    .Y(_1720_));
 sg13g2_nand2_1 _5508_ (.Y(_1721_),
    .A(_0422_),
    .B(net119));
 sg13g2_nand3_1 _5509_ (.B(net189),
    .C(net194),
    .A(net76),
    .Y(_1722_));
 sg13g2_a21oi_1 _5510_ (.A1(_1721_),
    .A2(_1722_),
    .Y(_1723_),
    .B1(_2600_));
 sg13g2_a21oi_1 _5511_ (.A1(_1160_),
    .A2(_3003_),
    .Y(_1724_),
    .B1(net138));
 sg13g2_nor4_1 _5512_ (.A(_1561_),
    .B(_1720_),
    .C(_1723_),
    .D(_1724_),
    .Y(_1725_));
 sg13g2_nand2_1 _5513_ (.Y(_1726_),
    .A(_1725_),
    .B(_2957_));
 sg13g2_inv_1 _5514_ (.Y(_1727_),
    .A(_1104_));
 sg13g2_o21ai_1 _5515_ (.B1(_2533_),
    .Y(_1728_),
    .A1(net98),
    .A2(_0942_));
 sg13g2_o21ai_1 _5516_ (.B1(_1728_),
    .Y(_1730_),
    .A1(_1727_),
    .A2(_2931_));
 sg13g2_o21ai_1 _5517_ (.B1(_2593_),
    .Y(_1731_),
    .A1(_0148_),
    .A2(_2574_));
 sg13g2_nor2_1 _5518_ (.A(_2494_),
    .B(net101),
    .Y(_1732_));
 sg13g2_a21oi_1 _5519_ (.A1(_1732_),
    .A2(_2649_),
    .Y(_1733_),
    .B1(net167));
 sg13g2_nand3_1 _5520_ (.B(_1731_),
    .C(_1733_),
    .A(_1730_),
    .Y(_1734_));
 sg13g2_nand3_1 _5521_ (.B(net112),
    .C(_1734_),
    .A(_1726_),
    .Y(_1735_));
 sg13g2_a21oi_1 _5522_ (.A1(_1109_),
    .A2(net65),
    .Y(_1736_),
    .B1(_1077_));
 sg13g2_o21ai_1 _5523_ (.B1(_2935_),
    .Y(_1737_),
    .A1(_2969_),
    .A2(_3029_));
 sg13g2_nand2_1 _5524_ (.Y(_1738_),
    .A(_1736_),
    .B(_1737_));
 sg13g2_nand2_1 _5525_ (.Y(_1739_),
    .A(_1738_),
    .B(_2559_));
 sg13g2_nand2_1 _5526_ (.Y(_1741_),
    .A(_2512_),
    .B(net37));
 sg13g2_o21ai_1 _5527_ (.B1(_1741_),
    .Y(_1742_),
    .A1(_2687_),
    .A2(_2906_));
 sg13g2_nor2_1 _5528_ (.A(_2351_),
    .B(net35),
    .Y(_1743_));
 sg13g2_nand2_1 _5529_ (.Y(_1744_),
    .A(_1742_),
    .B(_1743_));
 sg13g2_nor2_1 _5530_ (.A(_2923_),
    .B(_3029_),
    .Y(_1745_));
 sg13g2_nor3_1 _5531_ (.A(net168),
    .B(_2374_),
    .C(_1745_),
    .Y(_1746_));
 sg13g2_o21ai_1 _5532_ (.B1(_1746_),
    .Y(_1747_),
    .A1(_2642_),
    .A2(_0859_));
 sg13g2_nand3_1 _5533_ (.B(_1744_),
    .C(_1747_),
    .A(_1739_),
    .Y(_1748_));
 sg13g2_nand2_1 _5534_ (.Y(_1749_),
    .A(_1748_),
    .B(_2424_));
 sg13g2_nand2_1 _5535_ (.Y(_1750_),
    .A(_1735_),
    .B(_1749_));
 sg13g2_nor2_1 _5536_ (.A(net196),
    .B(_1750_),
    .Y(_1752_));
 sg13g2_nor2_1 _5537_ (.A(net155),
    .B(_2501_),
    .Y(_1753_));
 sg13g2_o21ai_1 _5538_ (.B1(_1054_),
    .Y(_1754_),
    .A1(_0795_),
    .A2(_0340_));
 sg13g2_a22oi_1 _5539_ (.Y(_1755_),
    .B1(_0165_),
    .B2(_1754_),
    .A2(_0949_),
    .A1(_1753_));
 sg13g2_nand3_1 _5540_ (.B(_1308_),
    .C(_0453_),
    .A(_2823_),
    .Y(_1756_));
 sg13g2_a21oi_1 _5541_ (.A1(_2239_),
    .A2(_2715_),
    .Y(_1757_),
    .B1(net124));
 sg13g2_nand2_1 _5542_ (.Y(_1758_),
    .A(_1756_),
    .B(_1757_));
 sg13g2_nand2_1 _5543_ (.Y(_1759_),
    .A(_1758_),
    .B(_1494_));
 sg13g2_nand2_1 _5544_ (.Y(_1760_),
    .A(_1759_),
    .B(_2596_));
 sg13g2_nand2_1 _5545_ (.Y(_1761_),
    .A(_1755_),
    .B(_1760_));
 sg13g2_nand2_1 _5546_ (.Y(_1763_),
    .A(_1761_),
    .B(_0728_));
 sg13g2_nor2b_1 _5547_ (.A(_1637_),
    .B_N(_0478_),
    .Y(_1764_));
 sg13g2_o21ai_1 _5548_ (.B1(_1764_),
    .Y(_1765_),
    .A1(net99),
    .A2(_0803_));
 sg13g2_a21oi_1 _5549_ (.A1(_1765_),
    .A2(_0959_),
    .Y(_1766_),
    .B1(net195));
 sg13g2_nand2_1 _5550_ (.Y(_1767_),
    .A(_1763_),
    .B(_1766_));
 sg13g2_a21oi_1 _5551_ (.A1(_2803_),
    .A2(_2989_),
    .Y(_1768_),
    .B1(net61));
 sg13g2_nand2_1 _5552_ (.Y(_1769_),
    .A(_0907_),
    .B(net88));
 sg13g2_nor2b_1 _5553_ (.A(_1125_),
    .B_N(_1769_),
    .Y(_1770_));
 sg13g2_nand2b_1 _5554_ (.Y(_1771_),
    .B(_1770_),
    .A_N(_1768_));
 sg13g2_nand2_1 _5555_ (.Y(_1772_),
    .A(_3019_),
    .B(_1370_));
 sg13g2_a21oi_1 _5556_ (.A1(_1772_),
    .A2(_1167_),
    .Y(_1774_),
    .B1(net116));
 sg13g2_nor2_1 _5557_ (.A(net33),
    .B(_1444_),
    .Y(_1775_));
 sg13g2_o21ai_1 _5558_ (.B1(net42),
    .Y(_1776_),
    .A1(_1775_),
    .A2(_2880_));
 sg13g2_nand4_1 _5559_ (.B(net24),
    .C(_2517_),
    .A(_0168_),
    .Y(_1777_),
    .D(net194));
 sg13g2_nand3_1 _5560_ (.B(_1776_),
    .C(_1777_),
    .A(_1774_),
    .Y(_1778_));
 sg13g2_a21oi_1 _5561_ (.A1(_1771_),
    .A2(_1778_),
    .Y(_1779_),
    .B1(net73));
 sg13g2_nor2_1 _5562_ (.A(net31),
    .B(_1197_),
    .Y(_1780_));
 sg13g2_o21ai_1 _5563_ (.B1(_0915_),
    .Y(_1781_),
    .A1(_2892_),
    .A2(_0209_));
 sg13g2_nand2_1 _5564_ (.Y(_1782_),
    .A(_1781_),
    .B(net123));
 sg13g2_a21oi_1 _5565_ (.A1(_0971_),
    .A2(net100),
    .Y(_1783_),
    .B1(net161));
 sg13g2_o21ai_1 _5566_ (.B1(net39),
    .Y(_1785_),
    .A1(_0527_),
    .A2(_2900_));
 sg13g2_nand2_1 _5567_ (.Y(_1786_),
    .A(_1514_),
    .B(net134));
 sg13g2_nand3_1 _5568_ (.B(_1785_),
    .C(_1786_),
    .A(_1783_),
    .Y(_1787_));
 sg13g2_o21ai_1 _5569_ (.B1(_1787_),
    .Y(_1788_),
    .A1(_1780_),
    .A2(_1782_));
 sg13g2_nor3_1 _5570_ (.A(_2678_),
    .B(_0483_),
    .C(_1727_),
    .Y(_1789_));
 sg13g2_nor3_1 _5571_ (.A(net197),
    .B(_1789_),
    .C(_1152_),
    .Y(_1790_));
 sg13g2_nand2_1 _5572_ (.Y(_1791_),
    .A(_1788_),
    .B(_1790_));
 sg13g2_nand2_1 _5573_ (.Y(_1792_),
    .A(_1791_),
    .B(net163));
 sg13g2_nor2_1 _5574_ (.A(_1779_),
    .B(_1792_),
    .Y(_1793_));
 sg13g2_nor2_1 _5575_ (.A(_1767_),
    .B(_1793_),
    .Y(_1794_));
 sg13g2_a21oi_1 _5576_ (.A1(_1719_),
    .A2(_1752_),
    .Y(_0020_),
    .B1(_1794_));
 sg13g2_buf_1 _5577_ (.A(ui_in[0]),
    .X(_1796_));
 sg13g2_buf_2 _5578_ (.A(ui_in[3]),
    .X(_1797_));
 sg13g2_buf_1 _5579_ (.A(_1797_),
    .X(_1798_));
 sg13g2_buf_1 _5580_ (.A(ui_in[2]),
    .X(_1799_));
 sg13g2_buf_1 _5581_ (.A(ui_in[1]),
    .X(_1800_));
 sg13g2_buf_1 _5582_ (.A(_1800_),
    .X(_1801_));
 sg13g2_inv_1 _5583_ (.Y(_1802_),
    .A(net216));
 sg13g2_nor2_1 _5584_ (.A(_1799_),
    .B(_1802_),
    .Y(_1803_));
 sg13g2_nor2_1 _5585_ (.A(net217),
    .B(_1803_),
    .Y(_1804_));
 sg13g2_inv_1 _5586_ (.Y(_1806_),
    .A(net218));
 sg13g2_nand2_1 _5587_ (.Y(_1807_),
    .A(_1806_),
    .B(net216));
 sg13g2_buf_1 _5588_ (.A(_1799_),
    .X(_1808_));
 sg13g2_nand2_1 _5589_ (.Y(_1809_),
    .A(_1807_),
    .B(net215));
 sg13g2_inv_1 _5590_ (.Y(_1810_),
    .A(_1797_));
 sg13g2_nand2_1 _5591_ (.Y(_1811_),
    .A(_1796_),
    .B(_1800_));
 sg13g2_buf_2 _5592_ (.A(_1811_),
    .X(_1812_));
 sg13g2_inv_1 _5593_ (.Y(_1813_),
    .A(_1812_));
 sg13g2_nor2_1 _5594_ (.A(net215),
    .B(_1813_),
    .Y(_1814_));
 sg13g2_nor2_1 _5595_ (.A(net214),
    .B(_1814_),
    .Y(_1815_));
 sg13g2_a22oi_1 _5596_ (.Y(_1817_),
    .B1(_1809_),
    .B2(_1815_),
    .A2(_1804_),
    .A1(net218));
 sg13g2_buf_1 _5597_ (.A(ui_in[4]),
    .X(_1818_));
 sg13g2_nor2_1 _5598_ (.A(_1818_),
    .B(net1),
    .Y(_1819_));
 sg13g2_buf_2 _5599_ (.A(_1819_),
    .X(_1820_));
 sg13g2_inv_1 _5600_ (.Y(_1821_),
    .A(_1820_));
 sg13g2_inv_1 _5601_ (.Y(_1822_),
    .A(net1));
 sg13g2_nor2_1 _5602_ (.A(_1818_),
    .B(_1822_),
    .Y(_1823_));
 sg13g2_buf_2 _5603_ (.A(_1823_),
    .X(_1824_));
 sg13g2_nor2_2 _5604_ (.A(net216),
    .B(net215),
    .Y(_1825_));
 sg13g2_nor2_2 _5605_ (.A(net214),
    .B(_1825_),
    .Y(_1826_));
 sg13g2_inv_1 _5606_ (.Y(_1828_),
    .A(_1799_));
 sg13g2_nor2_1 _5607_ (.A(net216),
    .B(_1828_),
    .Y(_1829_));
 sg13g2_nor2_2 _5608_ (.A(_1797_),
    .B(_1829_),
    .Y(_1830_));
 sg13g2_nor2_1 _5609_ (.A(net218),
    .B(_1799_),
    .Y(_1831_));
 sg13g2_inv_1 _5610_ (.Y(_1832_),
    .A(_1831_));
 sg13g2_o21ai_1 _5611_ (.B1(_1832_),
    .Y(_1833_),
    .A1(_1826_),
    .A2(_1830_));
 sg13g2_inv_1 _5612_ (.Y(_1834_),
    .A(_1818_));
 sg13g2_nor2_1 _5613_ (.A(net1),
    .B(_1834_),
    .Y(_1835_));
 sg13g2_buf_2 _5614_ (.A(_1835_),
    .X(_1836_));
 sg13g2_inv_1 _5615_ (.Y(_1837_),
    .A(_1836_));
 sg13g2_nor2_1 _5616_ (.A(_1831_),
    .B(_1803_),
    .Y(_1839_));
 sg13g2_nand2_1 _5617_ (.Y(_1840_),
    .A(_1796_),
    .B(_1808_));
 sg13g2_nand2_1 _5618_ (.Y(_1841_),
    .A(_1839_),
    .B(_1840_));
 sg13g2_nor2_1 _5619_ (.A(net217),
    .B(_1841_),
    .Y(_1842_));
 sg13g2_nor3_1 _5620_ (.A(_1826_),
    .B(net192),
    .C(_1842_),
    .Y(_1843_));
 sg13g2_a21oi_1 _5621_ (.A1(_1824_),
    .A2(_1833_),
    .Y(_1844_),
    .B1(_1843_));
 sg13g2_o21ai_1 _5622_ (.B1(_1844_),
    .Y(_0000_),
    .A1(_1817_),
    .A2(_1821_));
 sg13g2_nor2_1 _5623_ (.A(net218),
    .B(_1800_),
    .Y(_1845_));
 sg13g2_buf_2 _5624_ (.A(_1845_),
    .X(_1846_));
 sg13g2_nor2_1 _5625_ (.A(_1846_),
    .B(_1813_),
    .Y(_1847_));
 sg13g2_nand2_1 _5626_ (.Y(_1849_),
    .A(_1847_),
    .B(_1832_));
 sg13g2_buf_1 _5627_ (.A(_1828_),
    .X(_1850_));
 sg13g2_nor2_1 _5628_ (.A(_1797_),
    .B(net213),
    .Y(_1851_));
 sg13g2_a21oi_1 _5629_ (.A1(_1846_),
    .A2(net214),
    .Y(_1852_),
    .B1(_1851_));
 sg13g2_inv_1 _5630_ (.Y(_1853_),
    .A(_1852_));
 sg13g2_nand2_1 _5631_ (.Y(_1854_),
    .A(_1853_),
    .B(_1812_));
 sg13g2_o21ai_1 _5632_ (.B1(_1854_),
    .Y(_1855_),
    .A1(net214),
    .A2(_1849_));
 sg13g2_nand2_1 _5633_ (.Y(_1856_),
    .A(_1855_),
    .B(_1836_));
 sg13g2_nand2_1 _5634_ (.Y(_1857_),
    .A(_1839_),
    .B(_1797_));
 sg13g2_nand3_1 _5635_ (.B(_1807_),
    .C(_1824_),
    .A(_1857_),
    .Y(_1858_));
 sg13g2_inv_1 _5636_ (.Y(_1860_),
    .A(_1847_));
 sg13g2_nand2_1 _5637_ (.Y(_1861_),
    .A(_1860_),
    .B(_1850_));
 sg13g2_inv_1 _5638_ (.Y(_1862_),
    .A(_1846_));
 sg13g2_nand2_1 _5639_ (.Y(_1863_),
    .A(_1862_),
    .B(net215));
 sg13g2_a21oi_1 _5640_ (.A1(_1862_),
    .A2(net215),
    .Y(_1864_),
    .B1(net217));
 sg13g2_a21oi_1 _5641_ (.A1(_1861_),
    .A2(_1863_),
    .Y(_1865_),
    .B1(_1864_));
 sg13g2_nand2_1 _5642_ (.Y(_1866_),
    .A(_1865_),
    .B(_1820_));
 sg13g2_nand3_1 _5643_ (.B(_1858_),
    .C(_1866_),
    .A(_1856_),
    .Y(_0007_));
 sg13g2_buf_1 _5644_ (.A(net217),
    .X(_1867_));
 sg13g2_nor2_1 _5645_ (.A(net213),
    .B(_1860_),
    .Y(_1868_));
 sg13g2_nor2_1 _5646_ (.A(net217),
    .B(_1868_),
    .Y(_1870_));
 sg13g2_nand2_1 _5647_ (.Y(_1871_),
    .A(_1807_),
    .B(net213));
 sg13g2_nand2_1 _5648_ (.Y(_1872_),
    .A(net217),
    .B(net218));
 sg13g2_inv_1 _5649_ (.Y(_1873_),
    .A(_1872_));
 sg13g2_a221oi_1 _5650_ (.B2(_1871_),
    .C1(_1873_),
    .B1(_1870_),
    .A1(net212),
    .Y(_1874_),
    .A2(_1825_));
 sg13g2_nor2_1 _5651_ (.A(net216),
    .B(_1806_),
    .Y(_1875_));
 sg13g2_nor2_1 _5652_ (.A(net213),
    .B(_1875_),
    .Y(_1876_));
 sg13g2_nor2_1 _5653_ (.A(net215),
    .B(_1807_),
    .Y(_1877_));
 sg13g2_inv_1 _5654_ (.Y(_1878_),
    .A(_1877_));
 sg13g2_nand2_1 _5655_ (.Y(_1879_),
    .A(_1878_),
    .B(net212));
 sg13g2_nor2_1 _5656_ (.A(net215),
    .B(_1806_),
    .Y(_1881_));
 sg13g2_inv_1 _5657_ (.Y(_1882_),
    .A(_1830_));
 sg13g2_o21ai_1 _5658_ (.B1(_1824_),
    .Y(_1883_),
    .A1(_1881_),
    .A2(_1882_));
 sg13g2_o21ai_1 _5659_ (.B1(_1883_),
    .Y(_1884_),
    .A1(_1821_),
    .A2(_1853_));
 sg13g2_a22oi_1 _5660_ (.Y(_1885_),
    .B1(_1879_),
    .B2(_1884_),
    .A2(_1876_),
    .A1(_1820_));
 sg13g2_o21ai_1 _5661_ (.B1(_1885_),
    .Y(_0008_),
    .A1(net192),
    .A2(_1874_));
 sg13g2_nor2_1 _5662_ (.A(net213),
    .B(_1813_),
    .Y(_1886_));
 sg13g2_a21oi_1 _5663_ (.A1(_1860_),
    .A2(net213),
    .Y(_1887_),
    .B1(_1886_));
 sg13g2_inv_1 _5664_ (.Y(_1888_),
    .A(_1814_));
 sg13g2_nand2_1 _5665_ (.Y(_1889_),
    .A(_1801_),
    .B(_1808_));
 sg13g2_nand3_1 _5666_ (.B(_1889_),
    .C(_1824_),
    .A(_1888_),
    .Y(_1891_));
 sg13g2_o21ai_1 _5667_ (.B1(_1891_),
    .Y(_1892_),
    .A1(net192),
    .A2(_1887_));
 sg13g2_nand2_1 _5668_ (.Y(_1893_),
    .A(_1892_),
    .B(_1810_));
 sg13g2_nor2_2 _5669_ (.A(net214),
    .B(_1846_),
    .Y(_1894_));
 sg13g2_inv_1 _5670_ (.Y(_1895_),
    .A(_1824_));
 sg13g2_a21oi_1 _5671_ (.A1(_1895_),
    .A2(net192),
    .Y(_1896_),
    .B1(_1888_));
 sg13g2_nor2b_1 _5672_ (.A(_1881_),
    .B_N(_1889_),
    .Y(_1897_));
 sg13g2_inv_1 _5673_ (.Y(_1898_),
    .A(_1886_));
 sg13g2_a22oi_1 _5674_ (.Y(_1899_),
    .B1(_1804_),
    .B2(_1898_),
    .A2(_1867_),
    .A1(_1897_));
 sg13g2_a22oi_1 _5675_ (.Y(_1900_),
    .B1(_1820_),
    .B2(_1899_),
    .A2(_1896_),
    .A1(_1894_));
 sg13g2_nand2_1 _5676_ (.Y(_0009_),
    .A(_1893_),
    .B(_1900_));
 sg13g2_nor2_1 _5677_ (.A(net213),
    .B(_1812_),
    .Y(_1902_));
 sg13g2_inv_1 _5678_ (.Y(_1903_),
    .A(_1902_));
 sg13g2_a22oi_1 _5679_ (.Y(_1904_),
    .B1(_1830_),
    .B2(_1878_),
    .A2(net212),
    .A1(_1903_));
 sg13g2_nor2_1 _5680_ (.A(_1875_),
    .B(_1882_),
    .Y(_1905_));
 sg13g2_nand2_1 _5681_ (.Y(_1906_),
    .A(_1894_),
    .B(_1812_));
 sg13g2_nand2_1 _5682_ (.Y(_1907_),
    .A(_1797_),
    .B(_1799_));
 sg13g2_nand2_1 _5683_ (.Y(_1908_),
    .A(_1824_),
    .B(_1907_));
 sg13g2_inv_1 _5684_ (.Y(_1909_),
    .A(_1908_));
 sg13g2_nand2_1 _5685_ (.Y(_1910_),
    .A(_1906_),
    .B(_1909_));
 sg13g2_nor2_1 _5686_ (.A(_1905_),
    .B(_1910_),
    .Y(_1912_));
 sg13g2_nand3b_1 _5687_ (.B(net214),
    .C(net218),
    .Y(_1913_),
    .A_N(_1825_));
 sg13g2_a21oi_1 _5688_ (.A1(_1913_),
    .A2(_1906_),
    .Y(_1914_),
    .B1(_1821_));
 sg13g2_nor2_1 _5689_ (.A(_1912_),
    .B(_1914_),
    .Y(_1915_));
 sg13g2_o21ai_1 _5690_ (.B1(_1915_),
    .Y(_0010_),
    .A1(net192),
    .A2(_1904_));
 sg13g2_nand2_1 _5691_ (.Y(_1916_),
    .A(_1870_),
    .B(_1839_));
 sg13g2_nand3_1 _5692_ (.B(_1836_),
    .C(_1872_),
    .A(_1916_),
    .Y(_1917_));
 sg13g2_nor2_1 _5693_ (.A(_1821_),
    .B(_1830_),
    .Y(_1918_));
 sg13g2_nand2_1 _5694_ (.Y(_1919_),
    .A(_1826_),
    .B(_1812_));
 sg13g2_nor2_1 _5695_ (.A(_1894_),
    .B(_1908_),
    .Y(_1920_));
 sg13g2_a22oi_1 _5696_ (.Y(_1922_),
    .B1(_1849_),
    .B2(_1920_),
    .A2(_1919_),
    .A1(_1918_));
 sg13g2_nand2_1 _5697_ (.Y(_0011_),
    .A(_1917_),
    .B(_1922_));
 sg13g2_nand3_1 _5698_ (.B(_1818_),
    .C(_1906_),
    .A(_1854_),
    .Y(_1923_));
 sg13g2_nor2_1 _5699_ (.A(net216),
    .B(_1810_),
    .Y(_1924_));
 sg13g2_nand3b_1 _5700_ (.B(_1834_),
    .C(_1889_),
    .Y(_1925_),
    .A_N(_1924_));
 sg13g2_nand3_1 _5701_ (.B(_1822_),
    .C(_1925_),
    .A(_1923_),
    .Y(_1926_));
 sg13g2_o21ai_1 _5702_ (.B1(_1920_),
    .Y(_1927_),
    .A1(_1876_),
    .A2(_1852_));
 sg13g2_nand2_1 _5703_ (.Y(_0012_),
    .A(_1926_),
    .B(_1927_));
 sg13g2_nor3_1 _5704_ (.A(net212),
    .B(_1846_),
    .C(_1902_),
    .Y(_1928_));
 sg13g2_o21ai_1 _5705_ (.B1(_1836_),
    .Y(_1929_),
    .A1(_1902_),
    .A2(_1814_));
 sg13g2_a21oi_1 _5706_ (.A1(_1846_),
    .A2(_1867_),
    .Y(_1931_),
    .B1(_1895_));
 sg13g2_a22oi_1 _5707_ (.Y(_1932_),
    .B1(_1863_),
    .B2(_1931_),
    .A2(_1820_),
    .A1(_1826_));
 sg13g2_o21ai_1 _5708_ (.B1(_1932_),
    .Y(_0013_),
    .A1(_1928_),
    .A2(_1929_));
 sg13g2_inv_1 _5709_ (.Y(_1933_),
    .A(_1815_));
 sg13g2_nand3_1 _5710_ (.B(net214),
    .C(net213),
    .A(_1846_),
    .Y(_1934_));
 sg13g2_nand3_1 _5711_ (.B(_1836_),
    .C(_1934_),
    .A(_1933_),
    .Y(_1935_));
 sg13g2_o21ai_1 _5712_ (.B1(_1935_),
    .Y(_0014_),
    .A1(_1864_),
    .A2(_1908_));
 sg13g2_o21ai_1 _5713_ (.B1(_1908_),
    .Y(_0015_),
    .A1(net192),
    .A2(_1933_));
 sg13g2_nor2_1 _5714_ (.A(_1798_),
    .B(_1902_),
    .Y(_1936_));
 sg13g2_inv_1 _5715_ (.Y(_1937_),
    .A(_1857_));
 sg13g2_a22oi_1 _5716_ (.Y(_1939_),
    .B1(_1898_),
    .B2(_1937_),
    .A2(_1878_),
    .A1(_1936_));
 sg13g2_nor2_1 _5717_ (.A(net218),
    .B(_1850_),
    .Y(_1940_));
 sg13g2_o21ai_1 _5718_ (.B1(_1909_),
    .Y(_1941_),
    .A1(_1940_),
    .A2(_1924_));
 sg13g2_xor2_1 _5719_ (.B(net216),
    .A(_1798_),
    .X(_1942_));
 sg13g2_nand3_1 _5720_ (.B(_1942_),
    .C(_1822_),
    .A(_1863_),
    .Y(_1943_));
 sg13g2_nand3_1 _5721_ (.B(_1943_),
    .C(net192),
    .A(_1941_),
    .Y(_1944_));
 sg13g2_o21ai_1 _5722_ (.B1(_1944_),
    .Y(_0001_),
    .A1(net192),
    .A2(_1939_));
 sg13g2_inv_1 _5723_ (.Y(_1945_),
    .A(_1803_));
 sg13g2_nand2_1 _5724_ (.Y(_1946_),
    .A(_1945_),
    .B(net218));
 sg13g2_a21oi_1 _5725_ (.A1(_1946_),
    .A2(_1830_),
    .Y(_1947_),
    .B1(_1873_));
 sg13g2_a21oi_1 _5726_ (.A1(_1809_),
    .A2(_1945_),
    .Y(_1949_),
    .B1(net212));
 sg13g2_a21oi_1 _5727_ (.A1(_1894_),
    .A2(_1889_),
    .Y(_1950_),
    .B1(_1837_));
 sg13g2_o21ai_1 _5728_ (.B1(_1950_),
    .Y(_1951_),
    .A1(net212),
    .A2(_1868_));
 sg13g2_o21ai_1 _5729_ (.B1(_1951_),
    .Y(_1952_),
    .A1(_1910_),
    .A2(_1949_));
 sg13g2_a21oi_1 _5730_ (.A1(_1820_),
    .A2(_1947_),
    .Y(_0002_),
    .B1(_1952_));
 sg13g2_nor2_1 _5731_ (.A(net217),
    .B(_1840_),
    .Y(_1953_));
 sg13g2_nor2_1 _5732_ (.A(_1857_),
    .B(_1868_),
    .Y(_1954_));
 sg13g2_o21ai_1 _5733_ (.B1(_1836_),
    .Y(_1955_),
    .A1(_1953_),
    .A2(_1954_));
 sg13g2_nor2_1 _5734_ (.A(_1853_),
    .B(_1937_),
    .Y(_1956_));
 sg13g2_o21ai_1 _5735_ (.B1(_1820_),
    .Y(_1957_),
    .A1(_1940_),
    .A2(_1956_));
 sg13g2_o21ai_1 _5736_ (.B1(_1920_),
    .Y(_1959_),
    .A1(_1813_),
    .A2(_1882_));
 sg13g2_nand3_1 _5737_ (.B(_1957_),
    .C(_1959_),
    .A(_1955_),
    .Y(_0003_));
 sg13g2_nand2b_1 _5738_ (.Y(_1960_),
    .B(_1870_),
    .A_N(_1825_));
 sg13g2_nand3_1 _5739_ (.B(_1834_),
    .C(_1857_),
    .A(_1960_),
    .Y(_1961_));
 sg13g2_a21oi_1 _5740_ (.A1(_1841_),
    .A2(net217),
    .Y(_1962_),
    .B1(_1851_));
 sg13g2_a21oi_1 _5741_ (.A1(_1962_),
    .A2(_1818_),
    .Y(_1963_),
    .B1(net1));
 sg13g2_nand2_1 _5742_ (.Y(_1964_),
    .A(_1961_),
    .B(_1963_));
 sg13g2_nand2_1 _5743_ (.Y(_1965_),
    .A(_1853_),
    .B(_1809_));
 sg13g2_o21ai_1 _5744_ (.B1(net212),
    .Y(_1966_),
    .A1(net215),
    .A2(_1812_));
 sg13g2_nand3_1 _5745_ (.B(_1824_),
    .C(_1966_),
    .A(_1965_),
    .Y(_1967_));
 sg13g2_nand2_1 _5746_ (.Y(_0004_),
    .A(_1964_),
    .B(_1967_));
 sg13g2_o21ai_1 _5747_ (.B1(net214),
    .Y(_1969_),
    .A1(net216),
    .A2(_1840_));
 sg13g2_nor2b_1 _5748_ (.A(_1894_),
    .B_N(_1969_),
    .Y(_1970_));
 sg13g2_nor2_1 _5749_ (.A(_1801_),
    .B(_1881_),
    .Y(_1971_));
 sg13g2_nand2_1 _5750_ (.Y(_1972_),
    .A(_1820_),
    .B(_1907_));
 sg13g2_inv_1 _5751_ (.Y(_1973_),
    .A(_1972_));
 sg13g2_a22oi_1 _5752_ (.Y(_1974_),
    .B1(_1973_),
    .B2(_1969_),
    .A2(_1971_),
    .A1(_1909_));
 sg13g2_o21ai_1 _5753_ (.B1(_1974_),
    .Y(_0005_),
    .A1(_1837_),
    .A2(_1970_));
 sg13g2_nand3_1 _5754_ (.B(_1846_),
    .C(net212),
    .A(_1836_),
    .Y(_1975_));
 sg13g2_o21ai_1 _5755_ (.B1(_1975_),
    .Y(_0006_),
    .A1(_1895_),
    .A2(_1965_));
 sg13g2_nand2_1 _5756_ (.Y(_1977_),
    .A(_2239_),
    .B(net120));
 sg13g2_nand2_1 _5757_ (.Y(_1978_),
    .A(_3031_),
    .B(_1977_));
 sg13g2_a21oi_1 _5758_ (.A1(_1978_),
    .A2(_0234_),
    .Y(_1979_),
    .B1(net66));
 sg13g2_nand2_1 _5759_ (.Y(_1980_),
    .A(_0359_),
    .B(_0422_));
 sg13g2_o21ai_1 _5760_ (.B1(_1980_),
    .Y(_1981_),
    .A1(_0110_),
    .A2(_2961_));
 sg13g2_nand2_1 _5761_ (.Y(_1982_),
    .A(_1981_),
    .B(net105));
 sg13g2_nor3_1 _5762_ (.A(net203),
    .B(net64),
    .C(_2550_),
    .Y(_1983_));
 sg13g2_nand2_1 _5763_ (.Y(_1984_),
    .A(_2890_),
    .B(_1983_));
 sg13g2_nand2_1 _5764_ (.Y(_1985_),
    .A(_0333_),
    .B(_3026_));
 sg13g2_nand2_1 _5765_ (.Y(_1986_),
    .A(_1985_),
    .B(_0600_));
 sg13g2_nand3_1 _5766_ (.B(_1984_),
    .C(_1986_),
    .A(_1982_),
    .Y(_1988_));
 sg13g2_nor2_1 _5767_ (.A(_1979_),
    .B(_1988_),
    .Y(_1989_));
 sg13g2_nand2_1 _5768_ (.Y(_1990_),
    .A(_0100_),
    .B(_0921_));
 sg13g2_nor2b_1 _5769_ (.A(_1159_),
    .B_N(_2605_),
    .Y(_1991_));
 sg13g2_nand2_1 _5770_ (.Y(_1992_),
    .A(net86),
    .B(net125));
 sg13g2_nand2_1 _5771_ (.Y(_1993_),
    .A(_1991_),
    .B(_1992_));
 sg13g2_a22oi_1 _5772_ (.Y(_1994_),
    .B1(net25),
    .B2(_1993_),
    .A2(net32),
    .A1(_1990_));
 sg13g2_o21ai_1 _5773_ (.B1(_0542_),
    .Y(_1995_),
    .A1(_2758_),
    .A2(net59));
 sg13g2_nand2_1 _5774_ (.Y(_1996_),
    .A(_1995_),
    .B(net26));
 sg13g2_nand2_1 _5775_ (.Y(_1997_),
    .A(_1994_),
    .B(_1996_));
 sg13g2_nand2_1 _5776_ (.Y(_1999_),
    .A(_1997_),
    .B(net117));
 sg13g2_a21oi_1 _5777_ (.A1(_1989_),
    .A2(_1999_),
    .Y(_2000_),
    .B1(_0729_));
 sg13g2_nand3b_1 _5778_ (.B(_1446_),
    .C(net90),
    .Y(_2001_),
    .A_N(_2461_));
 sg13g2_nand3_1 _5779_ (.B(net141),
    .C(net49),
    .A(_0224_),
    .Y(_2002_));
 sg13g2_nand3_1 _5780_ (.B(_2002_),
    .C(net169),
    .A(_2001_),
    .Y(_2003_));
 sg13g2_a22oi_1 _5781_ (.Y(_2004_),
    .B1(net79),
    .B2(net141),
    .A2(net119),
    .A1(net153));
 sg13g2_o21ai_1 _5782_ (.B1(_2004_),
    .Y(_2005_),
    .A1(net102),
    .A2(net34));
 sg13g2_nand2_1 _5783_ (.Y(_2006_),
    .A(_2005_),
    .B(net129));
 sg13g2_nor2b_1 _5784_ (.A(_2003_),
    .B_N(_2006_),
    .Y(_2007_));
 sg13g2_nand2b_1 _5785_ (.Y(_2008_),
    .B(_0182_),
    .A_N(_1697_));
 sg13g2_nand2_1 _5786_ (.Y(_2010_),
    .A(_1463_),
    .B(_2585_));
 sg13g2_nand2_1 _5787_ (.Y(_2011_),
    .A(_2010_),
    .B(_2910_));
 sg13g2_nor2_1 _5788_ (.A(net23),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_a21oi_1 _5789_ (.A1(_2008_),
    .A2(net25),
    .Y(_2013_),
    .B1(_2012_));
 sg13g2_nand2_1 _5790_ (.Y(_2014_),
    .A(_2007_),
    .B(_2013_));
 sg13g2_a21oi_1 _5791_ (.A1(_2403_),
    .A2(_1160_),
    .Y(_2015_),
    .B1(net40));
 sg13g2_nor2_1 _5792_ (.A(net62),
    .B(_2900_),
    .Y(_2016_));
 sg13g2_a21oi_1 _5793_ (.A1(_2016_),
    .A2(_2933_),
    .Y(_2017_),
    .B1(net203));
 sg13g2_nor2b_1 _5794_ (.A(_2015_),
    .B_N(_2017_),
    .Y(_2018_));
 sg13g2_nand3_1 _5795_ (.B(net102),
    .C(net38),
    .A(net57),
    .Y(_2019_));
 sg13g2_nand2_1 _5796_ (.Y(_2021_),
    .A(_2019_),
    .B(_2514_));
 sg13g2_nand2_1 _5797_ (.Y(_2022_),
    .A(_2021_),
    .B(net25));
 sg13g2_o21ai_1 _5798_ (.B1(_2402_),
    .Y(_2023_),
    .A1(_1478_),
    .A2(_2501_));
 sg13g2_nand2_1 _5799_ (.Y(_2024_),
    .A(_2023_),
    .B(_2845_));
 sg13g2_nand2_1 _5800_ (.Y(_2025_),
    .A(_2024_),
    .B(net53));
 sg13g2_nand3_1 _5801_ (.B(_2022_),
    .C(_2025_),
    .A(_2018_),
    .Y(_2026_));
 sg13g2_nand3_1 _5802_ (.B(_2026_),
    .C(_2598_),
    .A(_2014_),
    .Y(_2027_));
 sg13g2_nand2_1 _5803_ (.Y(_2028_),
    .A(_2027_),
    .B(net195));
 sg13g2_nor2_1 _5804_ (.A(_2000_),
    .B(_2028_),
    .Y(_2029_));
 sg13g2_nand3_1 _5805_ (.B(_1197_),
    .C(net69),
    .A(_0704_),
    .Y(_2030_));
 sg13g2_nand2_1 _5806_ (.Y(_2032_),
    .A(_2030_),
    .B(_2556_));
 sg13g2_nand3_1 _5807_ (.B(_0782_),
    .C(_2526_),
    .A(_3048_),
    .Y(_2033_));
 sg13g2_nand2_1 _5808_ (.Y(_2034_),
    .A(_2033_),
    .B(net129));
 sg13g2_nand2_1 _5809_ (.Y(_2035_),
    .A(_2766_),
    .B(_1653_));
 sg13g2_nand2_1 _5810_ (.Y(_2036_),
    .A(_2035_),
    .B(net39));
 sg13g2_nand2_1 _5811_ (.Y(_2037_),
    .A(_2034_),
    .B(_2036_));
 sg13g2_nor2_1 _5812_ (.A(_2032_),
    .B(_2037_),
    .Y(_2038_));
 sg13g2_nor2_1 _5813_ (.A(net118),
    .B(_2038_),
    .Y(_2039_));
 sg13g2_a21oi_1 _5814_ (.A1(_2893_),
    .A2(_0100_),
    .Y(_2040_),
    .B1(net23));
 sg13g2_a21oi_1 _5815_ (.A1(_1425_),
    .A2(_2541_),
    .Y(_2041_),
    .B1(net31));
 sg13g2_nand2_1 _5816_ (.Y(_2043_),
    .A(_0234_),
    .B(_2961_));
 sg13g2_nand2_1 _5817_ (.Y(_2044_),
    .A(_2043_),
    .B(net110));
 sg13g2_nand2_1 _5818_ (.Y(_2045_),
    .A(_1114_),
    .B(_0617_));
 sg13g2_nand2_1 _5819_ (.Y(_2046_),
    .A(_2045_),
    .B(net134));
 sg13g2_nand2_1 _5820_ (.Y(_2047_),
    .A(_2044_),
    .B(_2046_));
 sg13g2_nor3_1 _5821_ (.A(_2040_),
    .B(_2041_),
    .C(_2047_),
    .Y(_2048_));
 sg13g2_nor2_1 _5822_ (.A(net63),
    .B(_2048_),
    .Y(_2049_));
 sg13g2_nor2_1 _5823_ (.A(_2039_),
    .B(_2049_),
    .Y(_2050_));
 sg13g2_nand3_1 _5824_ (.B(_3048_),
    .C(_2526_),
    .A(_0622_),
    .Y(_2051_));
 sg13g2_nand2_1 _5825_ (.Y(_2052_),
    .A(_2051_),
    .B(net129));
 sg13g2_nand2_1 _5826_ (.Y(_2054_),
    .A(_0318_),
    .B(_2617_));
 sg13g2_nand2_1 _5827_ (.Y(_2055_),
    .A(_2054_),
    .B(net39));
 sg13g2_nand2_1 _5828_ (.Y(_2056_),
    .A(_2052_),
    .B(_2055_));
 sg13g2_nor2_1 _5829_ (.A(net64),
    .B(_1169_),
    .Y(_2057_));
 sg13g2_nand2_1 _5830_ (.Y(_2058_),
    .A(_2057_),
    .B(_2797_));
 sg13g2_nor2_1 _5831_ (.A(net62),
    .B(_0346_),
    .Y(_2059_));
 sg13g2_nand2_1 _5832_ (.Y(_2060_),
    .A(_2834_),
    .B(net77));
 sg13g2_nand2_1 _5833_ (.Y(_2061_),
    .A(_2059_),
    .B(_2060_));
 sg13g2_nand3_1 _5834_ (.B(_2061_),
    .C(net167),
    .A(_2058_),
    .Y(_2062_));
 sg13g2_nor2_1 _5835_ (.A(_2056_),
    .B(_2062_),
    .Y(_2063_));
 sg13g2_nor2_1 _5836_ (.A(net166),
    .B(_2063_),
    .Y(_2065_));
 sg13g2_nand2_1 _5837_ (.Y(_2066_),
    .A(_2614_),
    .B(net84));
 sg13g2_nand2_1 _5838_ (.Y(_2067_),
    .A(_2674_),
    .B(_2992_));
 sg13g2_a21oi_1 _5839_ (.A1(_0958_),
    .A2(_2067_),
    .Y(_2068_),
    .B1(net81));
 sg13g2_o21ai_1 _5840_ (.B1(_2068_),
    .Y(_2069_),
    .A1(_2756_),
    .A2(_2066_));
 sg13g2_nand2_1 _5841_ (.Y(_2070_),
    .A(_0556_),
    .B(net92));
 sg13g2_nor2_1 _5842_ (.A(net151),
    .B(_2745_),
    .Y(_2071_));
 sg13g2_nand2_1 _5843_ (.Y(_2072_),
    .A(_2070_),
    .B(_2071_));
 sg13g2_nand2_1 _5844_ (.Y(_2073_),
    .A(_1104_),
    .B(_0833_));
 sg13g2_nand2_1 _5845_ (.Y(_2074_),
    .A(_2072_),
    .B(_2073_));
 sg13g2_nand2_1 _5846_ (.Y(_2076_),
    .A(_2074_),
    .B(net123));
 sg13g2_nand2_1 _5847_ (.Y(_2077_),
    .A(_2076_),
    .B(net35));
 sg13g2_nand2_1 _5848_ (.Y(_2078_),
    .A(_2069_),
    .B(_2077_));
 sg13g2_nand2_1 _5849_ (.Y(_2079_),
    .A(_2065_),
    .B(_2078_));
 sg13g2_nand2_1 _5850_ (.Y(_2080_),
    .A(_2050_),
    .B(_2079_));
 sg13g2_nand2_1 _5851_ (.Y(_2081_),
    .A(_2080_),
    .B(net132));
 sg13g2_a21oi_1 _5852_ (.A1(_0999_),
    .A2(_1574_),
    .Y(_2082_),
    .B1(_2716_));
 sg13g2_nand2_1 _5853_ (.Y(_2083_),
    .A(_1165_),
    .B(_1589_));
 sg13g2_nand2_1 _5854_ (.Y(_2084_),
    .A(_2082_),
    .B(_2083_));
 sg13g2_a21oi_1 _5855_ (.A1(_1318_),
    .A2(_1559_),
    .Y(_2085_),
    .B1(_2384_));
 sg13g2_a21oi_1 _5856_ (.A1(_2898_),
    .A2(_2010_),
    .Y(_2087_),
    .B1(_2085_));
 sg13g2_nand2_1 _5857_ (.Y(_2088_),
    .A(_2084_),
    .B(_2087_));
 sg13g2_nand2_1 _5858_ (.Y(_2089_),
    .A(_2088_),
    .B(_2665_));
 sg13g2_a21oi_1 _5859_ (.A1(_2394_),
    .A2(_0387_),
    .Y(_2090_),
    .B1(_0868_));
 sg13g2_nand3_1 _5860_ (.B(_2071_),
    .C(net113),
    .A(_1178_),
    .Y(_2091_));
 sg13g2_nand2_1 _5861_ (.Y(_2092_),
    .A(_2091_),
    .B(_2557_));
 sg13g2_nor2_1 _5862_ (.A(net41),
    .B(_1158_),
    .Y(_2093_));
 sg13g2_a22oi_1 _5863_ (.Y(_2094_),
    .B1(_0332_),
    .B2(_2093_),
    .A2(_2842_),
    .A1(_2577_));
 sg13g2_nand2_1 _5864_ (.Y(_2095_),
    .A(_0302_),
    .B(_2637_));
 sg13g2_a21oi_1 _5865_ (.A1(_2094_),
    .A2(_2095_),
    .Y(_2096_),
    .B1(_0118_));
 sg13g2_nor3_1 _5866_ (.A(_2090_),
    .B(_2092_),
    .C(_2096_),
    .Y(_2098_));
 sg13g2_a21oi_1 _5867_ (.A1(_2089_),
    .A2(_2098_),
    .Y(_2099_),
    .B1(net200));
 sg13g2_nor2_1 _5868_ (.A(net148),
    .B(_2392_),
    .Y(_2100_));
 sg13g2_nor3_1 _5869_ (.A(net149),
    .B(_2203_),
    .C(_2100_),
    .Y(_2101_));
 sg13g2_a21oi_1 _5870_ (.A1(_2101_),
    .A2(_2625_),
    .Y(_2102_),
    .B1(net81));
 sg13g2_nand3_1 _5871_ (.B(_3043_),
    .C(net84),
    .A(_2797_),
    .Y(_2103_));
 sg13g2_nand2_1 _5872_ (.Y(_2104_),
    .A(_2102_),
    .B(_2103_));
 sg13g2_nand2_1 _5873_ (.Y(_2105_),
    .A(_0223_),
    .B(_1407_));
 sg13g2_nand2_1 _5874_ (.Y(_2106_),
    .A(_2105_),
    .B(net26));
 sg13g2_nand2_1 _5875_ (.Y(_2107_),
    .A(_2019_),
    .B(_2970_));
 sg13g2_nand2_1 _5876_ (.Y(_2109_),
    .A(_2107_),
    .B(net70));
 sg13g2_nand3_1 _5877_ (.B(_2106_),
    .C(_2109_),
    .A(_2104_),
    .Y(_2110_));
 sg13g2_nand2_1 _5878_ (.Y(_2111_),
    .A(_2110_),
    .B(net83));
 sg13g2_inv_1 _5879_ (.Y(_2112_),
    .A(_0154_));
 sg13g2_nand2_1 _5880_ (.Y(_2113_),
    .A(_1204_),
    .B(_2506_));
 sg13g2_nand3_1 _5881_ (.B(net84),
    .C(_1991_),
    .A(_2113_),
    .Y(_2114_));
 sg13g2_nand2_1 _5882_ (.Y(_2115_),
    .A(_2114_),
    .B(net22));
 sg13g2_a21oi_1 _5883_ (.A1(_0221_),
    .A2(_2112_),
    .Y(_2116_),
    .B1(_2115_));
 sg13g2_a21oi_1 _5884_ (.A1(_0167_),
    .A2(_0387_),
    .Y(_2117_),
    .B1(net160));
 sg13g2_a21oi_1 _5885_ (.A1(net139),
    .A2(_1162_),
    .Y(_2118_),
    .B1(net142));
 sg13g2_nand3_1 _5886_ (.B(net206),
    .C(net119),
    .A(net30),
    .Y(_2120_));
 sg13g2_nand3_1 _5887_ (.B(_2118_),
    .C(_2120_),
    .A(_2548_),
    .Y(_2121_));
 sg13g2_a21oi_1 _5888_ (.A1(_2117_),
    .A2(_2121_),
    .Y(_2122_),
    .B1(net166));
 sg13g2_nor2b_1 _5889_ (.A(_2116_),
    .B_N(_2122_),
    .Y(_2123_));
 sg13g2_nand2_1 _5890_ (.Y(_2124_),
    .A(_2111_),
    .B(_2123_));
 sg13g2_nand2_1 _5891_ (.Y(_2125_),
    .A(_1056_),
    .B(_2688_));
 sg13g2_nor2_1 _5892_ (.A(_2125_),
    .B(_0324_),
    .Y(_2126_));
 sg13g2_nand3_1 _5893_ (.B(_0471_),
    .C(_2516_),
    .A(_0174_),
    .Y(_2127_));
 sg13g2_nand2_1 _5894_ (.Y(_2128_),
    .A(_2127_),
    .B(_1372_));
 sg13g2_nor2_1 _5895_ (.A(_2126_),
    .B(_2128_),
    .Y(_2129_));
 sg13g2_a22oi_1 _5896_ (.Y(_2131_),
    .B1(_2544_),
    .B2(_1097_),
    .A2(_0951_),
    .A1(net43));
 sg13g2_nand3_1 _5897_ (.B(net47),
    .C(net75),
    .A(_2571_),
    .Y(_2132_));
 sg13g2_inv_1 _5898_ (.Y(_2133_),
    .A(_0748_));
 sg13g2_a21oi_1 _5899_ (.A1(_2131_),
    .A2(_2132_),
    .Y(_2134_),
    .B1(_2133_));
 sg13g2_nor2_1 _5900_ (.A(_2129_),
    .B(_2134_),
    .Y(_2135_));
 sg13g2_a21oi_1 _5901_ (.A1(_0716_),
    .A2(_2651_),
    .Y(_2136_),
    .B1(_0483_));
 sg13g2_nand3_1 _5902_ (.B(_1171_),
    .C(_2653_),
    .A(_0285_),
    .Y(_2137_));
 sg13g2_nand2_1 _5903_ (.Y(_2138_),
    .A(_2136_),
    .B(_2137_));
 sg13g2_nand2_1 _5904_ (.Y(_2139_),
    .A(_2797_),
    .B(_3043_));
 sg13g2_nand2_1 _5905_ (.Y(_2140_),
    .A(_2139_),
    .B(_0600_));
 sg13g2_nand2_1 _5906_ (.Y(_2142_),
    .A(_2138_),
    .B(_2140_));
 sg13g2_nand3_1 _5907_ (.B(_2719_),
    .C(_0604_),
    .A(_2010_),
    .Y(_2143_));
 sg13g2_nor2b_1 _5908_ (.A(_2142_),
    .B_N(_2143_),
    .Y(_2144_));
 sg13g2_nand2_1 _5909_ (.Y(_2145_),
    .A(_2135_),
    .B(_2144_));
 sg13g2_nand2_1 _5910_ (.Y(_2146_),
    .A(_2145_),
    .B(_0728_));
 sg13g2_a221oi_1 _5911_ (.B2(_0958_),
    .C1(_0960_),
    .B1(_2943_),
    .A1(_0977_),
    .Y(_2147_),
    .A2(_1083_));
 sg13g2_nor2_1 _5912_ (.A(_2695_),
    .B(_2147_),
    .Y(_2148_));
 sg13g2_nand2_1 _5913_ (.Y(_2149_),
    .A(_2146_),
    .B(_2148_));
 sg13g2_a21oi_1 _5914_ (.A1(_2099_),
    .A2(_2124_),
    .Y(_2150_),
    .B1(_2149_));
 sg13g2_a21oi_1 _5915_ (.A1(_2029_),
    .A2(_2081_),
    .Y(_0016_),
    .B1(_2150_));
 sg13g2_buf_2 _5916_ (.A(\clk_picker.counter[9] ),
    .X(_2152_));
 sg13g2_nor3_1 _5917_ (.A(_2152_),
    .B(\clk_picker.counter[10] ),
    .C(\clk_picker.counter[11] ),
    .Y(_2153_));
 sg13g2_inv_1 _5918_ (.Y(_2154_),
    .A(\clk_picker.counter[7] ));
 sg13g2_inv_1 _5919_ (.Y(_2155_),
    .A(\clk_picker.counter[8] ));
 sg13g2_nand3_1 _5920_ (.B(_2154_),
    .C(_2155_),
    .A(_2153_),
    .Y(_2156_));
 sg13g2_buf_1 _5921_ (.A(\clk_picker.counter[17] ),
    .X(_2157_));
 sg13g2_nand2_1 _5922_ (.Y(_2158_),
    .A(\clk_picker.counter[12] ),
    .B(\clk_picker.counter[13] ));
 sg13g2_inv_1 _5923_ (.Y(_2159_),
    .A(_2158_));
 sg13g2_nand2_1 _5924_ (.Y(_2160_),
    .A(\clk_picker.counter[14] ),
    .B(\clk_picker.counter[15] ));
 sg13g2_inv_1 _5925_ (.Y(_2161_),
    .A(_2160_));
 sg13g2_nand4_1 _5926_ (.B(_2157_),
    .C(_2159_),
    .A(_2156_),
    .Y(_2163_),
    .D(_2161_));
 sg13g2_inv_1 _5927_ (.Y(_2164_),
    .A(\clk_picker.counter[18] ));
 sg13g2_nand2_1 _5928_ (.Y(_2165_),
    .A(\clk_picker.counter[16] ),
    .B(_2157_));
 sg13g2_nand3_1 _5929_ (.B(_2164_),
    .C(_2165_),
    .A(_2163_),
    .Y(_2166_));
 sg13g2_inv_1 _5930_ (.Y(_2167_),
    .A(\clk_picker.counter[20] ));
 sg13g2_inv_1 _5931_ (.Y(_2168_),
    .A(\clk_picker.counter[23] ));
 sg13g2_nand2_1 _5932_ (.Y(_2169_),
    .A(\clk_picker.counter[21] ),
    .B(\clk_picker.counter[22] ));
 sg13g2_nor3_1 _5933_ (.A(_2167_),
    .B(_2168_),
    .C(_2169_),
    .Y(_2170_));
 sg13g2_nand4_1 _5934_ (.B(\clk_picker.counter[19] ),
    .C(\clk_picker.counter[25] ),
    .A(_2166_),
    .Y(_2171_),
    .D(_2170_));
 sg13g2_nand2_1 _5935_ (.Y(_2172_),
    .A(\clk_picker.counter[24] ),
    .B(\clk_picker.counter[25] ));
 sg13g2_nand2_1 _5936_ (.Y(_2174_),
    .A(_2171_),
    .B(_2172_));
 sg13g2_nand2_1 _5937_ (.Y(_2175_),
    .A(_2174_),
    .B(_0030_));
 sg13g2_nand3_1 _5938_ (.B(\clk_picker.clk_slow ),
    .C(_2172_),
    .A(_2171_),
    .Y(_2176_));
 sg13g2_buf_1 _5939_ (.A(rst_n),
    .X(_2177_));
 sg13g2_inv_2 _5940_ (.Y(_2178_),
    .A(_2177_));
 sg13g2_buf_1 _5941_ (.A(_2178_),
    .X(_2179_));
 sg13g2_a21oi_1 _5942_ (.A1(_2175_),
    .A2(_2176_),
    .Y(_0040_),
    .B1(_2179_));
 sg13g2_nand3_1 _5943_ (.B(_2177_),
    .C(_2172_),
    .A(_2171_),
    .Y(_2180_));
 sg13g2_buf_2 _5944_ (.A(_2180_),
    .X(_2181_));
 sg13g2_buf_1 _5945_ (.A(_2181_),
    .X(_2182_));
 sg13g2_nor2b_1 _5946_ (.A(net21),
    .B_N(_0039_),
    .Y(_0041_));
 sg13g2_inv_1 _5947_ (.Y(_2184_),
    .A(\clk_picker.counter[10] ));
 sg13g2_inv_1 _5948_ (.Y(_2185_),
    .A(\clk_picker.counter[5] ));
 sg13g2_inv_1 _5949_ (.Y(_2186_),
    .A(\clk_picker.counter[6] ));
 sg13g2_nand2_1 _5950_ (.Y(_2187_),
    .A(\clk_picker.counter[1] ),
    .B(\clk_picker.counter[0] ));
 sg13g2_nor2b_1 _5951_ (.A(_2187_),
    .B_N(\clk_picker.counter[2] ),
    .Y(_2188_));
 sg13g2_and2_1 _5952_ (.A(_2188_),
    .B(\clk_picker.counter[3] ),
    .X(_2189_));
 sg13g2_buf_8 _5953_ (.A(_2189_),
    .X(_2190_));
 sg13g2_nand2_1 _5954_ (.Y(_2191_),
    .A(_2190_),
    .B(\clk_picker.counter[4] ));
 sg13g2_nor3_1 _5955_ (.A(_2185_),
    .B(_2186_),
    .C(_2191_),
    .Y(_2192_));
 sg13g2_nand2_1 _5956_ (.Y(_2194_),
    .A(_2192_),
    .B(\clk_picker.counter[7] ));
 sg13g2_nor2_2 _5957_ (.A(_2155_),
    .B(_2194_),
    .Y(_2195_));
 sg13g2_nand2_1 _5958_ (.Y(_2196_),
    .A(_2195_),
    .B(_2152_));
 sg13g2_xnor2_1 _5959_ (.Y(_2197_),
    .A(_2184_),
    .B(_2196_));
 sg13g2_buf_1 _5960_ (.A(_2181_),
    .X(_2198_));
 sg13g2_nor2_1 _5961_ (.A(_2197_),
    .B(net20),
    .Y(_0042_));
 sg13g2_inv_1 _5962_ (.Y(_2199_),
    .A(_2152_));
 sg13g2_nor4_1 _5963_ (.A(_2154_),
    .B(_2155_),
    .C(_2199_),
    .D(_2184_),
    .Y(_2200_));
 sg13g2_inv_1 _5964_ (.Y(_2201_),
    .A(_2200_));
 sg13g2_nor4_2 _5965_ (.A(_2185_),
    .B(_2186_),
    .C(_2201_),
    .Y(_2202_),
    .D(_2191_));
 sg13g2_xnor2_1 _5966_ (.Y(_2204_),
    .A(\clk_picker.counter[11] ),
    .B(_2202_));
 sg13g2_nor2_1 _5967_ (.A(_2204_),
    .B(net20),
    .Y(_0043_));
 sg13g2_inv_1 _5968_ (.Y(_2205_),
    .A(\clk_picker.counter[12] ));
 sg13g2_inv_2 _5969_ (.Y(_2206_),
    .A(_2194_));
 sg13g2_inv_1 _5970_ (.Y(_2207_),
    .A(\clk_picker.counter[11] ));
 sg13g2_nor4_1 _5971_ (.A(_2155_),
    .B(_2199_),
    .C(_2184_),
    .D(_2207_),
    .Y(_2208_));
 sg13g2_nand2_1 _5972_ (.Y(_2209_),
    .A(_2206_),
    .B(_2208_));
 sg13g2_xnor2_1 _5973_ (.Y(_2210_),
    .A(_2205_),
    .B(_2209_));
 sg13g2_nor2_1 _5974_ (.A(_2210_),
    .B(_2198_),
    .Y(_0044_));
 sg13g2_inv_1 _5975_ (.Y(_2211_),
    .A(\clk_picker.counter[13] ));
 sg13g2_nor4_1 _5976_ (.A(_2199_),
    .B(_2184_),
    .C(_2207_),
    .D(_2205_),
    .Y(_2213_));
 sg13g2_nand2_1 _5977_ (.Y(_2214_),
    .A(_2195_),
    .B(_2213_));
 sg13g2_xnor2_1 _5978_ (.Y(_2215_),
    .A(_2211_),
    .B(_2214_));
 sg13g2_nor2_1 _5979_ (.A(_2215_),
    .B(net20),
    .Y(_0045_));
 sg13g2_nor3_1 _5980_ (.A(_2184_),
    .B(_2207_),
    .C(_2158_),
    .Y(_2216_));
 sg13g2_inv_1 _5981_ (.Y(_2217_),
    .A(_2216_));
 sg13g2_nor2_1 _5982_ (.A(_2217_),
    .B(_2196_),
    .Y(_2218_));
 sg13g2_xnor2_1 _5983_ (.Y(_2219_),
    .A(\clk_picker.counter[14] ),
    .B(_2218_));
 sg13g2_nor2_1 _5984_ (.A(net21),
    .B(_2219_),
    .Y(_0046_));
 sg13g2_inv_1 _5985_ (.Y(_2220_),
    .A(\clk_picker.counter[15] ));
 sg13g2_inv_1 _5986_ (.Y(_2222_),
    .A(\clk_picker.counter[14] ));
 sg13g2_nor4_1 _5987_ (.A(_2207_),
    .B(_2205_),
    .C(_2211_),
    .D(_2222_),
    .Y(_2223_));
 sg13g2_nand2_1 _5988_ (.Y(_2224_),
    .A(_2202_),
    .B(_2223_));
 sg13g2_xnor2_1 _5989_ (.Y(_2225_),
    .A(_2220_),
    .B(_2224_));
 sg13g2_nor2_1 _5990_ (.A(_2225_),
    .B(net20),
    .Y(_0047_));
 sg13g2_nand2_1 _5991_ (.Y(_2226_),
    .A(_2159_),
    .B(_2161_));
 sg13g2_nor2_1 _5992_ (.A(_2226_),
    .B(_2209_),
    .Y(_2227_));
 sg13g2_xnor2_1 _5993_ (.Y(_2228_),
    .A(\clk_picker.counter[16] ),
    .B(_2227_));
 sg13g2_nor2_1 _5994_ (.A(_2228_),
    .B(net20),
    .Y(_0048_));
 sg13g2_inv_1 _5995_ (.Y(_2229_),
    .A(\clk_picker.counter[16] ));
 sg13g2_nor4_1 _5996_ (.A(_2211_),
    .B(_2222_),
    .C(_2220_),
    .D(_2229_),
    .Y(_2231_));
 sg13g2_nor2b_1 _5997_ (.A(_2214_),
    .B_N(_2231_),
    .Y(_2232_));
 sg13g2_xnor2_1 _5998_ (.Y(_2233_),
    .A(_2157_),
    .B(_2232_));
 sg13g2_nor2_1 _5999_ (.A(_2233_),
    .B(net20),
    .Y(_0049_));
 sg13g2_nor2_1 _6000_ (.A(_2165_),
    .B(_2160_),
    .Y(_2234_));
 sg13g2_nand2_1 _6001_ (.Y(_2235_),
    .A(_2218_),
    .B(_2234_));
 sg13g2_xnor2_1 _6002_ (.Y(_2236_),
    .A(_2164_),
    .B(_2235_));
 sg13g2_nor2_1 _6003_ (.A(net21),
    .B(_2236_),
    .Y(_0050_));
 sg13g2_inv_1 _6004_ (.Y(_2237_),
    .A(\clk_picker.counter[19] ));
 sg13g2_inv_1 _6005_ (.Y(_2238_),
    .A(_2157_));
 sg13g2_nor4_1 _6006_ (.A(_2220_),
    .B(_2229_),
    .C(_2238_),
    .D(_2164_),
    .Y(_2240_));
 sg13g2_nand3_1 _6007_ (.B(_2223_),
    .C(_2240_),
    .A(_2202_),
    .Y(_2241_));
 sg13g2_xnor2_1 _6008_ (.Y(_2242_),
    .A(_2237_),
    .B(_2241_));
 sg13g2_nor2_1 _6009_ (.A(_2242_),
    .B(net20),
    .Y(_0051_));
 sg13g2_inv_1 _6010_ (.Y(_2243_),
    .A(_2187_));
 sg13g2_nor2_1 _6011_ (.A(\clk_picker.counter[1] ),
    .B(\clk_picker.counter[0] ),
    .Y(_2244_));
 sg13g2_nor3_1 _6012_ (.A(_2243_),
    .B(_2244_),
    .C(_2182_),
    .Y(_0052_));
 sg13g2_nand2_1 _6013_ (.Y(_2245_),
    .A(\clk_picker.counter[18] ),
    .B(\clk_picker.counter[19] ));
 sg13g2_nor2_1 _6014_ (.A(_2165_),
    .B(_2245_),
    .Y(_2246_));
 sg13g2_nand2_1 _6015_ (.Y(_2247_),
    .A(_2227_),
    .B(_2246_));
 sg13g2_xnor2_1 _6016_ (.Y(_2249_),
    .A(_2167_),
    .B(_2247_));
 sg13g2_nor2_1 _6017_ (.A(net21),
    .B(_2249_),
    .Y(_0053_));
 sg13g2_inv_1 _6018_ (.Y(_2250_),
    .A(\clk_picker.counter[21] ));
 sg13g2_nor4_1 _6019_ (.A(_2238_),
    .B(_2164_),
    .C(_2237_),
    .D(_2167_),
    .Y(_2251_));
 sg13g2_nand2_1 _6020_ (.Y(_2252_),
    .A(_2232_),
    .B(_2251_));
 sg13g2_xnor2_1 _6021_ (.Y(_2253_),
    .A(_2250_),
    .B(_2252_));
 sg13g2_nor2_1 _6022_ (.A(net21),
    .B(_2253_),
    .Y(_0054_));
 sg13g2_nor2_1 _6023_ (.A(_2185_),
    .B(_2191_),
    .Y(_2254_));
 sg13g2_nor3_1 _6024_ (.A(_2167_),
    .B(_2250_),
    .C(_2245_),
    .Y(_2255_));
 sg13g2_nand4_1 _6025_ (.B(\clk_picker.counter[7] ),
    .C(\clk_picker.counter[8] ),
    .A(\clk_picker.counter[6] ),
    .Y(_2256_),
    .D(_2152_));
 sg13g2_nor2_1 _6026_ (.A(_2256_),
    .B(_2217_),
    .Y(_2258_));
 sg13g2_nand4_1 _6027_ (.B(_2255_),
    .C(_2258_),
    .A(_2254_),
    .Y(_2259_),
    .D(_2234_));
 sg13g2_xor2_1 _6028_ (.B(_2259_),
    .A(\clk_picker.counter[22] ),
    .X(_2260_));
 sg13g2_nor2_1 _6029_ (.A(_2260_),
    .B(_2198_),
    .Y(_0055_));
 sg13g2_nand2b_1 _6030_ (.Y(_2261_),
    .B(_2251_),
    .A_N(_2169_));
 sg13g2_nor4_1 _6031_ (.A(_2220_),
    .B(_2229_),
    .C(_2261_),
    .D(_2224_),
    .Y(_2262_));
 sg13g2_xnor2_1 _6032_ (.Y(_2263_),
    .A(\clk_picker.counter[23] ),
    .B(_2262_));
 sg13g2_nor2_1 _6033_ (.A(net21),
    .B(_2263_),
    .Y(_0056_));
 sg13g2_inv_1 _6034_ (.Y(_2264_),
    .A(\clk_picker.counter[24] ));
 sg13g2_nand3_1 _6035_ (.B(_2170_),
    .C(_2246_),
    .A(_2227_),
    .Y(_2265_));
 sg13g2_xnor2_1 _6036_ (.Y(_2267_),
    .A(_2264_),
    .B(_2265_));
 sg13g2_nor2_1 _6037_ (.A(net21),
    .B(_2267_),
    .Y(_0057_));
 sg13g2_nor3_1 _6038_ (.A(_2168_),
    .B(_2264_),
    .C(_2261_),
    .Y(_2268_));
 sg13g2_a21oi_1 _6039_ (.A1(_2232_),
    .A2(_2268_),
    .Y(_2269_),
    .B1(\clk_picker.counter[25] ));
 sg13g2_nor2_1 _6040_ (.A(_2269_),
    .B(net20),
    .Y(_0058_));
 sg13g2_nor2_1 _6041_ (.A(\clk_picker.counter[2] ),
    .B(_2243_),
    .Y(_2270_));
 sg13g2_nor3_1 _6042_ (.A(_2188_),
    .B(_2270_),
    .C(_2181_),
    .Y(_0059_));
 sg13g2_nor2_1 _6043_ (.A(\clk_picker.counter[3] ),
    .B(_2188_),
    .Y(_2271_));
 sg13g2_nor3_1 _6044_ (.A(_2190_),
    .B(_2271_),
    .C(_2181_),
    .Y(_0060_));
 sg13g2_xnor2_1 _6045_ (.Y(_2272_),
    .A(\clk_picker.counter[4] ),
    .B(_2190_));
 sg13g2_nor2_1 _6046_ (.A(_2272_),
    .B(net21),
    .Y(_0061_));
 sg13g2_a21oi_1 _6047_ (.A1(_2190_),
    .A2(\clk_picker.counter[4] ),
    .Y(_2274_),
    .B1(\clk_picker.counter[5] ));
 sg13g2_nor3_1 _6048_ (.A(_2254_),
    .B(_2274_),
    .C(_2181_),
    .Y(_0062_));
 sg13g2_nor2_1 _6049_ (.A(\clk_picker.counter[6] ),
    .B(_2254_),
    .Y(_2275_));
 sg13g2_nor3_1 _6050_ (.A(_2192_),
    .B(_2275_),
    .C(_2181_),
    .Y(_0063_));
 sg13g2_nor2_1 _6051_ (.A(\clk_picker.counter[7] ),
    .B(_2192_),
    .Y(_2276_));
 sg13g2_nor3_1 _6052_ (.A(_2206_),
    .B(_2276_),
    .C(_2181_),
    .Y(_0064_));
 sg13g2_nor2_1 _6053_ (.A(\clk_picker.counter[8] ),
    .B(_2206_),
    .Y(_2277_));
 sg13g2_nor3_1 _6054_ (.A(_2195_),
    .B(_2277_),
    .C(_2181_),
    .Y(_0065_));
 sg13g2_xnor2_1 _6055_ (.Y(_2278_),
    .A(_2152_),
    .B(_2195_));
 sg13g2_nor2_1 _6056_ (.A(_2278_),
    .B(_2182_),
    .Y(_0066_));
 sg13g2_nor2_1 _6057_ (.A(net2),
    .B(\transformer_1.started ),
    .Y(_2280_));
 sg13g2_buf_1 _6058_ (.A(_2280_),
    .X(_2281_));
 sg13g2_nor2_1 _6059_ (.A(_0031_),
    .B(net191),
    .Y(_2282_));
 sg13g2_nor3_1 _6060_ (.A(net2),
    .B(\transformer_1.started ),
    .C(\line_mapper_1.pointer_addr[10] ),
    .Y(_2283_));
 sg13g2_or2_1 _6061_ (.X(_2284_),
    .B(\chars_remaining[1] ),
    .A(\chars_remaining[2] ));
 sg13g2_nor2_1 _6062_ (.A(\chars_remaining[0] ),
    .B(_2284_),
    .Y(_2285_));
 sg13g2_inv_1 _6063_ (.Y(_2286_),
    .A(_2285_));
 sg13g2_nor4_2 _6064_ (.A(\chars_remaining[5] ),
    .B(\chars_remaining[4] ),
    .C(\chars_remaining[3] ),
    .Y(_2287_),
    .D(_2286_));
 sg13g2_nand2b_1 _6065_ (.Y(_2288_),
    .B(_2287_),
    .A_N(\chars_remaining[6] ));
 sg13g2_inv_1 _6066_ (.Y(_2290_),
    .A(\chars_remaining[8] ));
 sg13g2_nand2b_1 _6067_ (.Y(_2291_),
    .B(_2290_),
    .A_N(\chars_remaining[7] ));
 sg13g2_nor2_1 _6068_ (.A(\chars_remaining[9] ),
    .B(_2291_),
    .Y(_2292_));
 sg13g2_nor2b_1 _6069_ (.A(_2288_),
    .B_N(_2292_),
    .Y(_2293_));
 sg13g2_nor2b_1 _6070_ (.A(net191),
    .B_N(_2293_),
    .Y(_2294_));
 sg13g2_buf_1 _6071_ (.A(_2294_),
    .X(_2295_));
 sg13g2_nor4_1 _6072_ (.A(net211),
    .B(_2282_),
    .C(_2283_),
    .D(net19),
    .Y(_0067_));
 sg13g2_buf_1 _6073_ (.A(net191),
    .X(_2296_));
 sg13g2_xnor2_1 _6074_ (.Y(_2297_),
    .A(\chars_remaining[1] ),
    .B(\chars_remaining[0] ));
 sg13g2_nor2_1 _6075_ (.A(_2281_),
    .B(_2293_),
    .Y(_2298_));
 sg13g2_buf_2 _6076_ (.A(_2298_),
    .X(_2300_));
 sg13g2_buf_1 _6077_ (.A(_2300_),
    .X(_2301_));
 sg13g2_a22oi_1 _6078_ (.Y(_2302_),
    .B1(_2297_),
    .B2(net18),
    .A2(net159),
    .A1(\line_mapper_1.pointer_addr[11] ));
 sg13g2_nor2_1 _6079_ (.A(net211),
    .B(_2302_),
    .Y(_0068_));
 sg13g2_o21ai_1 _6080_ (.B1(\chars_remaining[2] ),
    .Y(_2303_),
    .A1(\chars_remaining[1] ),
    .A2(\chars_remaining[0] ));
 sg13g2_nand2_1 _6081_ (.Y(_2304_),
    .A(_2286_),
    .B(_2303_));
 sg13g2_a22oi_1 _6082_ (.Y(_2305_),
    .B1(_2304_),
    .B2(net18),
    .A2(net159),
    .A1(\line_mapper_1.pointer_addr[12] ));
 sg13g2_nor2_1 _6083_ (.A(net211),
    .B(_2305_),
    .Y(_0069_));
 sg13g2_nor2_1 _6084_ (.A(\chars_remaining[3] ),
    .B(_2286_),
    .Y(_2306_));
 sg13g2_nor2b_1 _6085_ (.A(_2285_),
    .B_N(\chars_remaining[3] ),
    .Y(_2307_));
 sg13g2_o21ai_1 _6086_ (.B1(_2300_),
    .Y(_2309_),
    .A1(_2306_),
    .A2(_2307_));
 sg13g2_nand2_1 _6087_ (.Y(_2310_),
    .A(net159),
    .B(\line_mapper_1.pointer_addr[13] ));
 sg13g2_a21oi_1 _6088_ (.A1(_2309_),
    .A2(_2310_),
    .Y(_0070_),
    .B1(net211));
 sg13g2_xor2_1 _6089_ (.B(_2306_),
    .A(\chars_remaining[4] ),
    .X(_2311_));
 sg13g2_a22oi_1 _6090_ (.Y(_2312_),
    .B1(_2311_),
    .B2(net18),
    .A2(net159),
    .A1(\line_mapper_1.pointer_addr[14] ));
 sg13g2_nor2_1 _6091_ (.A(net211),
    .B(_2312_),
    .Y(_0071_));
 sg13g2_nor3_1 _6092_ (.A(\chars_remaining[4] ),
    .B(\chars_remaining[3] ),
    .C(_2284_),
    .Y(_2313_));
 sg13g2_nand2_1 _6093_ (.Y(_2314_),
    .A(_2313_),
    .B(_0031_));
 sg13g2_xnor2_1 _6094_ (.Y(_2315_),
    .A(\chars_remaining[5] ),
    .B(_2314_));
 sg13g2_a22oi_1 _6095_ (.Y(_2316_),
    .B1(_2315_),
    .B2(net18),
    .A2(_2296_),
    .A1(\line_mapper_1.pointer_addr[15] ));
 sg13g2_nor2_1 _6096_ (.A(_2179_),
    .B(_2316_),
    .Y(_0072_));
 sg13g2_nor2_1 _6097_ (.A(_2178_),
    .B(_2281_),
    .Y(_2318_));
 sg13g2_inv_1 _6098_ (.Y(_2319_),
    .A(_2318_));
 sg13g2_xnor2_1 _6099_ (.Y(_2320_),
    .A(\chars_remaining[6] ),
    .B(_2287_));
 sg13g2_nor3_1 _6100_ (.A(_2319_),
    .B(_2293_),
    .C(_2320_),
    .Y(_0073_));
 sg13g2_or3_1 _6101_ (.A(\chars_remaining[7] ),
    .B(_2292_),
    .C(_2288_),
    .X(_2321_));
 sg13g2_buf_1 _6102_ (.A(_2321_),
    .X(_2322_));
 sg13g2_nand2_1 _6103_ (.Y(_2323_),
    .A(_2288_),
    .B(\chars_remaining[7] ));
 sg13g2_a21oi_1 _6104_ (.A1(_2322_),
    .A2(_2323_),
    .Y(_0074_),
    .B1(_2319_));
 sg13g2_o21ai_1 _6105_ (.B1(_2318_),
    .Y(_2324_),
    .A1(_2290_),
    .A2(_2322_));
 sg13g2_a21oi_1 _6106_ (.A1(_2290_),
    .A2(_2322_),
    .Y(_0075_),
    .B1(_2324_));
 sg13g2_inv_1 _6107_ (.Y(_2326_),
    .A(\chars_remaining[9] ));
 sg13g2_nor2_1 _6108_ (.A(_2291_),
    .B(_2288_),
    .Y(_2327_));
 sg13g2_nor3_1 _6109_ (.A(_2326_),
    .B(_2319_),
    .C(_2327_),
    .Y(_0076_));
 sg13g2_a22oi_1 _6110_ (.Y(_2328_),
    .B1(_1260_),
    .B2(net19),
    .A2(net159),
    .A1(\line_mapper_1.pointer_addr[0] ));
 sg13g2_a21oi_1 _6111_ (.A1(net18),
    .A2(_1162_),
    .Y(_2329_),
    .B1(net211));
 sg13g2_nand2_1 _6112_ (.Y(_0077_),
    .A(_2328_),
    .B(_2329_));
 sg13g2_a22oi_1 _6113_ (.Y(_2330_),
    .B1(net119),
    .B2(net19),
    .A2(_2300_),
    .A1(_2684_));
 sg13g2_a21oi_1 _6114_ (.A1(net159),
    .A2(\line_mapper_1.pointer_addr[1] ),
    .Y(_2331_),
    .B1(net211));
 sg13g2_nand2_1 _6115_ (.Y(_0078_),
    .A(_2330_),
    .B(_2331_));
 sg13g2_nand2_1 _6116_ (.Y(_2333_),
    .A(net19),
    .B(_1435_));
 sg13g2_nand2_1 _6117_ (.Y(_2334_),
    .A(net18),
    .B(_0258_));
 sg13g2_a21oi_1 _6118_ (.A1(net159),
    .A2(\line_mapper_1.pointer_addr[2] ),
    .Y(_2335_),
    .B1(_2178_));
 sg13g2_nand3_1 _6119_ (.B(_2334_),
    .C(_2335_),
    .A(_2333_),
    .Y(_0079_));
 sg13g2_nor2_1 _6120_ (.A(_1162_),
    .B(_2603_),
    .Y(_2336_));
 sg13g2_xnor2_1 _6121_ (.Y(_2337_),
    .A(net30),
    .B(_2336_));
 sg13g2_a22oi_1 _6122_ (.Y(_2338_),
    .B1(net33),
    .B2(net19),
    .A2(_2337_),
    .A1(_2300_));
 sg13g2_a21oi_1 _6123_ (.A1(_2296_),
    .A2(\line_mapper_1.pointer_addr[3] ),
    .Y(_2339_),
    .B1(_2178_));
 sg13g2_nand2_1 _6124_ (.Y(_0080_),
    .A(_2338_),
    .B(_2339_));
 sg13g2_nand2_1 _6125_ (.Y(_2340_),
    .A(net19),
    .B(_2419_));
 sg13g2_xnor2_1 _6126_ (.Y(_2342_),
    .A(_3023_),
    .B(_0598_));
 sg13g2_nand2_1 _6127_ (.Y(_2343_),
    .A(_2301_),
    .B(_2342_));
 sg13g2_a21oi_1 _6128_ (.A1(net191),
    .A2(\line_mapper_1.pointer_addr[4] ),
    .Y(_2344_),
    .B1(_2178_));
 sg13g2_nand3_1 _6129_ (.B(_2343_),
    .C(_2344_),
    .A(_2340_),
    .Y(_0081_));
 sg13g2_nor2_1 _6130_ (.A(_1998_),
    .B(_2020_),
    .Y(_2345_));
 sg13g2_inv_1 _6131_ (.Y(_2346_),
    .A(_2345_));
 sg13g2_nor2_1 _6132_ (.A(net75),
    .B(_2346_),
    .Y(_2347_));
 sg13g2_nand2_1 _6133_ (.Y(_2348_),
    .A(_2346_),
    .B(_2733_));
 sg13g2_nand3b_1 _6134_ (.B(_2300_),
    .C(_2348_),
    .Y(_2349_),
    .A_N(_2347_));
 sg13g2_nand2_1 _6135_ (.Y(_2350_),
    .A(net19),
    .B(net130));
 sg13g2_a21oi_1 _6136_ (.A1(net191),
    .A2(\line_mapper_1.pointer_addr[5] ),
    .Y(_2352_),
    .B1(_2178_));
 sg13g2_nand3_1 _6137_ (.B(_2350_),
    .C(_2352_),
    .A(_2349_),
    .Y(_0082_));
 sg13g2_nand2_1 _6138_ (.Y(_2353_),
    .A(_2295_),
    .B(net117));
 sg13g2_xnor2_1 _6139_ (.Y(_2354_),
    .A(net83),
    .B(_2347_));
 sg13g2_nand2_1 _6140_ (.Y(_2355_),
    .A(_2301_),
    .B(_2354_));
 sg13g2_a21oi_1 _6141_ (.A1(net191),
    .A2(\line_mapper_1.pointer_addr[6] ),
    .Y(_2356_),
    .B1(_2178_));
 sg13g2_nand3_1 _6142_ (.B(_2355_),
    .C(_2356_),
    .A(_2353_),
    .Y(_0083_));
 sg13g2_nand2_1 _6143_ (.Y(_2357_),
    .A(_1537_),
    .B(_2336_));
 sg13g2_xnor2_1 _6144_ (.Y(_2358_),
    .A(net164),
    .B(_2357_));
 sg13g2_a22oi_1 _6145_ (.Y(_2359_),
    .B1(net164),
    .B2(_2295_),
    .A2(_2358_),
    .A1(_2300_));
 sg13g2_a21oi_1 _6146_ (.A1(net159),
    .A2(\line_mapper_1.pointer_addr[7] ),
    .Y(_2361_),
    .B1(_2178_));
 sg13g2_nand2_1 _6147_ (.Y(_0084_),
    .A(_2359_),
    .B(_2361_));
 sg13g2_a22oi_1 _6148_ (.Y(_2362_),
    .B1(net200),
    .B2(net19),
    .A2(net191),
    .A1(\line_mapper_1.pointer_addr[8] ));
 sg13g2_nand2_1 _6149_ (.Y(_2363_),
    .A(_2347_),
    .B(_2559_));
 sg13g2_nor2_1 _6150_ (.A(net170),
    .B(_2363_),
    .Y(_2364_));
 sg13g2_nand2_1 _6151_ (.Y(_2365_),
    .A(_2363_),
    .B(net163));
 sg13g2_nand3b_1 _6152_ (.B(_2300_),
    .C(_2365_),
    .Y(_2366_),
    .A_N(_2364_));
 sg13g2_nand3_1 _6153_ (.B(_2177_),
    .C(_2366_),
    .A(_2362_),
    .Y(_0085_));
 sg13g2_a22oi_1 _6154_ (.Y(_2367_),
    .B1(net196),
    .B2(_2294_),
    .A2(net191),
    .A1(\line_mapper_1.pointer_addr[9] ));
 sg13g2_xnor2_1 _6155_ (.Y(_2368_),
    .A(net195),
    .B(_2364_));
 sg13g2_nand2_1 _6156_ (.Y(_2370_),
    .A(net18),
    .B(_2368_));
 sg13g2_nand3_1 _6157_ (.B(_2177_),
    .C(_2370_),
    .A(_2367_),
    .Y(_0086_));
 sg13g2_inv_1 _6158_ (.Y(_2371_),
    .A(\transformer_1.started ));
 sg13g2_a21oi_1 _6159_ (.A1(net18),
    .A2(_2371_),
    .Y(_0087_),
    .B1(net211));
 sg13g2_mux2_1 _6160_ (.A0(\clk_picker.clk_slow ),
    .A1(clknet_2_1__leaf_clk),
    .S(net3),
    .X(clk_buffered));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _6163__221 (.L_HI(net221));
 sg13g2_buf_1 _6163_ (.A(net221),
    .X(uio_oe[0]));
 sg13g2_buf_1 _6164_ (.A(net222),
    .X(uio_oe[1]));
 sg13g2_buf_1 _6165_ (.A(net223),
    .X(uio_oe[2]));
 sg13g2_buf_1 _6166_ (.A(net224),
    .X(uio_oe[3]));
 sg13g2_buf_1 _6167_ (.A(net225),
    .X(uio_oe[4]));
 sg13g2_buf_1 _6168_ (.A(net226),
    .X(uio_oe[5]));
 sg13g2_buf_1 _6169_ (.A(net227),
    .X(uio_oe[6]));
 sg13g2_buf_1 _6170_ (.A(net228),
    .X(uio_oe[7]));
 sg13g2_buf_1 _6171_ (.A(net219),
    .X(uio_out[7]));
 sg13g2_buf_1 _6172_ (.A(net220),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \clk_picker.clk_slow$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net229),
    .D(_0040_),
    .Q_N(_0030_),
    .Q(\clk_picker.clk_slow ));
 sg13g2_dfrbp_1 \clk_picker.counter[0]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net230),
    .D(_0041_),
    .Q_N(_0039_),
    .Q(\clk_picker.counter[0] ));
 sg13g2_dfrbp_1 \clk_picker.counter[10]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net231),
    .D(_0042_),
    .Q_N(_3087_),
    .Q(\clk_picker.counter[10] ));
 sg13g2_dfrbp_1 \clk_picker.counter[11]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net232),
    .D(_0043_),
    .Q_N(_3086_),
    .Q(\clk_picker.counter[11] ));
 sg13g2_dfrbp_1 \clk_picker.counter[12]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net233),
    .D(_0044_),
    .Q_N(_3085_),
    .Q(\clk_picker.counter[12] ));
 sg13g2_dfrbp_1 \clk_picker.counter[13]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net234),
    .D(_0045_),
    .Q_N(_3084_),
    .Q(\clk_picker.counter[13] ));
 sg13g2_dfrbp_1 \clk_picker.counter[14]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net235),
    .D(_0046_),
    .Q_N(_3083_),
    .Q(\clk_picker.counter[14] ));
 sg13g2_dfrbp_1 \clk_picker.counter[15]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net236),
    .D(_0047_),
    .Q_N(_3082_),
    .Q(\clk_picker.counter[15] ));
 sg13g2_dfrbp_1 \clk_picker.counter[16]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net237),
    .D(_0048_),
    .Q_N(_3081_),
    .Q(\clk_picker.counter[16] ));
 sg13g2_dfrbp_1 \clk_picker.counter[17]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net238),
    .D(_0049_),
    .Q_N(_3080_),
    .Q(\clk_picker.counter[17] ));
 sg13g2_dfrbp_1 \clk_picker.counter[18]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net239),
    .D(_0050_),
    .Q_N(_3079_),
    .Q(\clk_picker.counter[18] ));
 sg13g2_dfrbp_1 \clk_picker.counter[19]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net240),
    .D(_0051_),
    .Q_N(_3078_),
    .Q(\clk_picker.counter[19] ));
 sg13g2_dfrbp_1 \clk_picker.counter[1]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net241),
    .D(_0052_),
    .Q_N(_3077_),
    .Q(\clk_picker.counter[1] ));
 sg13g2_dfrbp_1 \clk_picker.counter[20]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net242),
    .D(_0053_),
    .Q_N(_3076_),
    .Q(\clk_picker.counter[20] ));
 sg13g2_dfrbp_1 \clk_picker.counter[21]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net243),
    .D(_0054_),
    .Q_N(_3075_),
    .Q(\clk_picker.counter[21] ));
 sg13g2_dfrbp_1 \clk_picker.counter[22]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net244),
    .D(_0055_),
    .Q_N(_3074_),
    .Q(\clk_picker.counter[22] ));
 sg13g2_dfrbp_1 \clk_picker.counter[23]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net245),
    .D(_0056_),
    .Q_N(_3073_),
    .Q(\clk_picker.counter[23] ));
 sg13g2_dfrbp_1 \clk_picker.counter[24]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net246),
    .D(_0057_),
    .Q_N(_3072_),
    .Q(\clk_picker.counter[24] ));
 sg13g2_dfrbp_1 \clk_picker.counter[25]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net247),
    .D(_0058_),
    .Q_N(_3071_),
    .Q(\clk_picker.counter[25] ));
 sg13g2_dfrbp_1 \clk_picker.counter[2]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net248),
    .D(_0059_),
    .Q_N(_3070_),
    .Q(\clk_picker.counter[2] ));
 sg13g2_dfrbp_1 \clk_picker.counter[3]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net249),
    .D(_0060_),
    .Q_N(_3069_),
    .Q(\clk_picker.counter[3] ));
 sg13g2_dfrbp_1 \clk_picker.counter[4]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net250),
    .D(_0061_),
    .Q_N(_3068_),
    .Q(\clk_picker.counter[4] ));
 sg13g2_dfrbp_1 \clk_picker.counter[5]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net251),
    .D(_0062_),
    .Q_N(_3067_),
    .Q(\clk_picker.counter[5] ));
 sg13g2_dfrbp_1 \clk_picker.counter[6]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net252),
    .D(_0063_),
    .Q_N(_3066_),
    .Q(\clk_picker.counter[6] ));
 sg13g2_dfrbp_1 \clk_picker.counter[7]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net253),
    .D(_0064_),
    .Q_N(_3065_),
    .Q(\clk_picker.counter[7] ));
 sg13g2_dfrbp_1 \clk_picker.counter[8]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net254),
    .D(_0065_),
    .Q_N(_3064_),
    .Q(\clk_picker.counter[8] ));
 sg13g2_dfrbp_1 \clk_picker.counter[9]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net255),
    .D(_0066_),
    .Q_N(_3088_),
    .Q(\clk_picker.counter[9] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[0]$_DFF_P_  (.CLK(clknet_3_0_0_clk_buffered),
    .RESET_B(net256),
    .D(_0000_),
    .Q_N(_3089_),
    .Q(\line_mapper_1.pointer_addr[0] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[10]$_DFF_P_  (.CLK(clknet_3_1_0_clk_buffered),
    .RESET_B(net257),
    .D(_0001_),
    .Q_N(_3090_),
    .Q(\line_mapper_1.pointer_addr[10] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[11]$_DFF_P_  (.CLK(clknet_3_3_0_clk_buffered),
    .RESET_B(net258),
    .D(_0002_),
    .Q_N(_3091_),
    .Q(\line_mapper_1.pointer_addr[11] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[12]$_DFF_P_  (.CLK(clknet_3_3_0_clk_buffered),
    .RESET_B(net259),
    .D(_0003_),
    .Q_N(_3092_),
    .Q(\line_mapper_1.pointer_addr[12] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[13]$_DFF_P_  (.CLK(clknet_3_2_0_clk_buffered),
    .RESET_B(net260),
    .D(_0004_),
    .Q_N(_3093_),
    .Q(\line_mapper_1.pointer_addr[13] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[14]$_DFF_P_  (.CLK(clknet_3_3_0_clk_buffered),
    .RESET_B(net261),
    .D(_0005_),
    .Q_N(_3094_),
    .Q(\line_mapper_1.pointer_addr[14] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[15]$_DFF_P_  (.CLK(clknet_3_1_0_clk_buffered),
    .RESET_B(net262),
    .D(_0006_),
    .Q_N(_3095_),
    .Q(\line_mapper_1.pointer_addr[15] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[1]$_DFF_P_  (.CLK(clknet_3_0_0_clk_buffered),
    .RESET_B(net263),
    .D(_0007_),
    .Q_N(_3096_),
    .Q(\line_mapper_1.pointer_addr[1] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[2]$_DFF_P_  (.CLK(clknet_3_0_0_clk_buffered),
    .RESET_B(net264),
    .D(_0008_),
    .Q_N(_3097_),
    .Q(\line_mapper_1.pointer_addr[2] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[3]$_DFF_P_  (.CLK(clknet_3_1_0_clk_buffered),
    .RESET_B(net265),
    .D(_0009_),
    .Q_N(_3098_),
    .Q(\line_mapper_1.pointer_addr[3] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[4]$_DFF_P_  (.CLK(clknet_3_0_0_clk_buffered),
    .RESET_B(net266),
    .D(_0010_),
    .Q_N(_3099_),
    .Q(\line_mapper_1.pointer_addr[4] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[5]$_DFF_P_  (.CLK(clknet_3_0_0_clk_buffered),
    .RESET_B(net267),
    .D(_0011_),
    .Q_N(_3100_),
    .Q(\line_mapper_1.pointer_addr[5] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[6]$_DFF_P_  (.CLK(clknet_3_1_0_clk_buffered),
    .RESET_B(net268),
    .D(_0012_),
    .Q_N(_3101_),
    .Q(\line_mapper_1.pointer_addr[6] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[7]$_DFF_P_  (.CLK(clknet_3_0_0_clk_buffered),
    .RESET_B(net269),
    .D(_0013_),
    .Q_N(_3102_),
    .Q(\line_mapper_1.pointer_addr[7] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[8]$_DFF_P_  (.CLK(clknet_3_0_0_clk_buffered),
    .RESET_B(net270),
    .D(_0014_),
    .Q_N(_3103_),
    .Q(\line_mapper_1.pointer_addr[8] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[9]$_DFF_P_  (.CLK(clknet_3_1_0_clk_buffered),
    .RESET_B(net271),
    .D(_0015_),
    .Q_N(_3104_),
    .Q(\line_mapper_1.pointer_addr[9] ));
 sg13g2_dfrbp_1 \memory_1.dout[0]$_DFF_P_  (.CLK(clknet_3_2_0_clk_buffered),
    .RESET_B(net272),
    .D(_0016_),
    .Q_N(_3105_),
    .Q(net11));
 sg13g2_dfrbp_1 \memory_1.dout[10]$_DFF_P_  (.CLK(clknet_3_2_0_clk_buffered),
    .RESET_B(net273),
    .D(_0029_),
    .Q_N(_3106_),
    .Q(net6));
 sg13g2_dfrbp_1 \memory_1.dout[11]$_DFF_P_  (.CLK(clknet_3_2_0_clk_buffered),
    .RESET_B(net274),
    .D(_0017_),
    .Q_N(_3107_),
    .Q(net7));
 sg13g2_dfrbp_1 \memory_1.dout[12]$_DFF_P_  (.CLK(clknet_3_7_0_clk_buffered),
    .RESET_B(net275),
    .D(_0018_),
    .Q_N(_3108_),
    .Q(net8));
 sg13g2_dfrbp_1 \memory_1.dout[13]$_DFF_P_  (.CLK(clknet_3_7_0_clk_buffered),
    .RESET_B(net276),
    .D(_0019_),
    .Q_N(_3109_),
    .Q(net9));
 sg13g2_dfrbp_1 \memory_1.dout[14]$_DFF_P_  (.CLK(clknet_3_7_0_clk_buffered),
    .RESET_B(net277),
    .D(_0020_),
    .Q_N(_3110_),
    .Q(net10));
 sg13g2_dfrbp_1 \memory_1.dout[1]$_DFF_P_  (.CLK(clknet_3_3_0_clk_buffered),
    .RESET_B(net278),
    .D(_0021_),
    .Q_N(_3111_),
    .Q(net12));
 sg13g2_dfrbp_1 \memory_1.dout[2]$_DFF_P_  (.CLK(clknet_3_2_0_clk_buffered),
    .RESET_B(net279),
    .D(_0022_),
    .Q_N(_3112_),
    .Q(net13));
 sg13g2_dfrbp_1 \memory_1.dout[3]$_DFF_P_  (.CLK(clknet_3_2_0_clk_buffered),
    .RESET_B(net280),
    .D(_0023_),
    .Q_N(_3113_),
    .Q(net14));
 sg13g2_dfrbp_1 \memory_1.dout[4]$_DFF_P_  (.CLK(clknet_3_2_0_clk_buffered),
    .RESET_B(net281),
    .D(_0024_),
    .Q_N(_3114_),
    .Q(net15));
 sg13g2_dfrbp_1 \memory_1.dout[5]$_DFF_P_  (.CLK(clknet_3_3_0_clk_buffered),
    .RESET_B(net282),
    .D(_0025_),
    .Q_N(_3115_),
    .Q(net16));
 sg13g2_dfrbp_1 \memory_1.dout[6]$_DFF_P_  (.CLK(clknet_3_7_0_clk_buffered),
    .RESET_B(net283),
    .D(_0026_),
    .Q_N(_3116_),
    .Q(net17));
 sg13g2_dfrbp_1 \memory_1.dout[8]$_DFF_P_  (.CLK(clknet_3_7_0_clk_buffered),
    .RESET_B(net284),
    .D(_0027_),
    .Q_N(_3117_),
    .Q(net4));
 sg13g2_dfrbp_1 \memory_1.dout[9]$_DFF_P_  (.CLK(clknet_3_3_0_clk_buffered),
    .RESET_B(net285),
    .D(_0028_),
    .Q_N(_3063_),
    .Q(net5));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[0]$_SDFFE_PN0P_  (.CLK(clknet_3_6_0_clk_buffered),
    .RESET_B(net286),
    .D(_0067_),
    .Q_N(_0031_),
    .Q(\chars_remaining[0] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[1]$_SDFFE_PN0P_  (.CLK(clknet_3_6_0_clk_buffered),
    .RESET_B(net287),
    .D(_0068_),
    .Q_N(_3062_),
    .Q(\chars_remaining[1] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[2]$_SDFFE_PN0P_  (.CLK(clknet_3_6_0_clk_buffered),
    .RESET_B(net288),
    .D(_0069_),
    .Q_N(_3061_),
    .Q(\chars_remaining[2] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[3]$_SDFFE_PN0P_  (.CLK(clknet_3_6_0_clk_buffered),
    .RESET_B(net289),
    .D(_0070_),
    .Q_N(_3060_),
    .Q(\chars_remaining[3] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[4]$_SDFFE_PN0P_  (.CLK(clknet_3_6_0_clk_buffered),
    .RESET_B(net290),
    .D(_0071_),
    .Q_N(_3059_),
    .Q(\chars_remaining[4] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[5]$_SDFFE_PN0P_  (.CLK(clknet_3_4_0_clk_buffered),
    .RESET_B(net291),
    .D(_0072_),
    .Q_N(_3058_),
    .Q(\chars_remaining[5] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[6]$_SDFFE_PN0P_  (.CLK(clknet_3_7_0_clk_buffered),
    .RESET_B(net292),
    .D(_0073_),
    .Q_N(_3057_),
    .Q(\chars_remaining[6] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[7]$_SDFFE_PN0P_  (.CLK(clknet_3_4_0_clk_buffered),
    .RESET_B(net293),
    .D(_0074_),
    .Q_N(_3056_),
    .Q(\chars_remaining[7] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[8]$_SDFFE_PN0P_  (.CLK(clknet_3_4_0_clk_buffered),
    .RESET_B(net294),
    .D(_0075_),
    .Q_N(_3055_),
    .Q(\chars_remaining[8] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[9]$_SDFFE_PN0P_  (.CLK(clknet_3_4_0_clk_buffered),
    .RESET_B(net295),
    .D(_0076_),
    .Q_N(_3054_),
    .Q(\chars_remaining[9] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[0]$_SDFFE_PN1P_  (.CLK(clknet_3_4_0_clk_buffered),
    .RESET_B(net296),
    .D(_0077_),
    .Q_N(_0032_),
    .Q(\mem_addr[0] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[1]$_SDFFE_PN1P_  (.CLK(clknet_3_5_0_clk_buffered),
    .RESET_B(net297),
    .D(_0078_),
    .Q_N(_0038_),
    .Q(\mem_addr[1] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[2]$_SDFFE_PN1P_  (.CLK(clknet_3_5_0_clk_buffered),
    .RESET_B(net298),
    .D(_0079_),
    .Q_N(_0037_),
    .Q(\mem_addr[2] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[3]$_SDFFE_PN1P_  (.CLK(clknet_3_5_0_clk_buffered),
    .RESET_B(net299),
    .D(_0080_),
    .Q_N(_0036_),
    .Q(\mem_addr[3] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[4]$_SDFFE_PN1P_  (.CLK(clknet_3_5_0_clk_buffered),
    .RESET_B(net300),
    .D(_0081_),
    .Q_N(_0035_),
    .Q(\mem_addr[4] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[5]$_SDFFE_PN1P_  (.CLK(clknet_3_5_0_clk_buffered),
    .RESET_B(net301),
    .D(_0082_),
    .Q_N(_0034_),
    .Q(\mem_addr[5] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[6]$_SDFFE_PN1P_  (.CLK(clknet_3_5_0_clk_buffered),
    .RESET_B(net302),
    .D(_0083_),
    .Q_N(_0033_),
    .Q(\mem_addr[6] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[7]$_SDFFE_PN1P_  (.CLK(clknet_3_4_0_clk_buffered),
    .RESET_B(net303),
    .D(_0084_),
    .Q_N(_3053_),
    .Q(\mem_addr[7] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[8]$_SDFFE_PN1P_  (.CLK(clknet_3_1_0_clk_buffered),
    .RESET_B(net304),
    .D(_0085_),
    .Q_N(_3052_),
    .Q(\mem_addr[8] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[9]$_SDFFE_PN1P_  (.CLK(clknet_3_4_0_clk_buffered),
    .RESET_B(net305),
    .D(_0086_),
    .Q_N(_3051_),
    .Q(\memory_1.mem_addr[9] ));
 sg13g2_dfrbp_1 \transformer_1.started$_SDFFE_PN0P_  (.CLK(clknet_3_6_0_clk_buffered),
    .RESET_B(net306),
    .D(_0087_),
    .Q_N(_3050_),
    .Q(\transformer_1.started ));
 sg13g2_buf_1 input1 (.A(ui_in[5]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[6]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[7]),
    .X(net3));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[0]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[1]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[2]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[3]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[4]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[5]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[6]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_2 fanout18 (.A(_2301_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_2295_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_2198_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_2182_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0521_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0294_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_3023_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_2991_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_2968_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_2844_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_2774_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_2512_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_2416_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_2384_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0334_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0326_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0181_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0163_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0110_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_3022_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_2997_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_2990_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_2963_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_2905_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_2895_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_2795_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_2778_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_2753_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_2733_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_2684_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2680_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_2615_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_2593_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_2589_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_2583_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2569_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2533_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2510_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_2506_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2503_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2491_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_2475_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_2415_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_2408_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_2383_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_2375_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1107_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0532_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0338_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0161_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0090_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_2935_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_2882_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_2860_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_2826_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2785_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2782_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_2732_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_2729_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_2728_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_2716_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_2711_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_2699_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_2689_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_2673_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_2665_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_2654_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_2649_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_2628_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_2603_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_2568_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_2518_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_2513_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_2509_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_2505_),
    .X(net92));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(_2490_));
 sg13g2_buf_2 fanout94 (.A(_2487_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_2458_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_2452_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_2449_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_2435_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_2419_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_2413_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_2407_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_2402_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_2387_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_2382_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_2053_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_1838_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_1707_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1631_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1522_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1347_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0856_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0728_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0511_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0220_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0165_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_3040_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_2957_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_2816_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_2808_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_2769_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_2749_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_2704_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_2698_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_2688_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_2682_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_2669_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_2664_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_2653_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_2626_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_2601_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_2596_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_2566_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_2554_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_2552_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_2508_),
    .X(net135));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(_2495_));
 sg13g2_buf_2 fanout137 (.A(_2477_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_2445_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_2442_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_2437_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_2426_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_2418_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_2401_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_2399_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_2390_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_2386_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_2360_),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(_2257_));
 sg13g2_buf_2 fanout149 (.A(_2173_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_1696_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_1555_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_1511_),
    .X(net152));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(_1435_));
 sg13g2_buf_2 fanout154 (.A(_1020_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0976_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_0910_),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(_0845_));
 sg13g2_buf_2 fanout158 (.A(_0757_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_2296_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_0483_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_3039_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_2760_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_2738_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_2736_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_2696_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_2646_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_2619_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_2600_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_2595_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_2565_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_2544_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_2517_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_2480_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_2417_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_2351_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_2193_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_2162_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_1773_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_1751_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_1685_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_1588_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_1544_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_1424_),
    .X(net183));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(_1282_));
 sg13g2_buf_2 fanout185 (.A(_1260_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_1249_),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(_1009_));
 sg13g2_buf_2 fanout188 (.A(_0834_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_0790_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_0746_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_2281_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_1837_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_0602_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_0530_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_2695_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_2610_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_2557_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_2543_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_2516_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_2424_),
    .X(net200));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(_1848_));
 sg13g2_buf_2 fanout202 (.A(_1740_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_1380_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_1205_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_0998_),
    .X(net205));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(_0943_));
 sg13g2_buf_2 fanout207 (.A(_0889_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_0867_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_1369_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_1053_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_2179_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_1867_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_1850_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_1810_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_1808_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_1801_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_1798_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_1796_),
    .X(net218));
 sg13g2_tielo _6171__219 (.L_LO(net219));
 sg13g2_tielo _6172__220 (.L_LO(net220));
 sg13g2_tiehi _6164__222 (.L_HI(net222));
 sg13g2_tiehi _6165__223 (.L_HI(net223));
 sg13g2_tiehi _6166__224 (.L_HI(net224));
 sg13g2_tiehi _6167__225 (.L_HI(net225));
 sg13g2_tiehi _6168__226 (.L_HI(net226));
 sg13g2_tiehi _6169__227 (.L_HI(net227));
 sg13g2_tiehi _6170__228 (.L_HI(net228));
 sg13g2_tiehi \clk_picker.clk_slow$_SDFFE_PN0P__229  (.L_HI(net229));
 sg13g2_tiehi \clk_picker.counter[0]$_SDFF_PN0__230  (.L_HI(net230));
 sg13g2_tiehi \clk_picker.counter[10]$_SDFF_PN0__231  (.L_HI(net231));
 sg13g2_tiehi \clk_picker.counter[11]$_SDFF_PN0__232  (.L_HI(net232));
 sg13g2_tiehi \clk_picker.counter[12]$_SDFF_PN0__233  (.L_HI(net233));
 sg13g2_tiehi \clk_picker.counter[13]$_SDFF_PN0__234  (.L_HI(net234));
 sg13g2_tiehi \clk_picker.counter[14]$_SDFF_PN0__235  (.L_HI(net235));
 sg13g2_tiehi \clk_picker.counter[15]$_SDFF_PN0__236  (.L_HI(net236));
 sg13g2_tiehi \clk_picker.counter[16]$_SDFF_PN0__237  (.L_HI(net237));
 sg13g2_tiehi \clk_picker.counter[17]$_SDFF_PN0__238  (.L_HI(net238));
 sg13g2_tiehi \clk_picker.counter[18]$_SDFF_PN0__239  (.L_HI(net239));
 sg13g2_tiehi \clk_picker.counter[19]$_SDFF_PN0__240  (.L_HI(net240));
 sg13g2_tiehi \clk_picker.counter[1]$_SDFF_PN0__241  (.L_HI(net241));
 sg13g2_tiehi \clk_picker.counter[20]$_SDFF_PN0__242  (.L_HI(net242));
 sg13g2_tiehi \clk_picker.counter[21]$_SDFF_PN0__243  (.L_HI(net243));
 sg13g2_tiehi \clk_picker.counter[22]$_SDFF_PN0__244  (.L_HI(net244));
 sg13g2_tiehi \clk_picker.counter[23]$_SDFF_PN0__245  (.L_HI(net245));
 sg13g2_tiehi \clk_picker.counter[24]$_SDFF_PN0__246  (.L_HI(net246));
 sg13g2_tiehi \clk_picker.counter[25]$_SDFF_PN0__247  (.L_HI(net247));
 sg13g2_tiehi \clk_picker.counter[2]$_SDFF_PN0__248  (.L_HI(net248));
 sg13g2_tiehi \clk_picker.counter[3]$_SDFF_PN0__249  (.L_HI(net249));
 sg13g2_tiehi \clk_picker.counter[4]$_SDFF_PN0__250  (.L_HI(net250));
 sg13g2_tiehi \clk_picker.counter[5]$_SDFF_PN0__251  (.L_HI(net251));
 sg13g2_tiehi \clk_picker.counter[6]$_SDFF_PN0__252  (.L_HI(net252));
 sg13g2_tiehi \clk_picker.counter[7]$_SDFF_PN0__253  (.L_HI(net253));
 sg13g2_tiehi \clk_picker.counter[8]$_SDFF_PN0__254  (.L_HI(net254));
 sg13g2_tiehi \clk_picker.counter[9]$_SDFF_PN0__255  (.L_HI(net255));
 sg13g2_tiehi \line_mapper_1.pointer_addr[0]$_DFF_P__256  (.L_HI(net256));
 sg13g2_tiehi \line_mapper_1.pointer_addr[10]$_DFF_P__257  (.L_HI(net257));
 sg13g2_tiehi \line_mapper_1.pointer_addr[11]$_DFF_P__258  (.L_HI(net258));
 sg13g2_tiehi \line_mapper_1.pointer_addr[12]$_DFF_P__259  (.L_HI(net259));
 sg13g2_tiehi \line_mapper_1.pointer_addr[13]$_DFF_P__260  (.L_HI(net260));
 sg13g2_tiehi \line_mapper_1.pointer_addr[14]$_DFF_P__261  (.L_HI(net261));
 sg13g2_tiehi \line_mapper_1.pointer_addr[15]$_DFF_P__262  (.L_HI(net262));
 sg13g2_tiehi \line_mapper_1.pointer_addr[1]$_DFF_P__263  (.L_HI(net263));
 sg13g2_tiehi \line_mapper_1.pointer_addr[2]$_DFF_P__264  (.L_HI(net264));
 sg13g2_tiehi \line_mapper_1.pointer_addr[3]$_DFF_P__265  (.L_HI(net265));
 sg13g2_tiehi \line_mapper_1.pointer_addr[4]$_DFF_P__266  (.L_HI(net266));
 sg13g2_tiehi \line_mapper_1.pointer_addr[5]$_DFF_P__267  (.L_HI(net267));
 sg13g2_tiehi \line_mapper_1.pointer_addr[6]$_DFF_P__268  (.L_HI(net268));
 sg13g2_tiehi \line_mapper_1.pointer_addr[7]$_DFF_P__269  (.L_HI(net269));
 sg13g2_tiehi \line_mapper_1.pointer_addr[8]$_DFF_P__270  (.L_HI(net270));
 sg13g2_tiehi \line_mapper_1.pointer_addr[9]$_DFF_P__271  (.L_HI(net271));
 sg13g2_tiehi \memory_1.dout[0]$_DFF_P__272  (.L_HI(net272));
 sg13g2_tiehi \memory_1.dout[10]$_DFF_P__273  (.L_HI(net273));
 sg13g2_tiehi \memory_1.dout[11]$_DFF_P__274  (.L_HI(net274));
 sg13g2_tiehi \memory_1.dout[12]$_DFF_P__275  (.L_HI(net275));
 sg13g2_tiehi \memory_1.dout[13]$_DFF_P__276  (.L_HI(net276));
 sg13g2_tiehi \memory_1.dout[14]$_DFF_P__277  (.L_HI(net277));
 sg13g2_tiehi \memory_1.dout[1]$_DFF_P__278  (.L_HI(net278));
 sg13g2_tiehi \memory_1.dout[2]$_DFF_P__279  (.L_HI(net279));
 sg13g2_tiehi \memory_1.dout[3]$_DFF_P__280  (.L_HI(net280));
 sg13g2_tiehi \memory_1.dout[4]$_DFF_P__281  (.L_HI(net281));
 sg13g2_tiehi \memory_1.dout[5]$_DFF_P__282  (.L_HI(net282));
 sg13g2_tiehi \memory_1.dout[6]$_DFF_P__283  (.L_HI(net283));
 sg13g2_tiehi \memory_1.dout[8]$_DFF_P__284  (.L_HI(net284));
 sg13g2_tiehi \memory_1.dout[9]$_DFF_P__285  (.L_HI(net285));
 sg13g2_tiehi \transformer_1.chars_remaining[0]$_SDFFE_PN0P__286  (.L_HI(net286));
 sg13g2_tiehi \transformer_1.chars_remaining[1]$_SDFFE_PN0P__287  (.L_HI(net287));
 sg13g2_tiehi \transformer_1.chars_remaining[2]$_SDFFE_PN0P__288  (.L_HI(net288));
 sg13g2_tiehi \transformer_1.chars_remaining[3]$_SDFFE_PN0P__289  (.L_HI(net289));
 sg13g2_tiehi \transformer_1.chars_remaining[4]$_SDFFE_PN0P__290  (.L_HI(net290));
 sg13g2_tiehi \transformer_1.chars_remaining[5]$_SDFFE_PN0P__291  (.L_HI(net291));
 sg13g2_tiehi \transformer_1.chars_remaining[6]$_SDFFE_PN0P__292  (.L_HI(net292));
 sg13g2_tiehi \transformer_1.chars_remaining[7]$_SDFFE_PN0P__293  (.L_HI(net293));
 sg13g2_tiehi \transformer_1.chars_remaining[8]$_SDFFE_PN0P__294  (.L_HI(net294));
 sg13g2_tiehi \transformer_1.chars_remaining[9]$_SDFFE_PN0P__295  (.L_HI(net295));
 sg13g2_tiehi \transformer_1.mem_addr[0]$_SDFFE_PN1P__296  (.L_HI(net296));
 sg13g2_tiehi \transformer_1.mem_addr[1]$_SDFFE_PN1P__297  (.L_HI(net297));
 sg13g2_tiehi \transformer_1.mem_addr[2]$_SDFFE_PN1P__298  (.L_HI(net298));
 sg13g2_tiehi \transformer_1.mem_addr[3]$_SDFFE_PN1P__299  (.L_HI(net299));
 sg13g2_tiehi \transformer_1.mem_addr[4]$_SDFFE_PN1P__300  (.L_HI(net300));
 sg13g2_tiehi \transformer_1.mem_addr[5]$_SDFFE_PN1P__301  (.L_HI(net301));
 sg13g2_tiehi \transformer_1.mem_addr[6]$_SDFFE_PN1P__302  (.L_HI(net302));
 sg13g2_tiehi \transformer_1.mem_addr[7]$_SDFFE_PN1P__303  (.L_HI(net303));
 sg13g2_tiehi \transformer_1.mem_addr[8]$_SDFFE_PN1P__304  (.L_HI(net304));
 sg13g2_tiehi \transformer_1.mem_addr[9]$_SDFFE_PN1P__305  (.L_HI(net305));
 sg13g2_tiehi \transformer_1.started$_SDFFE_PN0P__306  (.L_HI(net306));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_buf_4 clkbuf_level_0_1_10_clk (.X(clknet_level_0_1_10_clk),
    .A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkbuf_level_1_1_11_clk (.X(clknet_level_1_1_11_clk),
    .A(clknet_level_0_1_10_clk));
 sg13g2_buf_4 clkbuf_level_2_1_12_clk (.X(clknet_level_2_1_12_clk),
    .A(clknet_level_1_1_11_clk));
 sg13g2_buf_4 clkbuf_level_0_1_23_clk (.X(clknet_level_0_1_23_clk),
    .A(clknet_2_1__leaf_clk));
 sg13g2_buf_4 clkbuf_level_1_1_24_clk (.X(clknet_level_1_1_24_clk),
    .A(clknet_level_0_1_23_clk));
 sg13g2_buf_4 clkbuf_level_2_1_25_clk (.X(clknet_level_2_1_25_clk),
    .A(clknet_level_1_1_24_clk));
 sg13g2_buf_4 clkbuf_level_0_1_36_clk (.X(clknet_level_0_1_36_clk),
    .A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkbuf_level_1_1_37_clk (.X(clknet_level_1_1_37_clk),
    .A(clknet_level_0_1_36_clk));
 sg13g2_buf_4 clkbuf_level_2_1_38_clk (.X(clknet_level_2_1_38_clk),
    .A(clknet_level_1_1_37_clk));
 sg13g2_buf_4 clkbuf_level_0_1_49_clk (.X(clknet_level_0_1_49_clk),
    .A(clknet_2_3__leaf_clk));
 sg13g2_buf_4 clkbuf_level_1_1_410_clk (.X(clknet_level_1_1_410_clk),
    .A(clknet_level_0_1_49_clk));
 sg13g2_buf_4 clkbuf_level_2_1_411_clk (.X(clknet_level_2_1_411_clk),
    .A(clknet_level_1_1_410_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_2_3__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_buffered (.A(clk_buffered),
    .X(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_0_0_clk_buffered (.X(clknet_3_0_0_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_1_0_clk_buffered (.X(clknet_3_1_0_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_2_0_clk_buffered (.X(clknet_3_2_0_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_3_0_clk_buffered (.X(clknet_3_3_0_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_4_0_clk_buffered (.X(clknet_3_4_0_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_5_0_clk_buffered (.X(clknet_3_5_0_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_6_0_clk_buffered (.X(clknet_3_6_0_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_7_0_clk_buffered (.X(clknet_3_7_0_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_inv_1 clkload3 (.A(clknet_3_1_0_clk_buffered));
 sg13g2_inv_1 clkload4 (.A(clknet_3_3_0_clk_buffered));
 sg13g2_inv_1 clkload5 (.A(clknet_3_5_0_clk_buffered));
 sg13g2_inv_1 clkload6 (.A(clknet_3_6_0_clk_buffered));
 sg13g2_inv_1 clkload7 (.A(clknet_3_7_0_clk_buffered));
 sg13g2_antennanp ANTENNA_1 (.A(_0019_));
 sg13g2_antennanp ANTENNA_2 (.A(_0020_));
 sg13g2_antennanp ANTENNA_3 (.A(_0025_));
 sg13g2_antennanp ANTENNA_4 (.A(_0272_));
 sg13g2_antennanp ANTENNA_5 (.A(_0278_));
 sg13g2_antennanp ANTENNA_6 (.A(_0278_));
 sg13g2_antennanp ANTENNA_7 (.A(_0278_));
 sg13g2_antennanp ANTENNA_8 (.A(_0334_));
 sg13g2_antennanp ANTENNA_9 (.A(_0334_));
 sg13g2_antennanp ANTENNA_10 (.A(_0334_));
 sg13g2_antennanp ANTENNA_11 (.A(_0334_));
 sg13g2_antennanp ANTENNA_12 (.A(_0474_));
 sg13g2_antennanp ANTENNA_13 (.A(_0915_));
 sg13g2_antennanp ANTENNA_14 (.A(_0915_));
 sg13g2_antennanp ANTENNA_15 (.A(_0915_));
 sg13g2_antennanp ANTENNA_16 (.A(_1697_));
 sg13g2_antennanp ANTENNA_17 (.A(_1697_));
 sg13g2_antennanp ANTENNA_18 (.A(_1697_));
 sg13g2_antennanp ANTENNA_19 (.A(_2797_));
 sg13g2_antennanp ANTENNA_20 (.A(_2797_));
 sg13g2_antennanp ANTENNA_21 (.A(_2797_));
 sg13g2_antennanp ANTENNA_22 (.A(_2797_));
 sg13g2_antennanp ANTENNA_23 (.A(_2797_));
 sg13g2_antennanp ANTENNA_24 (.A(_2797_));
 sg13g2_antennanp ANTENNA_25 (.A(_2797_));
 sg13g2_antennanp ANTENNA_26 (.A(_2797_));
 sg13g2_antennanp ANTENNA_27 (.A(_2797_));
 sg13g2_antennanp ANTENNA_28 (.A(_2797_));
 sg13g2_antennanp ANTENNA_29 (.A(_2797_));
 sg13g2_antennanp ANTENNA_30 (.A(_0019_));
 sg13g2_antennanp ANTENNA_31 (.A(_0019_));
 sg13g2_antennanp ANTENNA_32 (.A(_0025_));
 sg13g2_antennanp ANTENNA_33 (.A(_0025_));
 sg13g2_antennanp ANTENNA_34 (.A(_0272_));
 sg13g2_antennanp ANTENNA_35 (.A(_0915_));
 sg13g2_antennanp ANTENNA_36 (.A(_0915_));
 sg13g2_antennanp ANTENNA_37 (.A(_0915_));
 sg13g2_antennanp ANTENNA_38 (.A(_1697_));
 sg13g2_antennanp ANTENNA_39 (.A(_1697_));
 sg13g2_antennanp ANTENNA_40 (.A(_2797_));
 sg13g2_antennanp ANTENNA_41 (.A(_2797_));
 sg13g2_antennanp ANTENNA_42 (.A(_2797_));
 sg13g2_antennanp ANTENNA_43 (.A(_2797_));
 sg13g2_antennanp ANTENNA_44 (.A(_2797_));
 sg13g2_antennanp ANTENNA_45 (.A(_2797_));
 sg13g2_antennanp ANTENNA_46 (.A(_2797_));
 sg13g2_antennanp ANTENNA_47 (.A(_2797_));
 sg13g2_antennanp ANTENNA_48 (.A(_2797_));
 sg13g2_antennanp ANTENNA_49 (.A(_2797_));
 sg13g2_antennanp ANTENNA_50 (.A(_2797_));
 sg13g2_antennanp ANTENNA_51 (.A(_0019_));
 sg13g2_antennanp ANTENNA_52 (.A(_0019_));
 sg13g2_antennanp ANTENNA_53 (.A(_0272_));
 sg13g2_antennanp ANTENNA_54 (.A(_0915_));
 sg13g2_antennanp ANTENNA_55 (.A(_0915_));
 sg13g2_antennanp ANTENNA_56 (.A(_0915_));
 sg13g2_antennanp ANTENNA_57 (.A(_1697_));
 sg13g2_antennanp ANTENNA_58 (.A(_1697_));
 sg13g2_antennanp ANTENNA_59 (.A(_2797_));
 sg13g2_antennanp ANTENNA_60 (.A(_2797_));
 sg13g2_antennanp ANTENNA_61 (.A(_2797_));
 sg13g2_antennanp ANTENNA_62 (.A(_2797_));
 sg13g2_antennanp ANTENNA_63 (.A(_2797_));
 sg13g2_antennanp ANTENNA_64 (.A(_2797_));
 sg13g2_antennanp ANTENNA_65 (.A(_2797_));
 sg13g2_antennanp ANTENNA_66 (.A(_2797_));
 sg13g2_antennanp ANTENNA_67 (.A(_2797_));
 sg13g2_antennanp ANTENNA_68 (.A(_2797_));
 sg13g2_antennanp ANTENNA_69 (.A(_2797_));
 sg13g2_antennanp ANTENNA_70 (.A(_0019_));
 sg13g2_antennanp ANTENNA_71 (.A(_0019_));
 sg13g2_antennanp ANTENNA_72 (.A(_0272_));
 sg13g2_antennanp ANTENNA_73 (.A(_0915_));
 sg13g2_antennanp ANTENNA_74 (.A(_0915_));
 sg13g2_antennanp ANTENNA_75 (.A(_0915_));
 sg13g2_antennanp ANTENNA_76 (.A(_1697_));
 sg13g2_antennanp ANTENNA_77 (.A(_1697_));
 sg13g2_antennanp ANTENNA_78 (.A(_2797_));
 sg13g2_antennanp ANTENNA_79 (.A(_2797_));
 sg13g2_antennanp ANTENNA_80 (.A(_2797_));
 sg13g2_antennanp ANTENNA_81 (.A(_2797_));
 sg13g2_antennanp ANTENNA_82 (.A(_2797_));
 sg13g2_antennanp ANTENNA_83 (.A(_2797_));
 sg13g2_antennanp ANTENNA_84 (.A(_2797_));
 sg13g2_antennanp ANTENNA_85 (.A(_2797_));
 sg13g2_antennanp ANTENNA_86 (.A(_2797_));
 sg13g2_antennanp ANTENNA_87 (.A(_2797_));
 sg13g2_antennanp ANTENNA_88 (.A(_2797_));
 sg13g2_antennanp ANTENNA_89 (.A(_0019_));
 sg13g2_antennanp ANTENNA_90 (.A(_0019_));
 sg13g2_antennanp ANTENNA_91 (.A(_0272_));
 sg13g2_antennanp ANTENNA_92 (.A(_1697_));
 sg13g2_antennanp ANTENNA_93 (.A(_1697_));
 sg13g2_antennanp ANTENNA_94 (.A(_2797_));
 sg13g2_antennanp ANTENNA_95 (.A(_2797_));
 sg13g2_antennanp ANTENNA_96 (.A(_2797_));
 sg13g2_antennanp ANTENNA_97 (.A(_2797_));
 sg13g2_antennanp ANTENNA_98 (.A(_2797_));
 sg13g2_antennanp ANTENNA_99 (.A(_2797_));
 sg13g2_antennanp ANTENNA_100 (.A(_2797_));
 sg13g2_antennanp ANTENNA_101 (.A(_2797_));
 sg13g2_antennanp ANTENNA_102 (.A(_2797_));
 sg13g2_antennanp ANTENNA_103 (.A(_2797_));
 sg13g2_antennanp ANTENNA_104 (.A(_2797_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_fill_2 FILLER_0_875 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_fill_2 FILLER_1_875 ();
 sg13g2_fill_1 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_fill_2 FILLER_2_875 ();
 sg13g2_fill_1 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_fill_2 FILLER_3_875 ();
 sg13g2_fill_1 FILLER_3_877 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_fill_2 FILLER_4_875 ();
 sg13g2_fill_1 FILLER_4_877 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_decap_8 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_5_868 ();
 sg13g2_fill_2 FILLER_5_875 ();
 sg13g2_fill_1 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_decap_8 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_6_868 ();
 sg13g2_fill_2 FILLER_6_875 ();
 sg13g2_fill_1 FILLER_6_877 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_fill_2 FILLER_7_875 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_fill_2 FILLER_8_875 ();
 sg13g2_fill_1 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_fill_2 FILLER_9_875 ();
 sg13g2_fill_1 FILLER_9_877 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_868 ();
 sg13g2_fill_2 FILLER_10_875 ();
 sg13g2_fill_1 FILLER_10_877 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_566 ();
 sg13g2_decap_8 FILLER_11_573 ();
 sg13g2_decap_8 FILLER_11_593 ();
 sg13g2_decap_8 FILLER_11_600 ();
 sg13g2_decap_8 FILLER_11_607 ();
 sg13g2_fill_1 FILLER_11_614 ();
 sg13g2_decap_8 FILLER_11_628 ();
 sg13g2_decap_8 FILLER_11_635 ();
 sg13g2_decap_8 FILLER_11_642 ();
 sg13g2_decap_8 FILLER_11_649 ();
 sg13g2_decap_8 FILLER_11_656 ();
 sg13g2_decap_8 FILLER_11_663 ();
 sg13g2_decap_8 FILLER_11_670 ();
 sg13g2_decap_8 FILLER_11_677 ();
 sg13g2_decap_8 FILLER_11_684 ();
 sg13g2_decap_8 FILLER_11_691 ();
 sg13g2_decap_8 FILLER_11_698 ();
 sg13g2_decap_8 FILLER_11_705 ();
 sg13g2_decap_8 FILLER_11_712 ();
 sg13g2_decap_8 FILLER_11_719 ();
 sg13g2_decap_8 FILLER_11_726 ();
 sg13g2_decap_8 FILLER_11_733 ();
 sg13g2_decap_8 FILLER_11_740 ();
 sg13g2_decap_8 FILLER_11_747 ();
 sg13g2_decap_8 FILLER_11_754 ();
 sg13g2_decap_8 FILLER_11_761 ();
 sg13g2_decap_8 FILLER_11_768 ();
 sg13g2_decap_8 FILLER_11_775 ();
 sg13g2_decap_8 FILLER_11_782 ();
 sg13g2_decap_8 FILLER_11_789 ();
 sg13g2_decap_8 FILLER_11_796 ();
 sg13g2_decap_8 FILLER_11_803 ();
 sg13g2_decap_8 FILLER_11_810 ();
 sg13g2_decap_8 FILLER_11_817 ();
 sg13g2_decap_8 FILLER_11_824 ();
 sg13g2_decap_8 FILLER_11_831 ();
 sg13g2_decap_8 FILLER_11_838 ();
 sg13g2_decap_8 FILLER_11_845 ();
 sg13g2_decap_8 FILLER_11_852 ();
 sg13g2_decap_8 FILLER_11_859 ();
 sg13g2_decap_8 FILLER_11_866 ();
 sg13g2_decap_4 FILLER_11_873 ();
 sg13g2_fill_1 FILLER_11_877 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_fill_1 FILLER_12_392 ();
 sg13g2_fill_1 FILLER_12_432 ();
 sg13g2_decap_8 FILLER_12_446 ();
 sg13g2_decap_8 FILLER_12_453 ();
 sg13g2_decap_8 FILLER_12_460 ();
 sg13g2_decap_8 FILLER_12_467 ();
 sg13g2_fill_1 FILLER_12_474 ();
 sg13g2_decap_4 FILLER_12_488 ();
 sg13g2_fill_1 FILLER_12_492 ();
 sg13g2_decap_8 FILLER_12_510 ();
 sg13g2_decap_8 FILLER_12_517 ();
 sg13g2_decap_8 FILLER_12_524 ();
 sg13g2_decap_4 FILLER_12_531 ();
 sg13g2_fill_1 FILLER_12_535 ();
 sg13g2_decap_8 FILLER_12_541 ();
 sg13g2_fill_2 FILLER_12_548 ();
 sg13g2_decap_8 FILLER_12_562 ();
 sg13g2_decap_4 FILLER_12_569 ();
 sg13g2_fill_1 FILLER_12_573 ();
 sg13g2_decap_8 FILLER_12_579 ();
 sg13g2_decap_8 FILLER_12_586 ();
 sg13g2_decap_8 FILLER_12_593 ();
 sg13g2_decap_8 FILLER_12_600 ();
 sg13g2_decap_8 FILLER_12_620 ();
 sg13g2_decap_4 FILLER_12_627 ();
 sg13g2_fill_1 FILLER_12_631 ();
 sg13g2_decap_4 FILLER_12_645 ();
 sg13g2_fill_1 FILLER_12_649 ();
 sg13g2_decap_8 FILLER_12_654 ();
 sg13g2_decap_8 FILLER_12_661 ();
 sg13g2_decap_8 FILLER_12_668 ();
 sg13g2_decap_8 FILLER_12_675 ();
 sg13g2_fill_2 FILLER_12_682 ();
 sg13g2_fill_1 FILLER_12_684 ();
 sg13g2_fill_2 FILLER_12_702 ();
 sg13g2_fill_1 FILLER_12_708 ();
 sg13g2_decap_8 FILLER_12_722 ();
 sg13g2_decap_8 FILLER_12_729 ();
 sg13g2_decap_8 FILLER_12_736 ();
 sg13g2_decap_8 FILLER_12_743 ();
 sg13g2_decap_8 FILLER_12_750 ();
 sg13g2_decap_8 FILLER_12_757 ();
 sg13g2_decap_8 FILLER_12_764 ();
 sg13g2_decap_8 FILLER_12_771 ();
 sg13g2_decap_8 FILLER_12_778 ();
 sg13g2_decap_8 FILLER_12_785 ();
 sg13g2_decap_8 FILLER_12_792 ();
 sg13g2_decap_8 FILLER_12_799 ();
 sg13g2_decap_8 FILLER_12_806 ();
 sg13g2_decap_8 FILLER_12_813 ();
 sg13g2_decap_8 FILLER_12_820 ();
 sg13g2_decap_8 FILLER_12_827 ();
 sg13g2_decap_8 FILLER_12_834 ();
 sg13g2_decap_8 FILLER_12_841 ();
 sg13g2_decap_8 FILLER_12_848 ();
 sg13g2_decap_8 FILLER_12_855 ();
 sg13g2_decap_8 FILLER_12_862 ();
 sg13g2_decap_8 FILLER_12_869 ();
 sg13g2_fill_2 FILLER_12_876 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_4 FILLER_13_441 ();
 sg13g2_fill_2 FILLER_13_445 ();
 sg13g2_decap_8 FILLER_13_464 ();
 sg13g2_decap_8 FILLER_13_471 ();
 sg13g2_decap_8 FILLER_13_478 ();
 sg13g2_decap_8 FILLER_13_485 ();
 sg13g2_decap_8 FILLER_13_492 ();
 sg13g2_decap_8 FILLER_13_499 ();
 sg13g2_decap_4 FILLER_13_506 ();
 sg13g2_decap_8 FILLER_13_515 ();
 sg13g2_decap_4 FILLER_13_522 ();
 sg13g2_decap_4 FILLER_13_531 ();
 sg13g2_decap_4 FILLER_13_540 ();
 sg13g2_fill_1 FILLER_13_544 ();
 sg13g2_fill_2 FILLER_13_549 ();
 sg13g2_decap_8 FILLER_13_563 ();
 sg13g2_decap_8 FILLER_13_570 ();
 sg13g2_decap_8 FILLER_13_577 ();
 sg13g2_decap_8 FILLER_13_584 ();
 sg13g2_decap_8 FILLER_13_591 ();
 sg13g2_decap_8 FILLER_13_598 ();
 sg13g2_decap_4 FILLER_13_605 ();
 sg13g2_fill_1 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_614 ();
 sg13g2_fill_1 FILLER_13_621 ();
 sg13g2_decap_8 FILLER_13_635 ();
 sg13g2_fill_2 FILLER_13_642 ();
 sg13g2_decap_8 FILLER_13_649 ();
 sg13g2_decap_8 FILLER_13_656 ();
 sg13g2_decap_8 FILLER_13_663 ();
 sg13g2_decap_8 FILLER_13_670 ();
 sg13g2_decap_8 FILLER_13_677 ();
 sg13g2_decap_8 FILLER_13_684 ();
 sg13g2_fill_2 FILLER_13_691 ();
 sg13g2_fill_1 FILLER_13_693 ();
 sg13g2_fill_2 FILLER_13_712 ();
 sg13g2_fill_2 FILLER_13_719 ();
 sg13g2_decap_8 FILLER_13_751 ();
 sg13g2_decap_8 FILLER_13_758 ();
 sg13g2_decap_8 FILLER_13_765 ();
 sg13g2_decap_8 FILLER_13_772 ();
 sg13g2_decap_8 FILLER_13_779 ();
 sg13g2_decap_8 FILLER_13_786 ();
 sg13g2_decap_8 FILLER_13_793 ();
 sg13g2_decap_8 FILLER_13_800 ();
 sg13g2_decap_8 FILLER_13_807 ();
 sg13g2_decap_8 FILLER_13_814 ();
 sg13g2_decap_8 FILLER_13_821 ();
 sg13g2_decap_8 FILLER_13_828 ();
 sg13g2_decap_8 FILLER_13_835 ();
 sg13g2_decap_8 FILLER_13_842 ();
 sg13g2_decap_8 FILLER_13_849 ();
 sg13g2_decap_8 FILLER_13_856 ();
 sg13g2_decap_8 FILLER_13_863 ();
 sg13g2_decap_8 FILLER_13_870 ();
 sg13g2_fill_1 FILLER_13_877 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_4 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_4 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_4 FILLER_14_359 ();
 sg13g2_fill_1 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_fill_1 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_fill_1 FILLER_14_391 ();
 sg13g2_fill_1 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_401 ();
 sg13g2_fill_2 FILLER_14_405 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_fill_1 FILLER_14_430 ();
 sg13g2_decap_8 FILLER_14_437 ();
 sg13g2_decap_8 FILLER_14_449 ();
 sg13g2_fill_1 FILLER_14_456 ();
 sg13g2_decap_8 FILLER_14_465 ();
 sg13g2_decap_8 FILLER_14_472 ();
 sg13g2_decap_8 FILLER_14_479 ();
 sg13g2_decap_8 FILLER_14_486 ();
 sg13g2_decap_8 FILLER_14_493 ();
 sg13g2_decap_8 FILLER_14_500 ();
 sg13g2_decap_8 FILLER_14_507 ();
 sg13g2_decap_8 FILLER_14_514 ();
 sg13g2_decap_4 FILLER_14_521 ();
 sg13g2_decap_8 FILLER_14_530 ();
 sg13g2_decap_4 FILLER_14_537 ();
 sg13g2_fill_1 FILLER_14_541 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_579 ();
 sg13g2_decap_8 FILLER_14_586 ();
 sg13g2_decap_8 FILLER_14_593 ();
 sg13g2_decap_8 FILLER_14_600 ();
 sg13g2_decap_8 FILLER_14_607 ();
 sg13g2_decap_4 FILLER_14_614 ();
 sg13g2_fill_2 FILLER_14_618 ();
 sg13g2_fill_1 FILLER_14_625 ();
 sg13g2_decap_8 FILLER_14_639 ();
 sg13g2_decap_8 FILLER_14_646 ();
 sg13g2_fill_2 FILLER_14_653 ();
 sg13g2_fill_1 FILLER_14_655 ();
 sg13g2_decap_8 FILLER_14_669 ();
 sg13g2_decap_8 FILLER_14_676 ();
 sg13g2_decap_8 FILLER_14_683 ();
 sg13g2_decap_8 FILLER_14_690 ();
 sg13g2_decap_8 FILLER_14_697 ();
 sg13g2_decap_4 FILLER_14_704 ();
 sg13g2_decap_4 FILLER_14_714 ();
 sg13g2_fill_2 FILLER_14_718 ();
 sg13g2_decap_8 FILLER_14_724 ();
 sg13g2_decap_8 FILLER_14_737 ();
 sg13g2_decap_8 FILLER_14_744 ();
 sg13g2_decap_8 FILLER_14_751 ();
 sg13g2_decap_8 FILLER_14_758 ();
 sg13g2_decap_8 FILLER_14_765 ();
 sg13g2_decap_8 FILLER_14_772 ();
 sg13g2_decap_8 FILLER_14_779 ();
 sg13g2_decap_8 FILLER_14_786 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_800 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_decap_8 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_821 ();
 sg13g2_decap_8 FILLER_14_828 ();
 sg13g2_decap_8 FILLER_14_835 ();
 sg13g2_decap_8 FILLER_14_842 ();
 sg13g2_decap_8 FILLER_14_849 ();
 sg13g2_decap_8 FILLER_14_856 ();
 sg13g2_decap_8 FILLER_14_863 ();
 sg13g2_decap_8 FILLER_14_870 ();
 sg13g2_fill_1 FILLER_14_877 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_202 ();
 sg13g2_decap_8 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_216 ();
 sg13g2_decap_8 FILLER_15_223 ();
 sg13g2_decap_4 FILLER_15_230 ();
 sg13g2_fill_1 FILLER_15_234 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_4 FILLER_15_259 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_decap_4 FILLER_15_276 ();
 sg13g2_fill_2 FILLER_15_280 ();
 sg13g2_decap_4 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_292 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_decap_4 FILLER_15_320 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_fill_2 FILLER_15_339 ();
 sg13g2_fill_1 FILLER_15_341 ();
 sg13g2_decap_4 FILLER_15_350 ();
 sg13g2_fill_1 FILLER_15_362 ();
 sg13g2_decap_4 FILLER_15_367 ();
 sg13g2_fill_2 FILLER_15_371 ();
 sg13g2_fill_2 FILLER_15_377 ();
 sg13g2_fill_1 FILLER_15_379 ();
 sg13g2_decap_4 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_fill_1 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_430 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_decap_4 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_474 ();
 sg13g2_decap_8 FILLER_15_481 ();
 sg13g2_fill_2 FILLER_15_488 ();
 sg13g2_fill_1 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_500 ();
 sg13g2_decap_8 FILLER_15_507 ();
 sg13g2_fill_2 FILLER_15_514 ();
 sg13g2_fill_1 FILLER_15_516 ();
 sg13g2_decap_4 FILLER_15_522 ();
 sg13g2_fill_1 FILLER_15_526 ();
 sg13g2_decap_4 FILLER_15_532 ();
 sg13g2_decap_4 FILLER_15_541 ();
 sg13g2_fill_2 FILLER_15_545 ();
 sg13g2_decap_8 FILLER_15_551 ();
 sg13g2_decap_8 FILLER_15_558 ();
 sg13g2_decap_8 FILLER_15_565 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_decap_8 FILLER_15_613 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_4 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_636 ();
 sg13g2_fill_2 FILLER_15_643 ();
 sg13g2_fill_2 FILLER_15_649 ();
 sg13g2_fill_1 FILLER_15_660 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_4 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_681 ();
 sg13g2_decap_8 FILLER_15_688 ();
 sg13g2_decap_4 FILLER_15_695 ();
 sg13g2_fill_2 FILLER_15_699 ();
 sg13g2_fill_1 FILLER_15_719 ();
 sg13g2_fill_1 FILLER_15_724 ();
 sg13g2_fill_2 FILLER_15_729 ();
 sg13g2_fill_1 FILLER_15_731 ();
 sg13g2_decap_8 FILLER_15_745 ();
 sg13g2_decap_8 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_759 ();
 sg13g2_decap_8 FILLER_15_766 ();
 sg13g2_decap_8 FILLER_15_773 ();
 sg13g2_decap_8 FILLER_15_780 ();
 sg13g2_decap_8 FILLER_15_787 ();
 sg13g2_decap_8 FILLER_15_794 ();
 sg13g2_decap_8 FILLER_15_801 ();
 sg13g2_decap_8 FILLER_15_808 ();
 sg13g2_decap_8 FILLER_15_815 ();
 sg13g2_decap_8 FILLER_15_822 ();
 sg13g2_decap_8 FILLER_15_829 ();
 sg13g2_decap_8 FILLER_15_836 ();
 sg13g2_decap_8 FILLER_15_843 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_decap_8 FILLER_15_857 ();
 sg13g2_decap_8 FILLER_15_864 ();
 sg13g2_decap_8 FILLER_15_871 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_4 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_169 ();
 sg13g2_decap_8 FILLER_16_176 ();
 sg13g2_decap_8 FILLER_16_183 ();
 sg13g2_decap_8 FILLER_16_190 ();
 sg13g2_decap_8 FILLER_16_197 ();
 sg13g2_decap_8 FILLER_16_204 ();
 sg13g2_fill_2 FILLER_16_211 ();
 sg13g2_decap_4 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_225 ();
 sg13g2_fill_2 FILLER_16_232 ();
 sg13g2_decap_8 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_decap_4 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_fill_2 FILLER_16_300 ();
 sg13g2_fill_1 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_4 FILLER_16_325 ();
 sg13g2_fill_2 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_4 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_4 FILLER_16_387 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_fill_1 FILLER_16_399 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_2 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_16_415 ();
 sg13g2_fill_1 FILLER_16_419 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_531 ();
 sg13g2_decap_4 FILLER_16_538 ();
 sg13g2_fill_2 FILLER_16_542 ();
 sg13g2_fill_2 FILLER_16_549 ();
 sg13g2_fill_1 FILLER_16_551 ();
 sg13g2_decap_8 FILLER_16_556 ();
 sg13g2_decap_8 FILLER_16_563 ();
 sg13g2_decap_8 FILLER_16_570 ();
 sg13g2_fill_1 FILLER_16_577 ();
 sg13g2_decap_4 FILLER_16_588 ();
 sg13g2_fill_2 FILLER_16_597 ();
 sg13g2_fill_1 FILLER_16_599 ();
 sg13g2_decap_8 FILLER_16_604 ();
 sg13g2_decap_8 FILLER_16_611 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_fill_2 FILLER_16_630 ();
 sg13g2_fill_1 FILLER_16_632 ();
 sg13g2_fill_2 FILLER_16_641 ();
 sg13g2_decap_8 FILLER_16_647 ();
 sg13g2_decap_8 FILLER_16_654 ();
 sg13g2_decap_8 FILLER_16_661 ();
 sg13g2_fill_1 FILLER_16_668 ();
 sg13g2_fill_1 FILLER_16_674 ();
 sg13g2_decap_8 FILLER_16_684 ();
 sg13g2_decap_8 FILLER_16_691 ();
 sg13g2_decap_8 FILLER_16_698 ();
 sg13g2_decap_4 FILLER_16_705 ();
 sg13g2_fill_2 FILLER_16_709 ();
 sg13g2_fill_2 FILLER_16_721 ();
 sg13g2_fill_1 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_decap_8 FILLER_16_753 ();
 sg13g2_decap_8 FILLER_16_760 ();
 sg13g2_decap_8 FILLER_16_767 ();
 sg13g2_decap_8 FILLER_16_774 ();
 sg13g2_decap_8 FILLER_16_781 ();
 sg13g2_decap_8 FILLER_16_788 ();
 sg13g2_decap_8 FILLER_16_795 ();
 sg13g2_decap_8 FILLER_16_802 ();
 sg13g2_decap_8 FILLER_16_809 ();
 sg13g2_decap_8 FILLER_16_816 ();
 sg13g2_decap_8 FILLER_16_823 ();
 sg13g2_decap_8 FILLER_16_830 ();
 sg13g2_decap_8 FILLER_16_837 ();
 sg13g2_decap_8 FILLER_16_844 ();
 sg13g2_decap_8 FILLER_16_851 ();
 sg13g2_decap_8 FILLER_16_858 ();
 sg13g2_decap_8 FILLER_16_865 ();
 sg13g2_decap_4 FILLER_16_872 ();
 sg13g2_fill_2 FILLER_16_876 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_163 ();
 sg13g2_decap_8 FILLER_17_169 ();
 sg13g2_decap_8 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_192 ();
 sg13g2_fill_2 FILLER_17_199 ();
 sg13g2_decap_4 FILLER_17_205 ();
 sg13g2_decap_8 FILLER_17_213 ();
 sg13g2_fill_2 FILLER_17_220 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_decap_8 FILLER_17_242 ();
 sg13g2_decap_8 FILLER_17_249 ();
 sg13g2_decap_4 FILLER_17_256 ();
 sg13g2_fill_1 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_decap_4 FILLER_17_278 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_4 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_302 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_315 ();
 sg13g2_fill_1 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_fill_2 FILLER_17_329 ();
 sg13g2_fill_1 FILLER_17_331 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_4 FILLER_17_392 ();
 sg13g2_fill_2 FILLER_17_396 ();
 sg13g2_decap_8 FILLER_17_412 ();
 sg13g2_decap_8 FILLER_17_419 ();
 sg13g2_fill_1 FILLER_17_426 ();
 sg13g2_fill_1 FILLER_17_433 ();
 sg13g2_decap_8 FILLER_17_438 ();
 sg13g2_decap_8 FILLER_17_445 ();
 sg13g2_decap_8 FILLER_17_452 ();
 sg13g2_fill_1 FILLER_17_459 ();
 sg13g2_decap_4 FILLER_17_464 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_fill_1 FILLER_17_497 ();
 sg13g2_fill_1 FILLER_17_506 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_fill_2 FILLER_17_539 ();
 sg13g2_decap_4 FILLER_17_545 ();
 sg13g2_fill_2 FILLER_17_549 ();
 sg13g2_decap_8 FILLER_17_556 ();
 sg13g2_decap_8 FILLER_17_563 ();
 sg13g2_decap_8 FILLER_17_570 ();
 sg13g2_fill_2 FILLER_17_577 ();
 sg13g2_decap_4 FILLER_17_584 ();
 sg13g2_decap_8 FILLER_17_592 ();
 sg13g2_decap_8 FILLER_17_605 ();
 sg13g2_decap_8 FILLER_17_612 ();
 sg13g2_decap_8 FILLER_17_619 ();
 sg13g2_decap_8 FILLER_17_626 ();
 sg13g2_decap_8 FILLER_17_642 ();
 sg13g2_decap_8 FILLER_17_649 ();
 sg13g2_decap_8 FILLER_17_656 ();
 sg13g2_decap_4 FILLER_17_663 ();
 sg13g2_fill_1 FILLER_17_667 ();
 sg13g2_decap_4 FILLER_17_677 ();
 sg13g2_decap_8 FILLER_17_685 ();
 sg13g2_decap_8 FILLER_17_692 ();
 sg13g2_decap_8 FILLER_17_699 ();
 sg13g2_decap_8 FILLER_17_706 ();
 sg13g2_fill_2 FILLER_17_713 ();
 sg13g2_fill_1 FILLER_17_715 ();
 sg13g2_fill_1 FILLER_17_731 ();
 sg13g2_decap_8 FILLER_17_736 ();
 sg13g2_decap_8 FILLER_17_743 ();
 sg13g2_decap_8 FILLER_17_750 ();
 sg13g2_decap_8 FILLER_17_757 ();
 sg13g2_decap_8 FILLER_17_764 ();
 sg13g2_decap_8 FILLER_17_771 ();
 sg13g2_decap_8 FILLER_17_778 ();
 sg13g2_decap_8 FILLER_17_785 ();
 sg13g2_decap_8 FILLER_17_792 ();
 sg13g2_decap_8 FILLER_17_799 ();
 sg13g2_decap_8 FILLER_17_806 ();
 sg13g2_decap_8 FILLER_17_813 ();
 sg13g2_decap_8 FILLER_17_820 ();
 sg13g2_decap_8 FILLER_17_827 ();
 sg13g2_decap_8 FILLER_17_834 ();
 sg13g2_decap_8 FILLER_17_841 ();
 sg13g2_decap_8 FILLER_17_848 ();
 sg13g2_decap_8 FILLER_17_855 ();
 sg13g2_decap_8 FILLER_17_862 ();
 sg13g2_decap_8 FILLER_17_869 ();
 sg13g2_fill_2 FILLER_17_876 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_182 ();
 sg13g2_fill_2 FILLER_18_187 ();
 sg13g2_fill_1 FILLER_18_193 ();
 sg13g2_decap_4 FILLER_18_198 ();
 sg13g2_fill_2 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_decap_4 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_4 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_290 ();
 sg13g2_decap_4 FILLER_18_297 ();
 sg13g2_fill_2 FILLER_18_309 ();
 sg13g2_fill_1 FILLER_18_311 ();
 sg13g2_decap_4 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_4 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_decap_4 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_fill_2 FILLER_18_411 ();
 sg13g2_fill_1 FILLER_18_413 ();
 sg13g2_fill_1 FILLER_18_418 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_decap_8 FILLER_18_430 ();
 sg13g2_decap_4 FILLER_18_437 ();
 sg13g2_decap_8 FILLER_18_445 ();
 sg13g2_fill_1 FILLER_18_452 ();
 sg13g2_fill_2 FILLER_18_457 ();
 sg13g2_fill_2 FILLER_18_463 ();
 sg13g2_fill_2 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_475 ();
 sg13g2_fill_2 FILLER_18_482 ();
 sg13g2_decap_4 FILLER_18_493 ();
 sg13g2_fill_1 FILLER_18_497 ();
 sg13g2_fill_1 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_517 ();
 sg13g2_decap_8 FILLER_18_524 ();
 sg13g2_decap_4 FILLER_18_531 ();
 sg13g2_decap_8 FILLER_18_540 ();
 sg13g2_decap_8 FILLER_18_547 ();
 sg13g2_fill_2 FILLER_18_554 ();
 sg13g2_fill_1 FILLER_18_556 ();
 sg13g2_decap_8 FILLER_18_565 ();
 sg13g2_decap_4 FILLER_18_572 ();
 sg13g2_fill_2 FILLER_18_576 ();
 sg13g2_decap_4 FILLER_18_582 ();
 sg13g2_decap_8 FILLER_18_592 ();
 sg13g2_decap_8 FILLER_18_599 ();
 sg13g2_fill_2 FILLER_18_606 ();
 sg13g2_decap_8 FILLER_18_611 ();
 sg13g2_decap_8 FILLER_18_618 ();
 sg13g2_decap_8 FILLER_18_625 ();
 sg13g2_decap_8 FILLER_18_632 ();
 sg13g2_decap_8 FILLER_18_639 ();
 sg13g2_decap_8 FILLER_18_646 ();
 sg13g2_decap_8 FILLER_18_653 ();
 sg13g2_decap_8 FILLER_18_660 ();
 sg13g2_decap_4 FILLER_18_671 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_fill_1 FILLER_18_721 ();
 sg13g2_fill_2 FILLER_18_727 ();
 sg13g2_decap_8 FILLER_18_733 ();
 sg13g2_decap_8 FILLER_18_740 ();
 sg13g2_decap_8 FILLER_18_747 ();
 sg13g2_decap_8 FILLER_18_754 ();
 sg13g2_decap_8 FILLER_18_761 ();
 sg13g2_decap_8 FILLER_18_768 ();
 sg13g2_decap_8 FILLER_18_775 ();
 sg13g2_decap_8 FILLER_18_782 ();
 sg13g2_decap_8 FILLER_18_789 ();
 sg13g2_decap_8 FILLER_18_796 ();
 sg13g2_decap_8 FILLER_18_803 ();
 sg13g2_decap_8 FILLER_18_810 ();
 sg13g2_decap_8 FILLER_18_817 ();
 sg13g2_decap_8 FILLER_18_824 ();
 sg13g2_decap_8 FILLER_18_831 ();
 sg13g2_decap_8 FILLER_18_838 ();
 sg13g2_decap_8 FILLER_18_845 ();
 sg13g2_decap_8 FILLER_18_852 ();
 sg13g2_decap_8 FILLER_18_859 ();
 sg13g2_decap_8 FILLER_18_866 ();
 sg13g2_decap_4 FILLER_18_873 ();
 sg13g2_fill_1 FILLER_18_877 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_fill_2 FILLER_19_140 ();
 sg13g2_fill_2 FILLER_19_146 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_decap_4 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_185 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_decap_4 FILLER_19_212 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_230 ();
 sg13g2_decap_4 FILLER_19_237 ();
 sg13g2_fill_2 FILLER_19_241 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_4 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_fill_1 FILLER_19_298 ();
 sg13g2_fill_2 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_353 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_fill_1 FILLER_19_397 ();
 sg13g2_decap_8 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_411 ();
 sg13g2_fill_1 FILLER_19_422 ();
 sg13g2_decap_8 FILLER_19_432 ();
 sg13g2_decap_8 FILLER_19_439 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_fill_2 FILLER_19_462 ();
 sg13g2_fill_1 FILLER_19_464 ();
 sg13g2_fill_1 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_474 ();
 sg13g2_decap_8 FILLER_19_481 ();
 sg13g2_decap_8 FILLER_19_492 ();
 sg13g2_decap_8 FILLER_19_499 ();
 sg13g2_decap_8 FILLER_19_506 ();
 sg13g2_decap_8 FILLER_19_513 ();
 sg13g2_fill_2 FILLER_19_520 ();
 sg13g2_fill_1 FILLER_19_522 ();
 sg13g2_decap_8 FILLER_19_541 ();
 sg13g2_decap_8 FILLER_19_548 ();
 sg13g2_decap_8 FILLER_19_555 ();
 sg13g2_decap_4 FILLER_19_566 ();
 sg13g2_fill_1 FILLER_19_570 ();
 sg13g2_decap_8 FILLER_19_575 ();
 sg13g2_decap_8 FILLER_19_582 ();
 sg13g2_decap_8 FILLER_19_589 ();
 sg13g2_decap_8 FILLER_19_596 ();
 sg13g2_fill_1 FILLER_19_603 ();
 sg13g2_decap_8 FILLER_19_621 ();
 sg13g2_decap_8 FILLER_19_628 ();
 sg13g2_decap_8 FILLER_19_635 ();
 sg13g2_decap_8 FILLER_19_642 ();
 sg13g2_decap_8 FILLER_19_649 ();
 sg13g2_fill_2 FILLER_19_656 ();
 sg13g2_fill_1 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_677 ();
 sg13g2_decap_8 FILLER_19_684 ();
 sg13g2_decap_8 FILLER_19_691 ();
 sg13g2_decap_8 FILLER_19_698 ();
 sg13g2_decap_4 FILLER_19_705 ();
 sg13g2_decap_8 FILLER_19_713 ();
 sg13g2_decap_4 FILLER_19_720 ();
 sg13g2_fill_2 FILLER_19_724 ();
 sg13g2_decap_8 FILLER_19_731 ();
 sg13g2_decap_8 FILLER_19_738 ();
 sg13g2_decap_8 FILLER_19_745 ();
 sg13g2_decap_8 FILLER_19_752 ();
 sg13g2_decap_8 FILLER_19_759 ();
 sg13g2_decap_8 FILLER_19_766 ();
 sg13g2_decap_8 FILLER_19_773 ();
 sg13g2_decap_8 FILLER_19_780 ();
 sg13g2_decap_8 FILLER_19_787 ();
 sg13g2_decap_8 FILLER_19_794 ();
 sg13g2_decap_8 FILLER_19_801 ();
 sg13g2_decap_8 FILLER_19_808 ();
 sg13g2_decap_8 FILLER_19_815 ();
 sg13g2_decap_8 FILLER_19_822 ();
 sg13g2_decap_8 FILLER_19_829 ();
 sg13g2_decap_8 FILLER_19_836 ();
 sg13g2_decap_8 FILLER_19_843 ();
 sg13g2_decap_8 FILLER_19_850 ();
 sg13g2_decap_8 FILLER_19_857 ();
 sg13g2_decap_8 FILLER_19_864 ();
 sg13g2_decap_8 FILLER_19_871 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_118 ();
 sg13g2_decap_8 FILLER_20_125 ();
 sg13g2_decap_8 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_146 ();
 sg13g2_decap_8 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_fill_2 FILLER_20_166 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_decap_4 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_decap_4 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_195 ();
 sg13g2_decap_4 FILLER_20_206 ();
 sg13g2_decap_8 FILLER_20_215 ();
 sg13g2_decap_8 FILLER_20_234 ();
 sg13g2_decap_4 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_fill_2 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_338 ();
 sg13g2_decap_4 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_fill_2 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_4 FILLER_20_417 ();
 sg13g2_fill_1 FILLER_20_425 ();
 sg13g2_decap_8 FILLER_20_432 ();
 sg13g2_fill_1 FILLER_20_439 ();
 sg13g2_decap_8 FILLER_20_443 ();
 sg13g2_decap_8 FILLER_20_450 ();
 sg13g2_decap_8 FILLER_20_457 ();
 sg13g2_fill_2 FILLER_20_464 ();
 sg13g2_fill_1 FILLER_20_466 ();
 sg13g2_decap_8 FILLER_20_471 ();
 sg13g2_fill_1 FILLER_20_478 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_500 ();
 sg13g2_decap_8 FILLER_20_507 ();
 sg13g2_decap_8 FILLER_20_514 ();
 sg13g2_fill_2 FILLER_20_521 ();
 sg13g2_fill_1 FILLER_20_523 ();
 sg13g2_decap_8 FILLER_20_528 ();
 sg13g2_fill_1 FILLER_20_535 ();
 sg13g2_decap_4 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_562 ();
 sg13g2_decap_4 FILLER_20_569 ();
 sg13g2_fill_2 FILLER_20_573 ();
 sg13g2_decap_8 FILLER_20_585 ();
 sg13g2_decap_8 FILLER_20_592 ();
 sg13g2_fill_2 FILLER_20_599 ();
 sg13g2_fill_1 FILLER_20_601 ();
 sg13g2_decap_4 FILLER_20_611 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_fill_2 FILLER_20_658 ();
 sg13g2_fill_1 FILLER_20_660 ();
 sg13g2_decap_4 FILLER_20_669 ();
 sg13g2_fill_2 FILLER_20_673 ();
 sg13g2_decap_4 FILLER_20_679 ();
 sg13g2_fill_1 FILLER_20_683 ();
 sg13g2_decap_8 FILLER_20_692 ();
 sg13g2_decap_4 FILLER_20_699 ();
 sg13g2_fill_1 FILLER_20_703 ();
 sg13g2_decap_8 FILLER_20_709 ();
 sg13g2_decap_8 FILLER_20_716 ();
 sg13g2_decap_8 FILLER_20_723 ();
 sg13g2_decap_8 FILLER_20_730 ();
 sg13g2_decap_8 FILLER_20_737 ();
 sg13g2_decap_8 FILLER_20_744 ();
 sg13g2_fill_1 FILLER_20_751 ();
 sg13g2_decap_8 FILLER_20_757 ();
 sg13g2_decap_8 FILLER_20_764 ();
 sg13g2_decap_8 FILLER_20_771 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_decap_8 FILLER_20_785 ();
 sg13g2_decap_8 FILLER_20_792 ();
 sg13g2_decap_8 FILLER_20_799 ();
 sg13g2_decap_8 FILLER_20_806 ();
 sg13g2_decap_8 FILLER_20_813 ();
 sg13g2_decap_8 FILLER_20_820 ();
 sg13g2_decap_8 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_decap_8 FILLER_20_841 ();
 sg13g2_decap_8 FILLER_20_848 ();
 sg13g2_decap_8 FILLER_20_855 ();
 sg13g2_decap_8 FILLER_20_862 ();
 sg13g2_decap_8 FILLER_20_869 ();
 sg13g2_fill_2 FILLER_20_876 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_4 FILLER_21_84 ();
 sg13g2_fill_1 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_93 ();
 sg13g2_decap_4 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_118 ();
 sg13g2_decap_8 FILLER_21_125 ();
 sg13g2_decap_8 FILLER_21_132 ();
 sg13g2_decap_8 FILLER_21_139 ();
 sg13g2_decap_4 FILLER_21_146 ();
 sg13g2_decap_4 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_decap_4 FILLER_21_164 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_fill_2 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_206 ();
 sg13g2_fill_2 FILLER_21_224 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_2 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_8 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_270 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_decap_4 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_329 ();
 sg13g2_decap_4 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_decap_4 FILLER_21_351 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_370 ();
 sg13g2_decap_8 FILLER_21_377 ();
 sg13g2_fill_2 FILLER_21_384 ();
 sg13g2_fill_1 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_4 FILLER_21_399 ();
 sg13g2_decap_4 FILLER_21_409 ();
 sg13g2_fill_2 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_21_430 ();
 sg13g2_decap_8 FILLER_21_437 ();
 sg13g2_decap_8 FILLER_21_444 ();
 sg13g2_decap_8 FILLER_21_451 ();
 sg13g2_decap_4 FILLER_21_458 ();
 sg13g2_fill_2 FILLER_21_462 ();
 sg13g2_decap_4 FILLER_21_468 ();
 sg13g2_fill_1 FILLER_21_472 ();
 sg13g2_decap_8 FILLER_21_479 ();
 sg13g2_decap_8 FILLER_21_486 ();
 sg13g2_fill_2 FILLER_21_493 ();
 sg13g2_fill_1 FILLER_21_495 ();
 sg13g2_decap_8 FILLER_21_500 ();
 sg13g2_fill_2 FILLER_21_507 ();
 sg13g2_fill_1 FILLER_21_509 ();
 sg13g2_decap_8 FILLER_21_514 ();
 sg13g2_fill_2 FILLER_21_521 ();
 sg13g2_fill_1 FILLER_21_523 ();
 sg13g2_decap_8 FILLER_21_535 ();
 sg13g2_decap_8 FILLER_21_549 ();
 sg13g2_fill_2 FILLER_21_556 ();
 sg13g2_fill_1 FILLER_21_558 ();
 sg13g2_fill_2 FILLER_21_564 ();
 sg13g2_decap_8 FILLER_21_572 ();
 sg13g2_decap_8 FILLER_21_579 ();
 sg13g2_decap_8 FILLER_21_586 ();
 sg13g2_decap_8 FILLER_21_593 ();
 sg13g2_decap_8 FILLER_21_600 ();
 sg13g2_decap_4 FILLER_21_607 ();
 sg13g2_fill_2 FILLER_21_611 ();
 sg13g2_decap_8 FILLER_21_617 ();
 sg13g2_decap_8 FILLER_21_624 ();
 sg13g2_decap_8 FILLER_21_631 ();
 sg13g2_decap_8 FILLER_21_638 ();
 sg13g2_decap_8 FILLER_21_645 ();
 sg13g2_decap_8 FILLER_21_652 ();
 sg13g2_decap_8 FILLER_21_659 ();
 sg13g2_fill_1 FILLER_21_666 ();
 sg13g2_decap_4 FILLER_21_672 ();
 sg13g2_fill_1 FILLER_21_676 ();
 sg13g2_fill_2 FILLER_21_685 ();
 sg13g2_fill_1 FILLER_21_687 ();
 sg13g2_fill_1 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_698 ();
 sg13g2_fill_1 FILLER_21_705 ();
 sg13g2_decap_8 FILLER_21_710 ();
 sg13g2_decap_8 FILLER_21_717 ();
 sg13g2_fill_1 FILLER_21_724 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_21_868 ();
 sg13g2_fill_2 FILLER_21_875 ();
 sg13g2_fill_1 FILLER_21_877 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_86 ();
 sg13g2_decap_4 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_99 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_decap_4 FILLER_22_119 ();
 sg13g2_fill_1 FILLER_22_123 ();
 sg13g2_decap_4 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_132 ();
 sg13g2_fill_2 FILLER_22_139 ();
 sg13g2_decap_8 FILLER_22_150 ();
 sg13g2_decap_8 FILLER_22_157 ();
 sg13g2_fill_1 FILLER_22_164 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_191 ();
 sg13g2_decap_4 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_fill_2 FILLER_22_228 ();
 sg13g2_fill_1 FILLER_22_230 ();
 sg13g2_decap_8 FILLER_22_239 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_decap_8 FILLER_22_271 ();
 sg13g2_decap_8 FILLER_22_278 ();
 sg13g2_fill_2 FILLER_22_285 ();
 sg13g2_decap_4 FILLER_22_295 ();
 sg13g2_fill_1 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_fill_2 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_332 ();
 sg13g2_decap_8 FILLER_22_339 ();
 sg13g2_decap_4 FILLER_22_346 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_fill_2 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_4 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_405 ();
 sg13g2_decap_4 FILLER_22_412 ();
 sg13g2_fill_1 FILLER_22_416 ();
 sg13g2_decap_8 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_22_435 ();
 sg13g2_decap_8 FILLER_22_442 ();
 sg13g2_decap_4 FILLER_22_455 ();
 sg13g2_fill_1 FILLER_22_459 ();
 sg13g2_decap_8 FILLER_22_465 ();
 sg13g2_decap_8 FILLER_22_472 ();
 sg13g2_decap_8 FILLER_22_479 ();
 sg13g2_fill_2 FILLER_22_486 ();
 sg13g2_fill_1 FILLER_22_492 ();
 sg13g2_fill_2 FILLER_22_502 ();
 sg13g2_fill_1 FILLER_22_504 ();
 sg13g2_fill_2 FILLER_22_509 ();
 sg13g2_decap_8 FILLER_22_519 ();
 sg13g2_decap_8 FILLER_22_526 ();
 sg13g2_decap_8 FILLER_22_533 ();
 sg13g2_fill_2 FILLER_22_540 ();
 sg13g2_fill_1 FILLER_22_542 ();
 sg13g2_decap_8 FILLER_22_557 ();
 sg13g2_decap_8 FILLER_22_564 ();
 sg13g2_decap_4 FILLER_22_571 ();
 sg13g2_fill_2 FILLER_22_575 ();
 sg13g2_decap_8 FILLER_22_585 ();
 sg13g2_fill_2 FILLER_22_592 ();
 sg13g2_decap_4 FILLER_22_602 ();
 sg13g2_fill_1 FILLER_22_610 ();
 sg13g2_decap_4 FILLER_22_615 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_4 FILLER_22_634 ();
 sg13g2_decap_8 FILLER_22_642 ();
 sg13g2_decap_4 FILLER_22_649 ();
 sg13g2_fill_2 FILLER_22_653 ();
 sg13g2_decap_8 FILLER_22_663 ();
 sg13g2_decap_8 FILLER_22_670 ();
 sg13g2_decap_4 FILLER_22_677 ();
 sg13g2_decap_4 FILLER_22_686 ();
 sg13g2_decap_4 FILLER_22_696 ();
 sg13g2_fill_2 FILLER_22_700 ();
 sg13g2_fill_1 FILLER_22_706 ();
 sg13g2_decap_8 FILLER_22_712 ();
 sg13g2_decap_8 FILLER_22_719 ();
 sg13g2_fill_2 FILLER_22_726 ();
 sg13g2_fill_1 FILLER_22_734 ();
 sg13g2_fill_2 FILLER_22_747 ();
 sg13g2_fill_1 FILLER_22_749 ();
 sg13g2_fill_1 FILLER_22_754 ();
 sg13g2_decap_8 FILLER_22_759 ();
 sg13g2_decap_8 FILLER_22_766 ();
 sg13g2_decap_8 FILLER_22_773 ();
 sg13g2_decap_8 FILLER_22_780 ();
 sg13g2_decap_8 FILLER_22_787 ();
 sg13g2_decap_8 FILLER_22_794 ();
 sg13g2_decap_8 FILLER_22_801 ();
 sg13g2_decap_8 FILLER_22_808 ();
 sg13g2_decap_8 FILLER_22_815 ();
 sg13g2_decap_8 FILLER_22_822 ();
 sg13g2_decap_8 FILLER_22_829 ();
 sg13g2_decap_8 FILLER_22_836 ();
 sg13g2_decap_8 FILLER_22_843 ();
 sg13g2_decap_8 FILLER_22_850 ();
 sg13g2_decap_8 FILLER_22_857 ();
 sg13g2_decap_8 FILLER_22_864 ();
 sg13g2_decap_8 FILLER_22_871 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_4 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_decap_4 FILLER_23_107 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_121 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_4 FILLER_23_175 ();
 sg13g2_fill_2 FILLER_23_179 ();
 sg13g2_decap_4 FILLER_23_189 ();
 sg13g2_fill_2 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_212 ();
 sg13g2_decap_4 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_237 ();
 sg13g2_fill_1 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_262 ();
 sg13g2_decap_8 FILLER_23_269 ();
 sg13g2_decap_8 FILLER_23_276 ();
 sg13g2_decap_4 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_337 ();
 sg13g2_fill_1 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_decap_4 FILLER_23_359 ();
 sg13g2_fill_2 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_4 FILLER_23_388 ();
 sg13g2_fill_1 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_decap_4 FILLER_23_408 ();
 sg13g2_fill_2 FILLER_23_412 ();
 sg13g2_decap_4 FILLER_23_422 ();
 sg13g2_fill_2 FILLER_23_437 ();
 sg13g2_decap_8 FILLER_23_452 ();
 sg13g2_decap_8 FILLER_23_463 ();
 sg13g2_decap_8 FILLER_23_470 ();
 sg13g2_fill_2 FILLER_23_481 ();
 sg13g2_fill_1 FILLER_23_483 ();
 sg13g2_fill_2 FILLER_23_493 ();
 sg13g2_decap_8 FILLER_23_499 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_fill_2 FILLER_23_526 ();
 sg13g2_decap_4 FILLER_23_533 ();
 sg13g2_fill_1 FILLER_23_537 ();
 sg13g2_fill_2 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_557 ();
 sg13g2_decap_8 FILLER_23_564 ();
 sg13g2_decap_8 FILLER_23_571 ();
 sg13g2_decap_8 FILLER_23_578 ();
 sg13g2_decap_4 FILLER_23_585 ();
 sg13g2_fill_2 FILLER_23_589 ();
 sg13g2_fill_2 FILLER_23_603 ();
 sg13g2_fill_1 FILLER_23_605 ();
 sg13g2_fill_1 FILLER_23_616 ();
 sg13g2_decap_4 FILLER_23_621 ();
 sg13g2_fill_2 FILLER_23_625 ();
 sg13g2_decap_4 FILLER_23_631 ();
 sg13g2_decap_8 FILLER_23_643 ();
 sg13g2_decap_4 FILLER_23_650 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_4 FILLER_23_672 ();
 sg13g2_fill_1 FILLER_23_676 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_decap_8 FILLER_23_690 ();
 sg13g2_decap_8 FILLER_23_697 ();
 sg13g2_decap_8 FILLER_23_704 ();
 sg13g2_fill_1 FILLER_23_711 ();
 sg13g2_decap_8 FILLER_23_715 ();
 sg13g2_decap_8 FILLER_23_722 ();
 sg13g2_fill_1 FILLER_23_729 ();
 sg13g2_fill_2 FILLER_23_743 ();
 sg13g2_fill_1 FILLER_23_745 ();
 sg13g2_fill_1 FILLER_23_754 ();
 sg13g2_decap_8 FILLER_23_760 ();
 sg13g2_decap_8 FILLER_23_767 ();
 sg13g2_decap_8 FILLER_23_774 ();
 sg13g2_decap_8 FILLER_23_781 ();
 sg13g2_decap_8 FILLER_23_788 ();
 sg13g2_decap_8 FILLER_23_795 ();
 sg13g2_decap_8 FILLER_23_802 ();
 sg13g2_decap_8 FILLER_23_809 ();
 sg13g2_decap_8 FILLER_23_816 ();
 sg13g2_decap_8 FILLER_23_823 ();
 sg13g2_decap_8 FILLER_23_830 ();
 sg13g2_decap_8 FILLER_23_837 ();
 sg13g2_decap_8 FILLER_23_844 ();
 sg13g2_decap_8 FILLER_23_851 ();
 sg13g2_decap_8 FILLER_23_858 ();
 sg13g2_decap_8 FILLER_23_865 ();
 sg13g2_decap_4 FILLER_23_872 ();
 sg13g2_fill_2 FILLER_23_876 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_4 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_decap_4 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_195 ();
 sg13g2_decap_4 FILLER_24_202 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_236 ();
 sg13g2_fill_2 FILLER_24_243 ();
 sg13g2_fill_1 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_285 ();
 sg13g2_decap_4 FILLER_24_290 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_fill_2 FILLER_24_319 ();
 sg13g2_fill_1 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_359 ();
 sg13g2_fill_1 FILLER_24_361 ();
 sg13g2_decap_4 FILLER_24_371 ();
 sg13g2_decap_4 FILLER_24_385 ();
 sg13g2_fill_2 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_24_409 ();
 sg13g2_decap_8 FILLER_24_423 ();
 sg13g2_fill_2 FILLER_24_430 ();
 sg13g2_fill_1 FILLER_24_432 ();
 sg13g2_decap_8 FILLER_24_437 ();
 sg13g2_decap_4 FILLER_24_444 ();
 sg13g2_fill_2 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_460 ();
 sg13g2_fill_2 FILLER_24_467 ();
 sg13g2_fill_2 FILLER_24_474 ();
 sg13g2_decap_8 FILLER_24_481 ();
 sg13g2_fill_2 FILLER_24_488 ();
 sg13g2_fill_1 FILLER_24_495 ();
 sg13g2_decap_8 FILLER_24_517 ();
 sg13g2_fill_1 FILLER_24_524 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_4 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_548 ();
 sg13g2_decap_4 FILLER_24_555 ();
 sg13g2_fill_1 FILLER_24_559 ();
 sg13g2_decap_4 FILLER_24_566 ();
 sg13g2_decap_8 FILLER_24_594 ();
 sg13g2_decap_8 FILLER_24_601 ();
 sg13g2_decap_4 FILLER_24_612 ();
 sg13g2_decap_4 FILLER_24_621 ();
 sg13g2_fill_2 FILLER_24_625 ();
 sg13g2_fill_1 FILLER_24_632 ();
 sg13g2_fill_1 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_653 ();
 sg13g2_decap_8 FILLER_24_660 ();
 sg13g2_decap_8 FILLER_24_667 ();
 sg13g2_decap_4 FILLER_24_674 ();
 sg13g2_decap_4 FILLER_24_684 ();
 sg13g2_fill_1 FILLER_24_688 ();
 sg13g2_decap_8 FILLER_24_697 ();
 sg13g2_decap_4 FILLER_24_704 ();
 sg13g2_decap_4 FILLER_24_712 ();
 sg13g2_fill_1 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_726 ();
 sg13g2_decap_8 FILLER_24_733 ();
 sg13g2_decap_8 FILLER_24_740 ();
 sg13g2_decap_8 FILLER_24_747 ();
 sg13g2_decap_8 FILLER_24_754 ();
 sg13g2_decap_8 FILLER_24_761 ();
 sg13g2_decap_8 FILLER_24_768 ();
 sg13g2_decap_8 FILLER_24_775 ();
 sg13g2_decap_8 FILLER_24_782 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_decap_8 FILLER_24_796 ();
 sg13g2_decap_8 FILLER_24_803 ();
 sg13g2_decap_8 FILLER_24_810 ();
 sg13g2_decap_8 FILLER_24_817 ();
 sg13g2_decap_8 FILLER_24_824 ();
 sg13g2_decap_8 FILLER_24_831 ();
 sg13g2_decap_8 FILLER_24_838 ();
 sg13g2_decap_8 FILLER_24_845 ();
 sg13g2_decap_8 FILLER_24_852 ();
 sg13g2_decap_8 FILLER_24_859 ();
 sg13g2_decap_8 FILLER_24_866 ();
 sg13g2_decap_4 FILLER_24_873 ();
 sg13g2_fill_1 FILLER_24_877 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_121 ();
 sg13g2_decap_8 FILLER_25_128 ();
 sg13g2_decap_4 FILLER_25_135 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_fill_1 FILLER_25_153 ();
 sg13g2_decap_8 FILLER_25_159 ();
 sg13g2_decap_4 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_decap_8 FILLER_25_185 ();
 sg13g2_decap_8 FILLER_25_192 ();
 sg13g2_decap_8 FILLER_25_199 ();
 sg13g2_decap_4 FILLER_25_206 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_decap_4 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_234 ();
 sg13g2_fill_2 FILLER_25_241 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_decap_4 FILLER_25_254 ();
 sg13g2_fill_1 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_278 ();
 sg13g2_decap_4 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_298 ();
 sg13g2_decap_8 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_decap_4 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_354 ();
 sg13g2_decap_4 FILLER_25_360 ();
 sg13g2_fill_1 FILLER_25_364 ();
 sg13g2_decap_4 FILLER_25_369 ();
 sg13g2_fill_2 FILLER_25_373 ();
 sg13g2_fill_1 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_414 ();
 sg13g2_fill_2 FILLER_25_430 ();
 sg13g2_decap_8 FILLER_25_436 ();
 sg13g2_decap_8 FILLER_25_443 ();
 sg13g2_decap_8 FILLER_25_460 ();
 sg13g2_decap_8 FILLER_25_467 ();
 sg13g2_decap_8 FILLER_25_474 ();
 sg13g2_decap_4 FILLER_25_481 ();
 sg13g2_fill_1 FILLER_25_485 ();
 sg13g2_decap_8 FILLER_25_491 ();
 sg13g2_decap_8 FILLER_25_498 ();
 sg13g2_decap_8 FILLER_25_505 ();
 sg13g2_decap_8 FILLER_25_512 ();
 sg13g2_decap_8 FILLER_25_519 ();
 sg13g2_decap_8 FILLER_25_526 ();
 sg13g2_decap_8 FILLER_25_533 ();
 sg13g2_decap_8 FILLER_25_540 ();
 sg13g2_decap_8 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_559 ();
 sg13g2_fill_1 FILLER_25_566 ();
 sg13g2_decap_4 FILLER_25_572 ();
 sg13g2_decap_4 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_611 ();
 sg13g2_decap_4 FILLER_25_618 ();
 sg13g2_fill_1 FILLER_25_622 ();
 sg13g2_decap_4 FILLER_25_628 ();
 sg13g2_fill_2 FILLER_25_632 ();
 sg13g2_decap_8 FILLER_25_638 ();
 sg13g2_decap_8 FILLER_25_645 ();
 sg13g2_decap_8 FILLER_25_652 ();
 sg13g2_decap_4 FILLER_25_659 ();
 sg13g2_fill_1 FILLER_25_663 ();
 sg13g2_decap_4 FILLER_25_669 ();
 sg13g2_fill_2 FILLER_25_673 ();
 sg13g2_decap_8 FILLER_25_689 ();
 sg13g2_decap_8 FILLER_25_696 ();
 sg13g2_decap_8 FILLER_25_703 ();
 sg13g2_decap_8 FILLER_25_710 ();
 sg13g2_fill_2 FILLER_25_717 ();
 sg13g2_decap_8 FILLER_25_723 ();
 sg13g2_fill_1 FILLER_25_730 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_decap_8 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_fill_2 FILLER_25_875 ();
 sg13g2_fill_1 FILLER_25_877 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_83 ();
 sg13g2_decap_8 FILLER_26_93 ();
 sg13g2_decap_8 FILLER_26_100 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_4 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_160 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_decap_4 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_230 ();
 sg13g2_decap_8 FILLER_26_237 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_fill_1 FILLER_26_315 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_fill_2 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_344 ();
 sg13g2_decap_4 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_364 ();
 sg13g2_decap_4 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_decap_8 FILLER_26_408 ();
 sg13g2_decap_4 FILLER_26_415 ();
 sg13g2_fill_1 FILLER_26_419 ();
 sg13g2_decap_4 FILLER_26_424 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_4 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_442 ();
 sg13g2_decap_8 FILLER_26_449 ();
 sg13g2_decap_8 FILLER_26_456 ();
 sg13g2_decap_8 FILLER_26_463 ();
 sg13g2_decap_8 FILLER_26_470 ();
 sg13g2_decap_8 FILLER_26_486 ();
 sg13g2_decap_8 FILLER_26_493 ();
 sg13g2_decap_4 FILLER_26_500 ();
 sg13g2_decap_8 FILLER_26_508 ();
 sg13g2_decap_4 FILLER_26_520 ();
 sg13g2_decap_8 FILLER_26_528 ();
 sg13g2_fill_2 FILLER_26_535 ();
 sg13g2_fill_2 FILLER_26_554 ();
 sg13g2_fill_2 FILLER_26_560 ();
 sg13g2_decap_4 FILLER_26_573 ();
 sg13g2_fill_1 FILLER_26_577 ();
 sg13g2_fill_2 FILLER_26_589 ();
 sg13g2_fill_2 FILLER_26_597 ();
 sg13g2_decap_8 FILLER_26_607 ();
 sg13g2_decap_8 FILLER_26_614 ();
 sg13g2_decap_4 FILLER_26_621 ();
 sg13g2_fill_2 FILLER_26_625 ();
 sg13g2_fill_2 FILLER_26_633 ();
 sg13g2_decap_8 FILLER_26_639 ();
 sg13g2_fill_1 FILLER_26_646 ();
 sg13g2_decap_8 FILLER_26_652 ();
 sg13g2_fill_1 FILLER_26_659 ();
 sg13g2_decap_4 FILLER_26_664 ();
 sg13g2_fill_2 FILLER_26_668 ();
 sg13g2_decap_8 FILLER_26_674 ();
 sg13g2_fill_1 FILLER_26_681 ();
 sg13g2_fill_2 FILLER_26_686 ();
 sg13g2_fill_1 FILLER_26_688 ();
 sg13g2_decap_4 FILLER_26_707 ();
 sg13g2_decap_4 FILLER_26_717 ();
 sg13g2_fill_2 FILLER_26_734 ();
 sg13g2_fill_1 FILLER_26_741 ();
 sg13g2_decap_8 FILLER_26_746 ();
 sg13g2_decap_8 FILLER_26_753 ();
 sg13g2_decap_8 FILLER_26_760 ();
 sg13g2_decap_8 FILLER_26_767 ();
 sg13g2_decap_8 FILLER_26_774 ();
 sg13g2_decap_8 FILLER_26_781 ();
 sg13g2_decap_8 FILLER_26_788 ();
 sg13g2_decap_8 FILLER_26_795 ();
 sg13g2_decap_8 FILLER_26_802 ();
 sg13g2_decap_8 FILLER_26_809 ();
 sg13g2_decap_8 FILLER_26_816 ();
 sg13g2_decap_8 FILLER_26_823 ();
 sg13g2_decap_8 FILLER_26_830 ();
 sg13g2_decap_8 FILLER_26_837 ();
 sg13g2_decap_8 FILLER_26_844 ();
 sg13g2_decap_8 FILLER_26_851 ();
 sg13g2_decap_8 FILLER_26_858 ();
 sg13g2_decap_8 FILLER_26_865 ();
 sg13g2_decap_4 FILLER_26_872 ();
 sg13g2_fill_2 FILLER_26_876 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_53 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_decap_8 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_107 ();
 sg13g2_decap_4 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_152 ();
 sg13g2_decap_4 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_163 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_4 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_decap_4 FILLER_27_185 ();
 sg13g2_decap_8 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_4 FILLER_27_287 ();
 sg13g2_fill_1 FILLER_27_291 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_4 FILLER_27_308 ();
 sg13g2_fill_2 FILLER_27_312 ();
 sg13g2_decap_4 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_4 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_4 FILLER_27_392 ();
 sg13g2_fill_2 FILLER_27_396 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_4 FILLER_27_436 ();
 sg13g2_fill_1 FILLER_27_440 ();
 sg13g2_fill_2 FILLER_27_444 ();
 sg13g2_fill_1 FILLER_27_446 ();
 sg13g2_decap_8 FILLER_27_452 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_fill_1 FILLER_27_474 ();
 sg13g2_decap_8 FILLER_27_484 ();
 sg13g2_decap_8 FILLER_27_491 ();
 sg13g2_decap_4 FILLER_27_498 ();
 sg13g2_fill_2 FILLER_27_502 ();
 sg13g2_decap_8 FILLER_27_507 ();
 sg13g2_fill_2 FILLER_27_514 ();
 sg13g2_decap_8 FILLER_27_521 ();
 sg13g2_fill_2 FILLER_27_528 ();
 sg13g2_fill_1 FILLER_27_530 ();
 sg13g2_decap_4 FILLER_27_536 ();
 sg13g2_fill_2 FILLER_27_540 ();
 sg13g2_fill_2 FILLER_27_546 ();
 sg13g2_fill_1 FILLER_27_558 ();
 sg13g2_fill_2 FILLER_27_563 ();
 sg13g2_fill_1 FILLER_27_565 ();
 sg13g2_decap_8 FILLER_27_570 ();
 sg13g2_fill_2 FILLER_27_577 ();
 sg13g2_fill_1 FILLER_27_579 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_4 FILLER_27_623 ();
 sg13g2_decap_4 FILLER_27_631 ();
 sg13g2_decap_8 FILLER_27_641 ();
 sg13g2_fill_1 FILLER_27_648 ();
 sg13g2_decap_4 FILLER_27_653 ();
 sg13g2_fill_2 FILLER_27_666 ();
 sg13g2_fill_1 FILLER_27_668 ();
 sg13g2_fill_1 FILLER_27_674 ();
 sg13g2_decap_8 FILLER_27_681 ();
 sg13g2_fill_1 FILLER_27_688 ();
 sg13g2_fill_2 FILLER_27_698 ();
 sg13g2_decap_8 FILLER_27_712 ();
 sg13g2_fill_1 FILLER_27_719 ();
 sg13g2_fill_1 FILLER_27_724 ();
 sg13g2_decap_8 FILLER_27_729 ();
 sg13g2_fill_1 FILLER_27_736 ();
 sg13g2_fill_1 FILLER_27_741 ();
 sg13g2_decap_8 FILLER_27_751 ();
 sg13g2_decap_8 FILLER_27_758 ();
 sg13g2_decap_8 FILLER_27_765 ();
 sg13g2_decap_8 FILLER_27_772 ();
 sg13g2_decap_8 FILLER_27_779 ();
 sg13g2_decap_8 FILLER_27_786 ();
 sg13g2_decap_8 FILLER_27_793 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_8 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_fill_1 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_4 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_73 ();
 sg13g2_decap_4 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_decap_4 FILLER_28_93 ();
 sg13g2_decap_8 FILLER_28_101 ();
 sg13g2_decap_8 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_4 FILLER_28_252 ();
 sg13g2_decap_4 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_decap_8 FILLER_28_279 ();
 sg13g2_decap_8 FILLER_28_286 ();
 sg13g2_decap_8 FILLER_28_293 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_decap_4 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_28_340 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_decap_4 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_4 FILLER_28_399 ();
 sg13g2_fill_1 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_409 ();
 sg13g2_decap_8 FILLER_28_430 ();
 sg13g2_fill_2 FILLER_28_437 ();
 sg13g2_fill_2 FILLER_28_444 ();
 sg13g2_fill_1 FILLER_28_446 ();
 sg13g2_fill_1 FILLER_28_472 ();
 sg13g2_decap_8 FILLER_28_477 ();
 sg13g2_decap_4 FILLER_28_484 ();
 sg13g2_fill_1 FILLER_28_488 ();
 sg13g2_decap_4 FILLER_28_493 ();
 sg13g2_fill_2 FILLER_28_497 ();
 sg13g2_fill_1 FILLER_28_504 ();
 sg13g2_decap_4 FILLER_28_514 ();
 sg13g2_decap_4 FILLER_28_523 ();
 sg13g2_fill_1 FILLER_28_527 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_fill_1 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_544 ();
 sg13g2_decap_8 FILLER_28_551 ();
 sg13g2_decap_8 FILLER_28_558 ();
 sg13g2_fill_2 FILLER_28_565 ();
 sg13g2_decap_8 FILLER_28_576 ();
 sg13g2_decap_8 FILLER_28_583 ();
 sg13g2_fill_2 FILLER_28_590 ();
 sg13g2_decap_8 FILLER_28_600 ();
 sg13g2_decap_8 FILLER_28_607 ();
 sg13g2_decap_8 FILLER_28_614 ();
 sg13g2_fill_2 FILLER_28_621 ();
 sg13g2_decap_8 FILLER_28_626 ();
 sg13g2_fill_1 FILLER_28_633 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_4 FILLER_28_658 ();
 sg13g2_fill_2 FILLER_28_666 ();
 sg13g2_fill_1 FILLER_28_668 ();
 sg13g2_decap_8 FILLER_28_673 ();
 sg13g2_decap_8 FILLER_28_680 ();
 sg13g2_fill_2 FILLER_28_687 ();
 sg13g2_fill_2 FILLER_28_693 ();
 sg13g2_fill_1 FILLER_28_695 ();
 sg13g2_decap_8 FILLER_28_701 ();
 sg13g2_fill_2 FILLER_28_708 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_4 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_737 ();
 sg13g2_decap_8 FILLER_28_744 ();
 sg13g2_decap_8 FILLER_28_751 ();
 sg13g2_decap_8 FILLER_28_758 ();
 sg13g2_decap_8 FILLER_28_765 ();
 sg13g2_decap_8 FILLER_28_772 ();
 sg13g2_decap_8 FILLER_28_779 ();
 sg13g2_decap_8 FILLER_28_786 ();
 sg13g2_decap_8 FILLER_28_793 ();
 sg13g2_decap_8 FILLER_28_800 ();
 sg13g2_decap_8 FILLER_28_807 ();
 sg13g2_decap_8 FILLER_28_814 ();
 sg13g2_decap_8 FILLER_28_821 ();
 sg13g2_decap_8 FILLER_28_828 ();
 sg13g2_decap_8 FILLER_28_835 ();
 sg13g2_decap_8 FILLER_28_842 ();
 sg13g2_decap_8 FILLER_28_849 ();
 sg13g2_decap_8 FILLER_28_856 ();
 sg13g2_decap_8 FILLER_28_863 ();
 sg13g2_decap_8 FILLER_28_870 ();
 sg13g2_fill_1 FILLER_28_877 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_79 ();
 sg13g2_fill_1 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_85 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_fill_1 FILLER_29_100 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_4 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_decap_8 FILLER_29_121 ();
 sg13g2_decap_8 FILLER_29_128 ();
 sg13g2_decap_4 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_157 ();
 sg13g2_fill_2 FILLER_29_164 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_decap_4 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_decap_4 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_225 ();
 sg13g2_decap_4 FILLER_29_232 ();
 sg13g2_fill_1 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_269 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_282 ();
 sg13g2_decap_4 FILLER_29_289 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_300 ();
 sg13g2_fill_2 FILLER_29_307 ();
 sg13g2_decap_4 FILLER_29_313 ();
 sg13g2_fill_1 FILLER_29_321 ();
 sg13g2_fill_2 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_fill_1 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_4 FILLER_29_358 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_4 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_424 ();
 sg13g2_fill_1 FILLER_29_431 ();
 sg13g2_fill_1 FILLER_29_451 ();
 sg13g2_decap_8 FILLER_29_456 ();
 sg13g2_decap_4 FILLER_29_463 ();
 sg13g2_decap_8 FILLER_29_481 ();
 sg13g2_fill_2 FILLER_29_488 ();
 sg13g2_decap_8 FILLER_29_502 ();
 sg13g2_decap_8 FILLER_29_509 ();
 sg13g2_fill_1 FILLER_29_516 ();
 sg13g2_decap_4 FILLER_29_522 ();
 sg13g2_fill_1 FILLER_29_526 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_4 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_562 ();
 sg13g2_decap_4 FILLER_29_569 ();
 sg13g2_fill_2 FILLER_29_573 ();
 sg13g2_decap_4 FILLER_29_581 ();
 sg13g2_fill_2 FILLER_29_585 ();
 sg13g2_decap_8 FILLER_29_600 ();
 sg13g2_fill_2 FILLER_29_607 ();
 sg13g2_decap_8 FILLER_29_614 ();
 sg13g2_fill_2 FILLER_29_621 ();
 sg13g2_fill_1 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_628 ();
 sg13g2_fill_1 FILLER_29_635 ();
 sg13g2_decap_4 FILLER_29_657 ();
 sg13g2_decap_8 FILLER_29_670 ();
 sg13g2_decap_8 FILLER_29_677 ();
 sg13g2_decap_8 FILLER_29_684 ();
 sg13g2_decap_4 FILLER_29_691 ();
 sg13g2_fill_2 FILLER_29_695 ();
 sg13g2_fill_2 FILLER_29_700 ();
 sg13g2_fill_1 FILLER_29_702 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_4 FILLER_29_728 ();
 sg13g2_fill_2 FILLER_29_732 ();
 sg13g2_decap_4 FILLER_29_738 ();
 sg13g2_fill_1 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_748 ();
 sg13g2_decap_8 FILLER_29_755 ();
 sg13g2_decap_8 FILLER_29_762 ();
 sg13g2_decap_8 FILLER_29_769 ();
 sg13g2_decap_8 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_783 ();
 sg13g2_decap_8 FILLER_29_790 ();
 sg13g2_decap_8 FILLER_29_797 ();
 sg13g2_decap_8 FILLER_29_804 ();
 sg13g2_decap_8 FILLER_29_811 ();
 sg13g2_decap_8 FILLER_29_818 ();
 sg13g2_decap_8 FILLER_29_825 ();
 sg13g2_decap_8 FILLER_29_832 ();
 sg13g2_decap_8 FILLER_29_839 ();
 sg13g2_decap_8 FILLER_29_846 ();
 sg13g2_decap_8 FILLER_29_853 ();
 sg13g2_decap_8 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_29_867 ();
 sg13g2_decap_4 FILLER_29_874 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_67 ();
 sg13g2_decap_4 FILLER_30_74 ();
 sg13g2_fill_1 FILLER_30_87 ();
 sg13g2_fill_2 FILLER_30_92 ();
 sg13g2_fill_1 FILLER_30_94 ();
 sg13g2_decap_8 FILLER_30_100 ();
 sg13g2_decap_8 FILLER_30_107 ();
 sg13g2_decap_8 FILLER_30_114 ();
 sg13g2_decap_4 FILLER_30_121 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_fill_2 FILLER_30_135 ();
 sg13g2_fill_1 FILLER_30_137 ();
 sg13g2_decap_8 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_150 ();
 sg13g2_decap_4 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_173 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_decap_4 FILLER_30_214 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_251 ();
 sg13g2_decap_8 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_decap_8 FILLER_30_276 ();
 sg13g2_decap_8 FILLER_30_283 ();
 sg13g2_decap_8 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_302 ();
 sg13g2_decap_4 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_decap_8 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_decap_4 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_4 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_4 FILLER_30_412 ();
 sg13g2_fill_1 FILLER_30_416 ();
 sg13g2_fill_1 FILLER_30_427 ();
 sg13g2_decap_4 FILLER_30_433 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_466 ();
 sg13g2_decap_8 FILLER_30_473 ();
 sg13g2_decap_8 FILLER_30_480 ();
 sg13g2_decap_8 FILLER_30_487 ();
 sg13g2_decap_8 FILLER_30_494 ();
 sg13g2_decap_4 FILLER_30_501 ();
 sg13g2_fill_2 FILLER_30_510 ();
 sg13g2_fill_1 FILLER_30_521 ();
 sg13g2_fill_2 FILLER_30_530 ();
 sg13g2_decap_8 FILLER_30_536 ();
 sg13g2_decap_8 FILLER_30_543 ();
 sg13g2_fill_2 FILLER_30_550 ();
 sg13g2_decap_8 FILLER_30_558 ();
 sg13g2_fill_2 FILLER_30_565 ();
 sg13g2_fill_1 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_576 ();
 sg13g2_decap_4 FILLER_30_583 ();
 sg13g2_fill_2 FILLER_30_591 ();
 sg13g2_fill_1 FILLER_30_593 ();
 sg13g2_decap_4 FILLER_30_604 ();
 sg13g2_fill_2 FILLER_30_608 ();
 sg13g2_fill_2 FILLER_30_615 ();
 sg13g2_fill_1 FILLER_30_637 ();
 sg13g2_decap_4 FILLER_30_648 ();
 sg13g2_fill_2 FILLER_30_652 ();
 sg13g2_decap_4 FILLER_30_659 ();
 sg13g2_fill_2 FILLER_30_663 ();
 sg13g2_decap_8 FILLER_30_669 ();
 sg13g2_decap_4 FILLER_30_676 ();
 sg13g2_decap_8 FILLER_30_684 ();
 sg13g2_decap_8 FILLER_30_691 ();
 sg13g2_decap_4 FILLER_30_698 ();
 sg13g2_fill_1 FILLER_30_702 ();
 sg13g2_decap_8 FILLER_30_711 ();
 sg13g2_decap_8 FILLER_30_718 ();
 sg13g2_fill_1 FILLER_30_725 ();
 sg13g2_decap_4 FILLER_30_731 ();
 sg13g2_fill_1 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_decap_8 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_30_868 ();
 sg13g2_fill_2 FILLER_30_875 ();
 sg13g2_fill_1 FILLER_30_877 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_fill_2 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_102 ();
 sg13g2_decap_4 FILLER_31_109 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_decap_8 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_129 ();
 sg13g2_fill_1 FILLER_31_136 ();
 sg13g2_decap_4 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_151 ();
 sg13g2_fill_2 FILLER_31_158 ();
 sg13g2_decap_8 FILLER_31_165 ();
 sg13g2_decap_4 FILLER_31_172 ();
 sg13g2_decap_4 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_205 ();
 sg13g2_decap_4 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_decap_8 FILLER_31_221 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_decap_8 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_264 ();
 sg13g2_decap_4 FILLER_31_271 ();
 sg13g2_decap_8 FILLER_31_279 ();
 sg13g2_decap_8 FILLER_31_286 ();
 sg13g2_fill_2 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_fill_1 FILLER_31_315 ();
 sg13g2_fill_1 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_decap_8 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_365 ();
 sg13g2_decap_4 FILLER_31_372 ();
 sg13g2_fill_1 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_4 FILLER_31_388 ();
 sg13g2_fill_1 FILLER_31_392 ();
 sg13g2_fill_1 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_1 FILLER_31_410 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_fill_1 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_474 ();
 sg13g2_fill_2 FILLER_31_481 ();
 sg13g2_decap_8 FILLER_31_492 ();
 sg13g2_fill_2 FILLER_31_499 ();
 sg13g2_fill_1 FILLER_31_501 ();
 sg13g2_decap_4 FILLER_31_508 ();
 sg13g2_fill_2 FILLER_31_525 ();
 sg13g2_fill_1 FILLER_31_527 ();
 sg13g2_fill_1 FILLER_31_537 ();
 sg13g2_decap_8 FILLER_31_544 ();
 sg13g2_decap_8 FILLER_31_551 ();
 sg13g2_decap_8 FILLER_31_558 ();
 sg13g2_fill_2 FILLER_31_565 ();
 sg13g2_decap_4 FILLER_31_572 ();
 sg13g2_fill_1 FILLER_31_576 ();
 sg13g2_decap_4 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_590 ();
 sg13g2_decap_4 FILLER_31_601 ();
 sg13g2_fill_2 FILLER_31_610 ();
 sg13g2_fill_1 FILLER_31_625 ();
 sg13g2_fill_1 FILLER_31_630 ();
 sg13g2_fill_2 FILLER_31_640 ();
 sg13g2_decap_8 FILLER_31_648 ();
 sg13g2_fill_1 FILLER_31_655 ();
 sg13g2_decap_4 FILLER_31_665 ();
 sg13g2_fill_1 FILLER_31_669 ();
 sg13g2_decap_8 FILLER_31_676 ();
 sg13g2_decap_4 FILLER_31_683 ();
 sg13g2_fill_1 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_698 ();
 sg13g2_decap_8 FILLER_31_705 ();
 sg13g2_decap_8 FILLER_31_712 ();
 sg13g2_decap_8 FILLER_31_719 ();
 sg13g2_decap_4 FILLER_31_726 ();
 sg13g2_fill_2 FILLER_31_730 ();
 sg13g2_fill_1 FILLER_31_745 ();
 sg13g2_fill_1 FILLER_31_751 ();
 sg13g2_decap_8 FILLER_31_758 ();
 sg13g2_decap_8 FILLER_31_765 ();
 sg13g2_decap_8 FILLER_31_772 ();
 sg13g2_decap_8 FILLER_31_779 ();
 sg13g2_decap_8 FILLER_31_786 ();
 sg13g2_decap_8 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_800 ();
 sg13g2_decap_8 FILLER_31_807 ();
 sg13g2_decap_8 FILLER_31_814 ();
 sg13g2_decap_8 FILLER_31_821 ();
 sg13g2_decap_8 FILLER_31_828 ();
 sg13g2_decap_8 FILLER_31_835 ();
 sg13g2_decap_8 FILLER_31_842 ();
 sg13g2_decap_8 FILLER_31_849 ();
 sg13g2_decap_8 FILLER_31_856 ();
 sg13g2_decap_8 FILLER_31_863 ();
 sg13g2_decap_8 FILLER_31_870 ();
 sg13g2_fill_1 FILLER_31_877 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_85 ();
 sg13g2_decap_8 FILLER_32_96 ();
 sg13g2_decap_8 FILLER_32_107 ();
 sg13g2_decap_8 FILLER_32_114 ();
 sg13g2_decap_8 FILLER_32_121 ();
 sg13g2_decap_4 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_decap_8 FILLER_32_142 ();
 sg13g2_fill_1 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_160 ();
 sg13g2_decap_8 FILLER_32_167 ();
 sg13g2_decap_8 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_4 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_253 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_269 ();
 sg13g2_decap_4 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_312 ();
 sg13g2_decap_4 FILLER_32_326 ();
 sg13g2_fill_2 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_fill_1 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_4 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_421 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_fill_1 FILLER_32_430 ();
 sg13g2_decap_8 FILLER_32_436 ();
 sg13g2_fill_2 FILLER_32_443 ();
 sg13g2_decap_4 FILLER_32_454 ();
 sg13g2_fill_2 FILLER_32_458 ();
 sg13g2_fill_1 FILLER_32_468 ();
 sg13g2_fill_2 FILLER_32_488 ();
 sg13g2_fill_1 FILLER_32_490 ();
 sg13g2_decap_8 FILLER_32_496 ();
 sg13g2_decap_8 FILLER_32_503 ();
 sg13g2_decap_8 FILLER_32_514 ();
 sg13g2_decap_4 FILLER_32_521 ();
 sg13g2_fill_1 FILLER_32_525 ();
 sg13g2_decap_8 FILLER_32_534 ();
 sg13g2_decap_8 FILLER_32_545 ();
 sg13g2_decap_8 FILLER_32_552 ();
 sg13g2_decap_8 FILLER_32_559 ();
 sg13g2_decap_8 FILLER_32_566 ();
 sg13g2_fill_1 FILLER_32_573 ();
 sg13g2_fill_2 FILLER_32_577 ();
 sg13g2_fill_1 FILLER_32_579 ();
 sg13g2_fill_2 FILLER_32_590 ();
 sg13g2_decap_8 FILLER_32_596 ();
 sg13g2_fill_2 FILLER_32_603 ();
 sg13g2_decap_8 FILLER_32_609 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_decap_4 FILLER_32_630 ();
 sg13g2_fill_1 FILLER_32_634 ();
 sg13g2_decap_8 FILLER_32_639 ();
 sg13g2_decap_8 FILLER_32_646 ();
 sg13g2_fill_1 FILLER_32_653 ();
 sg13g2_decap_8 FILLER_32_659 ();
 sg13g2_decap_8 FILLER_32_666 ();
 sg13g2_decap_8 FILLER_32_673 ();
 sg13g2_decap_8 FILLER_32_680 ();
 sg13g2_decap_8 FILLER_32_687 ();
 sg13g2_decap_4 FILLER_32_694 ();
 sg13g2_fill_2 FILLER_32_698 ();
 sg13g2_fill_2 FILLER_32_705 ();
 sg13g2_fill_1 FILLER_32_707 ();
 sg13g2_decap_8 FILLER_32_712 ();
 sg13g2_decap_8 FILLER_32_719 ();
 sg13g2_decap_4 FILLER_32_730 ();
 sg13g2_fill_1 FILLER_32_734 ();
 sg13g2_decap_4 FILLER_32_739 ();
 sg13g2_fill_1 FILLER_32_747 ();
 sg13g2_decap_8 FILLER_32_752 ();
 sg13g2_fill_2 FILLER_32_759 ();
 sg13g2_fill_1 FILLER_32_761 ();
 sg13g2_decap_8 FILLER_32_766 ();
 sg13g2_decap_8 FILLER_32_773 ();
 sg13g2_decap_8 FILLER_32_780 ();
 sg13g2_decap_8 FILLER_32_787 ();
 sg13g2_decap_8 FILLER_32_794 ();
 sg13g2_decap_8 FILLER_32_801 ();
 sg13g2_decap_8 FILLER_32_808 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_decap_8 FILLER_32_822 ();
 sg13g2_decap_8 FILLER_32_829 ();
 sg13g2_decap_8 FILLER_32_836 ();
 sg13g2_decap_8 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_850 ();
 sg13g2_decap_8 FILLER_32_857 ();
 sg13g2_decap_8 FILLER_32_864 ();
 sg13g2_decap_8 FILLER_32_871 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_fill_2 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_100 ();
 sg13g2_decap_8 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_114 ();
 sg13g2_decap_8 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_128 ();
 sg13g2_decap_8 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_157 ();
 sg13g2_decap_4 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_fill_2 FILLER_33_205 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_decap_8 FILLER_33_227 ();
 sg13g2_decap_8 FILLER_33_234 ();
 sg13g2_decap_8 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_253 ();
 sg13g2_decap_8 FILLER_33_260 ();
 sg13g2_decap_8 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_274 ();
 sg13g2_decap_4 FILLER_33_279 ();
 sg13g2_decap_4 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_4 FILLER_33_354 ();
 sg13g2_decap_4 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_4 FILLER_33_415 ();
 sg13g2_fill_2 FILLER_33_419 ();
 sg13g2_decap_8 FILLER_33_426 ();
 sg13g2_decap_8 FILLER_33_433 ();
 sg13g2_decap_8 FILLER_33_440 ();
 sg13g2_decap_8 FILLER_33_447 ();
 sg13g2_decap_8 FILLER_33_454 ();
 sg13g2_decap_8 FILLER_33_461 ();
 sg13g2_decap_8 FILLER_33_468 ();
 sg13g2_decap_8 FILLER_33_475 ();
 sg13g2_decap_8 FILLER_33_482 ();
 sg13g2_decap_8 FILLER_33_489 ();
 sg13g2_decap_8 FILLER_33_496 ();
 sg13g2_decap_8 FILLER_33_503 ();
 sg13g2_decap_4 FILLER_33_510 ();
 sg13g2_fill_2 FILLER_33_514 ();
 sg13g2_decap_4 FILLER_33_520 ();
 sg13g2_fill_2 FILLER_33_524 ();
 sg13g2_decap_8 FILLER_33_535 ();
 sg13g2_fill_2 FILLER_33_542 ();
 sg13g2_fill_1 FILLER_33_544 ();
 sg13g2_decap_8 FILLER_33_554 ();
 sg13g2_decap_8 FILLER_33_561 ();
 sg13g2_decap_4 FILLER_33_568 ();
 sg13g2_decap_8 FILLER_33_590 ();
 sg13g2_decap_8 FILLER_33_597 ();
 sg13g2_decap_4 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_623 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_fill_2 FILLER_33_637 ();
 sg13g2_fill_2 FILLER_33_645 ();
 sg13g2_fill_1 FILLER_33_647 ();
 sg13g2_decap_4 FILLER_33_661 ();
 sg13g2_decap_8 FILLER_33_668 ();
 sg13g2_decap_8 FILLER_33_675 ();
 sg13g2_decap_8 FILLER_33_696 ();
 sg13g2_decap_8 FILLER_33_703 ();
 sg13g2_decap_8 FILLER_33_710 ();
 sg13g2_decap_4 FILLER_33_717 ();
 sg13g2_fill_2 FILLER_33_721 ();
 sg13g2_decap_4 FILLER_33_732 ();
 sg13g2_decap_8 FILLER_33_745 ();
 sg13g2_decap_8 FILLER_33_752 ();
 sg13g2_decap_4 FILLER_33_759 ();
 sg13g2_decap_8 FILLER_33_768 ();
 sg13g2_decap_8 FILLER_33_775 ();
 sg13g2_decap_8 FILLER_33_782 ();
 sg13g2_decap_8 FILLER_33_789 ();
 sg13g2_decap_8 FILLER_33_796 ();
 sg13g2_decap_8 FILLER_33_803 ();
 sg13g2_decap_8 FILLER_33_810 ();
 sg13g2_decap_8 FILLER_33_817 ();
 sg13g2_decap_8 FILLER_33_824 ();
 sg13g2_decap_8 FILLER_33_831 ();
 sg13g2_decap_8 FILLER_33_838 ();
 sg13g2_decap_8 FILLER_33_845 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_decap_8 FILLER_33_859 ();
 sg13g2_decap_8 FILLER_33_866 ();
 sg13g2_decap_4 FILLER_33_873 ();
 sg13g2_fill_1 FILLER_33_877 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_63 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_decap_8 FILLER_34_72 ();
 sg13g2_decap_8 FILLER_34_79 ();
 sg13g2_decap_4 FILLER_34_86 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_decap_8 FILLER_34_94 ();
 sg13g2_decap_8 FILLER_34_101 ();
 sg13g2_decap_8 FILLER_34_108 ();
 sg13g2_decap_4 FILLER_34_115 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_137 ();
 sg13g2_decap_8 FILLER_34_143 ();
 sg13g2_fill_2 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_152 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_168 ();
 sg13g2_fill_1 FILLER_34_178 ();
 sg13g2_decap_8 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_200 ();
 sg13g2_fill_2 FILLER_34_207 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_fill_2 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_decap_4 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_288 ();
 sg13g2_decap_8 FILLER_34_295 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_fill_1 FILLER_34_304 ();
 sg13g2_fill_2 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_316 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_4 FILLER_34_357 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_fill_1 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_fill_2 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_415 ();
 sg13g2_decap_8 FILLER_34_422 ();
 sg13g2_decap_8 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_34_436 ();
 sg13g2_decap_4 FILLER_34_443 ();
 sg13g2_fill_2 FILLER_34_447 ();
 sg13g2_fill_2 FILLER_34_467 ();
 sg13g2_fill_1 FILLER_34_473 ();
 sg13g2_decap_4 FILLER_34_482 ();
 sg13g2_fill_2 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_496 ();
 sg13g2_decap_8 FILLER_34_503 ();
 sg13g2_decap_4 FILLER_34_510 ();
 sg13g2_fill_1 FILLER_34_514 ();
 sg13g2_decap_4 FILLER_34_519 ();
 sg13g2_fill_1 FILLER_34_523 ();
 sg13g2_fill_1 FILLER_34_529 ();
 sg13g2_fill_1 FILLER_34_543 ();
 sg13g2_decap_8 FILLER_34_548 ();
 sg13g2_decap_8 FILLER_34_555 ();
 sg13g2_decap_8 FILLER_34_562 ();
 sg13g2_decap_4 FILLER_34_569 ();
 sg13g2_fill_2 FILLER_34_573 ();
 sg13g2_decap_8 FILLER_34_586 ();
 sg13g2_decap_8 FILLER_34_593 ();
 sg13g2_fill_2 FILLER_34_600 ();
 sg13g2_fill_2 FILLER_34_606 ();
 sg13g2_decap_4 FILLER_34_613 ();
 sg13g2_fill_2 FILLER_34_617 ();
 sg13g2_decap_8 FILLER_34_623 ();
 sg13g2_fill_2 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_636 ();
 sg13g2_fill_2 FILLER_34_643 ();
 sg13g2_fill_2 FILLER_34_649 ();
 sg13g2_fill_1 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_656 ();
 sg13g2_decap_8 FILLER_34_663 ();
 sg13g2_decap_8 FILLER_34_670 ();
 sg13g2_decap_8 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_691 ();
 sg13g2_decap_8 FILLER_34_698 ();
 sg13g2_decap_8 FILLER_34_709 ();
 sg13g2_decap_8 FILLER_34_716 ();
 sg13g2_fill_2 FILLER_34_723 ();
 sg13g2_fill_1 FILLER_34_725 ();
 sg13g2_decap_4 FILLER_34_732 ();
 sg13g2_fill_2 FILLER_34_736 ();
 sg13g2_fill_1 FILLER_34_742 ();
 sg13g2_decap_4 FILLER_34_750 ();
 sg13g2_fill_1 FILLER_34_754 ();
 sg13g2_decap_8 FILLER_34_759 ();
 sg13g2_decap_8 FILLER_34_766 ();
 sg13g2_decap_8 FILLER_34_773 ();
 sg13g2_decap_8 FILLER_34_780 ();
 sg13g2_decap_8 FILLER_34_787 ();
 sg13g2_decap_8 FILLER_34_794 ();
 sg13g2_decap_8 FILLER_34_801 ();
 sg13g2_decap_8 FILLER_34_808 ();
 sg13g2_decap_8 FILLER_34_815 ();
 sg13g2_decap_8 FILLER_34_822 ();
 sg13g2_decap_8 FILLER_34_829 ();
 sg13g2_decap_8 FILLER_34_836 ();
 sg13g2_decap_8 FILLER_34_843 ();
 sg13g2_decap_8 FILLER_34_850 ();
 sg13g2_decap_8 FILLER_34_857 ();
 sg13g2_decap_8 FILLER_34_864 ();
 sg13g2_decap_8 FILLER_34_871 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_72 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_88 ();
 sg13g2_fill_2 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_104 ();
 sg13g2_decap_8 FILLER_35_111 ();
 sg13g2_decap_4 FILLER_35_130 ();
 sg13g2_decap_4 FILLER_35_139 ();
 sg13g2_fill_2 FILLER_35_143 ();
 sg13g2_decap_4 FILLER_35_150 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_decap_4 FILLER_35_182 ();
 sg13g2_fill_2 FILLER_35_186 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_decap_4 FILLER_35_206 ();
 sg13g2_decap_8 FILLER_35_220 ();
 sg13g2_decap_8 FILLER_35_227 ();
 sg13g2_fill_2 FILLER_35_234 ();
 sg13g2_decap_4 FILLER_35_240 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_decap_8 FILLER_35_257 ();
 sg13g2_decap_4 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_decap_8 FILLER_35_275 ();
 sg13g2_decap_8 FILLER_35_286 ();
 sg13g2_decap_8 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_308 ();
 sg13g2_decap_4 FILLER_35_327 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_decap_4 FILLER_35_337 ();
 sg13g2_decap_4 FILLER_35_349 ();
 sg13g2_fill_2 FILLER_35_353 ();
 sg13g2_fill_2 FILLER_35_359 ();
 sg13g2_fill_2 FILLER_35_370 ();
 sg13g2_decap_4 FILLER_35_376 ();
 sg13g2_fill_2 FILLER_35_385 ();
 sg13g2_fill_1 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_1 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_35_417 ();
 sg13g2_decap_8 FILLER_35_436 ();
 sg13g2_decap_8 FILLER_35_443 ();
 sg13g2_decap_8 FILLER_35_450 ();
 sg13g2_decap_8 FILLER_35_457 ();
 sg13g2_decap_4 FILLER_35_464 ();
 sg13g2_decap_8 FILLER_35_473 ();
 sg13g2_decap_4 FILLER_35_480 ();
 sg13g2_decap_8 FILLER_35_489 ();
 sg13g2_decap_8 FILLER_35_496 ();
 sg13g2_decap_8 FILLER_35_507 ();
 sg13g2_decap_8 FILLER_35_514 ();
 sg13g2_fill_2 FILLER_35_521 ();
 sg13g2_decap_8 FILLER_35_532 ();
 sg13g2_fill_2 FILLER_35_539 ();
 sg13g2_fill_1 FILLER_35_541 ();
 sg13g2_decap_8 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_decap_8 FILLER_35_560 ();
 sg13g2_decap_4 FILLER_35_567 ();
 sg13g2_decap_4 FILLER_35_579 ();
 sg13g2_fill_1 FILLER_35_583 ();
 sg13g2_decap_4 FILLER_35_601 ();
 sg13g2_fill_1 FILLER_35_605 ();
 sg13g2_fill_2 FILLER_35_611 ();
 sg13g2_decap_8 FILLER_35_617 ();
 sg13g2_decap_8 FILLER_35_624 ();
 sg13g2_decap_8 FILLER_35_631 ();
 sg13g2_decap_4 FILLER_35_638 ();
 sg13g2_decap_8 FILLER_35_650 ();
 sg13g2_decap_4 FILLER_35_657 ();
 sg13g2_decap_8 FILLER_35_666 ();
 sg13g2_decap_8 FILLER_35_673 ();
 sg13g2_decap_8 FILLER_35_680 ();
 sg13g2_decap_8 FILLER_35_687 ();
 sg13g2_fill_1 FILLER_35_694 ();
 sg13g2_decap_4 FILLER_35_699 ();
 sg13g2_fill_2 FILLER_35_703 ();
 sg13g2_decap_8 FILLER_35_710 ();
 sg13g2_fill_1 FILLER_35_717 ();
 sg13g2_decap_4 FILLER_35_722 ();
 sg13g2_fill_1 FILLER_35_726 ();
 sg13g2_fill_2 FILLER_35_731 ();
 sg13g2_fill_1 FILLER_35_733 ();
 sg13g2_decap_8 FILLER_35_743 ();
 sg13g2_fill_2 FILLER_35_750 ();
 sg13g2_decap_4 FILLER_35_761 ();
 sg13g2_fill_1 FILLER_35_765 ();
 sg13g2_decap_8 FILLER_35_779 ();
 sg13g2_decap_8 FILLER_35_786 ();
 sg13g2_decap_8 FILLER_35_793 ();
 sg13g2_decap_8 FILLER_35_800 ();
 sg13g2_decap_8 FILLER_35_807 ();
 sg13g2_decap_8 FILLER_35_814 ();
 sg13g2_decap_8 FILLER_35_821 ();
 sg13g2_decap_8 FILLER_35_828 ();
 sg13g2_decap_8 FILLER_35_835 ();
 sg13g2_decap_8 FILLER_35_842 ();
 sg13g2_decap_8 FILLER_35_849 ();
 sg13g2_decap_8 FILLER_35_856 ();
 sg13g2_decap_8 FILLER_35_863 ();
 sg13g2_decap_8 FILLER_35_870 ();
 sg13g2_fill_1 FILLER_35_877 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_60 ();
 sg13g2_fill_2 FILLER_36_85 ();
 sg13g2_fill_1 FILLER_36_87 ();
 sg13g2_decap_8 FILLER_36_97 ();
 sg13g2_fill_2 FILLER_36_104 ();
 sg13g2_fill_1 FILLER_36_106 ();
 sg13g2_decap_4 FILLER_36_111 ();
 sg13g2_fill_1 FILLER_36_134 ();
 sg13g2_decap_8 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_decap_8 FILLER_36_160 ();
 sg13g2_decap_8 FILLER_36_167 ();
 sg13g2_decap_8 FILLER_36_174 ();
 sg13g2_decap_8 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_decap_4 FILLER_36_219 ();
 sg13g2_decap_4 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_239 ();
 sg13g2_decap_8 FILLER_36_264 ();
 sg13g2_decap_4 FILLER_36_271 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_288 ();
 sg13g2_decap_8 FILLER_36_295 ();
 sg13g2_decap_4 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_337 ();
 sg13g2_decap_8 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_351 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_decap_4 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_4 FILLER_36_401 ();
 sg13g2_fill_2 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_36_412 ();
 sg13g2_decap_8 FILLER_36_419 ();
 sg13g2_decap_4 FILLER_36_426 ();
 sg13g2_fill_2 FILLER_36_430 ();
 sg13g2_decap_8 FILLER_36_437 ();
 sg13g2_decap_4 FILLER_36_444 ();
 sg13g2_fill_1 FILLER_36_448 ();
 sg13g2_decap_8 FILLER_36_457 ();
 sg13g2_decap_8 FILLER_36_464 ();
 sg13g2_decap_8 FILLER_36_471 ();
 sg13g2_decap_8 FILLER_36_478 ();
 sg13g2_decap_8 FILLER_36_489 ();
 sg13g2_decap_8 FILLER_36_496 ();
 sg13g2_decap_8 FILLER_36_503 ();
 sg13g2_decap_8 FILLER_36_510 ();
 sg13g2_decap_8 FILLER_36_517 ();
 sg13g2_decap_8 FILLER_36_524 ();
 sg13g2_fill_2 FILLER_36_531 ();
 sg13g2_decap_8 FILLER_36_538 ();
 sg13g2_fill_2 FILLER_36_545 ();
 sg13g2_fill_1 FILLER_36_547 ();
 sg13g2_decap_8 FILLER_36_552 ();
 sg13g2_decap_8 FILLER_36_559 ();
 sg13g2_decap_8 FILLER_36_566 ();
 sg13g2_decap_8 FILLER_36_573 ();
 sg13g2_decap_4 FILLER_36_580 ();
 sg13g2_fill_1 FILLER_36_584 ();
 sg13g2_decap_4 FILLER_36_598 ();
 sg13g2_decap_4 FILLER_36_616 ();
 sg13g2_fill_1 FILLER_36_620 ();
 sg13g2_fill_2 FILLER_36_636 ();
 sg13g2_fill_2 FILLER_36_644 ();
 sg13g2_fill_2 FILLER_36_651 ();
 sg13g2_decap_8 FILLER_36_657 ();
 sg13g2_decap_4 FILLER_36_664 ();
 sg13g2_fill_1 FILLER_36_668 ();
 sg13g2_decap_8 FILLER_36_673 ();
 sg13g2_decap_8 FILLER_36_680 ();
 sg13g2_decap_8 FILLER_36_687 ();
 sg13g2_fill_1 FILLER_36_694 ();
 sg13g2_fill_1 FILLER_36_710 ();
 sg13g2_fill_1 FILLER_36_720 ();
 sg13g2_decap_4 FILLER_36_726 ();
 sg13g2_fill_2 FILLER_36_730 ();
 sg13g2_decap_4 FILLER_36_738 ();
 sg13g2_fill_2 FILLER_36_742 ();
 sg13g2_fill_1 FILLER_36_749 ();
 sg13g2_decap_8 FILLER_36_755 ();
 sg13g2_decap_8 FILLER_36_762 ();
 sg13g2_decap_8 FILLER_36_769 ();
 sg13g2_decap_8 FILLER_36_776 ();
 sg13g2_decap_8 FILLER_36_783 ();
 sg13g2_decap_8 FILLER_36_790 ();
 sg13g2_decap_8 FILLER_36_797 ();
 sg13g2_decap_8 FILLER_36_804 ();
 sg13g2_decap_8 FILLER_36_811 ();
 sg13g2_decap_8 FILLER_36_818 ();
 sg13g2_decap_8 FILLER_36_825 ();
 sg13g2_decap_8 FILLER_36_832 ();
 sg13g2_decap_8 FILLER_36_839 ();
 sg13g2_decap_8 FILLER_36_846 ();
 sg13g2_decap_8 FILLER_36_853 ();
 sg13g2_decap_8 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_36_867 ();
 sg13g2_decap_4 FILLER_36_874 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_4 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_60 ();
 sg13g2_fill_1 FILLER_37_66 ();
 sg13g2_fill_2 FILLER_37_87 ();
 sg13g2_fill_2 FILLER_37_93 ();
 sg13g2_fill_1 FILLER_37_95 ();
 sg13g2_decap_8 FILLER_37_99 ();
 sg13g2_decap_8 FILLER_37_106 ();
 sg13g2_fill_2 FILLER_37_113 ();
 sg13g2_fill_1 FILLER_37_115 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_4 FILLER_37_189 ();
 sg13g2_decap_4 FILLER_37_198 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_decap_8 FILLER_37_216 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_decap_4 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_234 ();
 sg13g2_decap_4 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_fill_2 FILLER_37_253 ();
 sg13g2_fill_2 FILLER_37_265 ();
 sg13g2_decap_4 FILLER_37_283 ();
 sg13g2_decap_8 FILLER_37_291 ();
 sg13g2_decap_8 FILLER_37_298 ();
 sg13g2_decap_8 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_4 FILLER_37_353 ();
 sg13g2_fill_1 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_8 FILLER_37_403 ();
 sg13g2_decap_8 FILLER_37_410 ();
 sg13g2_decap_8 FILLER_37_417 ();
 sg13g2_fill_1 FILLER_37_428 ();
 sg13g2_decap_4 FILLER_37_434 ();
 sg13g2_fill_2 FILLER_37_438 ();
 sg13g2_decap_4 FILLER_37_445 ();
 sg13g2_fill_2 FILLER_37_449 ();
 sg13g2_decap_8 FILLER_37_463 ();
 sg13g2_decap_8 FILLER_37_470 ();
 sg13g2_decap_8 FILLER_37_477 ();
 sg13g2_fill_2 FILLER_37_484 ();
 sg13g2_fill_1 FILLER_37_486 ();
 sg13g2_decap_8 FILLER_37_491 ();
 sg13g2_fill_2 FILLER_37_498 ();
 sg13g2_decap_8 FILLER_37_515 ();
 sg13g2_decap_8 FILLER_37_522 ();
 sg13g2_decap_8 FILLER_37_534 ();
 sg13g2_fill_2 FILLER_37_541 ();
 sg13g2_fill_1 FILLER_37_543 ();
 sg13g2_decap_8 FILLER_37_548 ();
 sg13g2_decap_8 FILLER_37_555 ();
 sg13g2_decap_4 FILLER_37_562 ();
 sg13g2_fill_2 FILLER_37_576 ();
 sg13g2_fill_1 FILLER_37_578 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_fill_2 FILLER_37_602 ();
 sg13g2_fill_2 FILLER_37_609 ();
 sg13g2_fill_1 FILLER_37_611 ();
 sg13g2_fill_2 FILLER_37_617 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_fill_1 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_643 ();
 sg13g2_decap_4 FILLER_37_658 ();
 sg13g2_fill_1 FILLER_37_662 ();
 sg13g2_decap_8 FILLER_37_674 ();
 sg13g2_decap_8 FILLER_37_681 ();
 sg13g2_decap_8 FILLER_37_688 ();
 sg13g2_decap_4 FILLER_37_695 ();
 sg13g2_decap_8 FILLER_37_713 ();
 sg13g2_decap_8 FILLER_37_720 ();
 sg13g2_decap_8 FILLER_37_727 ();
 sg13g2_decap_8 FILLER_37_734 ();
 sg13g2_decap_4 FILLER_37_746 ();
 sg13g2_fill_1 FILLER_37_750 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_decap_8 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_37_868 ();
 sg13g2_fill_2 FILLER_37_875 ();
 sg13g2_fill_1 FILLER_37_877 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_4 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_67 ();
 sg13g2_fill_2 FILLER_38_78 ();
 sg13g2_decap_4 FILLER_38_86 ();
 sg13g2_fill_1 FILLER_38_90 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_97 ();
 sg13g2_decap_8 FILLER_38_111 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_128 ();
 sg13g2_decap_4 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_146 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_decap_8 FILLER_38_158 ();
 sg13g2_decap_8 FILLER_38_165 ();
 sg13g2_fill_2 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_174 ();
 sg13g2_decap_4 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_fill_1 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_226 ();
 sg13g2_decap_4 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_258 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_decap_8 FILLER_38_288 ();
 sg13g2_decap_8 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_302 ();
 sg13g2_fill_2 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_fill_1 FILLER_38_363 ();
 sg13g2_decap_4 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_fill_2 FILLER_38_413 ();
 sg13g2_decap_4 FILLER_38_419 ();
 sg13g2_fill_1 FILLER_38_423 ();
 sg13g2_decap_4 FILLER_38_428 ();
 sg13g2_fill_1 FILLER_38_450 ();
 sg13g2_decap_8 FILLER_38_454 ();
 sg13g2_decap_8 FILLER_38_461 ();
 sg13g2_decap_8 FILLER_38_468 ();
 sg13g2_decap_8 FILLER_38_475 ();
 sg13g2_decap_8 FILLER_38_482 ();
 sg13g2_decap_8 FILLER_38_489 ();
 sg13g2_fill_1 FILLER_38_496 ();
 sg13g2_decap_4 FILLER_38_505 ();
 sg13g2_fill_2 FILLER_38_509 ();
 sg13g2_decap_8 FILLER_38_521 ();
 sg13g2_decap_8 FILLER_38_528 ();
 sg13g2_decap_8 FILLER_38_535 ();
 sg13g2_decap_4 FILLER_38_542 ();
 sg13g2_fill_1 FILLER_38_546 ();
 sg13g2_decap_4 FILLER_38_552 ();
 sg13g2_fill_2 FILLER_38_556 ();
 sg13g2_decap_8 FILLER_38_562 ();
 sg13g2_decap_8 FILLER_38_569 ();
 sg13g2_decap_8 FILLER_38_576 ();
 sg13g2_decap_8 FILLER_38_588 ();
 sg13g2_decap_8 FILLER_38_595 ();
 sg13g2_decap_4 FILLER_38_602 ();
 sg13g2_fill_2 FILLER_38_615 ();
 sg13g2_decap_8 FILLER_38_622 ();
 sg13g2_decap_4 FILLER_38_629 ();
 sg13g2_decap_4 FILLER_38_641 ();
 sg13g2_fill_2 FILLER_38_645 ();
 sg13g2_decap_8 FILLER_38_652 ();
 sg13g2_decap_8 FILLER_38_659 ();
 sg13g2_decap_4 FILLER_38_666 ();
 sg13g2_fill_2 FILLER_38_670 ();
 sg13g2_decap_8 FILLER_38_682 ();
 sg13g2_decap_4 FILLER_38_689 ();
 sg13g2_fill_2 FILLER_38_693 ();
 sg13g2_decap_4 FILLER_38_700 ();
 sg13g2_fill_1 FILLER_38_704 ();
 sg13g2_decap_8 FILLER_38_708 ();
 sg13g2_decap_4 FILLER_38_715 ();
 sg13g2_fill_1 FILLER_38_719 ();
 sg13g2_fill_1 FILLER_38_725 ();
 sg13g2_fill_1 FILLER_38_731 ();
 sg13g2_decap_8 FILLER_38_736 ();
 sg13g2_fill_1 FILLER_38_743 ();
 sg13g2_decap_4 FILLER_38_753 ();
 sg13g2_decap_8 FILLER_38_762 ();
 sg13g2_decap_8 FILLER_38_769 ();
 sg13g2_fill_1 FILLER_38_776 ();
 sg13g2_decap_8 FILLER_38_782 ();
 sg13g2_decap_8 FILLER_38_789 ();
 sg13g2_decap_8 FILLER_38_796 ();
 sg13g2_decap_8 FILLER_38_803 ();
 sg13g2_decap_8 FILLER_38_810 ();
 sg13g2_decap_8 FILLER_38_817 ();
 sg13g2_decap_8 FILLER_38_824 ();
 sg13g2_decap_8 FILLER_38_831 ();
 sg13g2_decap_8 FILLER_38_838 ();
 sg13g2_decap_8 FILLER_38_845 ();
 sg13g2_decap_8 FILLER_38_852 ();
 sg13g2_decap_8 FILLER_38_859 ();
 sg13g2_decap_8 FILLER_38_866 ();
 sg13g2_decap_4 FILLER_38_873 ();
 sg13g2_fill_1 FILLER_38_877 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_4 FILLER_39_49 ();
 sg13g2_fill_2 FILLER_39_53 ();
 sg13g2_fill_1 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_76 ();
 sg13g2_fill_1 FILLER_39_83 ();
 sg13g2_fill_1 FILLER_39_89 ();
 sg13g2_decap_4 FILLER_39_95 ();
 sg13g2_fill_1 FILLER_39_99 ();
 sg13g2_fill_1 FILLER_39_115 ();
 sg13g2_decap_8 FILLER_39_121 ();
 sg13g2_fill_1 FILLER_39_128 ();
 sg13g2_decap_8 FILLER_39_144 ();
 sg13g2_fill_2 FILLER_39_151 ();
 sg13g2_fill_1 FILLER_39_153 ();
 sg13g2_decap_8 FILLER_39_163 ();
 sg13g2_fill_1 FILLER_39_170 ();
 sg13g2_decap_8 FILLER_39_183 ();
 sg13g2_decap_8 FILLER_39_190 ();
 sg13g2_decap_8 FILLER_39_197 ();
 sg13g2_decap_8 FILLER_39_204 ();
 sg13g2_decap_8 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_227 ();
 sg13g2_fill_2 FILLER_39_234 ();
 sg13g2_fill_2 FILLER_39_241 ();
 sg13g2_fill_1 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_249 ();
 sg13g2_fill_1 FILLER_39_251 ();
 sg13g2_fill_1 FILLER_39_256 ();
 sg13g2_fill_1 FILLER_39_266 ();
 sg13g2_fill_1 FILLER_39_272 ();
 sg13g2_fill_2 FILLER_39_278 ();
 sg13g2_decap_8 FILLER_39_285 ();
 sg13g2_fill_2 FILLER_39_292 ();
 sg13g2_decap_8 FILLER_39_304 ();
 sg13g2_fill_2 FILLER_39_311 ();
 sg13g2_decap_4 FILLER_39_316 ();
 sg13g2_fill_1 FILLER_39_320 ();
 sg13g2_decap_8 FILLER_39_330 ();
 sg13g2_decap_8 FILLER_39_337 ();
 sg13g2_decap_8 FILLER_39_344 ();
 sg13g2_decap_8 FILLER_39_351 ();
 sg13g2_fill_2 FILLER_39_358 ();
 sg13g2_decap_4 FILLER_39_370 ();
 sg13g2_fill_1 FILLER_39_379 ();
 sg13g2_fill_2 FILLER_39_385 ();
 sg13g2_fill_2 FILLER_39_392 ();
 sg13g2_fill_2 FILLER_39_399 ();
 sg13g2_decap_4 FILLER_39_411 ();
 sg13g2_fill_2 FILLER_39_415 ();
 sg13g2_fill_1 FILLER_39_422 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_4 FILLER_39_434 ();
 sg13g2_fill_1 FILLER_39_438 ();
 sg13g2_decap_4 FILLER_39_444 ();
 sg13g2_decap_8 FILLER_39_452 ();
 sg13g2_decap_4 FILLER_39_459 ();
 sg13g2_fill_2 FILLER_39_463 ();
 sg13g2_decap_8 FILLER_39_470 ();
 sg13g2_decap_8 FILLER_39_477 ();
 sg13g2_decap_4 FILLER_39_484 ();
 sg13g2_fill_2 FILLER_39_488 ();
 sg13g2_decap_8 FILLER_39_499 ();
 sg13g2_fill_2 FILLER_39_506 ();
 sg13g2_fill_1 FILLER_39_508 ();
 sg13g2_decap_4 FILLER_39_515 ();
 sg13g2_decap_8 FILLER_39_537 ();
 sg13g2_fill_2 FILLER_39_544 ();
 sg13g2_fill_2 FILLER_39_551 ();
 sg13g2_decap_4 FILLER_39_558 ();
 sg13g2_fill_1 FILLER_39_562 ();
 sg13g2_decap_8 FILLER_39_568 ();
 sg13g2_fill_1 FILLER_39_575 ();
 sg13g2_fill_2 FILLER_39_581 ();
 sg13g2_fill_2 FILLER_39_590 ();
 sg13g2_fill_1 FILLER_39_592 ();
 sg13g2_decap_4 FILLER_39_597 ();
 sg13g2_decap_8 FILLER_39_608 ();
 sg13g2_decap_8 FILLER_39_615 ();
 sg13g2_decap_8 FILLER_39_622 ();
 sg13g2_decap_8 FILLER_39_629 ();
 sg13g2_fill_2 FILLER_39_636 ();
 sg13g2_decap_4 FILLER_39_642 ();
 sg13g2_fill_1 FILLER_39_646 ();
 sg13g2_decap_8 FILLER_39_652 ();
 sg13g2_decap_8 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_672 ();
 sg13g2_decap_8 FILLER_39_679 ();
 sg13g2_decap_4 FILLER_39_686 ();
 sg13g2_fill_1 FILLER_39_690 ();
 sg13g2_decap_4 FILLER_39_701 ();
 sg13g2_fill_1 FILLER_39_705 ();
 sg13g2_fill_2 FILLER_39_738 ();
 sg13g2_fill_2 FILLER_39_748 ();
 sg13g2_fill_1 FILLER_39_750 ();
 sg13g2_fill_2 FILLER_39_756 ();
 sg13g2_decap_4 FILLER_39_769 ();
 sg13g2_fill_1 FILLER_39_773 ();
 sg13g2_decap_4 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_788 ();
 sg13g2_decap_8 FILLER_39_795 ();
 sg13g2_decap_8 FILLER_39_802 ();
 sg13g2_decap_8 FILLER_39_809 ();
 sg13g2_decap_8 FILLER_39_816 ();
 sg13g2_decap_8 FILLER_39_823 ();
 sg13g2_decap_8 FILLER_39_830 ();
 sg13g2_decap_8 FILLER_39_837 ();
 sg13g2_decap_8 FILLER_39_844 ();
 sg13g2_decap_8 FILLER_39_851 ();
 sg13g2_decap_8 FILLER_39_858 ();
 sg13g2_decap_8 FILLER_39_865 ();
 sg13g2_decap_4 FILLER_39_872 ();
 sg13g2_fill_2 FILLER_39_876 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_4 FILLER_40_70 ();
 sg13g2_fill_2 FILLER_40_74 ();
 sg13g2_decap_8 FILLER_40_80 ();
 sg13g2_decap_8 FILLER_40_87 ();
 sg13g2_decap_8 FILLER_40_99 ();
 sg13g2_fill_1 FILLER_40_106 ();
 sg13g2_decap_8 FILLER_40_116 ();
 sg13g2_decap_8 FILLER_40_123 ();
 sg13g2_decap_8 FILLER_40_130 ();
 sg13g2_decap_8 FILLER_40_137 ();
 sg13g2_decap_8 FILLER_40_144 ();
 sg13g2_fill_1 FILLER_40_151 ();
 sg13g2_decap_8 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_164 ();
 sg13g2_fill_1 FILLER_40_166 ();
 sg13g2_decap_4 FILLER_40_171 ();
 sg13g2_decap_8 FILLER_40_192 ();
 sg13g2_decap_8 FILLER_40_199 ();
 sg13g2_decap_8 FILLER_40_206 ();
 sg13g2_decap_8 FILLER_40_213 ();
 sg13g2_decap_8 FILLER_40_220 ();
 sg13g2_decap_8 FILLER_40_227 ();
 sg13g2_decap_8 FILLER_40_234 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_4 FILLER_40_252 ();
 sg13g2_fill_1 FILLER_40_256 ();
 sg13g2_decap_4 FILLER_40_261 ();
 sg13g2_decap_8 FILLER_40_269 ();
 sg13g2_decap_8 FILLER_40_276 ();
 sg13g2_decap_8 FILLER_40_283 ();
 sg13g2_decap_8 FILLER_40_290 ();
 sg13g2_decap_8 FILLER_40_297 ();
 sg13g2_decap_8 FILLER_40_307 ();
 sg13g2_decap_8 FILLER_40_314 ();
 sg13g2_decap_8 FILLER_40_321 ();
 sg13g2_decap_8 FILLER_40_328 ();
 sg13g2_decap_8 FILLER_40_335 ();
 sg13g2_decap_8 FILLER_40_342 ();
 sg13g2_decap_8 FILLER_40_349 ();
 sg13g2_decap_8 FILLER_40_356 ();
 sg13g2_decap_8 FILLER_40_363 ();
 sg13g2_decap_8 FILLER_40_382 ();
 sg13g2_fill_1 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_395 ();
 sg13g2_fill_1 FILLER_40_402 ();
 sg13g2_decap_8 FILLER_40_411 ();
 sg13g2_fill_2 FILLER_40_418 ();
 sg13g2_decap_4 FILLER_40_424 ();
 sg13g2_fill_2 FILLER_40_428 ();
 sg13g2_decap_4 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_456 ();
 sg13g2_fill_1 FILLER_40_463 ();
 sg13g2_fill_2 FILLER_40_469 ();
 sg13g2_fill_1 FILLER_40_471 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_fill_2 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_505 ();
 sg13g2_decap_8 FILLER_40_512 ();
 sg13g2_decap_4 FILLER_40_524 ();
 sg13g2_fill_2 FILLER_40_528 ();
 sg13g2_fill_2 FILLER_40_534 ();
 sg13g2_fill_1 FILLER_40_536 ();
 sg13g2_fill_1 FILLER_40_543 ();
 sg13g2_decap_8 FILLER_40_549 ();
 sg13g2_decap_4 FILLER_40_556 ();
 sg13g2_fill_1 FILLER_40_560 ();
 sg13g2_decap_4 FILLER_40_570 ();
 sg13g2_fill_2 FILLER_40_579 ();
 sg13g2_fill_2 FILLER_40_586 ();
 sg13g2_fill_1 FILLER_40_592 ();
 sg13g2_fill_1 FILLER_40_597 ();
 sg13g2_decap_8 FILLER_40_602 ();
 sg13g2_decap_8 FILLER_40_609 ();
 sg13g2_decap_8 FILLER_40_616 ();
 sg13g2_fill_2 FILLER_40_627 ();
 sg13g2_fill_1 FILLER_40_629 ();
 sg13g2_fill_1 FILLER_40_635 ();
 sg13g2_fill_1 FILLER_40_651 ();
 sg13g2_fill_1 FILLER_40_657 ();
 sg13g2_fill_1 FILLER_40_663 ();
 sg13g2_fill_1 FILLER_40_669 ();
 sg13g2_decap_4 FILLER_40_674 ();
 sg13g2_decap_8 FILLER_40_683 ();
 sg13g2_decap_4 FILLER_40_690 ();
 sg13g2_fill_1 FILLER_40_698 ();
 sg13g2_decap_8 FILLER_40_707 ();
 sg13g2_fill_2 FILLER_40_714 ();
 sg13g2_fill_1 FILLER_40_724 ();
 sg13g2_decap_8 FILLER_40_735 ();
 sg13g2_decap_8 FILLER_40_750 ();
 sg13g2_decap_8 FILLER_40_757 ();
 sg13g2_decap_8 FILLER_40_764 ();
 sg13g2_decap_8 FILLER_40_771 ();
 sg13g2_decap_8 FILLER_40_786 ();
 sg13g2_decap_8 FILLER_40_793 ();
 sg13g2_decap_8 FILLER_40_800 ();
 sg13g2_decap_8 FILLER_40_807 ();
 sg13g2_decap_8 FILLER_40_814 ();
 sg13g2_decap_8 FILLER_40_821 ();
 sg13g2_decap_8 FILLER_40_828 ();
 sg13g2_decap_8 FILLER_40_835 ();
 sg13g2_decap_8 FILLER_40_842 ();
 sg13g2_decap_8 FILLER_40_849 ();
 sg13g2_decap_8 FILLER_40_856 ();
 sg13g2_decap_8 FILLER_40_863 ();
 sg13g2_decap_8 FILLER_40_870 ();
 sg13g2_fill_1 FILLER_40_877 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_4 FILLER_41_49 ();
 sg13g2_fill_1 FILLER_41_53 ();
 sg13g2_decap_8 FILLER_41_58 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_decap_4 FILLER_41_75 ();
 sg13g2_fill_2 FILLER_41_79 ();
 sg13g2_decap_8 FILLER_41_86 ();
 sg13g2_decap_8 FILLER_41_93 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_fill_1 FILLER_41_122 ();
 sg13g2_decap_4 FILLER_41_127 ();
 sg13g2_fill_1 FILLER_41_131 ();
 sg13g2_decap_4 FILLER_41_137 ();
 sg13g2_fill_2 FILLER_41_153 ();
 sg13g2_decap_8 FILLER_41_159 ();
 sg13g2_decap_8 FILLER_41_166 ();
 sg13g2_fill_1 FILLER_41_173 ();
 sg13g2_decap_4 FILLER_41_187 ();
 sg13g2_decap_8 FILLER_41_195 ();
 sg13g2_decap_8 FILLER_41_202 ();
 sg13g2_decap_4 FILLER_41_209 ();
 sg13g2_fill_2 FILLER_41_213 ();
 sg13g2_decap_8 FILLER_41_227 ();
 sg13g2_decap_8 FILLER_41_234 ();
 sg13g2_decap_8 FILLER_41_241 ();
 sg13g2_decap_8 FILLER_41_248 ();
 sg13g2_decap_4 FILLER_41_255 ();
 sg13g2_fill_2 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_265 ();
 sg13g2_decap_8 FILLER_41_272 ();
 sg13g2_decap_8 FILLER_41_279 ();
 sg13g2_decap_8 FILLER_41_286 ();
 sg13g2_fill_1 FILLER_41_305 ();
 sg13g2_decap_8 FILLER_41_311 ();
 sg13g2_fill_2 FILLER_41_318 ();
 sg13g2_decap_8 FILLER_41_325 ();
 sg13g2_decap_4 FILLER_41_332 ();
 sg13g2_decap_8 FILLER_41_341 ();
 sg13g2_decap_8 FILLER_41_348 ();
 sg13g2_fill_2 FILLER_41_355 ();
 sg13g2_fill_1 FILLER_41_357 ();
 sg13g2_fill_2 FILLER_41_367 ();
 sg13g2_fill_1 FILLER_41_382 ();
 sg13g2_fill_2 FILLER_41_386 ();
 sg13g2_decap_4 FILLER_41_395 ();
 sg13g2_fill_2 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_41_412 ();
 sg13g2_decap_8 FILLER_41_424 ();
 sg13g2_decap_8 FILLER_41_431 ();
 sg13g2_fill_2 FILLER_41_438 ();
 sg13g2_decap_8 FILLER_41_453 ();
 sg13g2_fill_1 FILLER_41_460 ();
 sg13g2_decap_8 FILLER_41_466 ();
 sg13g2_decap_8 FILLER_41_473 ();
 sg13g2_fill_2 FILLER_41_480 ();
 sg13g2_fill_1 FILLER_41_482 ();
 sg13g2_fill_1 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_503 ();
 sg13g2_fill_2 FILLER_41_510 ();
 sg13g2_fill_1 FILLER_41_512 ();
 sg13g2_fill_2 FILLER_41_517 ();
 sg13g2_fill_2 FILLER_41_523 ();
 sg13g2_decap_4 FILLER_41_534 ();
 sg13g2_decap_4 FILLER_41_548 ();
 sg13g2_fill_2 FILLER_41_552 ();
 sg13g2_decap_8 FILLER_41_558 ();
 sg13g2_decap_8 FILLER_41_565 ();
 sg13g2_decap_8 FILLER_41_572 ();
 sg13g2_decap_8 FILLER_41_579 ();
 sg13g2_fill_2 FILLER_41_586 ();
 sg13g2_decap_8 FILLER_41_592 ();
 sg13g2_decap_4 FILLER_41_599 ();
 sg13g2_fill_1 FILLER_41_603 ();
 sg13g2_fill_2 FILLER_41_608 ();
 sg13g2_fill_1 FILLER_41_610 ();
 sg13g2_fill_2 FILLER_41_615 ();
 sg13g2_fill_1 FILLER_41_623 ();
 sg13g2_decap_8 FILLER_41_640 ();
 sg13g2_decap_8 FILLER_41_647 ();
 sg13g2_decap_8 FILLER_41_654 ();
 sg13g2_decap_4 FILLER_41_661 ();
 sg13g2_fill_1 FILLER_41_665 ();
 sg13g2_decap_4 FILLER_41_670 ();
 sg13g2_decap_8 FILLER_41_677 ();
 sg13g2_fill_2 FILLER_41_687 ();
 sg13g2_decap_8 FILLER_41_692 ();
 sg13g2_decap_8 FILLER_41_699 ();
 sg13g2_decap_8 FILLER_41_706 ();
 sg13g2_fill_2 FILLER_41_713 ();
 sg13g2_fill_2 FILLER_41_718 ();
 sg13g2_fill_1 FILLER_41_720 ();
 sg13g2_fill_1 FILLER_41_726 ();
 sg13g2_decap_8 FILLER_41_734 ();
 sg13g2_decap_4 FILLER_41_741 ();
 sg13g2_decap_4 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_759 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_fill_2 FILLER_41_773 ();
 sg13g2_fill_2 FILLER_41_783 ();
 sg13g2_decap_8 FILLER_41_789 ();
 sg13g2_decap_8 FILLER_41_796 ();
 sg13g2_decap_8 FILLER_41_803 ();
 sg13g2_decap_8 FILLER_41_810 ();
 sg13g2_decap_8 FILLER_41_817 ();
 sg13g2_decap_8 FILLER_41_824 ();
 sg13g2_decap_8 FILLER_41_831 ();
 sg13g2_decap_8 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_845 ();
 sg13g2_decap_8 FILLER_41_852 ();
 sg13g2_decap_8 FILLER_41_859 ();
 sg13g2_decap_8 FILLER_41_866 ();
 sg13g2_decap_4 FILLER_41_873 ();
 sg13g2_fill_1 FILLER_41_877 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_fill_2 FILLER_42_49 ();
 sg13g2_fill_1 FILLER_42_51 ();
 sg13g2_decap_8 FILLER_42_61 ();
 sg13g2_fill_1 FILLER_42_68 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_102 ();
 sg13g2_fill_2 FILLER_42_109 ();
 sg13g2_fill_1 FILLER_42_116 ();
 sg13g2_fill_2 FILLER_42_126 ();
 sg13g2_decap_4 FILLER_42_132 ();
 sg13g2_decap_8 FILLER_42_145 ();
 sg13g2_decap_8 FILLER_42_152 ();
 sg13g2_decap_8 FILLER_42_159 ();
 sg13g2_decap_8 FILLER_42_166 ();
 sg13g2_decap_4 FILLER_42_173 ();
 sg13g2_fill_2 FILLER_42_177 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_fill_1 FILLER_42_196 ();
 sg13g2_decap_4 FILLER_42_206 ();
 sg13g2_fill_1 FILLER_42_210 ();
 sg13g2_fill_1 FILLER_42_220 ();
 sg13g2_decap_8 FILLER_42_226 ();
 sg13g2_decap_8 FILLER_42_233 ();
 sg13g2_decap_8 FILLER_42_240 ();
 sg13g2_fill_1 FILLER_42_247 ();
 sg13g2_decap_8 FILLER_42_256 ();
 sg13g2_decap_8 FILLER_42_263 ();
 sg13g2_decap_8 FILLER_42_270 ();
 sg13g2_fill_2 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_decap_8 FILLER_42_284 ();
 sg13g2_decap_4 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_299 ();
 sg13g2_decap_8 FILLER_42_309 ();
 sg13g2_decap_8 FILLER_42_316 ();
 sg13g2_decap_8 FILLER_42_323 ();
 sg13g2_decap_4 FILLER_42_330 ();
 sg13g2_fill_2 FILLER_42_334 ();
 sg13g2_fill_1 FILLER_42_340 ();
 sg13g2_fill_2 FILLER_42_350 ();
 sg13g2_fill_1 FILLER_42_352 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_fill_2 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_376 ();
 sg13g2_decap_8 FILLER_42_383 ();
 sg13g2_decap_8 FILLER_42_390 ();
 sg13g2_decap_8 FILLER_42_397 ();
 sg13g2_decap_8 FILLER_42_404 ();
 sg13g2_decap_8 FILLER_42_411 ();
 sg13g2_decap_8 FILLER_42_418 ();
 sg13g2_decap_8 FILLER_42_425 ();
 sg13g2_decap_8 FILLER_42_432 ();
 sg13g2_decap_8 FILLER_42_439 ();
 sg13g2_decap_8 FILLER_42_446 ();
 sg13g2_decap_8 FILLER_42_453 ();
 sg13g2_fill_2 FILLER_42_460 ();
 sg13g2_fill_1 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_decap_8 FILLER_42_511 ();
 sg13g2_decap_8 FILLER_42_518 ();
 sg13g2_fill_2 FILLER_42_525 ();
 sg13g2_decap_4 FILLER_42_532 ();
 sg13g2_decap_4 FILLER_42_541 ();
 sg13g2_decap_8 FILLER_42_549 ();
 sg13g2_decap_8 FILLER_42_556 ();
 sg13g2_decap_8 FILLER_42_563 ();
 sg13g2_decap_4 FILLER_42_570 ();
 sg13g2_decap_4 FILLER_42_580 ();
 sg13g2_fill_2 FILLER_42_584 ();
 sg13g2_fill_2 FILLER_42_598 ();
 sg13g2_fill_1 FILLER_42_610 ();
 sg13g2_decap_4 FILLER_42_615 ();
 sg13g2_fill_2 FILLER_42_619 ();
 sg13g2_decap_8 FILLER_42_631 ();
 sg13g2_fill_2 FILLER_42_638 ();
 sg13g2_decap_8 FILLER_42_650 ();
 sg13g2_decap_8 FILLER_42_657 ();
 sg13g2_decap_8 FILLER_42_664 ();
 sg13g2_fill_2 FILLER_42_671 ();
 sg13g2_fill_1 FILLER_42_673 ();
 sg13g2_fill_2 FILLER_42_677 ();
 sg13g2_fill_1 FILLER_42_679 ();
 sg13g2_decap_8 FILLER_42_694 ();
 sg13g2_fill_1 FILLER_42_701 ();
 sg13g2_decap_8 FILLER_42_706 ();
 sg13g2_decap_8 FILLER_42_713 ();
 sg13g2_decap_4 FILLER_42_720 ();
 sg13g2_decap_4 FILLER_42_728 ();
 sg13g2_fill_2 FILLER_42_732 ();
 sg13g2_decap_8 FILLER_42_743 ();
 sg13g2_decap_8 FILLER_42_750 ();
 sg13g2_fill_2 FILLER_42_757 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_fill_2 FILLER_42_777 ();
 sg13g2_fill_1 FILLER_42_779 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_decap_8 FILLER_42_790 ();
 sg13g2_decap_8 FILLER_42_797 ();
 sg13g2_decap_8 FILLER_42_804 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_846 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_decap_8 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_42_867 ();
 sg13g2_decap_4 FILLER_42_874 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_4 FILLER_43_49 ();
 sg13g2_fill_1 FILLER_43_53 ();
 sg13g2_decap_8 FILLER_43_58 ();
 sg13g2_decap_8 FILLER_43_65 ();
 sg13g2_decap_8 FILLER_43_72 ();
 sg13g2_decap_8 FILLER_43_79 ();
 sg13g2_decap_8 FILLER_43_86 ();
 sg13g2_decap_8 FILLER_43_93 ();
 sg13g2_decap_8 FILLER_43_100 ();
 sg13g2_decap_4 FILLER_43_107 ();
 sg13g2_decap_8 FILLER_43_115 ();
 sg13g2_decap_8 FILLER_43_122 ();
 sg13g2_decap_4 FILLER_43_129 ();
 sg13g2_fill_1 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_142 ();
 sg13g2_decap_8 FILLER_43_149 ();
 sg13g2_decap_8 FILLER_43_156 ();
 sg13g2_decap_8 FILLER_43_163 ();
 sg13g2_decap_8 FILLER_43_170 ();
 sg13g2_decap_4 FILLER_43_177 ();
 sg13g2_fill_1 FILLER_43_181 ();
 sg13g2_decap_4 FILLER_43_186 ();
 sg13g2_fill_2 FILLER_43_190 ();
 sg13g2_decap_4 FILLER_43_211 ();
 sg13g2_fill_2 FILLER_43_215 ();
 sg13g2_decap_4 FILLER_43_222 ();
 sg13g2_fill_2 FILLER_43_226 ();
 sg13g2_decap_4 FILLER_43_232 ();
 sg13g2_fill_2 FILLER_43_236 ();
 sg13g2_decap_4 FILLER_43_242 ();
 sg13g2_fill_2 FILLER_43_246 ();
 sg13g2_decap_8 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_264 ();
 sg13g2_decap_8 FILLER_43_278 ();
 sg13g2_decap_8 FILLER_43_285 ();
 sg13g2_fill_2 FILLER_43_292 ();
 sg13g2_fill_1 FILLER_43_294 ();
 sg13g2_fill_1 FILLER_43_300 ();
 sg13g2_fill_1 FILLER_43_305 ();
 sg13g2_decap_4 FILLER_43_310 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_4 FILLER_43_357 ();
 sg13g2_fill_2 FILLER_43_361 ();
 sg13g2_decap_8 FILLER_43_367 ();
 sg13g2_decap_8 FILLER_43_374 ();
 sg13g2_decap_8 FILLER_43_381 ();
 sg13g2_decap_4 FILLER_43_388 ();
 sg13g2_fill_2 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_403 ();
 sg13g2_decap_4 FILLER_43_410 ();
 sg13g2_fill_1 FILLER_43_414 ();
 sg13g2_decap_4 FILLER_43_419 ();
 sg13g2_decap_8 FILLER_43_428 ();
 sg13g2_decap_8 FILLER_43_435 ();
 sg13g2_decap_4 FILLER_43_442 ();
 sg13g2_decap_8 FILLER_43_451 ();
 sg13g2_decap_8 FILLER_43_458 ();
 sg13g2_fill_2 FILLER_43_465 ();
 sg13g2_fill_1 FILLER_43_467 ();
 sg13g2_fill_2 FILLER_43_482 ();
 sg13g2_fill_1 FILLER_43_484 ();
 sg13g2_decap_8 FILLER_43_498 ();
 sg13g2_decap_8 FILLER_43_505 ();
 sg13g2_decap_8 FILLER_43_512 ();
 sg13g2_decap_8 FILLER_43_519 ();
 sg13g2_decap_8 FILLER_43_526 ();
 sg13g2_decap_8 FILLER_43_533 ();
 sg13g2_decap_8 FILLER_43_540 ();
 sg13g2_decap_4 FILLER_43_547 ();
 sg13g2_decap_8 FILLER_43_556 ();
 sg13g2_fill_2 FILLER_43_563 ();
 sg13g2_decap_8 FILLER_43_570 ();
 sg13g2_fill_1 FILLER_43_577 ();
 sg13g2_fill_2 FILLER_43_588 ();
 sg13g2_fill_2 FILLER_43_594 ();
 sg13g2_decap_8 FILLER_43_606 ();
 sg13g2_decap_8 FILLER_43_613 ();
 sg13g2_decap_8 FILLER_43_620 ();
 sg13g2_fill_1 FILLER_43_627 ();
 sg13g2_fill_1 FILLER_43_637 ();
 sg13g2_fill_2 FILLER_43_642 ();
 sg13g2_decap_8 FILLER_43_648 ();
 sg13g2_fill_2 FILLER_43_655 ();
 sg13g2_decap_8 FILLER_43_662 ();
 sg13g2_fill_1 FILLER_43_673 ();
 sg13g2_fill_2 FILLER_43_678 ();
 sg13g2_fill_1 FILLER_43_680 ();
 sg13g2_fill_2 FILLER_43_686 ();
 sg13g2_fill_1 FILLER_43_688 ();
 sg13g2_decap_4 FILLER_43_699 ();
 sg13g2_fill_2 FILLER_43_703 ();
 sg13g2_decap_8 FILLER_43_710 ();
 sg13g2_decap_8 FILLER_43_717 ();
 sg13g2_decap_4 FILLER_43_724 ();
 sg13g2_fill_1 FILLER_43_734 ();
 sg13g2_decap_8 FILLER_43_744 ();
 sg13g2_decap_4 FILLER_43_751 ();
 sg13g2_fill_1 FILLER_43_755 ();
 sg13g2_decap_8 FILLER_43_762 ();
 sg13g2_decap_8 FILLER_43_769 ();
 sg13g2_fill_2 FILLER_43_776 ();
 sg13g2_fill_1 FILLER_43_778 ();
 sg13g2_decap_8 FILLER_43_783 ();
 sg13g2_decap_8 FILLER_43_790 ();
 sg13g2_decap_8 FILLER_43_797 ();
 sg13g2_decap_8 FILLER_43_804 ();
 sg13g2_decap_8 FILLER_43_811 ();
 sg13g2_decap_8 FILLER_43_818 ();
 sg13g2_decap_8 FILLER_43_825 ();
 sg13g2_decap_8 FILLER_43_832 ();
 sg13g2_decap_8 FILLER_43_839 ();
 sg13g2_decap_8 FILLER_43_846 ();
 sg13g2_decap_8 FILLER_43_853 ();
 sg13g2_decap_8 FILLER_43_860 ();
 sg13g2_decap_8 FILLER_43_867 ();
 sg13g2_decap_4 FILLER_43_874 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_4 FILLER_44_49 ();
 sg13g2_fill_2 FILLER_44_66 ();
 sg13g2_decap_4 FILLER_44_73 ();
 sg13g2_decap_4 FILLER_44_81 ();
 sg13g2_decap_8 FILLER_44_89 ();
 sg13g2_decap_8 FILLER_44_96 ();
 sg13g2_decap_8 FILLER_44_103 ();
 sg13g2_fill_1 FILLER_44_110 ();
 sg13g2_fill_2 FILLER_44_125 ();
 sg13g2_fill_1 FILLER_44_132 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_fill_2 FILLER_44_147 ();
 sg13g2_fill_1 FILLER_44_149 ();
 sg13g2_decap_8 FILLER_44_155 ();
 sg13g2_decap_8 FILLER_44_162 ();
 sg13g2_decap_4 FILLER_44_169 ();
 sg13g2_decap_4 FILLER_44_190 ();
 sg13g2_fill_1 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_208 ();
 sg13g2_decap_8 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_222 ();
 sg13g2_decap_8 FILLER_44_229 ();
 sg13g2_decap_8 FILLER_44_244 ();
 sg13g2_decap_4 FILLER_44_251 ();
 sg13g2_decap_4 FILLER_44_260 ();
 sg13g2_fill_1 FILLER_44_264 ();
 sg13g2_decap_4 FILLER_44_269 ();
 sg13g2_fill_1 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_279 ();
 sg13g2_fill_2 FILLER_44_286 ();
 sg13g2_fill_1 FILLER_44_288 ();
 sg13g2_fill_1 FILLER_44_293 ();
 sg13g2_fill_2 FILLER_44_299 ();
 sg13g2_fill_1 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_307 ();
 sg13g2_fill_2 FILLER_44_314 ();
 sg13g2_decap_8 FILLER_44_324 ();
 sg13g2_decap_8 FILLER_44_331 ();
 sg13g2_decap_8 FILLER_44_338 ();
 sg13g2_decap_8 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_368 ();
 sg13g2_decap_8 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_4 FILLER_44_396 ();
 sg13g2_fill_2 FILLER_44_400 ();
 sg13g2_fill_1 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_44_428 ();
 sg13g2_fill_2 FILLER_44_444 ();
 sg13g2_decap_8 FILLER_44_454 ();
 sg13g2_decap_8 FILLER_44_461 ();
 sg13g2_decap_8 FILLER_44_468 ();
 sg13g2_decap_4 FILLER_44_492 ();
 sg13g2_fill_1 FILLER_44_496 ();
 sg13g2_decap_8 FILLER_44_505 ();
 sg13g2_decap_8 FILLER_44_512 ();
 sg13g2_decap_8 FILLER_44_519 ();
 sg13g2_decap_8 FILLER_44_526 ();
 sg13g2_fill_1 FILLER_44_539 ();
 sg13g2_decap_8 FILLER_44_546 ();
 sg13g2_decap_8 FILLER_44_553 ();
 sg13g2_decap_4 FILLER_44_560 ();
 sg13g2_fill_1 FILLER_44_564 ();
 sg13g2_decap_8 FILLER_44_574 ();
 sg13g2_decap_8 FILLER_44_581 ();
 sg13g2_fill_2 FILLER_44_594 ();
 sg13g2_decap_4 FILLER_44_601 ();
 sg13g2_decap_8 FILLER_44_611 ();
 sg13g2_decap_8 FILLER_44_618 ();
 sg13g2_decap_8 FILLER_44_629 ();
 sg13g2_decap_8 FILLER_44_636 ();
 sg13g2_decap_8 FILLER_44_643 ();
 sg13g2_decap_4 FILLER_44_650 ();
 sg13g2_fill_2 FILLER_44_662 ();
 sg13g2_decap_4 FILLER_44_669 ();
 sg13g2_fill_2 FILLER_44_673 ();
 sg13g2_decap_8 FILLER_44_690 ();
 sg13g2_decap_8 FILLER_44_697 ();
 sg13g2_decap_4 FILLER_44_704 ();
 sg13g2_fill_1 FILLER_44_708 ();
 sg13g2_decap_8 FILLER_44_713 ();
 sg13g2_decap_4 FILLER_44_720 ();
 sg13g2_fill_2 FILLER_44_724 ();
 sg13g2_fill_2 FILLER_44_731 ();
 sg13g2_fill_1 FILLER_44_738 ();
 sg13g2_decap_8 FILLER_44_747 ();
 sg13g2_decap_8 FILLER_44_754 ();
 sg13g2_decap_8 FILLER_44_761 ();
 sg13g2_decap_8 FILLER_44_768 ();
 sg13g2_decap_8 FILLER_44_775 ();
 sg13g2_decap_8 FILLER_44_782 ();
 sg13g2_decap_8 FILLER_44_789 ();
 sg13g2_decap_8 FILLER_44_796 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_decap_8 FILLER_44_810 ();
 sg13g2_decap_8 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_decap_8 FILLER_44_831 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_decap_8 FILLER_44_859 ();
 sg13g2_decap_8 FILLER_44_866 ();
 sg13g2_decap_4 FILLER_44_873 ();
 sg13g2_fill_1 FILLER_44_877 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_4 FILLER_45_49 ();
 sg13g2_fill_2 FILLER_45_53 ();
 sg13g2_fill_1 FILLER_45_59 ();
 sg13g2_fill_1 FILLER_45_64 ();
 sg13g2_fill_1 FILLER_45_69 ();
 sg13g2_fill_2 FILLER_45_74 ();
 sg13g2_fill_1 FILLER_45_76 ();
 sg13g2_fill_1 FILLER_45_82 ();
 sg13g2_fill_2 FILLER_45_87 ();
 sg13g2_decap_8 FILLER_45_93 ();
 sg13g2_decap_8 FILLER_45_100 ();
 sg13g2_decap_8 FILLER_45_107 ();
 sg13g2_decap_4 FILLER_45_114 ();
 sg13g2_fill_1 FILLER_45_118 ();
 sg13g2_decap_8 FILLER_45_127 ();
 sg13g2_decap_8 FILLER_45_134 ();
 sg13g2_decap_8 FILLER_45_141 ();
 sg13g2_fill_1 FILLER_45_148 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_4 FILLER_45_161 ();
 sg13g2_decap_4 FILLER_45_168 ();
 sg13g2_fill_1 FILLER_45_172 ();
 sg13g2_fill_2 FILLER_45_178 ();
 sg13g2_decap_8 FILLER_45_184 ();
 sg13g2_decap_8 FILLER_45_199 ();
 sg13g2_fill_2 FILLER_45_206 ();
 sg13g2_fill_1 FILLER_45_208 ();
 sg13g2_decap_8 FILLER_45_214 ();
 sg13g2_decap_8 FILLER_45_221 ();
 sg13g2_decap_8 FILLER_45_228 ();
 sg13g2_decap_8 FILLER_45_240 ();
 sg13g2_decap_8 FILLER_45_247 ();
 sg13g2_decap_8 FILLER_45_254 ();
 sg13g2_fill_2 FILLER_45_261 ();
 sg13g2_fill_1 FILLER_45_263 ();
 sg13g2_decap_8 FILLER_45_268 ();
 sg13g2_decap_8 FILLER_45_275 ();
 sg13g2_decap_8 FILLER_45_282 ();
 sg13g2_fill_2 FILLER_45_289 ();
 sg13g2_fill_1 FILLER_45_291 ();
 sg13g2_decap_4 FILLER_45_297 ();
 sg13g2_fill_2 FILLER_45_301 ();
 sg13g2_fill_2 FILLER_45_312 ();
 sg13g2_decap_8 FILLER_45_327 ();
 sg13g2_decap_8 FILLER_45_334 ();
 sg13g2_decap_8 FILLER_45_341 ();
 sg13g2_decap_8 FILLER_45_348 ();
 sg13g2_decap_4 FILLER_45_355 ();
 sg13g2_fill_1 FILLER_45_359 ();
 sg13g2_fill_1 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_370 ();
 sg13g2_decap_4 FILLER_45_377 ();
 sg13g2_fill_1 FILLER_45_381 ();
 sg13g2_decap_8 FILLER_45_390 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_45_417 ();
 sg13g2_fill_1 FILLER_45_424 ();
 sg13g2_decap_8 FILLER_45_429 ();
 sg13g2_decap_4 FILLER_45_436 ();
 sg13g2_fill_1 FILLER_45_440 ();
 sg13g2_decap_8 FILLER_45_445 ();
 sg13g2_decap_8 FILLER_45_456 ();
 sg13g2_fill_1 FILLER_45_463 ();
 sg13g2_decap_4 FILLER_45_473 ();
 sg13g2_fill_1 FILLER_45_477 ();
 sg13g2_decap_8 FILLER_45_482 ();
 sg13g2_decap_8 FILLER_45_489 ();
 sg13g2_decap_4 FILLER_45_496 ();
 sg13g2_fill_2 FILLER_45_500 ();
 sg13g2_decap_4 FILLER_45_507 ();
 sg13g2_fill_1 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_517 ();
 sg13g2_decap_4 FILLER_45_524 ();
 sg13g2_fill_1 FILLER_45_528 ();
 sg13g2_decap_4 FILLER_45_534 ();
 sg13g2_fill_2 FILLER_45_538 ();
 sg13g2_decap_8 FILLER_45_548 ();
 sg13g2_fill_2 FILLER_45_555 ();
 sg13g2_fill_1 FILLER_45_557 ();
 sg13g2_decap_8 FILLER_45_570 ();
 sg13g2_decap_8 FILLER_45_577 ();
 sg13g2_decap_8 FILLER_45_584 ();
 sg13g2_decap_8 FILLER_45_591 ();
 sg13g2_decap_8 FILLER_45_598 ();
 sg13g2_decap_8 FILLER_45_605 ();
 sg13g2_decap_8 FILLER_45_612 ();
 sg13g2_fill_2 FILLER_45_619 ();
 sg13g2_decap_8 FILLER_45_625 ();
 sg13g2_decap_8 FILLER_45_632 ();
 sg13g2_fill_2 FILLER_45_639 ();
 sg13g2_fill_2 FILLER_45_650 ();
 sg13g2_decap_8 FILLER_45_656 ();
 sg13g2_decap_8 FILLER_45_663 ();
 sg13g2_decap_4 FILLER_45_670 ();
 sg13g2_fill_1 FILLER_45_674 ();
 sg13g2_decap_8 FILLER_45_679 ();
 sg13g2_decap_4 FILLER_45_686 ();
 sg13g2_fill_1 FILLER_45_690 ();
 sg13g2_decap_4 FILLER_45_695 ();
 sg13g2_decap_8 FILLER_45_703 ();
 sg13g2_decap_8 FILLER_45_710 ();
 sg13g2_decap_4 FILLER_45_717 ();
 sg13g2_fill_1 FILLER_45_721 ();
 sg13g2_fill_1 FILLER_45_728 ();
 sg13g2_decap_8 FILLER_45_743 ();
 sg13g2_decap_4 FILLER_45_750 ();
 sg13g2_decap_4 FILLER_45_772 ();
 sg13g2_decap_8 FILLER_45_780 ();
 sg13g2_decap_8 FILLER_45_787 ();
 sg13g2_decap_8 FILLER_45_794 ();
 sg13g2_decap_8 FILLER_45_801 ();
 sg13g2_decap_8 FILLER_45_808 ();
 sg13g2_decap_8 FILLER_45_815 ();
 sg13g2_decap_8 FILLER_45_822 ();
 sg13g2_decap_8 FILLER_45_829 ();
 sg13g2_decap_8 FILLER_45_836 ();
 sg13g2_decap_8 FILLER_45_843 ();
 sg13g2_decap_8 FILLER_45_850 ();
 sg13g2_decap_8 FILLER_45_857 ();
 sg13g2_decap_8 FILLER_45_864 ();
 sg13g2_decap_8 FILLER_45_871 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_fill_1 FILLER_46_63 ();
 sg13g2_fill_2 FILLER_46_72 ();
 sg13g2_fill_1 FILLER_46_74 ();
 sg13g2_fill_2 FILLER_46_83 ();
 sg13g2_fill_1 FILLER_46_85 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_fill_2 FILLER_46_126 ();
 sg13g2_fill_1 FILLER_46_128 ();
 sg13g2_decap_4 FILLER_46_133 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_150 ();
 sg13g2_decap_8 FILLER_46_157 ();
 sg13g2_decap_8 FILLER_46_164 ();
 sg13g2_decap_8 FILLER_46_171 ();
 sg13g2_decap_8 FILLER_46_178 ();
 sg13g2_decap_8 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_192 ();
 sg13g2_decap_8 FILLER_46_199 ();
 sg13g2_decap_8 FILLER_46_206 ();
 sg13g2_fill_2 FILLER_46_213 ();
 sg13g2_decap_8 FILLER_46_228 ();
 sg13g2_decap_8 FILLER_46_235 ();
 sg13g2_fill_2 FILLER_46_242 ();
 sg13g2_fill_1 FILLER_46_244 ();
 sg13g2_fill_1 FILLER_46_254 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_fill_1 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_299 ();
 sg13g2_decap_8 FILLER_46_306 ();
 sg13g2_decap_4 FILLER_46_313 ();
 sg13g2_fill_2 FILLER_46_317 ();
 sg13g2_decap_8 FILLER_46_324 ();
 sg13g2_decap_8 FILLER_46_331 ();
 sg13g2_decap_8 FILLER_46_338 ();
 sg13g2_decap_8 FILLER_46_345 ();
 sg13g2_decap_8 FILLER_46_352 ();
 sg13g2_decap_8 FILLER_46_359 ();
 sg13g2_fill_2 FILLER_46_366 ();
 sg13g2_fill_1 FILLER_46_377 ();
 sg13g2_decap_8 FILLER_46_383 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_fill_2 FILLER_46_409 ();
 sg13g2_fill_1 FILLER_46_411 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_4 FILLER_46_441 ();
 sg13g2_fill_2 FILLER_46_445 ();
 sg13g2_decap_8 FILLER_46_450 ();
 sg13g2_decap_8 FILLER_46_457 ();
 sg13g2_decap_4 FILLER_46_464 ();
 sg13g2_fill_1 FILLER_46_468 ();
 sg13g2_decap_8 FILLER_46_473 ();
 sg13g2_decap_4 FILLER_46_480 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_fill_2 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_545 ();
 sg13g2_decap_8 FILLER_46_552 ();
 sg13g2_fill_1 FILLER_46_559 ();
 sg13g2_fill_1 FILLER_46_565 ();
 sg13g2_decap_4 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_584 ();
 sg13g2_decap_8 FILLER_46_591 ();
 sg13g2_decap_8 FILLER_46_598 ();
 sg13g2_fill_2 FILLER_46_605 ();
 sg13g2_fill_1 FILLER_46_607 ();
 sg13g2_decap_8 FILLER_46_622 ();
 sg13g2_decap_8 FILLER_46_629 ();
 sg13g2_decap_8 FILLER_46_636 ();
 sg13g2_fill_2 FILLER_46_643 ();
 sg13g2_fill_1 FILLER_46_645 ();
 sg13g2_decap_8 FILLER_46_650 ();
 sg13g2_decap_8 FILLER_46_657 ();
 sg13g2_decap_8 FILLER_46_664 ();
 sg13g2_decap_4 FILLER_46_671 ();
 sg13g2_decap_8 FILLER_46_689 ();
 sg13g2_fill_1 FILLER_46_696 ();
 sg13g2_decap_8 FILLER_46_702 ();
 sg13g2_decap_4 FILLER_46_709 ();
 sg13g2_fill_1 FILLER_46_713 ();
 sg13g2_fill_2 FILLER_46_719 ();
 sg13g2_fill_1 FILLER_46_721 ();
 sg13g2_decap_4 FILLER_46_726 ();
 sg13g2_fill_2 FILLER_46_740 ();
 sg13g2_decap_4 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_757 ();
 sg13g2_decap_8 FILLER_46_764 ();
 sg13g2_fill_2 FILLER_46_771 ();
 sg13g2_fill_1 FILLER_46_773 ();
 sg13g2_decap_8 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_793 ();
 sg13g2_decap_8 FILLER_46_800 ();
 sg13g2_decap_8 FILLER_46_807 ();
 sg13g2_decap_8 FILLER_46_814 ();
 sg13g2_decap_8 FILLER_46_821 ();
 sg13g2_decap_8 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_835 ();
 sg13g2_decap_8 FILLER_46_842 ();
 sg13g2_decap_8 FILLER_46_849 ();
 sg13g2_decap_8 FILLER_46_856 ();
 sg13g2_decap_8 FILLER_46_863 ();
 sg13g2_decap_8 FILLER_46_870 ();
 sg13g2_fill_1 FILLER_46_877 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_4 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_60 ();
 sg13g2_fill_1 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_79 ();
 sg13g2_fill_2 FILLER_47_86 ();
 sg13g2_fill_1 FILLER_47_88 ();
 sg13g2_decap_8 FILLER_47_102 ();
 sg13g2_fill_2 FILLER_47_109 ();
 sg13g2_decap_8 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_122 ();
 sg13g2_decap_8 FILLER_47_127 ();
 sg13g2_decap_4 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_148 ();
 sg13g2_decap_8 FILLER_47_159 ();
 sg13g2_decap_8 FILLER_47_166 ();
 sg13g2_decap_8 FILLER_47_173 ();
 sg13g2_fill_1 FILLER_47_180 ();
 sg13g2_decap_4 FILLER_47_199 ();
 sg13g2_fill_1 FILLER_47_203 ();
 sg13g2_decap_4 FILLER_47_208 ();
 sg13g2_decap_8 FILLER_47_227 ();
 sg13g2_fill_2 FILLER_47_234 ();
 sg13g2_decap_4 FILLER_47_245 ();
 sg13g2_fill_2 FILLER_47_258 ();
 sg13g2_fill_1 FILLER_47_260 ();
 sg13g2_decap_8 FILLER_47_264 ();
 sg13g2_decap_8 FILLER_47_271 ();
 sg13g2_fill_2 FILLER_47_278 ();
 sg13g2_decap_4 FILLER_47_285 ();
 sg13g2_fill_2 FILLER_47_289 ();
 sg13g2_decap_8 FILLER_47_300 ();
 sg13g2_decap_4 FILLER_47_307 ();
 sg13g2_fill_1 FILLER_47_311 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_4 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_375 ();
 sg13g2_decap_8 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_47_389 ();
 sg13g2_decap_4 FILLER_47_396 ();
 sg13g2_fill_2 FILLER_47_400 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_fill_2 FILLER_47_425 ();
 sg13g2_fill_1 FILLER_47_443 ();
 sg13g2_fill_2 FILLER_47_449 ();
 sg13g2_fill_2 FILLER_47_455 ();
 sg13g2_decap_4 FILLER_47_460 ();
 sg13g2_fill_1 FILLER_47_464 ();
 sg13g2_decap_8 FILLER_47_470 ();
 sg13g2_fill_1 FILLER_47_477 ();
 sg13g2_decap_8 FILLER_47_481 ();
 sg13g2_decap_8 FILLER_47_488 ();
 sg13g2_decap_4 FILLER_47_495 ();
 sg13g2_decap_8 FILLER_47_503 ();
 sg13g2_fill_1 FILLER_47_510 ();
 sg13g2_decap_8 FILLER_47_517 ();
 sg13g2_fill_2 FILLER_47_524 ();
 sg13g2_fill_1 FILLER_47_526 ();
 sg13g2_fill_2 FILLER_47_536 ();
 sg13g2_fill_1 FILLER_47_538 ();
 sg13g2_fill_2 FILLER_47_544 ();
 sg13g2_decap_8 FILLER_47_550 ();
 sg13g2_fill_2 FILLER_47_557 ();
 sg13g2_fill_2 FILLER_47_576 ();
 sg13g2_decap_4 FILLER_47_586 ();
 sg13g2_fill_2 FILLER_47_590 ();
 sg13g2_decap_8 FILLER_47_600 ();
 sg13g2_decap_8 FILLER_47_607 ();
 sg13g2_decap_8 FILLER_47_614 ();
 sg13g2_fill_1 FILLER_47_621 ();
 sg13g2_decap_8 FILLER_47_627 ();
 sg13g2_decap_4 FILLER_47_634 ();
 sg13g2_decap_4 FILLER_47_646 ();
 sg13g2_decap_8 FILLER_47_655 ();
 sg13g2_decap_4 FILLER_47_662 ();
 sg13g2_fill_2 FILLER_47_666 ();
 sg13g2_fill_1 FILLER_47_682 ();
 sg13g2_fill_2 FILLER_47_691 ();
 sg13g2_fill_1 FILLER_47_697 ();
 sg13g2_fill_1 FILLER_47_707 ();
 sg13g2_fill_1 FILLER_47_713 ();
 sg13g2_decap_4 FILLER_47_718 ();
 sg13g2_fill_1 FILLER_47_722 ();
 sg13g2_decap_4 FILLER_47_735 ();
 sg13g2_decap_4 FILLER_47_754 ();
 sg13g2_fill_2 FILLER_47_758 ();
 sg13g2_decap_8 FILLER_47_764 ();
 sg13g2_decap_8 FILLER_47_771 ();
 sg13g2_decap_8 FILLER_47_778 ();
 sg13g2_decap_8 FILLER_47_785 ();
 sg13g2_decap_8 FILLER_47_792 ();
 sg13g2_decap_8 FILLER_47_799 ();
 sg13g2_decap_8 FILLER_47_806 ();
 sg13g2_decap_8 FILLER_47_813 ();
 sg13g2_decap_8 FILLER_47_820 ();
 sg13g2_decap_8 FILLER_47_827 ();
 sg13g2_decap_8 FILLER_47_834 ();
 sg13g2_decap_8 FILLER_47_841 ();
 sg13g2_decap_8 FILLER_47_848 ();
 sg13g2_decap_8 FILLER_47_855 ();
 sg13g2_decap_8 FILLER_47_862 ();
 sg13g2_decap_8 FILLER_47_869 ();
 sg13g2_fill_2 FILLER_47_876 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_fill_2 FILLER_48_70 ();
 sg13g2_decap_4 FILLER_48_80 ();
 sg13g2_decap_8 FILLER_48_88 ();
 sg13g2_decap_8 FILLER_48_95 ();
 sg13g2_decap_8 FILLER_48_102 ();
 sg13g2_decap_8 FILLER_48_109 ();
 sg13g2_decap_8 FILLER_48_116 ();
 sg13g2_decap_8 FILLER_48_123 ();
 sg13g2_fill_2 FILLER_48_130 ();
 sg13g2_fill_1 FILLER_48_132 ();
 sg13g2_decap_4 FILLER_48_140 ();
 sg13g2_fill_1 FILLER_48_154 ();
 sg13g2_fill_1 FILLER_48_159 ();
 sg13g2_decap_8 FILLER_48_165 ();
 sg13g2_fill_2 FILLER_48_172 ();
 sg13g2_fill_1 FILLER_48_174 ();
 sg13g2_fill_2 FILLER_48_179 ();
 sg13g2_fill_1 FILLER_48_181 ();
 sg13g2_decap_8 FILLER_48_187 ();
 sg13g2_decap_8 FILLER_48_194 ();
 sg13g2_decap_8 FILLER_48_201 ();
 sg13g2_fill_1 FILLER_48_208 ();
 sg13g2_decap_8 FILLER_48_218 ();
 sg13g2_fill_2 FILLER_48_225 ();
 sg13g2_fill_1 FILLER_48_227 ();
 sg13g2_decap_8 FILLER_48_233 ();
 sg13g2_decap_4 FILLER_48_245 ();
 sg13g2_fill_2 FILLER_48_254 ();
 sg13g2_fill_1 FILLER_48_256 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_fill_1 FILLER_48_264 ();
 sg13g2_decap_8 FILLER_48_279 ();
 sg13g2_decap_8 FILLER_48_286 ();
 sg13g2_fill_2 FILLER_48_293 ();
 sg13g2_fill_1 FILLER_48_300 ();
 sg13g2_decap_8 FILLER_48_306 ();
 sg13g2_decap_4 FILLER_48_313 ();
 sg13g2_fill_1 FILLER_48_317 ();
 sg13g2_decap_8 FILLER_48_323 ();
 sg13g2_decap_4 FILLER_48_330 ();
 sg13g2_decap_8 FILLER_48_349 ();
 sg13g2_decap_4 FILLER_48_356 ();
 sg13g2_fill_1 FILLER_48_360 ();
 sg13g2_decap_4 FILLER_48_365 ();
 sg13g2_fill_1 FILLER_48_369 ();
 sg13g2_decap_8 FILLER_48_374 ();
 sg13g2_decap_8 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_48_388 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_fill_1 FILLER_48_409 ();
 sg13g2_decap_8 FILLER_48_417 ();
 sg13g2_decap_8 FILLER_48_424 ();
 sg13g2_fill_2 FILLER_48_431 ();
 sg13g2_fill_1 FILLER_48_453 ();
 sg13g2_fill_2 FILLER_48_464 ();
 sg13g2_fill_1 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_482 ();
 sg13g2_fill_2 FILLER_48_489 ();
 sg13g2_fill_1 FILLER_48_491 ();
 sg13g2_decap_8 FILLER_48_505 ();
 sg13g2_decap_8 FILLER_48_512 ();
 sg13g2_decap_8 FILLER_48_519 ();
 sg13g2_decap_8 FILLER_48_526 ();
 sg13g2_fill_1 FILLER_48_537 ();
 sg13g2_decap_4 FILLER_48_541 ();
 sg13g2_decap_8 FILLER_48_549 ();
 sg13g2_decap_4 FILLER_48_556 ();
 sg13g2_decap_8 FILLER_48_568 ();
 sg13g2_decap_8 FILLER_48_575 ();
 sg13g2_decap_8 FILLER_48_582 ();
 sg13g2_decap_4 FILLER_48_589 ();
 sg13g2_fill_2 FILLER_48_593 ();
 sg13g2_decap_8 FILLER_48_599 ();
 sg13g2_decap_8 FILLER_48_606 ();
 sg13g2_fill_2 FILLER_48_618 ();
 sg13g2_fill_1 FILLER_48_620 ();
 sg13g2_decap_8 FILLER_48_634 ();
 sg13g2_decap_8 FILLER_48_641 ();
 sg13g2_decap_8 FILLER_48_648 ();
 sg13g2_decap_8 FILLER_48_655 ();
 sg13g2_decap_8 FILLER_48_662 ();
 sg13g2_decap_8 FILLER_48_669 ();
 sg13g2_decap_8 FILLER_48_676 ();
 sg13g2_decap_8 FILLER_48_683 ();
 sg13g2_fill_2 FILLER_48_690 ();
 sg13g2_fill_1 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_730 ();
 sg13g2_decap_8 FILLER_48_737 ();
 sg13g2_decap_8 FILLER_48_744 ();
 sg13g2_fill_1 FILLER_48_751 ();
 sg13g2_decap_4 FILLER_48_758 ();
 sg13g2_fill_1 FILLER_48_767 ();
 sg13g2_decap_8 FILLER_48_772 ();
 sg13g2_decap_8 FILLER_48_779 ();
 sg13g2_fill_2 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_801 ();
 sg13g2_decap_8 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_850 ();
 sg13g2_decap_8 FILLER_48_857 ();
 sg13g2_decap_8 FILLER_48_864 ();
 sg13g2_decap_8 FILLER_48_871 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_4 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_83 ();
 sg13g2_decap_4 FILLER_49_99 ();
 sg13g2_fill_1 FILLER_49_103 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_fill_2 FILLER_49_119 ();
 sg13g2_fill_1 FILLER_49_121 ();
 sg13g2_fill_1 FILLER_49_140 ();
 sg13g2_decap_4 FILLER_49_150 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_fill_1 FILLER_49_169 ();
 sg13g2_decap_8 FILLER_49_173 ();
 sg13g2_decap_4 FILLER_49_180 ();
 sg13g2_fill_1 FILLER_49_184 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_fill_2 FILLER_49_196 ();
 sg13g2_decap_4 FILLER_49_202 ();
 sg13g2_fill_1 FILLER_49_206 ();
 sg13g2_decap_8 FILLER_49_216 ();
 sg13g2_decap_8 FILLER_49_223 ();
 sg13g2_decap_8 FILLER_49_230 ();
 sg13g2_decap_8 FILLER_49_237 ();
 sg13g2_decap_8 FILLER_49_244 ();
 sg13g2_decap_8 FILLER_49_251 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_fill_2 FILLER_49_270 ();
 sg13g2_fill_1 FILLER_49_272 ();
 sg13g2_decap_8 FILLER_49_282 ();
 sg13g2_fill_2 FILLER_49_289 ();
 sg13g2_fill_1 FILLER_49_291 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_4 FILLER_49_315 ();
 sg13g2_fill_1 FILLER_49_319 ();
 sg13g2_decap_8 FILLER_49_324 ();
 sg13g2_fill_2 FILLER_49_331 ();
 sg13g2_decap_8 FILLER_49_338 ();
 sg13g2_fill_1 FILLER_49_345 ();
 sg13g2_fill_2 FILLER_49_351 ();
 sg13g2_fill_1 FILLER_49_353 ();
 sg13g2_fill_2 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_fill_1 FILLER_49_373 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_decap_8 FILLER_49_386 ();
 sg13g2_fill_2 FILLER_49_393 ();
 sg13g2_decap_4 FILLER_49_399 ();
 sg13g2_fill_1 FILLER_49_403 ();
 sg13g2_decap_4 FILLER_49_408 ();
 sg13g2_fill_1 FILLER_49_412 ();
 sg13g2_decap_8 FILLER_49_423 ();
 sg13g2_decap_8 FILLER_49_430 ();
 sg13g2_fill_1 FILLER_49_437 ();
 sg13g2_decap_8 FILLER_49_446 ();
 sg13g2_decap_4 FILLER_49_453 ();
 sg13g2_fill_1 FILLER_49_457 ();
 sg13g2_decap_4 FILLER_49_462 ();
 sg13g2_fill_2 FILLER_49_466 ();
 sg13g2_decap_8 FILLER_49_486 ();
 sg13g2_decap_8 FILLER_49_493 ();
 sg13g2_decap_8 FILLER_49_500 ();
 sg13g2_decap_8 FILLER_49_507 ();
 sg13g2_decap_8 FILLER_49_514 ();
 sg13g2_decap_8 FILLER_49_521 ();
 sg13g2_decap_8 FILLER_49_528 ();
 sg13g2_decap_4 FILLER_49_535 ();
 sg13g2_fill_2 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_545 ();
 sg13g2_decap_8 FILLER_49_552 ();
 sg13g2_decap_8 FILLER_49_559 ();
 sg13g2_decap_8 FILLER_49_566 ();
 sg13g2_decap_8 FILLER_49_573 ();
 sg13g2_fill_2 FILLER_49_588 ();
 sg13g2_fill_1 FILLER_49_590 ();
 sg13g2_decap_8 FILLER_49_601 ();
 sg13g2_decap_8 FILLER_49_608 ();
 sg13g2_fill_1 FILLER_49_615 ();
 sg13g2_fill_1 FILLER_49_626 ();
 sg13g2_decap_4 FILLER_49_635 ();
 sg13g2_decap_8 FILLER_49_648 ();
 sg13g2_decap_4 FILLER_49_655 ();
 sg13g2_decap_8 FILLER_49_666 ();
 sg13g2_decap_8 FILLER_49_673 ();
 sg13g2_decap_8 FILLER_49_680 ();
 sg13g2_decap_4 FILLER_49_687 ();
 sg13g2_fill_1 FILLER_49_691 ();
 sg13g2_decap_8 FILLER_49_698 ();
 sg13g2_decap_8 FILLER_49_705 ();
 sg13g2_fill_1 FILLER_49_712 ();
 sg13g2_decap_8 FILLER_49_718 ();
 sg13g2_decap_4 FILLER_49_725 ();
 sg13g2_decap_4 FILLER_49_738 ();
 sg13g2_fill_1 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_753 ();
 sg13g2_fill_2 FILLER_49_760 ();
 sg13g2_fill_1 FILLER_49_762 ();
 sg13g2_decap_8 FILLER_49_768 ();
 sg13g2_decap_8 FILLER_49_775 ();
 sg13g2_decap_4 FILLER_49_782 ();
 sg13g2_fill_1 FILLER_49_786 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_fill_2 FILLER_49_875 ();
 sg13g2_fill_1 FILLER_49_877 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_4 FILLER_50_49 ();
 sg13g2_fill_1 FILLER_50_53 ();
 sg13g2_decap_4 FILLER_50_74 ();
 sg13g2_fill_1 FILLER_50_78 ();
 sg13g2_decap_8 FILLER_50_83 ();
 sg13g2_decap_8 FILLER_50_94 ();
 sg13g2_decap_8 FILLER_50_101 ();
 sg13g2_decap_8 FILLER_50_108 ();
 sg13g2_decap_8 FILLER_50_115 ();
 sg13g2_decap_8 FILLER_50_122 ();
 sg13g2_decap_8 FILLER_50_129 ();
 sg13g2_decap_8 FILLER_50_141 ();
 sg13g2_fill_1 FILLER_50_148 ();
 sg13g2_decap_4 FILLER_50_153 ();
 sg13g2_fill_1 FILLER_50_157 ();
 sg13g2_fill_2 FILLER_50_162 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_decap_8 FILLER_50_189 ();
 sg13g2_decap_8 FILLER_50_196 ();
 sg13g2_fill_2 FILLER_50_203 ();
 sg13g2_fill_2 FILLER_50_215 ();
 sg13g2_decap_8 FILLER_50_232 ();
 sg13g2_decap_8 FILLER_50_239 ();
 sg13g2_decap_8 FILLER_50_246 ();
 sg13g2_decap_4 FILLER_50_253 ();
 sg13g2_decap_4 FILLER_50_263 ();
 sg13g2_fill_1 FILLER_50_271 ();
 sg13g2_fill_2 FILLER_50_277 ();
 sg13g2_decap_8 FILLER_50_291 ();
 sg13g2_fill_2 FILLER_50_298 ();
 sg13g2_fill_1 FILLER_50_300 ();
 sg13g2_decap_4 FILLER_50_305 ();
 sg13g2_decap_8 FILLER_50_313 ();
 sg13g2_decap_8 FILLER_50_320 ();
 sg13g2_decap_8 FILLER_50_327 ();
 sg13g2_decap_8 FILLER_50_334 ();
 sg13g2_decap_8 FILLER_50_341 ();
 sg13g2_decap_8 FILLER_50_348 ();
 sg13g2_decap_4 FILLER_50_355 ();
 sg13g2_fill_2 FILLER_50_359 ();
 sg13g2_decap_8 FILLER_50_366 ();
 sg13g2_decap_4 FILLER_50_373 ();
 sg13g2_fill_2 FILLER_50_377 ();
 sg13g2_decap_8 FILLER_50_384 ();
 sg13g2_decap_4 FILLER_50_391 ();
 sg13g2_decap_8 FILLER_50_400 ();
 sg13g2_decap_4 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_50_424 ();
 sg13g2_decap_8 FILLER_50_431 ();
 sg13g2_decap_8 FILLER_50_438 ();
 sg13g2_decap_8 FILLER_50_445 ();
 sg13g2_fill_2 FILLER_50_452 ();
 sg13g2_fill_1 FILLER_50_454 ();
 sg13g2_decap_8 FILLER_50_464 ();
 sg13g2_decap_8 FILLER_50_471 ();
 sg13g2_decap_8 FILLER_50_478 ();
 sg13g2_decap_8 FILLER_50_485 ();
 sg13g2_decap_8 FILLER_50_492 ();
 sg13g2_decap_8 FILLER_50_499 ();
 sg13g2_fill_2 FILLER_50_506 ();
 sg13g2_fill_1 FILLER_50_508 ();
 sg13g2_decap_8 FILLER_50_513 ();
 sg13g2_decap_8 FILLER_50_520 ();
 sg13g2_decap_8 FILLER_50_527 ();
 sg13g2_decap_8 FILLER_50_534 ();
 sg13g2_fill_1 FILLER_50_541 ();
 sg13g2_fill_1 FILLER_50_550 ();
 sg13g2_decap_8 FILLER_50_565 ();
 sg13g2_decap_8 FILLER_50_572 ();
 sg13g2_fill_2 FILLER_50_579 ();
 sg13g2_fill_1 FILLER_50_581 ();
 sg13g2_decap_8 FILLER_50_586 ();
 sg13g2_decap_8 FILLER_50_593 ();
 sg13g2_decap_8 FILLER_50_600 ();
 sg13g2_decap_8 FILLER_50_607 ();
 sg13g2_decap_8 FILLER_50_614 ();
 sg13g2_fill_2 FILLER_50_621 ();
 sg13g2_fill_1 FILLER_50_623 ();
 sg13g2_fill_1 FILLER_50_629 ();
 sg13g2_fill_2 FILLER_50_634 ();
 sg13g2_fill_1 FILLER_50_636 ();
 sg13g2_decap_4 FILLER_50_641 ();
 sg13g2_fill_2 FILLER_50_645 ();
 sg13g2_fill_2 FILLER_50_652 ();
 sg13g2_fill_1 FILLER_50_654 ();
 sg13g2_fill_2 FILLER_50_667 ();
 sg13g2_decap_8 FILLER_50_674 ();
 sg13g2_fill_1 FILLER_50_681 ();
 sg13g2_fill_2 FILLER_50_689 ();
 sg13g2_decap_4 FILLER_50_700 ();
 sg13g2_fill_1 FILLER_50_704 ();
 sg13g2_decap_8 FILLER_50_716 ();
 sg13g2_decap_4 FILLER_50_733 ();
 sg13g2_fill_1 FILLER_50_737 ();
 sg13g2_decap_4 FILLER_50_747 ();
 sg13g2_decap_8 FILLER_50_756 ();
 sg13g2_decap_8 FILLER_50_763 ();
 sg13g2_decap_8 FILLER_50_770 ();
 sg13g2_decap_8 FILLER_50_777 ();
 sg13g2_decap_8 FILLER_50_784 ();
 sg13g2_decap_8 FILLER_50_791 ();
 sg13g2_decap_8 FILLER_50_798 ();
 sg13g2_decap_8 FILLER_50_805 ();
 sg13g2_decap_8 FILLER_50_812 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_decap_8 FILLER_50_826 ();
 sg13g2_decap_8 FILLER_50_833 ();
 sg13g2_decap_8 FILLER_50_840 ();
 sg13g2_decap_8 FILLER_50_847 ();
 sg13g2_decap_8 FILLER_50_854 ();
 sg13g2_decap_8 FILLER_50_861 ();
 sg13g2_decap_8 FILLER_50_868 ();
 sg13g2_fill_2 FILLER_50_875 ();
 sg13g2_fill_1 FILLER_50_877 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_60 ();
 sg13g2_decap_4 FILLER_51_67 ();
 sg13g2_fill_2 FILLER_51_75 ();
 sg13g2_decap_4 FILLER_51_81 ();
 sg13g2_decap_8 FILLER_51_89 ();
 sg13g2_decap_8 FILLER_51_96 ();
 sg13g2_decap_8 FILLER_51_103 ();
 sg13g2_decap_8 FILLER_51_110 ();
 sg13g2_decap_8 FILLER_51_117 ();
 sg13g2_decap_8 FILLER_51_124 ();
 sg13g2_decap_8 FILLER_51_131 ();
 sg13g2_decap_8 FILLER_51_138 ();
 sg13g2_decap_4 FILLER_51_145 ();
 sg13g2_decap_8 FILLER_51_173 ();
 sg13g2_decap_8 FILLER_51_180 ();
 sg13g2_fill_2 FILLER_51_187 ();
 sg13g2_decap_8 FILLER_51_193 ();
 sg13g2_decap_8 FILLER_51_200 ();
 sg13g2_decap_4 FILLER_51_207 ();
 sg13g2_fill_2 FILLER_51_211 ();
 sg13g2_decap_8 FILLER_51_219 ();
 sg13g2_decap_4 FILLER_51_226 ();
 sg13g2_decap_8 FILLER_51_236 ();
 sg13g2_decap_8 FILLER_51_243 ();
 sg13g2_decap_8 FILLER_51_259 ();
 sg13g2_decap_4 FILLER_51_266 ();
 sg13g2_fill_2 FILLER_51_270 ();
 sg13g2_fill_2 FILLER_51_277 ();
 sg13g2_decap_8 FILLER_51_283 ();
 sg13g2_fill_2 FILLER_51_290 ();
 sg13g2_decap_8 FILLER_51_297 ();
 sg13g2_decap_4 FILLER_51_304 ();
 sg13g2_decap_4 FILLER_51_312 ();
 sg13g2_fill_1 FILLER_51_316 ();
 sg13g2_fill_1 FILLER_51_322 ();
 sg13g2_fill_2 FILLER_51_328 ();
 sg13g2_decap_4 FILLER_51_333 ();
 sg13g2_fill_2 FILLER_51_337 ();
 sg13g2_decap_4 FILLER_51_348 ();
 sg13g2_decap_8 FILLER_51_356 ();
 sg13g2_decap_8 FILLER_51_363 ();
 sg13g2_decap_8 FILLER_51_370 ();
 sg13g2_decap_8 FILLER_51_377 ();
 sg13g2_decap_8 FILLER_51_384 ();
 sg13g2_fill_2 FILLER_51_391 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_decap_8 FILLER_51_406 ();
 sg13g2_decap_8 FILLER_51_419 ();
 sg13g2_decap_8 FILLER_51_426 ();
 sg13g2_fill_2 FILLER_51_433 ();
 sg13g2_fill_1 FILLER_51_435 ();
 sg13g2_decap_8 FILLER_51_442 ();
 sg13g2_decap_8 FILLER_51_449 ();
 sg13g2_decap_8 FILLER_51_456 ();
 sg13g2_decap_8 FILLER_51_468 ();
 sg13g2_fill_2 FILLER_51_475 ();
 sg13g2_decap_4 FILLER_51_481 ();
 sg13g2_decap_8 FILLER_51_499 ();
 sg13g2_decap_8 FILLER_51_506 ();
 sg13g2_decap_8 FILLER_51_513 ();
 sg13g2_decap_8 FILLER_51_520 ();
 sg13g2_decap_8 FILLER_51_527 ();
 sg13g2_decap_8 FILLER_51_534 ();
 sg13g2_fill_1 FILLER_51_541 ();
 sg13g2_decap_4 FILLER_51_551 ();
 sg13g2_fill_1 FILLER_51_555 ();
 sg13g2_fill_2 FILLER_51_560 ();
 sg13g2_fill_1 FILLER_51_562 ();
 sg13g2_decap_8 FILLER_51_568 ();
 sg13g2_decap_8 FILLER_51_575 ();
 sg13g2_decap_8 FILLER_51_582 ();
 sg13g2_decap_8 FILLER_51_589 ();
 sg13g2_decap_8 FILLER_51_596 ();
 sg13g2_decap_8 FILLER_51_603 ();
 sg13g2_decap_8 FILLER_51_610 ();
 sg13g2_decap_8 FILLER_51_617 ();
 sg13g2_decap_8 FILLER_51_624 ();
 sg13g2_decap_8 FILLER_51_631 ();
 sg13g2_decap_8 FILLER_51_642 ();
 sg13g2_decap_8 FILLER_51_649 ();
 sg13g2_decap_4 FILLER_51_661 ();
 sg13g2_decap_4 FILLER_51_669 ();
 sg13g2_fill_1 FILLER_51_678 ();
 sg13g2_fill_1 FILLER_51_684 ();
 sg13g2_fill_2 FILLER_51_690 ();
 sg13g2_fill_1 FILLER_51_692 ();
 sg13g2_decap_8 FILLER_51_698 ();
 sg13g2_fill_1 FILLER_51_705 ();
 sg13g2_decap_8 FILLER_51_711 ();
 sg13g2_decap_8 FILLER_51_718 ();
 sg13g2_decap_8 FILLER_51_725 ();
 sg13g2_decap_8 FILLER_51_732 ();
 sg13g2_fill_2 FILLER_51_739 ();
 sg13g2_fill_1 FILLER_51_747 ();
 sg13g2_decap_8 FILLER_51_752 ();
 sg13g2_decap_8 FILLER_51_759 ();
 sg13g2_decap_8 FILLER_51_766 ();
 sg13g2_decap_8 FILLER_51_773 ();
 sg13g2_decap_8 FILLER_51_780 ();
 sg13g2_decap_8 FILLER_51_787 ();
 sg13g2_decap_8 FILLER_51_794 ();
 sg13g2_decap_8 FILLER_51_801 ();
 sg13g2_decap_8 FILLER_51_808 ();
 sg13g2_decap_8 FILLER_51_815 ();
 sg13g2_decap_8 FILLER_51_822 ();
 sg13g2_decap_8 FILLER_51_829 ();
 sg13g2_decap_8 FILLER_51_836 ();
 sg13g2_decap_8 FILLER_51_843 ();
 sg13g2_decap_8 FILLER_51_850 ();
 sg13g2_decap_8 FILLER_51_857 ();
 sg13g2_decap_8 FILLER_51_864 ();
 sg13g2_decap_8 FILLER_51_871 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_4 FILLER_52_28 ();
 sg13g2_fill_2 FILLER_52_32 ();
 sg13g2_fill_2 FILLER_52_57 ();
 sg13g2_decap_4 FILLER_52_63 ();
 sg13g2_fill_1 FILLER_52_67 ();
 sg13g2_decap_8 FILLER_52_79 ();
 sg13g2_fill_2 FILLER_52_90 ();
 sg13g2_fill_1 FILLER_52_92 ();
 sg13g2_decap_8 FILLER_52_97 ();
 sg13g2_fill_2 FILLER_52_113 ();
 sg13g2_fill_2 FILLER_52_119 ();
 sg13g2_fill_1 FILLER_52_121 ();
 sg13g2_decap_8 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_137 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_fill_2 FILLER_52_153 ();
 sg13g2_fill_1 FILLER_52_155 ();
 sg13g2_fill_1 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_172 ();
 sg13g2_decap_4 FILLER_52_183 ();
 sg13g2_fill_2 FILLER_52_187 ();
 sg13g2_decap_8 FILLER_52_193 ();
 sg13g2_fill_1 FILLER_52_200 ();
 sg13g2_decap_8 FILLER_52_204 ();
 sg13g2_decap_8 FILLER_52_211 ();
 sg13g2_decap_8 FILLER_52_223 ();
 sg13g2_decap_8 FILLER_52_230 ();
 sg13g2_decap_8 FILLER_52_237 ();
 sg13g2_decap_8 FILLER_52_244 ();
 sg13g2_fill_2 FILLER_52_251 ();
 sg13g2_fill_1 FILLER_52_253 ();
 sg13g2_fill_1 FILLER_52_259 ();
 sg13g2_fill_1 FILLER_52_265 ();
 sg13g2_decap_4 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_274 ();
 sg13g2_decap_4 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_286 ();
 sg13g2_decap_8 FILLER_52_291 ();
 sg13g2_decap_4 FILLER_52_298 ();
 sg13g2_fill_2 FILLER_52_306 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_fill_2 FILLER_52_318 ();
 sg13g2_decap_8 FILLER_52_325 ();
 sg13g2_decap_8 FILLER_52_332 ();
 sg13g2_decap_8 FILLER_52_339 ();
 sg13g2_decap_8 FILLER_52_346 ();
 sg13g2_decap_8 FILLER_52_353 ();
 sg13g2_fill_1 FILLER_52_360 ();
 sg13g2_decap_4 FILLER_52_365 ();
 sg13g2_fill_1 FILLER_52_369 ();
 sg13g2_fill_2 FILLER_52_374 ();
 sg13g2_decap_8 FILLER_52_382 ();
 sg13g2_decap_4 FILLER_52_389 ();
 sg13g2_fill_2 FILLER_52_393 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_fill_2 FILLER_52_406 ();
 sg13g2_fill_2 FILLER_52_422 ();
 sg13g2_fill_1 FILLER_52_424 ();
 sg13g2_fill_2 FILLER_52_430 ();
 sg13g2_decap_4 FILLER_52_438 ();
 sg13g2_fill_2 FILLER_52_446 ();
 sg13g2_fill_2 FILLER_52_453 ();
 sg13g2_decap_8 FILLER_52_460 ();
 sg13g2_decap_8 FILLER_52_467 ();
 sg13g2_decap_4 FILLER_52_474 ();
 sg13g2_decap_8 FILLER_52_486 ();
 sg13g2_fill_2 FILLER_52_493 ();
 sg13g2_decap_4 FILLER_52_500 ();
 sg13g2_decap_8 FILLER_52_517 ();
 sg13g2_fill_2 FILLER_52_524 ();
 sg13g2_decap_8 FILLER_52_531 ();
 sg13g2_decap_4 FILLER_52_538 ();
 sg13g2_decap_8 FILLER_52_546 ();
 sg13g2_fill_2 FILLER_52_553 ();
 sg13g2_fill_1 FILLER_52_555 ();
 sg13g2_fill_2 FILLER_52_560 ();
 sg13g2_decap_8 FILLER_52_577 ();
 sg13g2_decap_8 FILLER_52_584 ();
 sg13g2_fill_2 FILLER_52_591 ();
 sg13g2_decap_8 FILLER_52_601 ();
 sg13g2_fill_2 FILLER_52_608 ();
 sg13g2_fill_1 FILLER_52_615 ();
 sg13g2_decap_4 FILLER_52_620 ();
 sg13g2_fill_1 FILLER_52_624 ();
 sg13g2_decap_8 FILLER_52_634 ();
 sg13g2_decap_8 FILLER_52_641 ();
 sg13g2_decap_8 FILLER_52_654 ();
 sg13g2_decap_8 FILLER_52_661 ();
 sg13g2_decap_4 FILLER_52_668 ();
 sg13g2_decap_8 FILLER_52_676 ();
 sg13g2_fill_2 FILLER_52_683 ();
 sg13g2_fill_1 FILLER_52_685 ();
 sg13g2_decap_8 FILLER_52_691 ();
 sg13g2_fill_1 FILLER_52_698 ();
 sg13g2_decap_4 FILLER_52_705 ();
 sg13g2_decap_4 FILLER_52_715 ();
 sg13g2_fill_2 FILLER_52_719 ();
 sg13g2_decap_8 FILLER_52_725 ();
 sg13g2_decap_8 FILLER_52_732 ();
 sg13g2_fill_2 FILLER_52_743 ();
 sg13g2_decap_4 FILLER_52_749 ();
 sg13g2_fill_1 FILLER_52_753 ();
 sg13g2_fill_2 FILLER_52_763 ();
 sg13g2_decap_8 FILLER_52_769 ();
 sg13g2_decap_8 FILLER_52_776 ();
 sg13g2_decap_8 FILLER_52_783 ();
 sg13g2_decap_8 FILLER_52_790 ();
 sg13g2_decap_8 FILLER_52_797 ();
 sg13g2_decap_8 FILLER_52_804 ();
 sg13g2_decap_8 FILLER_52_811 ();
 sg13g2_decap_8 FILLER_52_818 ();
 sg13g2_decap_8 FILLER_52_825 ();
 sg13g2_decap_8 FILLER_52_832 ();
 sg13g2_decap_8 FILLER_52_839 ();
 sg13g2_decap_8 FILLER_52_846 ();
 sg13g2_decap_8 FILLER_52_853 ();
 sg13g2_decap_8 FILLER_52_860 ();
 sg13g2_decap_8 FILLER_52_867 ();
 sg13g2_decap_4 FILLER_52_874 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_53 ();
 sg13g2_decap_8 FILLER_53_60 ();
 sg13g2_decap_4 FILLER_53_67 ();
 sg13g2_fill_1 FILLER_53_71 ();
 sg13g2_decap_4 FILLER_53_76 ();
 sg13g2_decap_8 FILLER_53_88 ();
 sg13g2_fill_2 FILLER_53_95 ();
 sg13g2_decap_8 FILLER_53_106 ();
 sg13g2_decap_8 FILLER_53_113 ();
 sg13g2_fill_2 FILLER_53_124 ();
 sg13g2_fill_2 FILLER_53_135 ();
 sg13g2_decap_4 FILLER_53_141 ();
 sg13g2_fill_2 FILLER_53_145 ();
 sg13g2_fill_2 FILLER_53_157 ();
 sg13g2_fill_1 FILLER_53_159 ();
 sg13g2_fill_2 FILLER_53_164 ();
 sg13g2_fill_1 FILLER_53_166 ();
 sg13g2_decap_8 FILLER_53_171 ();
 sg13g2_decap_8 FILLER_53_178 ();
 sg13g2_decap_8 FILLER_53_185 ();
 sg13g2_decap_8 FILLER_53_192 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_decap_8 FILLER_53_225 ();
 sg13g2_decap_8 FILLER_53_232 ();
 sg13g2_decap_8 FILLER_53_239 ();
 sg13g2_decap_8 FILLER_53_246 ();
 sg13g2_decap_4 FILLER_53_253 ();
 sg13g2_fill_1 FILLER_53_262 ();
 sg13g2_decap_4 FILLER_53_272 ();
 sg13g2_fill_2 FILLER_53_279 ();
 sg13g2_fill_1 FILLER_53_281 ();
 sg13g2_decap_8 FILLER_53_287 ();
 sg13g2_decap_8 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_301 ();
 sg13g2_decap_4 FILLER_53_308 ();
 sg13g2_fill_1 FILLER_53_312 ();
 sg13g2_decap_8 FILLER_53_320 ();
 sg13g2_decap_8 FILLER_53_327 ();
 sg13g2_decap_8 FILLER_53_334 ();
 sg13g2_decap_8 FILLER_53_341 ();
 sg13g2_fill_1 FILLER_53_348 ();
 sg13g2_decap_8 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_361 ();
 sg13g2_decap_4 FILLER_53_366 ();
 sg13g2_decap_8 FILLER_53_380 ();
 sg13g2_decap_8 FILLER_53_387 ();
 sg13g2_decap_8 FILLER_53_424 ();
 sg13g2_decap_8 FILLER_53_431 ();
 sg13g2_decap_8 FILLER_53_438 ();
 sg13g2_decap_8 FILLER_53_445 ();
 sg13g2_decap_8 FILLER_53_452 ();
 sg13g2_decap_8 FILLER_53_459 ();
 sg13g2_decap_8 FILLER_53_466 ();
 sg13g2_fill_2 FILLER_53_473 ();
 sg13g2_decap_8 FILLER_53_484 ();
 sg13g2_decap_8 FILLER_53_491 ();
 sg13g2_decap_8 FILLER_53_498 ();
 sg13g2_decap_8 FILLER_53_505 ();
 sg13g2_decap_8 FILLER_53_512 ();
 sg13g2_decap_8 FILLER_53_519 ();
 sg13g2_decap_4 FILLER_53_526 ();
 sg13g2_fill_1 FILLER_53_530 ();
 sg13g2_fill_2 FILLER_53_537 ();
 sg13g2_fill_1 FILLER_53_548 ();
 sg13g2_fill_2 FILLER_53_566 ();
 sg13g2_fill_1 FILLER_53_568 ();
 sg13g2_decap_8 FILLER_53_574 ();
 sg13g2_decap_8 FILLER_53_581 ();
 sg13g2_fill_2 FILLER_53_588 ();
 sg13g2_decap_4 FILLER_53_598 ();
 sg13g2_fill_1 FILLER_53_602 ();
 sg13g2_decap_8 FILLER_53_608 ();
 sg13g2_decap_8 FILLER_53_615 ();
 sg13g2_decap_4 FILLER_53_622 ();
 sg13g2_fill_2 FILLER_53_626 ();
 sg13g2_fill_2 FILLER_53_635 ();
 sg13g2_fill_1 FILLER_53_637 ();
 sg13g2_decap_8 FILLER_53_642 ();
 sg13g2_fill_2 FILLER_53_649 ();
 sg13g2_fill_1 FILLER_53_651 ();
 sg13g2_decap_8 FILLER_53_657 ();
 sg13g2_decap_8 FILLER_53_664 ();
 sg13g2_fill_2 FILLER_53_671 ();
 sg13g2_fill_1 FILLER_53_673 ();
 sg13g2_decap_8 FILLER_53_693 ();
 sg13g2_decap_8 FILLER_53_705 ();
 sg13g2_fill_1 FILLER_53_712 ();
 sg13g2_decap_8 FILLER_53_717 ();
 sg13g2_decap_8 FILLER_53_724 ();
 sg13g2_decap_8 FILLER_53_731 ();
 sg13g2_decap_4 FILLER_53_738 ();
 sg13g2_fill_2 FILLER_53_742 ();
 sg13g2_decap_8 FILLER_53_752 ();
 sg13g2_decap_8 FILLER_53_759 ();
 sg13g2_decap_8 FILLER_53_766 ();
 sg13g2_decap_8 FILLER_53_773 ();
 sg13g2_decap_8 FILLER_53_780 ();
 sg13g2_decap_8 FILLER_53_787 ();
 sg13g2_decap_8 FILLER_53_794 ();
 sg13g2_decap_8 FILLER_53_801 ();
 sg13g2_decap_8 FILLER_53_808 ();
 sg13g2_decap_8 FILLER_53_815 ();
 sg13g2_decap_8 FILLER_53_822 ();
 sg13g2_decap_8 FILLER_53_829 ();
 sg13g2_decap_8 FILLER_53_836 ();
 sg13g2_decap_8 FILLER_53_843 ();
 sg13g2_decap_8 FILLER_53_850 ();
 sg13g2_decap_8 FILLER_53_857 ();
 sg13g2_decap_8 FILLER_53_864 ();
 sg13g2_decap_8 FILLER_53_871 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_4 FILLER_54_49 ();
 sg13g2_fill_2 FILLER_54_53 ();
 sg13g2_fill_1 FILLER_54_59 ();
 sg13g2_decap_4 FILLER_54_65 ();
 sg13g2_fill_2 FILLER_54_69 ();
 sg13g2_decap_4 FILLER_54_76 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_102 ();
 sg13g2_decap_8 FILLER_54_109 ();
 sg13g2_decap_8 FILLER_54_116 ();
 sg13g2_decap_8 FILLER_54_123 ();
 sg13g2_decap_8 FILLER_54_130 ();
 sg13g2_decap_8 FILLER_54_137 ();
 sg13g2_fill_2 FILLER_54_144 ();
 sg13g2_decap_8 FILLER_54_151 ();
 sg13g2_decap_8 FILLER_54_158 ();
 sg13g2_decap_8 FILLER_54_165 ();
 sg13g2_decap_4 FILLER_54_172 ();
 sg13g2_fill_2 FILLER_54_176 ();
 sg13g2_decap_4 FILLER_54_183 ();
 sg13g2_fill_2 FILLER_54_187 ();
 sg13g2_decap_4 FILLER_54_194 ();
 sg13g2_fill_1 FILLER_54_198 ();
 sg13g2_decap_8 FILLER_54_209 ();
 sg13g2_decap_4 FILLER_54_216 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_decap_8 FILLER_54_229 ();
 sg13g2_decap_8 FILLER_54_241 ();
 sg13g2_decap_8 FILLER_54_248 ();
 sg13g2_decap_4 FILLER_54_264 ();
 sg13g2_fill_1 FILLER_54_268 ();
 sg13g2_fill_2 FILLER_54_274 ();
 sg13g2_fill_1 FILLER_54_276 ();
 sg13g2_decap_8 FILLER_54_281 ();
 sg13g2_decap_8 FILLER_54_288 ();
 sg13g2_decap_8 FILLER_54_295 ();
 sg13g2_decap_8 FILLER_54_302 ();
 sg13g2_decap_8 FILLER_54_309 ();
 sg13g2_decap_4 FILLER_54_316 ();
 sg13g2_decap_8 FILLER_54_325 ();
 sg13g2_decap_8 FILLER_54_332 ();
 sg13g2_decap_8 FILLER_54_339 ();
 sg13g2_decap_8 FILLER_54_346 ();
 sg13g2_decap_8 FILLER_54_353 ();
 sg13g2_decap_8 FILLER_54_360 ();
 sg13g2_decap_4 FILLER_54_367 ();
 sg13g2_decap_8 FILLER_54_375 ();
 sg13g2_decap_4 FILLER_54_382 ();
 sg13g2_fill_1 FILLER_54_386 ();
 sg13g2_decap_8 FILLER_54_391 ();
 sg13g2_decap_4 FILLER_54_398 ();
 sg13g2_fill_1 FILLER_54_406 ();
 sg13g2_decap_8 FILLER_54_421 ();
 sg13g2_decap_4 FILLER_54_436 ();
 sg13g2_fill_2 FILLER_54_440 ();
 sg13g2_fill_2 FILLER_54_450 ();
 sg13g2_decap_4 FILLER_54_457 ();
 sg13g2_fill_1 FILLER_54_461 ();
 sg13g2_decap_8 FILLER_54_467 ();
 sg13g2_decap_8 FILLER_54_474 ();
 sg13g2_decap_8 FILLER_54_481 ();
 sg13g2_decap_8 FILLER_54_488 ();
 sg13g2_decap_8 FILLER_54_495 ();
 sg13g2_decap_8 FILLER_54_502 ();
 sg13g2_decap_4 FILLER_54_509 ();
 sg13g2_fill_2 FILLER_54_513 ();
 sg13g2_decap_4 FILLER_54_519 ();
 sg13g2_fill_1 FILLER_54_523 ();
 sg13g2_decap_8 FILLER_54_533 ();
 sg13g2_fill_1 FILLER_54_540 ();
 sg13g2_fill_2 FILLER_54_547 ();
 sg13g2_fill_1 FILLER_54_549 ();
 sg13g2_decap_8 FILLER_54_560 ();
 sg13g2_fill_2 FILLER_54_572 ();
 sg13g2_decap_8 FILLER_54_579 ();
 sg13g2_decap_8 FILLER_54_586 ();
 sg13g2_decap_8 FILLER_54_593 ();
 sg13g2_fill_1 FILLER_54_600 ();
 sg13g2_decap_8 FILLER_54_609 ();
 sg13g2_decap_8 FILLER_54_616 ();
 sg13g2_fill_2 FILLER_54_623 ();
 sg13g2_fill_1 FILLER_54_625 ();
 sg13g2_fill_1 FILLER_54_630 ();
 sg13g2_decap_8 FILLER_54_641 ();
 sg13g2_decap_4 FILLER_54_648 ();
 sg13g2_decap_8 FILLER_54_655 ();
 sg13g2_decap_4 FILLER_54_662 ();
 sg13g2_decap_8 FILLER_54_670 ();
 sg13g2_decap_8 FILLER_54_677 ();
 sg13g2_fill_1 FILLER_54_684 ();
 sg13g2_fill_2 FILLER_54_689 ();
 sg13g2_fill_1 FILLER_54_691 ();
 sg13g2_decap_4 FILLER_54_696 ();
 sg13g2_fill_1 FILLER_54_700 ();
 sg13g2_fill_1 FILLER_54_710 ();
 sg13g2_decap_8 FILLER_54_725 ();
 sg13g2_decap_8 FILLER_54_732 ();
 sg13g2_decap_4 FILLER_54_739 ();
 sg13g2_fill_2 FILLER_54_743 ();
 sg13g2_decap_8 FILLER_54_749 ();
 sg13g2_decap_8 FILLER_54_756 ();
 sg13g2_decap_8 FILLER_54_763 ();
 sg13g2_decap_8 FILLER_54_770 ();
 sg13g2_decap_8 FILLER_54_777 ();
 sg13g2_decap_8 FILLER_54_784 ();
 sg13g2_decap_8 FILLER_54_791 ();
 sg13g2_decap_8 FILLER_54_798 ();
 sg13g2_decap_8 FILLER_54_805 ();
 sg13g2_decap_8 FILLER_54_812 ();
 sg13g2_decap_8 FILLER_54_819 ();
 sg13g2_decap_8 FILLER_54_826 ();
 sg13g2_decap_8 FILLER_54_833 ();
 sg13g2_decap_8 FILLER_54_840 ();
 sg13g2_decap_8 FILLER_54_847 ();
 sg13g2_decap_8 FILLER_54_854 ();
 sg13g2_decap_8 FILLER_54_861 ();
 sg13g2_decap_8 FILLER_54_868 ();
 sg13g2_fill_2 FILLER_54_875 ();
 sg13g2_fill_1 FILLER_54_877 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_4 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_39 ();
 sg13g2_decap_8 FILLER_55_51 ();
 sg13g2_fill_1 FILLER_55_58 ();
 sg13g2_decap_4 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_72 ();
 sg13g2_fill_1 FILLER_55_79 ();
 sg13g2_decap_8 FILLER_55_85 ();
 sg13g2_decap_4 FILLER_55_92 ();
 sg13g2_decap_8 FILLER_55_101 ();
 sg13g2_decap_8 FILLER_55_108 ();
 sg13g2_decap_8 FILLER_55_115 ();
 sg13g2_decap_8 FILLER_55_122 ();
 sg13g2_decap_4 FILLER_55_134 ();
 sg13g2_fill_1 FILLER_55_138 ();
 sg13g2_fill_2 FILLER_55_143 ();
 sg13g2_fill_1 FILLER_55_145 ();
 sg13g2_decap_8 FILLER_55_155 ();
 sg13g2_decap_8 FILLER_55_162 ();
 sg13g2_decap_8 FILLER_55_169 ();
 sg13g2_decap_4 FILLER_55_176 ();
 sg13g2_fill_2 FILLER_55_189 ();
 sg13g2_decap_8 FILLER_55_195 ();
 sg13g2_fill_2 FILLER_55_202 ();
 sg13g2_fill_1 FILLER_55_204 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_4 FILLER_55_217 ();
 sg13g2_decap_8 FILLER_55_230 ();
 sg13g2_decap_8 FILLER_55_237 ();
 sg13g2_decap_4 FILLER_55_244 ();
 sg13g2_decap_8 FILLER_55_260 ();
 sg13g2_decap_4 FILLER_55_267 ();
 sg13g2_fill_1 FILLER_55_271 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_4 FILLER_55_287 ();
 sg13g2_fill_1 FILLER_55_291 ();
 sg13g2_fill_1 FILLER_55_296 ();
 sg13g2_decap_8 FILLER_55_301 ();
 sg13g2_decap_8 FILLER_55_308 ();
 sg13g2_fill_2 FILLER_55_315 ();
 sg13g2_fill_1 FILLER_55_317 ();
 sg13g2_decap_4 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_326 ();
 sg13g2_decap_8 FILLER_55_336 ();
 sg13g2_decap_8 FILLER_55_343 ();
 sg13g2_decap_8 FILLER_55_350 ();
 sg13g2_fill_2 FILLER_55_357 ();
 sg13g2_fill_1 FILLER_55_359 ();
 sg13g2_decap_8 FILLER_55_363 ();
 sg13g2_decap_8 FILLER_55_374 ();
 sg13g2_decap_4 FILLER_55_381 ();
 sg13g2_fill_2 FILLER_55_385 ();
 sg13g2_decap_4 FILLER_55_391 ();
 sg13g2_fill_2 FILLER_55_395 ();
 sg13g2_decap_4 FILLER_55_405 ();
 sg13g2_fill_2 FILLER_55_409 ();
 sg13g2_decap_8 FILLER_55_416 ();
 sg13g2_decap_4 FILLER_55_423 ();
 sg13g2_decap_8 FILLER_55_432 ();
 sg13g2_fill_2 FILLER_55_439 ();
 sg13g2_fill_1 FILLER_55_441 ();
 sg13g2_decap_4 FILLER_55_460 ();
 sg13g2_fill_2 FILLER_55_464 ();
 sg13g2_decap_8 FILLER_55_481 ();
 sg13g2_decap_4 FILLER_55_488 ();
 sg13g2_fill_1 FILLER_55_492 ();
 sg13g2_fill_2 FILLER_55_500 ();
 sg13g2_fill_1 FILLER_55_502 ();
 sg13g2_decap_8 FILLER_55_508 ();
 sg13g2_decap_8 FILLER_55_515 ();
 sg13g2_decap_8 FILLER_55_531 ();
 sg13g2_decap_8 FILLER_55_538 ();
 sg13g2_decap_4 FILLER_55_550 ();
 sg13g2_decap_4 FILLER_55_559 ();
 sg13g2_decap_8 FILLER_55_572 ();
 sg13g2_decap_4 FILLER_55_579 ();
 sg13g2_decap_4 FILLER_55_588 ();
 sg13g2_fill_1 FILLER_55_602 ();
 sg13g2_decap_8 FILLER_55_608 ();
 sg13g2_decap_8 FILLER_55_615 ();
 sg13g2_decap_8 FILLER_55_622 ();
 sg13g2_decap_8 FILLER_55_629 ();
 sg13g2_decap_8 FILLER_55_636 ();
 sg13g2_decap_8 FILLER_55_643 ();
 sg13g2_decap_4 FILLER_55_650 ();
 sg13g2_decap_4 FILLER_55_659 ();
 sg13g2_fill_1 FILLER_55_663 ();
 sg13g2_decap_8 FILLER_55_669 ();
 sg13g2_decap_8 FILLER_55_676 ();
 sg13g2_fill_2 FILLER_55_683 ();
 sg13g2_fill_1 FILLER_55_685 ();
 sg13g2_decap_8 FILLER_55_694 ();
 sg13g2_fill_1 FILLER_55_701 ();
 sg13g2_decap_4 FILLER_55_707 ();
 sg13g2_fill_2 FILLER_55_715 ();
 sg13g2_decap_8 FILLER_55_722 ();
 sg13g2_decap_4 FILLER_55_729 ();
 sg13g2_fill_1 FILLER_55_733 ();
 sg13g2_decap_4 FILLER_55_738 ();
 sg13g2_fill_1 FILLER_55_742 ();
 sg13g2_decap_8 FILLER_55_747 ();
 sg13g2_fill_2 FILLER_55_754 ();
 sg13g2_decap_8 FILLER_55_765 ();
 sg13g2_decap_8 FILLER_55_772 ();
 sg13g2_decap_8 FILLER_55_779 ();
 sg13g2_decap_8 FILLER_55_786 ();
 sg13g2_decap_8 FILLER_55_793 ();
 sg13g2_decap_8 FILLER_55_800 ();
 sg13g2_decap_8 FILLER_55_807 ();
 sg13g2_decap_8 FILLER_55_814 ();
 sg13g2_decap_8 FILLER_55_821 ();
 sg13g2_decap_8 FILLER_55_828 ();
 sg13g2_decap_8 FILLER_55_835 ();
 sg13g2_decap_8 FILLER_55_842 ();
 sg13g2_decap_8 FILLER_55_849 ();
 sg13g2_decap_8 FILLER_55_856 ();
 sg13g2_decap_8 FILLER_55_863 ();
 sg13g2_decap_8 FILLER_55_870 ();
 sg13g2_fill_1 FILLER_55_877 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_4 FILLER_56_28 ();
 sg13g2_fill_1 FILLER_56_32 ();
 sg13g2_decap_8 FILLER_56_37 ();
 sg13g2_decap_4 FILLER_56_44 ();
 sg13g2_fill_2 FILLER_56_48 ();
 sg13g2_decap_8 FILLER_56_54 ();
 sg13g2_fill_2 FILLER_56_61 ();
 sg13g2_fill_1 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_68 ();
 sg13g2_fill_1 FILLER_56_75 ();
 sg13g2_fill_1 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_90 ();
 sg13g2_decap_8 FILLER_56_102 ();
 sg13g2_fill_2 FILLER_56_109 ();
 sg13g2_decap_8 FILLER_56_120 ();
 sg13g2_fill_2 FILLER_56_127 ();
 sg13g2_fill_1 FILLER_56_129 ();
 sg13g2_decap_4 FILLER_56_134 ();
 sg13g2_fill_2 FILLER_56_138 ();
 sg13g2_fill_1 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_151 ();
 sg13g2_fill_2 FILLER_56_157 ();
 sg13g2_decap_4 FILLER_56_172 ();
 sg13g2_decap_8 FILLER_56_180 ();
 sg13g2_decap_4 FILLER_56_187 ();
 sg13g2_fill_1 FILLER_56_191 ();
 sg13g2_fill_1 FILLER_56_197 ();
 sg13g2_fill_1 FILLER_56_202 ();
 sg13g2_decap_8 FILLER_56_213 ();
 sg13g2_decap_4 FILLER_56_220 ();
 sg13g2_fill_1 FILLER_56_224 ();
 sg13g2_decap_8 FILLER_56_229 ();
 sg13g2_decap_8 FILLER_56_241 ();
 sg13g2_decap_8 FILLER_56_248 ();
 sg13g2_decap_4 FILLER_56_255 ();
 sg13g2_fill_1 FILLER_56_259 ();
 sg13g2_decap_8 FILLER_56_273 ();
 sg13g2_decap_8 FILLER_56_280 ();
 sg13g2_decap_4 FILLER_56_287 ();
 sg13g2_fill_2 FILLER_56_291 ();
 sg13g2_fill_1 FILLER_56_301 ();
 sg13g2_decap_8 FILLER_56_312 ();
 sg13g2_decap_4 FILLER_56_319 ();
 sg13g2_decap_4 FILLER_56_328 ();
 sg13g2_fill_2 FILLER_56_337 ();
 sg13g2_fill_2 FILLER_56_344 ();
 sg13g2_fill_2 FILLER_56_351 ();
 sg13g2_fill_1 FILLER_56_353 ();
 sg13g2_decap_8 FILLER_56_359 ();
 sg13g2_decap_4 FILLER_56_366 ();
 sg13g2_fill_1 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_375 ();
 sg13g2_fill_2 FILLER_56_382 ();
 sg13g2_decap_8 FILLER_56_400 ();
 sg13g2_decap_8 FILLER_56_407 ();
 sg13g2_decap_4 FILLER_56_414 ();
 sg13g2_decap_8 FILLER_56_422 ();
 sg13g2_decap_4 FILLER_56_429 ();
 sg13g2_fill_2 FILLER_56_433 ();
 sg13g2_decap_4 FILLER_56_444 ();
 sg13g2_decap_8 FILLER_56_452 ();
 sg13g2_decap_8 FILLER_56_463 ();
 sg13g2_decap_4 FILLER_56_470 ();
 sg13g2_fill_1 FILLER_56_479 ();
 sg13g2_decap_8 FILLER_56_485 ();
 sg13g2_fill_1 FILLER_56_492 ();
 sg13g2_decap_8 FILLER_56_508 ();
 sg13g2_decap_8 FILLER_56_515 ();
 sg13g2_fill_2 FILLER_56_527 ();
 sg13g2_fill_1 FILLER_56_529 ();
 sg13g2_decap_8 FILLER_56_533 ();
 sg13g2_fill_1 FILLER_56_540 ();
 sg13g2_decap_8 FILLER_56_558 ();
 sg13g2_decap_4 FILLER_56_565 ();
 sg13g2_fill_2 FILLER_56_569 ();
 sg13g2_decap_4 FILLER_56_580 ();
 sg13g2_decap_8 FILLER_56_600 ();
 sg13g2_decap_8 FILLER_56_607 ();
 sg13g2_decap_8 FILLER_56_614 ();
 sg13g2_decap_8 FILLER_56_621 ();
 sg13g2_decap_8 FILLER_56_628 ();
 sg13g2_decap_4 FILLER_56_635 ();
 sg13g2_fill_1 FILLER_56_639 ();
 sg13g2_decap_8 FILLER_56_644 ();
 sg13g2_fill_1 FILLER_56_651 ();
 sg13g2_decap_8 FILLER_56_655 ();
 sg13g2_decap_8 FILLER_56_662 ();
 sg13g2_decap_4 FILLER_56_669 ();
 sg13g2_decap_4 FILLER_56_678 ();
 sg13g2_fill_2 FILLER_56_682 ();
 sg13g2_fill_1 FILLER_56_688 ();
 sg13g2_fill_2 FILLER_56_718 ();
 sg13g2_decap_4 FILLER_56_727 ();
 sg13g2_decap_8 FILLER_56_735 ();
 sg13g2_decap_8 FILLER_56_742 ();
 sg13g2_decap_8 FILLER_56_758 ();
 sg13g2_decap_8 FILLER_56_765 ();
 sg13g2_decap_8 FILLER_56_772 ();
 sg13g2_decap_8 FILLER_56_779 ();
 sg13g2_decap_8 FILLER_56_786 ();
 sg13g2_decap_8 FILLER_56_793 ();
 sg13g2_decap_8 FILLER_56_800 ();
 sg13g2_decap_8 FILLER_56_807 ();
 sg13g2_decap_8 FILLER_56_814 ();
 sg13g2_decap_8 FILLER_56_821 ();
 sg13g2_decap_8 FILLER_56_828 ();
 sg13g2_decap_8 FILLER_56_835 ();
 sg13g2_decap_8 FILLER_56_842 ();
 sg13g2_decap_8 FILLER_56_849 ();
 sg13g2_decap_8 FILLER_56_856 ();
 sg13g2_decap_8 FILLER_56_863 ();
 sg13g2_decap_8 FILLER_56_870 ();
 sg13g2_fill_1 FILLER_56_877 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_4 FILLER_57_77 ();
 sg13g2_fill_1 FILLER_57_85 ();
 sg13g2_decap_4 FILLER_57_90 ();
 sg13g2_fill_1 FILLER_57_94 ();
 sg13g2_decap_8 FILLER_57_104 ();
 sg13g2_decap_8 FILLER_57_111 ();
 sg13g2_decap_8 FILLER_57_118 ();
 sg13g2_decap_8 FILLER_57_125 ();
 sg13g2_decap_4 FILLER_57_132 ();
 sg13g2_decap_8 FILLER_57_144 ();
 sg13g2_decap_4 FILLER_57_151 ();
 sg13g2_fill_1 FILLER_57_155 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_4 FILLER_57_168 ();
 sg13g2_fill_2 FILLER_57_172 ();
 sg13g2_decap_8 FILLER_57_179 ();
 sg13g2_decap_8 FILLER_57_186 ();
 sg13g2_decap_8 FILLER_57_193 ();
 sg13g2_fill_2 FILLER_57_200 ();
 sg13g2_decap_8 FILLER_57_207 ();
 sg13g2_decap_8 FILLER_57_214 ();
 sg13g2_fill_1 FILLER_57_221 ();
 sg13g2_decap_8 FILLER_57_226 ();
 sg13g2_decap_8 FILLER_57_233 ();
 sg13g2_decap_8 FILLER_57_240 ();
 sg13g2_decap_8 FILLER_57_247 ();
 sg13g2_decap_8 FILLER_57_254 ();
 sg13g2_decap_8 FILLER_57_261 ();
 sg13g2_decap_4 FILLER_57_268 ();
 sg13g2_decap_8 FILLER_57_276 ();
 sg13g2_decap_8 FILLER_57_283 ();
 sg13g2_fill_2 FILLER_57_290 ();
 sg13g2_fill_2 FILLER_57_295 ();
 sg13g2_decap_8 FILLER_57_310 ();
 sg13g2_decap_8 FILLER_57_317 ();
 sg13g2_fill_2 FILLER_57_324 ();
 sg13g2_fill_1 FILLER_57_338 ();
 sg13g2_decap_8 FILLER_57_344 ();
 sg13g2_decap_8 FILLER_57_351 ();
 sg13g2_decap_8 FILLER_57_358 ();
 sg13g2_decap_8 FILLER_57_365 ();
 sg13g2_decap_8 FILLER_57_372 ();
 sg13g2_decap_8 FILLER_57_379 ();
 sg13g2_fill_1 FILLER_57_386 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_57_406 ();
 sg13g2_fill_2 FILLER_57_413 ();
 sg13g2_fill_1 FILLER_57_415 ();
 sg13g2_decap_8 FILLER_57_420 ();
 sg13g2_decap_8 FILLER_57_427 ();
 sg13g2_decap_8 FILLER_57_434 ();
 sg13g2_decap_8 FILLER_57_445 ();
 sg13g2_decap_8 FILLER_57_452 ();
 sg13g2_decap_8 FILLER_57_459 ();
 sg13g2_decap_8 FILLER_57_466 ();
 sg13g2_decap_8 FILLER_57_478 ();
 sg13g2_decap_8 FILLER_57_485 ();
 sg13g2_decap_4 FILLER_57_492 ();
 sg13g2_decap_8 FILLER_57_505 ();
 sg13g2_decap_8 FILLER_57_512 ();
 sg13g2_decap_4 FILLER_57_519 ();
 sg13g2_fill_1 FILLER_57_523 ();
 sg13g2_decap_8 FILLER_57_529 ();
 sg13g2_fill_1 FILLER_57_536 ();
 sg13g2_decap_4 FILLER_57_541 ();
 sg13g2_decap_8 FILLER_57_549 ();
 sg13g2_decap_8 FILLER_57_556 ();
 sg13g2_decap_4 FILLER_57_563 ();
 sg13g2_fill_2 FILLER_57_567 ();
 sg13g2_fill_2 FILLER_57_573 ();
 sg13g2_decap_8 FILLER_57_579 ();
 sg13g2_decap_4 FILLER_57_586 ();
 sg13g2_fill_1 FILLER_57_590 ();
 sg13g2_decap_8 FILLER_57_596 ();
 sg13g2_decap_8 FILLER_57_603 ();
 sg13g2_decap_8 FILLER_57_610 ();
 sg13g2_decap_8 FILLER_57_617 ();
 sg13g2_decap_8 FILLER_57_624 ();
 sg13g2_fill_2 FILLER_57_631 ();
 sg13g2_fill_1 FILLER_57_633 ();
 sg13g2_decap_4 FILLER_57_638 ();
 sg13g2_decap_8 FILLER_57_651 ();
 sg13g2_decap_8 FILLER_57_658 ();
 sg13g2_decap_8 FILLER_57_665 ();
 sg13g2_decap_8 FILLER_57_672 ();
 sg13g2_decap_8 FILLER_57_679 ();
 sg13g2_fill_2 FILLER_57_686 ();
 sg13g2_fill_1 FILLER_57_688 ();
 sg13g2_decap_4 FILLER_57_694 ();
 sg13g2_fill_2 FILLER_57_698 ();
 sg13g2_decap_8 FILLER_57_704 ();
 sg13g2_fill_2 FILLER_57_711 ();
 sg13g2_fill_1 FILLER_57_713 ();
 sg13g2_fill_1 FILLER_57_722 ();
 sg13g2_decap_4 FILLER_57_728 ();
 sg13g2_decap_8 FILLER_57_737 ();
 sg13g2_decap_8 FILLER_57_744 ();
 sg13g2_decap_8 FILLER_57_751 ();
 sg13g2_decap_8 FILLER_57_758 ();
 sg13g2_decap_8 FILLER_57_765 ();
 sg13g2_decap_8 FILLER_57_772 ();
 sg13g2_decap_8 FILLER_57_779 ();
 sg13g2_decap_8 FILLER_57_786 ();
 sg13g2_decap_8 FILLER_57_793 ();
 sg13g2_decap_8 FILLER_57_800 ();
 sg13g2_decap_8 FILLER_57_807 ();
 sg13g2_decap_8 FILLER_57_814 ();
 sg13g2_decap_8 FILLER_57_821 ();
 sg13g2_decap_8 FILLER_57_828 ();
 sg13g2_decap_8 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_842 ();
 sg13g2_decap_8 FILLER_57_849 ();
 sg13g2_decap_8 FILLER_57_856 ();
 sg13g2_decap_8 FILLER_57_863 ();
 sg13g2_decap_8 FILLER_57_870 ();
 sg13g2_fill_1 FILLER_57_877 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_4 FILLER_58_56 ();
 sg13g2_fill_1 FILLER_58_69 ();
 sg13g2_decap_4 FILLER_58_74 ();
 sg13g2_decap_4 FILLER_58_82 ();
 sg13g2_fill_2 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_118 ();
 sg13g2_fill_2 FILLER_58_125 ();
 sg13g2_decap_8 FILLER_58_131 ();
 sg13g2_decap_8 FILLER_58_146 ();
 sg13g2_decap_4 FILLER_58_153 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_fill_1 FILLER_58_173 ();
 sg13g2_decap_4 FILLER_58_178 ();
 sg13g2_fill_1 FILLER_58_182 ();
 sg13g2_decap_4 FILLER_58_187 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_fill_1 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_208 ();
 sg13g2_decap_8 FILLER_58_215 ();
 sg13g2_decap_8 FILLER_58_222 ();
 sg13g2_decap_8 FILLER_58_229 ();
 sg13g2_decap_8 FILLER_58_236 ();
 sg13g2_fill_2 FILLER_58_243 ();
 sg13g2_fill_1 FILLER_58_249 ();
 sg13g2_decap_8 FILLER_58_255 ();
 sg13g2_decap_8 FILLER_58_262 ();
 sg13g2_fill_1 FILLER_58_269 ();
 sg13g2_decap_8 FILLER_58_274 ();
 sg13g2_fill_2 FILLER_58_281 ();
 sg13g2_fill_1 FILLER_58_283 ();
 sg13g2_decap_8 FILLER_58_288 ();
 sg13g2_decap_8 FILLER_58_295 ();
 sg13g2_decap_8 FILLER_58_302 ();
 sg13g2_decap_4 FILLER_58_313 ();
 sg13g2_fill_2 FILLER_58_326 ();
 sg13g2_fill_1 FILLER_58_328 ();
 sg13g2_decap_4 FILLER_58_334 ();
 sg13g2_decap_8 FILLER_58_342 ();
 sg13g2_decap_8 FILLER_58_349 ();
 sg13g2_decap_8 FILLER_58_356 ();
 sg13g2_decap_8 FILLER_58_368 ();
 sg13g2_decap_8 FILLER_58_375 ();
 sg13g2_decap_8 FILLER_58_382 ();
 sg13g2_decap_8 FILLER_58_389 ();
 sg13g2_decap_8 FILLER_58_396 ();
 sg13g2_decap_8 FILLER_58_403 ();
 sg13g2_decap_4 FILLER_58_410 ();
 sg13g2_fill_2 FILLER_58_414 ();
 sg13g2_decap_8 FILLER_58_420 ();
 sg13g2_decap_8 FILLER_58_431 ();
 sg13g2_fill_1 FILLER_58_438 ();
 sg13g2_decap_8 FILLER_58_443 ();
 sg13g2_fill_2 FILLER_58_450 ();
 sg13g2_decap_8 FILLER_58_456 ();
 sg13g2_decap_8 FILLER_58_463 ();
 sg13g2_decap_8 FILLER_58_470 ();
 sg13g2_decap_8 FILLER_58_477 ();
 sg13g2_decap_8 FILLER_58_484 ();
 sg13g2_fill_2 FILLER_58_491 ();
 sg13g2_decap_8 FILLER_58_498 ();
 sg13g2_decap_8 FILLER_58_505 ();
 sg13g2_decap_8 FILLER_58_512 ();
 sg13g2_decap_4 FILLER_58_519 ();
 sg13g2_fill_1 FILLER_58_523 ();
 sg13g2_decap_4 FILLER_58_528 ();
 sg13g2_fill_2 FILLER_58_532 ();
 sg13g2_decap_4 FILLER_58_538 ();
 sg13g2_decap_8 FILLER_58_551 ();
 sg13g2_decap_8 FILLER_58_558 ();
 sg13g2_decap_4 FILLER_58_565 ();
 sg13g2_decap_8 FILLER_58_574 ();
 sg13g2_decap_8 FILLER_58_581 ();
 sg13g2_decap_4 FILLER_58_588 ();
 sg13g2_fill_1 FILLER_58_592 ();
 sg13g2_decap_4 FILLER_58_601 ();
 sg13g2_fill_2 FILLER_58_605 ();
 sg13g2_decap_8 FILLER_58_613 ();
 sg13g2_decap_8 FILLER_58_620 ();
 sg13g2_fill_2 FILLER_58_627 ();
 sg13g2_fill_1 FILLER_58_629 ();
 sg13g2_decap_4 FILLER_58_634 ();
 sg13g2_fill_2 FILLER_58_648 ();
 sg13g2_decap_8 FILLER_58_656 ();
 sg13g2_decap_8 FILLER_58_663 ();
 sg13g2_fill_1 FILLER_58_675 ();
 sg13g2_decap_8 FILLER_58_680 ();
 sg13g2_decap_8 FILLER_58_687 ();
 sg13g2_decap_8 FILLER_58_694 ();
 sg13g2_decap_4 FILLER_58_701 ();
 sg13g2_decap_4 FILLER_58_710 ();
 sg13g2_fill_1 FILLER_58_714 ();
 sg13g2_decap_8 FILLER_58_719 ();
 sg13g2_decap_8 FILLER_58_726 ();
 sg13g2_decap_8 FILLER_58_733 ();
 sg13g2_decap_8 FILLER_58_740 ();
 sg13g2_decap_8 FILLER_58_747 ();
 sg13g2_decap_8 FILLER_58_754 ();
 sg13g2_decap_8 FILLER_58_761 ();
 sg13g2_decap_8 FILLER_58_768 ();
 sg13g2_decap_8 FILLER_58_775 ();
 sg13g2_decap_8 FILLER_58_782 ();
 sg13g2_decap_8 FILLER_58_789 ();
 sg13g2_decap_8 FILLER_58_796 ();
 sg13g2_decap_8 FILLER_58_803 ();
 sg13g2_decap_8 FILLER_58_810 ();
 sg13g2_decap_8 FILLER_58_817 ();
 sg13g2_decap_8 FILLER_58_824 ();
 sg13g2_decap_8 FILLER_58_831 ();
 sg13g2_decap_8 FILLER_58_838 ();
 sg13g2_decap_8 FILLER_58_845 ();
 sg13g2_decap_8 FILLER_58_852 ();
 sg13g2_decap_8 FILLER_58_859 ();
 sg13g2_decap_8 FILLER_58_866 ();
 sg13g2_decap_4 FILLER_58_873 ();
 sg13g2_fill_1 FILLER_58_877 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_67 ();
 sg13g2_fill_2 FILLER_59_74 ();
 sg13g2_fill_1 FILLER_59_76 ();
 sg13g2_decap_8 FILLER_59_87 ();
 sg13g2_fill_1 FILLER_59_94 ();
 sg13g2_decap_8 FILLER_59_99 ();
 sg13g2_decap_8 FILLER_59_106 ();
 sg13g2_decap_8 FILLER_59_113 ();
 sg13g2_decap_8 FILLER_59_120 ();
 sg13g2_decap_8 FILLER_59_127 ();
 sg13g2_decap_8 FILLER_59_134 ();
 sg13g2_decap_8 FILLER_59_141 ();
 sg13g2_decap_8 FILLER_59_148 ();
 sg13g2_decap_8 FILLER_59_160 ();
 sg13g2_decap_4 FILLER_59_167 ();
 sg13g2_fill_2 FILLER_59_171 ();
 sg13g2_decap_8 FILLER_59_178 ();
 sg13g2_decap_4 FILLER_59_185 ();
 sg13g2_fill_2 FILLER_59_189 ();
 sg13g2_fill_1 FILLER_59_195 ();
 sg13g2_decap_4 FILLER_59_210 ();
 sg13g2_decap_8 FILLER_59_218 ();
 sg13g2_fill_2 FILLER_59_225 ();
 sg13g2_decap_8 FILLER_59_231 ();
 sg13g2_decap_8 FILLER_59_243 ();
 sg13g2_decap_4 FILLER_59_262 ();
 sg13g2_decap_4 FILLER_59_274 ();
 sg13g2_fill_1 FILLER_59_278 ();
 sg13g2_decap_8 FILLER_59_288 ();
 sg13g2_fill_1 FILLER_59_295 ();
 sg13g2_fill_2 FILLER_59_301 ();
 sg13g2_decap_4 FILLER_59_307 ();
 sg13g2_fill_2 FILLER_59_315 ();
 sg13g2_fill_2 FILLER_59_326 ();
 sg13g2_decap_8 FILLER_59_333 ();
 sg13g2_decap_8 FILLER_59_340 ();
 sg13g2_decap_8 FILLER_59_347 ();
 sg13g2_decap_4 FILLER_59_354 ();
 sg13g2_fill_1 FILLER_59_358 ();
 sg13g2_fill_1 FILLER_59_368 ();
 sg13g2_fill_1 FILLER_59_373 ();
 sg13g2_decap_8 FILLER_59_379 ();
 sg13g2_decap_4 FILLER_59_386 ();
 sg13g2_fill_1 FILLER_59_390 ();
 sg13g2_fill_2 FILLER_59_404 ();
 sg13g2_decap_8 FILLER_59_409 ();
 sg13g2_decap_8 FILLER_59_416 ();
 sg13g2_fill_1 FILLER_59_423 ();
 sg13g2_decap_8 FILLER_59_428 ();
 sg13g2_decap_8 FILLER_59_435 ();
 sg13g2_decap_8 FILLER_59_442 ();
 sg13g2_decap_4 FILLER_59_449 ();
 sg13g2_fill_1 FILLER_59_461 ();
 sg13g2_decap_8 FILLER_59_466 ();
 sg13g2_decap_8 FILLER_59_473 ();
 sg13g2_decap_8 FILLER_59_480 ();
 sg13g2_decap_8 FILLER_59_487 ();
 sg13g2_fill_2 FILLER_59_508 ();
 sg13g2_fill_2 FILLER_59_515 ();
 sg13g2_decap_8 FILLER_59_526 ();
 sg13g2_fill_1 FILLER_59_533 ();
 sg13g2_decap_8 FILLER_59_538 ();
 sg13g2_fill_2 FILLER_59_545 ();
 sg13g2_decap_8 FILLER_59_552 ();
 sg13g2_decap_8 FILLER_59_559 ();
 sg13g2_fill_2 FILLER_59_566 ();
 sg13g2_decap_4 FILLER_59_577 ();
 sg13g2_fill_2 FILLER_59_590 ();
 sg13g2_fill_1 FILLER_59_592 ();
 sg13g2_decap_4 FILLER_59_597 ();
 sg13g2_fill_1 FILLER_59_601 ();
 sg13g2_decap_8 FILLER_59_611 ();
 sg13g2_decap_8 FILLER_59_618 ();
 sg13g2_decap_4 FILLER_59_625 ();
 sg13g2_decap_4 FILLER_59_634 ();
 sg13g2_decap_8 FILLER_59_647 ();
 sg13g2_decap_4 FILLER_59_654 ();
 sg13g2_decap_8 FILLER_59_662 ();
 sg13g2_fill_2 FILLER_59_669 ();
 sg13g2_decap_4 FILLER_59_679 ();
 sg13g2_fill_1 FILLER_59_683 ();
 sg13g2_decap_8 FILLER_59_689 ();
 sg13g2_decap_4 FILLER_59_696 ();
 sg13g2_fill_2 FILLER_59_700 ();
 sg13g2_decap_8 FILLER_59_706 ();
 sg13g2_decap_4 FILLER_59_713 ();
 sg13g2_decap_8 FILLER_59_732 ();
 sg13g2_decap_8 FILLER_59_739 ();
 sg13g2_decap_8 FILLER_59_746 ();
 sg13g2_decap_8 FILLER_59_753 ();
 sg13g2_decap_8 FILLER_59_760 ();
 sg13g2_decap_8 FILLER_59_767 ();
 sg13g2_decap_8 FILLER_59_774 ();
 sg13g2_decap_8 FILLER_59_781 ();
 sg13g2_decap_8 FILLER_59_788 ();
 sg13g2_decap_8 FILLER_59_795 ();
 sg13g2_decap_8 FILLER_59_802 ();
 sg13g2_decap_8 FILLER_59_809 ();
 sg13g2_decap_8 FILLER_59_816 ();
 sg13g2_decap_8 FILLER_59_823 ();
 sg13g2_decap_8 FILLER_59_830 ();
 sg13g2_decap_8 FILLER_59_837 ();
 sg13g2_decap_8 FILLER_59_844 ();
 sg13g2_decap_8 FILLER_59_851 ();
 sg13g2_decap_8 FILLER_59_858 ();
 sg13g2_decap_8 FILLER_59_865 ();
 sg13g2_decap_4 FILLER_59_872 ();
 sg13g2_fill_2 FILLER_59_876 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_4 FILLER_60_77 ();
 sg13g2_fill_2 FILLER_60_81 ();
 sg13g2_decap_8 FILLER_60_88 ();
 sg13g2_decap_8 FILLER_60_95 ();
 sg13g2_decap_8 FILLER_60_102 ();
 sg13g2_decap_8 FILLER_60_109 ();
 sg13g2_decap_4 FILLER_60_116 ();
 sg13g2_fill_2 FILLER_60_120 ();
 sg13g2_decap_8 FILLER_60_127 ();
 sg13g2_decap_8 FILLER_60_134 ();
 sg13g2_decap_8 FILLER_60_141 ();
 sg13g2_decap_4 FILLER_60_148 ();
 sg13g2_decap_8 FILLER_60_156 ();
 sg13g2_fill_2 FILLER_60_163 ();
 sg13g2_decap_4 FILLER_60_169 ();
 sg13g2_fill_1 FILLER_60_173 ();
 sg13g2_decap_8 FILLER_60_178 ();
 sg13g2_decap_8 FILLER_60_185 ();
 sg13g2_decap_4 FILLER_60_192 ();
 sg13g2_fill_1 FILLER_60_196 ();
 sg13g2_fill_1 FILLER_60_201 ();
 sg13g2_fill_1 FILLER_60_206 ();
 sg13g2_decap_4 FILLER_60_219 ();
 sg13g2_fill_2 FILLER_60_223 ();
 sg13g2_decap_8 FILLER_60_229 ();
 sg13g2_fill_2 FILLER_60_236 ();
 sg13g2_fill_2 FILLER_60_242 ();
 sg13g2_decap_8 FILLER_60_248 ();
 sg13g2_decap_8 FILLER_60_255 ();
 sg13g2_decap_8 FILLER_60_262 ();
 sg13g2_fill_2 FILLER_60_269 ();
 sg13g2_fill_1 FILLER_60_271 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_fill_2 FILLER_60_287 ();
 sg13g2_fill_1 FILLER_60_289 ();
 sg13g2_fill_2 FILLER_60_294 ();
 sg13g2_fill_2 FILLER_60_300 ();
 sg13g2_decap_4 FILLER_60_307 ();
 sg13g2_fill_1 FILLER_60_311 ();
 sg13g2_decap_4 FILLER_60_325 ();
 sg13g2_fill_1 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_334 ();
 sg13g2_decap_8 FILLER_60_341 ();
 sg13g2_decap_8 FILLER_60_348 ();
 sg13g2_decap_8 FILLER_60_355 ();
 sg13g2_decap_4 FILLER_60_362 ();
 sg13g2_decap_4 FILLER_60_371 ();
 sg13g2_fill_1 FILLER_60_375 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_2 FILLER_60_397 ();
 sg13g2_decap_8 FILLER_60_412 ();
 sg13g2_fill_2 FILLER_60_419 ();
 sg13g2_decap_8 FILLER_60_426 ();
 sg13g2_decap_4 FILLER_60_433 ();
 sg13g2_fill_2 FILLER_60_437 ();
 sg13g2_decap_8 FILLER_60_442 ();
 sg13g2_fill_1 FILLER_60_449 ();
 sg13g2_decap_4 FILLER_60_455 ();
 sg13g2_fill_2 FILLER_60_459 ();
 sg13g2_decap_8 FILLER_60_465 ();
 sg13g2_decap_4 FILLER_60_472 ();
 sg13g2_fill_2 FILLER_60_476 ();
 sg13g2_decap_4 FILLER_60_482 ();
 sg13g2_fill_1 FILLER_60_486 ();
 sg13g2_decap_4 FILLER_60_497 ();
 sg13g2_fill_2 FILLER_60_501 ();
 sg13g2_decap_8 FILLER_60_509 ();
 sg13g2_decap_4 FILLER_60_516 ();
 sg13g2_decap_8 FILLER_60_525 ();
 sg13g2_decap_8 FILLER_60_532 ();
 sg13g2_fill_2 FILLER_60_539 ();
 sg13g2_fill_1 FILLER_60_541 ();
 sg13g2_decap_4 FILLER_60_553 ();
 sg13g2_fill_2 FILLER_60_557 ();
 sg13g2_decap_4 FILLER_60_563 ();
 sg13g2_decap_8 FILLER_60_571 ();
 sg13g2_decap_8 FILLER_60_578 ();
 sg13g2_decap_4 FILLER_60_585 ();
 sg13g2_decap_8 FILLER_60_594 ();
 sg13g2_fill_2 FILLER_60_601 ();
 sg13g2_decap_8 FILLER_60_608 ();
 sg13g2_decap_8 FILLER_60_615 ();
 sg13g2_decap_4 FILLER_60_622 ();
 sg13g2_decap_8 FILLER_60_630 ();
 sg13g2_decap_8 FILLER_60_637 ();
 sg13g2_decap_4 FILLER_60_644 ();
 sg13g2_fill_2 FILLER_60_648 ();
 sg13g2_decap_8 FILLER_60_654 ();
 sg13g2_fill_1 FILLER_60_661 ();
 sg13g2_decap_8 FILLER_60_667 ();
 sg13g2_decap_8 FILLER_60_674 ();
 sg13g2_decap_4 FILLER_60_681 ();
 sg13g2_fill_1 FILLER_60_685 ();
 sg13g2_fill_2 FILLER_60_694 ();
 sg13g2_fill_1 FILLER_60_696 ();
 sg13g2_decap_8 FILLER_60_706 ();
 sg13g2_decap_4 FILLER_60_713 ();
 sg13g2_fill_1 FILLER_60_717 ();
 sg13g2_decap_8 FILLER_60_722 ();
 sg13g2_decap_8 FILLER_60_729 ();
 sg13g2_decap_8 FILLER_60_736 ();
 sg13g2_decap_4 FILLER_60_743 ();
 sg13g2_decap_8 FILLER_60_752 ();
 sg13g2_decap_8 FILLER_60_759 ();
 sg13g2_decap_8 FILLER_60_766 ();
 sg13g2_decap_8 FILLER_60_773 ();
 sg13g2_decap_8 FILLER_60_780 ();
 sg13g2_decap_8 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_794 ();
 sg13g2_decap_8 FILLER_60_801 ();
 sg13g2_decap_8 FILLER_60_808 ();
 sg13g2_decap_8 FILLER_60_815 ();
 sg13g2_decap_8 FILLER_60_822 ();
 sg13g2_decap_8 FILLER_60_829 ();
 sg13g2_decap_8 FILLER_60_836 ();
 sg13g2_decap_8 FILLER_60_843 ();
 sg13g2_decap_8 FILLER_60_850 ();
 sg13g2_decap_8 FILLER_60_857 ();
 sg13g2_decap_8 FILLER_60_864 ();
 sg13g2_decap_8 FILLER_60_871 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_4 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_170 ();
 sg13g2_decap_8 FILLER_61_177 ();
 sg13g2_decap_8 FILLER_61_184 ();
 sg13g2_decap_8 FILLER_61_191 ();
 sg13g2_fill_1 FILLER_61_198 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_4 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_218 ();
 sg13g2_decap_8 FILLER_61_225 ();
 sg13g2_decap_8 FILLER_61_232 ();
 sg13g2_decap_8 FILLER_61_239 ();
 sg13g2_decap_8 FILLER_61_246 ();
 sg13g2_decap_8 FILLER_61_253 ();
 sg13g2_decap_8 FILLER_61_273 ();
 sg13g2_decap_8 FILLER_61_280 ();
 sg13g2_decap_8 FILLER_61_287 ();
 sg13g2_fill_2 FILLER_61_294 ();
 sg13g2_fill_1 FILLER_61_296 ();
 sg13g2_decap_4 FILLER_61_305 ();
 sg13g2_fill_2 FILLER_61_309 ();
 sg13g2_decap_4 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_327 ();
 sg13g2_decap_8 FILLER_61_334 ();
 sg13g2_decap_8 FILLER_61_341 ();
 sg13g2_decap_8 FILLER_61_348 ();
 sg13g2_decap_8 FILLER_61_355 ();
 sg13g2_fill_1 FILLER_61_362 ();
 sg13g2_decap_8 FILLER_61_368 ();
 sg13g2_decap_8 FILLER_61_375 ();
 sg13g2_fill_1 FILLER_61_382 ();
 sg13g2_fill_1 FILLER_61_387 ();
 sg13g2_fill_1 FILLER_61_392 ();
 sg13g2_decap_4 FILLER_61_403 ();
 sg13g2_decap_8 FILLER_61_411 ();
 sg13g2_decap_4 FILLER_61_418 ();
 sg13g2_fill_1 FILLER_61_422 ();
 sg13g2_decap_8 FILLER_61_427 ();
 sg13g2_fill_1 FILLER_61_434 ();
 sg13g2_decap_4 FILLER_61_439 ();
 sg13g2_fill_1 FILLER_61_443 ();
 sg13g2_fill_2 FILLER_61_449 ();
 sg13g2_fill_1 FILLER_61_451 ();
 sg13g2_decap_4 FILLER_61_456 ();
 sg13g2_fill_1 FILLER_61_460 ();
 sg13g2_decap_8 FILLER_61_468 ();
 sg13g2_decap_8 FILLER_61_475 ();
 sg13g2_decap_4 FILLER_61_482 ();
 sg13g2_fill_2 FILLER_61_486 ();
 sg13g2_decap_8 FILLER_61_496 ();
 sg13g2_decap_8 FILLER_61_503 ();
 sg13g2_decap_8 FILLER_61_510 ();
 sg13g2_decap_8 FILLER_61_529 ();
 sg13g2_decap_8 FILLER_61_541 ();
 sg13g2_fill_1 FILLER_61_548 ();
 sg13g2_fill_1 FILLER_61_553 ();
 sg13g2_decap_8 FILLER_61_559 ();
 sg13g2_decap_8 FILLER_61_571 ();
 sg13g2_decap_8 FILLER_61_578 ();
 sg13g2_decap_8 FILLER_61_585 ();
 sg13g2_decap_8 FILLER_61_592 ();
 sg13g2_decap_8 FILLER_61_599 ();
 sg13g2_decap_8 FILLER_61_606 ();
 sg13g2_decap_8 FILLER_61_613 ();
 sg13g2_fill_2 FILLER_61_620 ();
 sg13g2_decap_8 FILLER_61_638 ();
 sg13g2_fill_2 FILLER_61_645 ();
 sg13g2_fill_1 FILLER_61_647 ();
 sg13g2_decap_8 FILLER_61_657 ();
 sg13g2_decap_4 FILLER_61_664 ();
 sg13g2_fill_1 FILLER_61_668 ();
 sg13g2_decap_8 FILLER_61_677 ();
 sg13g2_decap_8 FILLER_61_688 ();
 sg13g2_decap_8 FILLER_61_695 ();
 sg13g2_decap_8 FILLER_61_702 ();
 sg13g2_decap_8 FILLER_61_709 ();
 sg13g2_decap_8 FILLER_61_716 ();
 sg13g2_decap_8 FILLER_61_723 ();
 sg13g2_decap_8 FILLER_61_730 ();
 sg13g2_decap_8 FILLER_61_737 ();
 sg13g2_decap_8 FILLER_61_744 ();
 sg13g2_decap_8 FILLER_61_751 ();
 sg13g2_decap_8 FILLER_61_758 ();
 sg13g2_decap_8 FILLER_61_765 ();
 sg13g2_decap_8 FILLER_61_772 ();
 sg13g2_decap_8 FILLER_61_779 ();
 sg13g2_decap_8 FILLER_61_786 ();
 sg13g2_decap_8 FILLER_61_793 ();
 sg13g2_decap_8 FILLER_61_800 ();
 sg13g2_decap_8 FILLER_61_807 ();
 sg13g2_decap_8 FILLER_61_814 ();
 sg13g2_decap_8 FILLER_61_821 ();
 sg13g2_decap_8 FILLER_61_828 ();
 sg13g2_decap_8 FILLER_61_835 ();
 sg13g2_decap_8 FILLER_61_842 ();
 sg13g2_decap_8 FILLER_61_849 ();
 sg13g2_decap_8 FILLER_61_856 ();
 sg13g2_decap_8 FILLER_61_863 ();
 sg13g2_decap_8 FILLER_61_870 ();
 sg13g2_fill_1 FILLER_61_877 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_60 ();
 sg13g2_decap_8 FILLER_62_67 ();
 sg13g2_decap_8 FILLER_62_74 ();
 sg13g2_decap_8 FILLER_62_111 ();
 sg13g2_decap_8 FILLER_62_118 ();
 sg13g2_decap_8 FILLER_62_125 ();
 sg13g2_decap_8 FILLER_62_132 ();
 sg13g2_decap_8 FILLER_62_139 ();
 sg13g2_decap_8 FILLER_62_146 ();
 sg13g2_decap_8 FILLER_62_153 ();
 sg13g2_decap_8 FILLER_62_160 ();
 sg13g2_fill_1 FILLER_62_167 ();
 sg13g2_decap_8 FILLER_62_172 ();
 sg13g2_decap_8 FILLER_62_179 ();
 sg13g2_decap_8 FILLER_62_186 ();
 sg13g2_decap_8 FILLER_62_193 ();
 sg13g2_decap_8 FILLER_62_200 ();
 sg13g2_decap_8 FILLER_62_207 ();
 sg13g2_decap_8 FILLER_62_214 ();
 sg13g2_decap_8 FILLER_62_221 ();
 sg13g2_decap_8 FILLER_62_228 ();
 sg13g2_decap_8 FILLER_62_235 ();
 sg13g2_decap_8 FILLER_62_242 ();
 sg13g2_decap_8 FILLER_62_249 ();
 sg13g2_decap_8 FILLER_62_256 ();
 sg13g2_decap_8 FILLER_62_263 ();
 sg13g2_decap_8 FILLER_62_270 ();
 sg13g2_decap_8 FILLER_62_277 ();
 sg13g2_decap_8 FILLER_62_284 ();
 sg13g2_decap_8 FILLER_62_291 ();
 sg13g2_decap_8 FILLER_62_302 ();
 sg13g2_decap_8 FILLER_62_309 ();
 sg13g2_decap_4 FILLER_62_316 ();
 sg13g2_fill_1 FILLER_62_320 ();
 sg13g2_decap_8 FILLER_62_330 ();
 sg13g2_decap_8 FILLER_62_337 ();
 sg13g2_decap_8 FILLER_62_344 ();
 sg13g2_decap_8 FILLER_62_351 ();
 sg13g2_decap_4 FILLER_62_358 ();
 sg13g2_fill_2 FILLER_62_362 ();
 sg13g2_decap_8 FILLER_62_368 ();
 sg13g2_decap_8 FILLER_62_375 ();
 sg13g2_decap_4 FILLER_62_382 ();
 sg13g2_decap_8 FILLER_62_394 ();
 sg13g2_decap_8 FILLER_62_401 ();
 sg13g2_decap_8 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_fill_1 FILLER_62_434 ();
 sg13g2_decap_8 FILLER_62_439 ();
 sg13g2_decap_8 FILLER_62_446 ();
 sg13g2_decap_8 FILLER_62_453 ();
 sg13g2_decap_8 FILLER_62_460 ();
 sg13g2_decap_8 FILLER_62_467 ();
 sg13g2_decap_4 FILLER_62_474 ();
 sg13g2_fill_1 FILLER_62_483 ();
 sg13g2_decap_8 FILLER_62_492 ();
 sg13g2_decap_4 FILLER_62_499 ();
 sg13g2_fill_2 FILLER_62_503 ();
 sg13g2_decap_8 FILLER_62_518 ();
 sg13g2_decap_8 FILLER_62_525 ();
 sg13g2_decap_8 FILLER_62_532 ();
 sg13g2_decap_8 FILLER_62_539 ();
 sg13g2_decap_8 FILLER_62_568 ();
 sg13g2_decap_8 FILLER_62_575 ();
 sg13g2_decap_8 FILLER_62_582 ();
 sg13g2_decap_8 FILLER_62_589 ();
 sg13g2_fill_2 FILLER_62_596 ();
 sg13g2_decap_8 FILLER_62_602 ();
 sg13g2_fill_2 FILLER_62_609 ();
 sg13g2_fill_1 FILLER_62_611 ();
 sg13g2_decap_8 FILLER_62_616 ();
 sg13g2_decap_8 FILLER_62_623 ();
 sg13g2_decap_8 FILLER_62_630 ();
 sg13g2_decap_4 FILLER_62_637 ();
 sg13g2_fill_2 FILLER_62_641 ();
 sg13g2_decap_8 FILLER_62_648 ();
 sg13g2_decap_8 FILLER_62_655 ();
 sg13g2_decap_8 FILLER_62_662 ();
 sg13g2_decap_8 FILLER_62_669 ();
 sg13g2_decap_8 FILLER_62_676 ();
 sg13g2_decap_8 FILLER_62_683 ();
 sg13g2_decap_8 FILLER_62_690 ();
 sg13g2_decap_8 FILLER_62_697 ();
 sg13g2_decap_8 FILLER_62_704 ();
 sg13g2_decap_8 FILLER_62_711 ();
 sg13g2_decap_8 FILLER_62_718 ();
 sg13g2_decap_8 FILLER_62_725 ();
 sg13g2_decap_8 FILLER_62_732 ();
 sg13g2_decap_8 FILLER_62_739 ();
 sg13g2_decap_8 FILLER_62_746 ();
 sg13g2_decap_8 FILLER_62_753 ();
 sg13g2_decap_8 FILLER_62_760 ();
 sg13g2_decap_8 FILLER_62_767 ();
 sg13g2_decap_8 FILLER_62_774 ();
 sg13g2_decap_8 FILLER_62_781 ();
 sg13g2_decap_8 FILLER_62_788 ();
 sg13g2_decap_8 FILLER_62_795 ();
 sg13g2_decap_8 FILLER_62_802 ();
 sg13g2_decap_8 FILLER_62_809 ();
 sg13g2_decap_8 FILLER_62_816 ();
 sg13g2_decap_8 FILLER_62_823 ();
 sg13g2_decap_8 FILLER_62_830 ();
 sg13g2_decap_8 FILLER_62_837 ();
 sg13g2_decap_8 FILLER_62_844 ();
 sg13g2_decap_8 FILLER_62_851 ();
 sg13g2_decap_8 FILLER_62_858 ();
 sg13g2_decap_8 FILLER_62_865 ();
 sg13g2_decap_4 FILLER_62_872 ();
 sg13g2_fill_2 FILLER_62_876 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_fill_1 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_40 ();
 sg13g2_fill_2 FILLER_63_47 ();
 sg13g2_fill_1 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_76 ();
 sg13g2_decap_4 FILLER_63_83 ();
 sg13g2_fill_2 FILLER_63_87 ();
 sg13g2_decap_4 FILLER_63_93 ();
 sg13g2_fill_2 FILLER_63_97 ();
 sg13g2_decap_8 FILLER_63_125 ();
 sg13g2_decap_8 FILLER_63_132 ();
 sg13g2_decap_8 FILLER_63_139 ();
 sg13g2_fill_1 FILLER_63_146 ();
 sg13g2_decap_8 FILLER_63_151 ();
 sg13g2_decap_8 FILLER_63_158 ();
 sg13g2_decap_8 FILLER_63_165 ();
 sg13g2_decap_8 FILLER_63_172 ();
 sg13g2_decap_8 FILLER_63_179 ();
 sg13g2_decap_8 FILLER_63_186 ();
 sg13g2_decap_8 FILLER_63_193 ();
 sg13g2_decap_8 FILLER_63_200 ();
 sg13g2_decap_8 FILLER_63_207 ();
 sg13g2_decap_8 FILLER_63_214 ();
 sg13g2_decap_8 FILLER_63_221 ();
 sg13g2_decap_8 FILLER_63_228 ();
 sg13g2_decap_8 FILLER_63_235 ();
 sg13g2_decap_8 FILLER_63_242 ();
 sg13g2_decap_8 FILLER_63_249 ();
 sg13g2_decap_8 FILLER_63_256 ();
 sg13g2_decap_8 FILLER_63_263 ();
 sg13g2_decap_8 FILLER_63_270 ();
 sg13g2_decap_8 FILLER_63_277 ();
 sg13g2_decap_8 FILLER_63_284 ();
 sg13g2_decap_8 FILLER_63_291 ();
 sg13g2_decap_8 FILLER_63_298 ();
 sg13g2_decap_8 FILLER_63_305 ();
 sg13g2_decap_8 FILLER_63_312 ();
 sg13g2_decap_8 FILLER_63_319 ();
 sg13g2_decap_8 FILLER_63_326 ();
 sg13g2_fill_2 FILLER_63_333 ();
 sg13g2_fill_1 FILLER_63_335 ();
 sg13g2_decap_8 FILLER_63_344 ();
 sg13g2_decap_8 FILLER_63_351 ();
 sg13g2_decap_8 FILLER_63_358 ();
 sg13g2_fill_1 FILLER_63_365 ();
 sg13g2_decap_8 FILLER_63_370 ();
 sg13g2_decap_8 FILLER_63_377 ();
 sg13g2_decap_4 FILLER_63_384 ();
 sg13g2_fill_1 FILLER_63_388 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_decap_4 FILLER_63_427 ();
 sg13g2_fill_2 FILLER_63_431 ();
 sg13g2_decap_8 FILLER_63_441 ();
 sg13g2_decap_8 FILLER_63_448 ();
 sg13g2_decap_8 FILLER_63_455 ();
 sg13g2_decap_8 FILLER_63_462 ();
 sg13g2_decap_8 FILLER_63_469 ();
 sg13g2_fill_2 FILLER_63_476 ();
 sg13g2_fill_1 FILLER_63_478 ();
 sg13g2_decap_4 FILLER_63_483 ();
 sg13g2_decap_8 FILLER_63_490 ();
 sg13g2_decap_8 FILLER_63_497 ();
 sg13g2_decap_8 FILLER_63_504 ();
 sg13g2_decap_8 FILLER_63_511 ();
 sg13g2_decap_8 FILLER_63_518 ();
 sg13g2_decap_8 FILLER_63_525 ();
 sg13g2_decap_8 FILLER_63_532 ();
 sg13g2_fill_2 FILLER_63_539 ();
 sg13g2_decap_8 FILLER_63_545 ();
 sg13g2_decap_8 FILLER_63_552 ();
 sg13g2_decap_8 FILLER_63_559 ();
 sg13g2_decap_8 FILLER_63_566 ();
 sg13g2_decap_8 FILLER_63_573 ();
 sg13g2_decap_8 FILLER_63_580 ();
 sg13g2_decap_8 FILLER_63_587 ();
 sg13g2_decap_8 FILLER_63_625 ();
 sg13g2_decap_8 FILLER_63_632 ();
 sg13g2_decap_8 FILLER_63_639 ();
 sg13g2_fill_1 FILLER_63_646 ();
 sg13g2_decap_8 FILLER_63_651 ();
 sg13g2_decap_8 FILLER_63_658 ();
 sg13g2_decap_8 FILLER_63_665 ();
 sg13g2_decap_8 FILLER_63_672 ();
 sg13g2_decap_8 FILLER_63_679 ();
 sg13g2_decap_8 FILLER_63_686 ();
 sg13g2_decap_8 FILLER_63_693 ();
 sg13g2_decap_8 FILLER_63_700 ();
 sg13g2_decap_8 FILLER_63_707 ();
 sg13g2_decap_8 FILLER_63_714 ();
 sg13g2_decap_8 FILLER_63_721 ();
 sg13g2_decap_8 FILLER_63_728 ();
 sg13g2_decap_8 FILLER_63_735 ();
 sg13g2_decap_8 FILLER_63_742 ();
 sg13g2_decap_8 FILLER_63_749 ();
 sg13g2_decap_8 FILLER_63_756 ();
 sg13g2_decap_8 FILLER_63_763 ();
 sg13g2_decap_8 FILLER_63_770 ();
 sg13g2_decap_8 FILLER_63_777 ();
 sg13g2_decap_8 FILLER_63_784 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_decap_8 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_decap_8 FILLER_63_812 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_decap_8 FILLER_63_840 ();
 sg13g2_decap_8 FILLER_63_847 ();
 sg13g2_decap_8 FILLER_63_854 ();
 sg13g2_decap_8 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_63_868 ();
 sg13g2_fill_2 FILLER_63_875 ();
 sg13g2_fill_1 FILLER_63_877 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_fill_2 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_60 ();
 sg13g2_decap_8 FILLER_64_67 ();
 sg13g2_decap_8 FILLER_64_74 ();
 sg13g2_decap_8 FILLER_64_81 ();
 sg13g2_decap_8 FILLER_64_88 ();
 sg13g2_decap_8 FILLER_64_95 ();
 sg13g2_decap_8 FILLER_64_102 ();
 sg13g2_decap_8 FILLER_64_109 ();
 sg13g2_decap_8 FILLER_64_116 ();
 sg13g2_decap_8 FILLER_64_123 ();
 sg13g2_decap_8 FILLER_64_130 ();
 sg13g2_fill_2 FILLER_64_137 ();
 sg13g2_decap_4 FILLER_64_165 ();
 sg13g2_fill_1 FILLER_64_169 ();
 sg13g2_decap_8 FILLER_64_174 ();
 sg13g2_decap_8 FILLER_64_181 ();
 sg13g2_decap_8 FILLER_64_188 ();
 sg13g2_decap_8 FILLER_64_195 ();
 sg13g2_decap_8 FILLER_64_202 ();
 sg13g2_decap_8 FILLER_64_209 ();
 sg13g2_decap_8 FILLER_64_216 ();
 sg13g2_decap_8 FILLER_64_223 ();
 sg13g2_decap_8 FILLER_64_230 ();
 sg13g2_decap_8 FILLER_64_237 ();
 sg13g2_decap_8 FILLER_64_244 ();
 sg13g2_decap_8 FILLER_64_251 ();
 sg13g2_decap_8 FILLER_64_258 ();
 sg13g2_decap_8 FILLER_64_265 ();
 sg13g2_decap_8 FILLER_64_272 ();
 sg13g2_decap_8 FILLER_64_279 ();
 sg13g2_decap_8 FILLER_64_286 ();
 sg13g2_decap_8 FILLER_64_293 ();
 sg13g2_decap_8 FILLER_64_300 ();
 sg13g2_decap_8 FILLER_64_307 ();
 sg13g2_decap_8 FILLER_64_314 ();
 sg13g2_decap_8 FILLER_64_321 ();
 sg13g2_decap_8 FILLER_64_328 ();
 sg13g2_decap_8 FILLER_64_347 ();
 sg13g2_decap_8 FILLER_64_354 ();
 sg13g2_decap_8 FILLER_64_361 ();
 sg13g2_decap_8 FILLER_64_368 ();
 sg13g2_decap_8 FILLER_64_375 ();
 sg13g2_decap_8 FILLER_64_382 ();
 sg13g2_decap_8 FILLER_64_389 ();
 sg13g2_decap_8 FILLER_64_396 ();
 sg13g2_decap_8 FILLER_64_409 ();
 sg13g2_fill_2 FILLER_64_416 ();
 sg13g2_fill_1 FILLER_64_418 ();
 sg13g2_decap_4 FILLER_64_425 ();
 sg13g2_decap_8 FILLER_64_440 ();
 sg13g2_decap_4 FILLER_64_447 ();
 sg13g2_decap_4 FILLER_64_459 ();
 sg13g2_fill_1 FILLER_64_463 ();
 sg13g2_decap_8 FILLER_64_468 ();
 sg13g2_decap_8 FILLER_64_475 ();
 sg13g2_decap_8 FILLER_64_482 ();
 sg13g2_decap_8 FILLER_64_489 ();
 sg13g2_decap_8 FILLER_64_496 ();
 sg13g2_fill_2 FILLER_64_503 ();
 sg13g2_fill_1 FILLER_64_505 ();
 sg13g2_decap_8 FILLER_64_510 ();
 sg13g2_decap_8 FILLER_64_517 ();
 sg13g2_decap_8 FILLER_64_524 ();
 sg13g2_decap_8 FILLER_64_531 ();
 sg13g2_decap_8 FILLER_64_538 ();
 sg13g2_decap_4 FILLER_64_545 ();
 sg13g2_fill_2 FILLER_64_549 ();
 sg13g2_decap_8 FILLER_64_556 ();
 sg13g2_decap_8 FILLER_64_563 ();
 sg13g2_decap_8 FILLER_64_570 ();
 sg13g2_decap_8 FILLER_64_577 ();
 sg13g2_decap_8 FILLER_64_584 ();
 sg13g2_decap_8 FILLER_64_591 ();
 sg13g2_decap_8 FILLER_64_598 ();
 sg13g2_decap_8 FILLER_64_605 ();
 sg13g2_decap_8 FILLER_64_612 ();
 sg13g2_decap_8 FILLER_64_619 ();
 sg13g2_decap_8 FILLER_64_626 ();
 sg13g2_decap_8 FILLER_64_633 ();
 sg13g2_decap_8 FILLER_64_640 ();
 sg13g2_decap_8 FILLER_64_647 ();
 sg13g2_decap_8 FILLER_64_654 ();
 sg13g2_decap_8 FILLER_64_661 ();
 sg13g2_decap_8 FILLER_64_668 ();
 sg13g2_decap_8 FILLER_64_675 ();
 sg13g2_decap_8 FILLER_64_682 ();
 sg13g2_decap_8 FILLER_64_689 ();
 sg13g2_decap_8 FILLER_64_696 ();
 sg13g2_decap_8 FILLER_64_703 ();
 sg13g2_decap_8 FILLER_64_710 ();
 sg13g2_decap_8 FILLER_64_717 ();
 sg13g2_decap_8 FILLER_64_724 ();
 sg13g2_decap_8 FILLER_64_731 ();
 sg13g2_decap_8 FILLER_64_738 ();
 sg13g2_decap_8 FILLER_64_745 ();
 sg13g2_decap_8 FILLER_64_752 ();
 sg13g2_decap_8 FILLER_64_759 ();
 sg13g2_decap_8 FILLER_64_766 ();
 sg13g2_decap_8 FILLER_64_773 ();
 sg13g2_decap_8 FILLER_64_780 ();
 sg13g2_decap_8 FILLER_64_787 ();
 sg13g2_decap_8 FILLER_64_794 ();
 sg13g2_decap_8 FILLER_64_801 ();
 sg13g2_decap_8 FILLER_64_808 ();
 sg13g2_decap_8 FILLER_64_815 ();
 sg13g2_decap_8 FILLER_64_822 ();
 sg13g2_decap_8 FILLER_64_829 ();
 sg13g2_decap_8 FILLER_64_836 ();
 sg13g2_decap_8 FILLER_64_843 ();
 sg13g2_decap_8 FILLER_64_850 ();
 sg13g2_decap_8 FILLER_64_857 ();
 sg13g2_decap_8 FILLER_64_864 ();
 sg13g2_decap_8 FILLER_64_871 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_4 FILLER_65_42 ();
 sg13g2_fill_2 FILLER_65_46 ();
 sg13g2_decap_8 FILLER_65_74 ();
 sg13g2_decap_8 FILLER_65_81 ();
 sg13g2_decap_4 FILLER_65_88 ();
 sg13g2_fill_1 FILLER_65_92 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_4 FILLER_65_126 ();
 sg13g2_fill_2 FILLER_65_135 ();
 sg13g2_fill_1 FILLER_65_137 ();
 sg13g2_decap_8 FILLER_65_144 ();
 sg13g2_decap_8 FILLER_65_151 ();
 sg13g2_decap_4 FILLER_65_158 ();
 sg13g2_decap_8 FILLER_65_188 ();
 sg13g2_decap_8 FILLER_65_199 ();
 sg13g2_decap_8 FILLER_65_206 ();
 sg13g2_decap_8 FILLER_65_213 ();
 sg13g2_fill_1 FILLER_65_220 ();
 sg13g2_decap_8 FILLER_65_225 ();
 sg13g2_decap_8 FILLER_65_232 ();
 sg13g2_decap_8 FILLER_65_239 ();
 sg13g2_decap_8 FILLER_65_246 ();
 sg13g2_decap_8 FILLER_65_253 ();
 sg13g2_decap_8 FILLER_65_260 ();
 sg13g2_decap_8 FILLER_65_267 ();
 sg13g2_fill_2 FILLER_65_274 ();
 sg13g2_fill_1 FILLER_65_276 ();
 sg13g2_decap_8 FILLER_65_281 ();
 sg13g2_fill_2 FILLER_65_288 ();
 sg13g2_fill_1 FILLER_65_290 ();
 sg13g2_decap_8 FILLER_65_296 ();
 sg13g2_decap_8 FILLER_65_303 ();
 sg13g2_decap_8 FILLER_65_310 ();
 sg13g2_decap_8 FILLER_65_317 ();
 sg13g2_decap_4 FILLER_65_324 ();
 sg13g2_fill_1 FILLER_65_334 ();
 sg13g2_fill_2 FILLER_65_342 ();
 sg13g2_decap_8 FILLER_65_348 ();
 sg13g2_decap_8 FILLER_65_355 ();
 sg13g2_decap_8 FILLER_65_362 ();
 sg13g2_decap_8 FILLER_65_369 ();
 sg13g2_decap_4 FILLER_65_376 ();
 sg13g2_fill_1 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_65_409 ();
 sg13g2_fill_2 FILLER_65_416 ();
 sg13g2_fill_1 FILLER_65_418 ();
 sg13g2_decap_8 FILLER_65_423 ();
 sg13g2_fill_1 FILLER_65_430 ();
 sg13g2_decap_8 FILLER_65_436 ();
 sg13g2_decap_8 FILLER_65_443 ();
 sg13g2_fill_2 FILLER_65_459 ();
 sg13g2_fill_2 FILLER_65_466 ();
 sg13g2_decap_4 FILLER_65_494 ();
 sg13g2_fill_1 FILLER_65_498 ();
 sg13g2_decap_8 FILLER_65_551 ();
 sg13g2_decap_8 FILLER_65_558 ();
 sg13g2_decap_8 FILLER_65_565 ();
 sg13g2_decap_4 FILLER_65_572 ();
 sg13g2_fill_1 FILLER_65_576 ();
 sg13g2_decap_8 FILLER_65_590 ();
 sg13g2_fill_1 FILLER_65_597 ();
 sg13g2_decap_8 FILLER_65_628 ();
 sg13g2_decap_8 FILLER_65_635 ();
 sg13g2_decap_8 FILLER_65_642 ();
 sg13g2_decap_8 FILLER_65_649 ();
 sg13g2_decap_8 FILLER_65_656 ();
 sg13g2_decap_8 FILLER_65_663 ();
 sg13g2_decap_8 FILLER_65_670 ();
 sg13g2_fill_2 FILLER_65_677 ();
 sg13g2_fill_2 FILLER_65_684 ();
 sg13g2_fill_2 FILLER_65_690 ();
 sg13g2_fill_1 FILLER_65_692 ();
 sg13g2_decap_8 FILLER_65_705 ();
 sg13g2_decap_8 FILLER_65_712 ();
 sg13g2_decap_8 FILLER_65_719 ();
 sg13g2_decap_8 FILLER_65_726 ();
 sg13g2_decap_8 FILLER_65_733 ();
 sg13g2_decap_8 FILLER_65_740 ();
 sg13g2_decap_8 FILLER_65_747 ();
 sg13g2_decap_8 FILLER_65_754 ();
 sg13g2_fill_1 FILLER_65_761 ();
 sg13g2_decap_8 FILLER_65_775 ();
 sg13g2_decap_8 FILLER_65_782 ();
 sg13g2_decap_8 FILLER_65_789 ();
 sg13g2_decap_8 FILLER_65_796 ();
 sg13g2_decap_8 FILLER_65_803 ();
 sg13g2_decap_8 FILLER_65_810 ();
 sg13g2_decap_8 FILLER_65_817 ();
 sg13g2_decap_8 FILLER_65_824 ();
 sg13g2_decap_8 FILLER_65_831 ();
 sg13g2_decap_8 FILLER_65_838 ();
 sg13g2_decap_8 FILLER_65_845 ();
 sg13g2_decap_8 FILLER_65_852 ();
 sg13g2_decap_8 FILLER_65_859 ();
 sg13g2_decap_8 FILLER_65_866 ();
 sg13g2_decap_4 FILLER_65_873 ();
 sg13g2_fill_1 FILLER_65_877 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_4 FILLER_66_35 ();
 sg13g2_fill_2 FILLER_66_48 ();
 sg13g2_decap_8 FILLER_66_59 ();
 sg13g2_decap_8 FILLER_66_66 ();
 sg13g2_decap_8 FILLER_66_73 ();
 sg13g2_decap_8 FILLER_66_80 ();
 sg13g2_decap_8 FILLER_66_87 ();
 sg13g2_decap_8 FILLER_66_94 ();
 sg13g2_fill_1 FILLER_66_101 ();
 sg13g2_decap_8 FILLER_66_106 ();
 sg13g2_fill_1 FILLER_66_113 ();
 sg13g2_fill_2 FILLER_66_146 ();
 sg13g2_decap_8 FILLER_66_163 ();
 sg13g2_decap_8 FILLER_66_170 ();
 sg13g2_decap_8 FILLER_66_177 ();
 sg13g2_decap_4 FILLER_66_184 ();
 sg13g2_decap_8 FILLER_66_240 ();
 sg13g2_decap_8 FILLER_66_247 ();
 sg13g2_decap_8 FILLER_66_254 ();
 sg13g2_decap_8 FILLER_66_261 ();
 sg13g2_fill_2 FILLER_66_268 ();
 sg13g2_decap_8 FILLER_66_296 ();
 sg13g2_decap_8 FILLER_66_303 ();
 sg13g2_decap_8 FILLER_66_310 ();
 sg13g2_decap_8 FILLER_66_317 ();
 sg13g2_decap_8 FILLER_66_324 ();
 sg13g2_fill_2 FILLER_66_331 ();
 sg13g2_fill_1 FILLER_66_333 ();
 sg13g2_decap_4 FILLER_66_339 ();
 sg13g2_fill_2 FILLER_66_343 ();
 sg13g2_decap_8 FILLER_66_351 ();
 sg13g2_decap_8 FILLER_66_358 ();
 sg13g2_decap_8 FILLER_66_365 ();
 sg13g2_fill_1 FILLER_66_372 ();
 sg13g2_decap_4 FILLER_66_382 ();
 sg13g2_fill_2 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_393 ();
 sg13g2_decap_8 FILLER_66_400 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_66_415 ();
 sg13g2_fill_1 FILLER_66_430 ();
 sg13g2_fill_1 FILLER_66_435 ();
 sg13g2_fill_2 FILLER_66_441 ();
 sg13g2_decap_8 FILLER_66_447 ();
 sg13g2_decap_8 FILLER_66_454 ();
 sg13g2_decap_8 FILLER_66_461 ();
 sg13g2_decap_4 FILLER_66_468 ();
 sg13g2_fill_2 FILLER_66_472 ();
 sg13g2_decap_8 FILLER_66_478 ();
 sg13g2_decap_8 FILLER_66_485 ();
 sg13g2_decap_8 FILLER_66_492 ();
 sg13g2_decap_8 FILLER_66_499 ();
 sg13g2_decap_8 FILLER_66_506 ();
 sg13g2_decap_8 FILLER_66_513 ();
 sg13g2_decap_8 FILLER_66_520 ();
 sg13g2_decap_4 FILLER_66_527 ();
 sg13g2_fill_1 FILLER_66_531 ();
 sg13g2_decap_8 FILLER_66_536 ();
 sg13g2_decap_8 FILLER_66_543 ();
 sg13g2_decap_8 FILLER_66_550 ();
 sg13g2_decap_8 FILLER_66_557 ();
 sg13g2_decap_8 FILLER_66_564 ();
 sg13g2_decap_8 FILLER_66_571 ();
 sg13g2_decap_8 FILLER_66_578 ();
 sg13g2_decap_8 FILLER_66_585 ();
 sg13g2_decap_8 FILLER_66_592 ();
 sg13g2_fill_1 FILLER_66_599 ();
 sg13g2_decap_8 FILLER_66_630 ();
 sg13g2_decap_8 FILLER_66_637 ();
 sg13g2_fill_2 FILLER_66_644 ();
 sg13g2_fill_1 FILLER_66_646 ();
 sg13g2_fill_2 FILLER_66_673 ();
 sg13g2_fill_1 FILLER_66_675 ();
 sg13g2_fill_2 FILLER_66_702 ();
 sg13g2_fill_1 FILLER_66_704 ();
 sg13g2_fill_2 FILLER_66_731 ();
 sg13g2_decap_8 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_744 ();
 sg13g2_decap_8 FILLER_66_751 ();
 sg13g2_fill_1 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_799 ();
 sg13g2_decap_8 FILLER_66_806 ();
 sg13g2_decap_8 FILLER_66_813 ();
 sg13g2_decap_8 FILLER_66_820 ();
 sg13g2_decap_8 FILLER_66_827 ();
 sg13g2_decap_8 FILLER_66_834 ();
 sg13g2_decap_8 FILLER_66_841 ();
 sg13g2_decap_8 FILLER_66_848 ();
 sg13g2_decap_8 FILLER_66_855 ();
 sg13g2_decap_8 FILLER_66_862 ();
 sg13g2_decap_8 FILLER_66_869 ();
 sg13g2_fill_2 FILLER_66_876 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_fill_2 FILLER_67_35 ();
 sg13g2_fill_1 FILLER_67_37 ();
 sg13g2_fill_1 FILLER_67_56 ();
 sg13g2_decap_4 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_92 ();
 sg13g2_decap_4 FILLER_67_102 ();
 sg13g2_fill_2 FILLER_67_106 ();
 sg13g2_decap_4 FILLER_67_120 ();
 sg13g2_fill_1 FILLER_67_124 ();
 sg13g2_fill_1 FILLER_67_130 ();
 sg13g2_fill_1 FILLER_67_146 ();
 sg13g2_decap_8 FILLER_67_151 ();
 sg13g2_decap_8 FILLER_67_158 ();
 sg13g2_decap_8 FILLER_67_165 ();
 sg13g2_decap_8 FILLER_67_172 ();
 sg13g2_decap_8 FILLER_67_179 ();
 sg13g2_decap_8 FILLER_67_186 ();
 sg13g2_decap_8 FILLER_67_193 ();
 sg13g2_decap_8 FILLER_67_200 ();
 sg13g2_decap_8 FILLER_67_207 ();
 sg13g2_decap_8 FILLER_67_214 ();
 sg13g2_decap_8 FILLER_67_221 ();
 sg13g2_decap_8 FILLER_67_228 ();
 sg13g2_fill_2 FILLER_67_235 ();
 sg13g2_fill_2 FILLER_67_241 ();
 sg13g2_fill_1 FILLER_67_243 ();
 sg13g2_decap_8 FILLER_67_255 ();
 sg13g2_fill_2 FILLER_67_262 ();
 sg13g2_fill_1 FILLER_67_264 ();
 sg13g2_decap_8 FILLER_67_295 ();
 sg13g2_decap_8 FILLER_67_302 ();
 sg13g2_decap_8 FILLER_67_309 ();
 sg13g2_decap_8 FILLER_67_316 ();
 sg13g2_decap_8 FILLER_67_323 ();
 sg13g2_decap_8 FILLER_67_330 ();
 sg13g2_decap_8 FILLER_67_337 ();
 sg13g2_decap_8 FILLER_67_349 ();
 sg13g2_decap_8 FILLER_67_382 ();
 sg13g2_fill_2 FILLER_67_389 ();
 sg13g2_fill_2 FILLER_67_396 ();
 sg13g2_fill_1 FILLER_67_398 ();
 sg13g2_decap_8 FILLER_67_404 ();
 sg13g2_fill_2 FILLER_67_411 ();
 sg13g2_fill_1 FILLER_67_413 ();
 sg13g2_fill_2 FILLER_67_419 ();
 sg13g2_fill_1 FILLER_67_421 ();
 sg13g2_decap_8 FILLER_67_432 ();
 sg13g2_decap_8 FILLER_67_439 ();
 sg13g2_decap_8 FILLER_67_446 ();
 sg13g2_decap_8 FILLER_67_453 ();
 sg13g2_decap_8 FILLER_67_460 ();
 sg13g2_decap_8 FILLER_67_467 ();
 sg13g2_fill_1 FILLER_67_474 ();
 sg13g2_decap_8 FILLER_67_479 ();
 sg13g2_decap_8 FILLER_67_486 ();
 sg13g2_decap_8 FILLER_67_493 ();
 sg13g2_decap_8 FILLER_67_500 ();
 sg13g2_decap_8 FILLER_67_507 ();
 sg13g2_decap_8 FILLER_67_525 ();
 sg13g2_decap_8 FILLER_67_532 ();
 sg13g2_decap_8 FILLER_67_539 ();
 sg13g2_decap_8 FILLER_67_546 ();
 sg13g2_decap_8 FILLER_67_553 ();
 sg13g2_decap_8 FILLER_67_560 ();
 sg13g2_decap_8 FILLER_67_567 ();
 sg13g2_decap_8 FILLER_67_574 ();
 sg13g2_decap_8 FILLER_67_581 ();
 sg13g2_decap_8 FILLER_67_588 ();
 sg13g2_decap_8 FILLER_67_595 ();
 sg13g2_decap_8 FILLER_67_602 ();
 sg13g2_decap_8 FILLER_67_609 ();
 sg13g2_decap_8 FILLER_67_616 ();
 sg13g2_decap_8 FILLER_67_623 ();
 sg13g2_decap_8 FILLER_67_630 ();
 sg13g2_decap_8 FILLER_67_637 ();
 sg13g2_decap_8 FILLER_67_644 ();
 sg13g2_fill_2 FILLER_67_651 ();
 sg13g2_fill_1 FILLER_67_657 ();
 sg13g2_decap_8 FILLER_67_663 ();
 sg13g2_decap_8 FILLER_67_670 ();
 sg13g2_decap_4 FILLER_67_677 ();
 sg13g2_fill_2 FILLER_67_681 ();
 sg13g2_decap_8 FILLER_67_691 ();
 sg13g2_fill_2 FILLER_67_698 ();
 sg13g2_fill_1 FILLER_67_700 ();
 sg13g2_decap_4 FILLER_67_706 ();
 sg13g2_fill_2 FILLER_67_710 ();
 sg13g2_decap_4 FILLER_67_716 ();
 sg13g2_fill_1 FILLER_67_720 ();
 sg13g2_fill_1 FILLER_67_725 ();
 sg13g2_decap_8 FILLER_67_760 ();
 sg13g2_decap_8 FILLER_67_767 ();
 sg13g2_decap_4 FILLER_67_774 ();
 sg13g2_fill_1 FILLER_67_778 ();
 sg13g2_decap_8 FILLER_67_783 ();
 sg13g2_decap_8 FILLER_67_790 ();
 sg13g2_decap_8 FILLER_67_797 ();
 sg13g2_decap_8 FILLER_67_804 ();
 sg13g2_decap_8 FILLER_67_811 ();
 sg13g2_decap_8 FILLER_67_818 ();
 sg13g2_decap_8 FILLER_67_825 ();
 sg13g2_decap_8 FILLER_67_832 ();
 sg13g2_decap_8 FILLER_67_839 ();
 sg13g2_decap_8 FILLER_67_846 ();
 sg13g2_decap_8 FILLER_67_853 ();
 sg13g2_decap_8 FILLER_67_860 ();
 sg13g2_decap_8 FILLER_67_867 ();
 sg13g2_decap_4 FILLER_67_874 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_4 FILLER_68_28 ();
 sg13g2_fill_2 FILLER_68_32 ();
 sg13g2_fill_1 FILLER_68_41 ();
 sg13g2_fill_1 FILLER_68_55 ();
 sg13g2_decap_8 FILLER_68_80 ();
 sg13g2_decap_4 FILLER_68_87 ();
 sg13g2_fill_1 FILLER_68_94 ();
 sg13g2_fill_1 FILLER_68_111 ();
 sg13g2_decap_8 FILLER_68_159 ();
 sg13g2_decap_8 FILLER_68_166 ();
 sg13g2_decap_8 FILLER_68_173 ();
 sg13g2_decap_8 FILLER_68_180 ();
 sg13g2_decap_4 FILLER_68_187 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_decap_4 FILLER_68_224 ();
 sg13g2_fill_2 FILLER_68_228 ();
 sg13g2_decap_8 FILLER_68_256 ();
 sg13g2_decap_8 FILLER_68_263 ();
 sg13g2_decap_8 FILLER_68_278 ();
 sg13g2_decap_8 FILLER_68_285 ();
 sg13g2_decap_8 FILLER_68_292 ();
 sg13g2_decap_8 FILLER_68_299 ();
 sg13g2_decap_8 FILLER_68_306 ();
 sg13g2_fill_1 FILLER_68_313 ();
 sg13g2_decap_8 FILLER_68_318 ();
 sg13g2_fill_2 FILLER_68_325 ();
 sg13g2_decap_8 FILLER_68_337 ();
 sg13g2_decap_8 FILLER_68_344 ();
 sg13g2_decap_8 FILLER_68_351 ();
 sg13g2_decap_4 FILLER_68_358 ();
 sg13g2_fill_1 FILLER_68_362 ();
 sg13g2_decap_8 FILLER_68_367 ();
 sg13g2_fill_2 FILLER_68_379 ();
 sg13g2_fill_1 FILLER_68_381 ();
 sg13g2_decap_8 FILLER_68_386 ();
 sg13g2_decap_4 FILLER_68_393 ();
 sg13g2_fill_2 FILLER_68_397 ();
 sg13g2_decap_8 FILLER_68_403 ();
 sg13g2_decap_8 FILLER_68_410 ();
 sg13g2_decap_8 FILLER_68_417 ();
 sg13g2_fill_2 FILLER_68_424 ();
 sg13g2_decap_8 FILLER_68_430 ();
 sg13g2_fill_1 FILLER_68_437 ();
 sg13g2_decap_8 FILLER_68_443 ();
 sg13g2_decap_4 FILLER_68_450 ();
 sg13g2_fill_2 FILLER_68_454 ();
 sg13g2_decap_8 FILLER_68_487 ();
 sg13g2_decap_8 FILLER_68_494 ();
 sg13g2_decap_8 FILLER_68_501 ();
 sg13g2_decap_8 FILLER_68_508 ();
 sg13g2_decap_8 FILLER_68_515 ();
 sg13g2_decap_8 FILLER_68_522 ();
 sg13g2_decap_8 FILLER_68_529 ();
 sg13g2_decap_8 FILLER_68_536 ();
 sg13g2_decap_4 FILLER_68_543 ();
 sg13g2_fill_2 FILLER_68_547 ();
 sg13g2_decap_8 FILLER_68_553 ();
 sg13g2_decap_8 FILLER_68_560 ();
 sg13g2_decap_8 FILLER_68_567 ();
 sg13g2_fill_2 FILLER_68_574 ();
 sg13g2_fill_1 FILLER_68_576 ();
 sg13g2_decap_4 FILLER_68_581 ();
 sg13g2_fill_1 FILLER_68_585 ();
 sg13g2_decap_8 FILLER_68_590 ();
 sg13g2_decap_8 FILLER_68_597 ();
 sg13g2_decap_8 FILLER_68_604 ();
 sg13g2_decap_8 FILLER_68_611 ();
 sg13g2_decap_8 FILLER_68_618 ();
 sg13g2_decap_8 FILLER_68_625 ();
 sg13g2_decap_8 FILLER_68_632 ();
 sg13g2_decap_8 FILLER_68_639 ();
 sg13g2_decap_8 FILLER_68_646 ();
 sg13g2_decap_8 FILLER_68_653 ();
 sg13g2_decap_8 FILLER_68_660 ();
 sg13g2_decap_8 FILLER_68_667 ();
 sg13g2_decap_8 FILLER_68_674 ();
 sg13g2_decap_8 FILLER_68_681 ();
 sg13g2_decap_8 FILLER_68_688 ();
 sg13g2_decap_8 FILLER_68_695 ();
 sg13g2_decap_8 FILLER_68_702 ();
 sg13g2_decap_8 FILLER_68_709 ();
 sg13g2_decap_8 FILLER_68_716 ();
 sg13g2_fill_2 FILLER_68_723 ();
 sg13g2_decap_8 FILLER_68_733 ();
 sg13g2_decap_8 FILLER_68_740 ();
 sg13g2_decap_8 FILLER_68_747 ();
 sg13g2_decap_8 FILLER_68_754 ();
 sg13g2_decap_8 FILLER_68_761 ();
 sg13g2_decap_8 FILLER_68_768 ();
 sg13g2_decap_8 FILLER_68_775 ();
 sg13g2_decap_8 FILLER_68_782 ();
 sg13g2_decap_8 FILLER_68_789 ();
 sg13g2_decap_8 FILLER_68_796 ();
 sg13g2_decap_8 FILLER_68_803 ();
 sg13g2_decap_8 FILLER_68_810 ();
 sg13g2_decap_8 FILLER_68_817 ();
 sg13g2_decap_8 FILLER_68_824 ();
 sg13g2_decap_8 FILLER_68_831 ();
 sg13g2_decap_8 FILLER_68_838 ();
 sg13g2_decap_8 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_852 ();
 sg13g2_decap_8 FILLER_68_859 ();
 sg13g2_decap_8 FILLER_68_866 ();
 sg13g2_decap_4 FILLER_68_873 ();
 sg13g2_fill_1 FILLER_68_877 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_4 FILLER_69_28 ();
 sg13g2_fill_2 FILLER_69_59 ();
 sg13g2_decap_8 FILLER_69_66 ();
 sg13g2_decap_4 FILLER_69_73 ();
 sg13g2_decap_4 FILLER_69_82 ();
 sg13g2_decap_4 FILLER_69_96 ();
 sg13g2_decap_4 FILLER_69_108 ();
 sg13g2_fill_2 FILLER_69_116 ();
 sg13g2_fill_1 FILLER_69_123 ();
 sg13g2_decap_4 FILLER_69_128 ();
 sg13g2_fill_2 FILLER_69_132 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_168 ();
 sg13g2_decap_8 FILLER_69_175 ();
 sg13g2_decap_8 FILLER_69_182 ();
 sg13g2_decap_8 FILLER_69_189 ();
 sg13g2_decap_4 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_204 ();
 sg13g2_decap_8 FILLER_69_211 ();
 sg13g2_decap_8 FILLER_69_218 ();
 sg13g2_decap_8 FILLER_69_225 ();
 sg13g2_fill_1 FILLER_69_232 ();
 sg13g2_decap_8 FILLER_69_259 ();
 sg13g2_decap_8 FILLER_69_266 ();
 sg13g2_decap_8 FILLER_69_273 ();
 sg13g2_decap_8 FILLER_69_280 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_8 FILLER_69_294 ();
 sg13g2_decap_4 FILLER_69_301 ();
 sg13g2_fill_2 FILLER_69_305 ();
 sg13g2_fill_2 FILLER_69_338 ();
 sg13g2_fill_1 FILLER_69_340 ();
 sg13g2_decap_8 FILLER_69_345 ();
 sg13g2_fill_1 FILLER_69_352 ();
 sg13g2_decap_8 FILLER_69_357 ();
 sg13g2_fill_2 FILLER_69_364 ();
 sg13g2_fill_1 FILLER_69_366 ();
 sg13g2_fill_2 FILLER_69_381 ();
 sg13g2_decap_4 FILLER_69_388 ();
 sg13g2_decap_4 FILLER_69_396 ();
 sg13g2_fill_2 FILLER_69_400 ();
 sg13g2_decap_8 FILLER_69_406 ();
 sg13g2_decap_8 FILLER_69_413 ();
 sg13g2_decap_8 FILLER_69_420 ();
 sg13g2_decap_4 FILLER_69_427 ();
 sg13g2_fill_1 FILLER_69_431 ();
 sg13g2_decap_4 FILLER_69_458 ();
 sg13g2_fill_1 FILLER_69_462 ();
 sg13g2_decap_8 FILLER_69_467 ();
 sg13g2_decap_8 FILLER_69_474 ();
 sg13g2_decap_8 FILLER_69_481 ();
 sg13g2_decap_8 FILLER_69_488 ();
 sg13g2_decap_8 FILLER_69_495 ();
 sg13g2_decap_8 FILLER_69_502 ();
 sg13g2_decap_8 FILLER_69_509 ();
 sg13g2_decap_8 FILLER_69_516 ();
 sg13g2_decap_8 FILLER_69_523 ();
 sg13g2_decap_8 FILLER_69_530 ();
 sg13g2_decap_8 FILLER_69_537 ();
 sg13g2_decap_8 FILLER_69_544 ();
 sg13g2_decap_8 FILLER_69_603 ();
 sg13g2_decap_4 FILLER_69_610 ();
 sg13g2_fill_1 FILLER_69_614 ();
 sg13g2_decap_8 FILLER_69_619 ();
 sg13g2_decap_8 FILLER_69_626 ();
 sg13g2_decap_8 FILLER_69_633 ();
 sg13g2_decap_8 FILLER_69_640 ();
 sg13g2_decap_8 FILLER_69_647 ();
 sg13g2_decap_8 FILLER_69_654 ();
 sg13g2_decap_8 FILLER_69_661 ();
 sg13g2_decap_8 FILLER_69_668 ();
 sg13g2_decap_8 FILLER_69_675 ();
 sg13g2_decap_8 FILLER_69_682 ();
 sg13g2_decap_8 FILLER_69_689 ();
 sg13g2_decap_8 FILLER_69_696 ();
 sg13g2_decap_8 FILLER_69_703 ();
 sg13g2_fill_2 FILLER_69_710 ();
 sg13g2_fill_1 FILLER_69_712 ();
 sg13g2_decap_8 FILLER_69_737 ();
 sg13g2_decap_8 FILLER_69_744 ();
 sg13g2_fill_2 FILLER_69_751 ();
 sg13g2_decap_8 FILLER_69_793 ();
 sg13g2_decap_8 FILLER_69_800 ();
 sg13g2_decap_8 FILLER_69_807 ();
 sg13g2_decap_8 FILLER_69_814 ();
 sg13g2_decap_8 FILLER_69_821 ();
 sg13g2_decap_8 FILLER_69_828 ();
 sg13g2_decap_8 FILLER_69_835 ();
 sg13g2_decap_8 FILLER_69_842 ();
 sg13g2_decap_8 FILLER_69_849 ();
 sg13g2_decap_8 FILLER_69_856 ();
 sg13g2_decap_8 FILLER_69_863 ();
 sg13g2_decap_8 FILLER_69_870 ();
 sg13g2_fill_1 FILLER_69_877 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_28 ();
 sg13g2_fill_1 FILLER_70_30 ();
 sg13g2_fill_2 FILLER_70_39 ();
 sg13g2_fill_1 FILLER_70_41 ();
 sg13g2_fill_1 FILLER_70_45 ();
 sg13g2_decap_4 FILLER_70_63 ();
 sg13g2_fill_1 FILLER_70_67 ();
 sg13g2_decap_8 FILLER_70_72 ();
 sg13g2_decap_8 FILLER_70_86 ();
 sg13g2_fill_1 FILLER_70_97 ();
 sg13g2_decap_4 FILLER_70_102 ();
 sg13g2_fill_1 FILLER_70_106 ();
 sg13g2_decap_8 FILLER_70_115 ();
 sg13g2_fill_1 FILLER_70_122 ();
 sg13g2_decap_8 FILLER_70_129 ();
 sg13g2_decap_8 FILLER_70_136 ();
 sg13g2_fill_2 FILLER_70_143 ();
 sg13g2_decap_8 FILLER_70_149 ();
 sg13g2_decap_8 FILLER_70_156 ();
 sg13g2_decap_8 FILLER_70_163 ();
 sg13g2_decap_8 FILLER_70_170 ();
 sg13g2_decap_8 FILLER_70_177 ();
 sg13g2_decap_8 FILLER_70_184 ();
 sg13g2_decap_8 FILLER_70_191 ();
 sg13g2_decap_8 FILLER_70_198 ();
 sg13g2_decap_8 FILLER_70_205 ();
 sg13g2_decap_8 FILLER_70_212 ();
 sg13g2_decap_8 FILLER_70_219 ();
 sg13g2_decap_8 FILLER_70_226 ();
 sg13g2_decap_8 FILLER_70_233 ();
 sg13g2_fill_2 FILLER_70_240 ();
 sg13g2_decap_8 FILLER_70_246 ();
 sg13g2_decap_8 FILLER_70_253 ();
 sg13g2_decap_8 FILLER_70_260 ();
 sg13g2_decap_8 FILLER_70_267 ();
 sg13g2_decap_8 FILLER_70_274 ();
 sg13g2_decap_8 FILLER_70_281 ();
 sg13g2_decap_8 FILLER_70_288 ();
 sg13g2_decap_8 FILLER_70_295 ();
 sg13g2_decap_8 FILLER_70_302 ();
 sg13g2_decap_8 FILLER_70_309 ();
 sg13g2_decap_8 FILLER_70_316 ();
 sg13g2_decap_8 FILLER_70_323 ();
 sg13g2_decap_8 FILLER_70_330 ();
 sg13g2_decap_8 FILLER_70_337 ();
 sg13g2_decap_8 FILLER_70_344 ();
 sg13g2_fill_2 FILLER_70_351 ();
 sg13g2_decap_8 FILLER_70_359 ();
 sg13g2_decap_8 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_391 ();
 sg13g2_decap_8 FILLER_70_398 ();
 sg13g2_decap_4 FILLER_70_405 ();
 sg13g2_decap_8 FILLER_70_414 ();
 sg13g2_decap_8 FILLER_70_421 ();
 sg13g2_decap_8 FILLER_70_428 ();
 sg13g2_fill_2 FILLER_70_435 ();
 sg13g2_decap_8 FILLER_70_445 ();
 sg13g2_decap_8 FILLER_70_452 ();
 sg13g2_decap_8 FILLER_70_459 ();
 sg13g2_decap_8 FILLER_70_466 ();
 sg13g2_decap_8 FILLER_70_473 ();
 sg13g2_decap_8 FILLER_70_480 ();
 sg13g2_decap_8 FILLER_70_487 ();
 sg13g2_decap_8 FILLER_70_494 ();
 sg13g2_decap_8 FILLER_70_501 ();
 sg13g2_decap_4 FILLER_70_508 ();
 sg13g2_fill_2 FILLER_70_512 ();
 sg13g2_decap_8 FILLER_70_544 ();
 sg13g2_fill_2 FILLER_70_556 ();
 sg13g2_decap_8 FILLER_70_583 ();
 sg13g2_decap_8 FILLER_70_590 ();
 sg13g2_decap_8 FILLER_70_597 ();
 sg13g2_decap_8 FILLER_70_634 ();
 sg13g2_decap_8 FILLER_70_641 ();
 sg13g2_decap_4 FILLER_70_648 ();
 sg13g2_fill_1 FILLER_70_652 ();
 sg13g2_decap_8 FILLER_70_683 ();
 sg13g2_decap_8 FILLER_70_690 ();
 sg13g2_decap_8 FILLER_70_697 ();
 sg13g2_decap_8 FILLER_70_734 ();
 sg13g2_decap_8 FILLER_70_741 ();
 sg13g2_decap_4 FILLER_70_748 ();
 sg13g2_fill_1 FILLER_70_752 ();
 sg13g2_decap_8 FILLER_70_760 ();
 sg13g2_decap_8 FILLER_70_767 ();
 sg13g2_decap_8 FILLER_70_778 ();
 sg13g2_decap_8 FILLER_70_785 ();
 sg13g2_decap_8 FILLER_70_792 ();
 sg13g2_decap_8 FILLER_70_799 ();
 sg13g2_decap_8 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_813 ();
 sg13g2_decap_8 FILLER_70_820 ();
 sg13g2_decap_8 FILLER_70_827 ();
 sg13g2_decap_8 FILLER_70_834 ();
 sg13g2_decap_8 FILLER_70_841 ();
 sg13g2_decap_8 FILLER_70_848 ();
 sg13g2_decap_8 FILLER_70_855 ();
 sg13g2_decap_8 FILLER_70_862 ();
 sg13g2_decap_8 FILLER_70_869 ();
 sg13g2_fill_2 FILLER_70_876 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_fill_2 FILLER_71_35 ();
 sg13g2_fill_1 FILLER_71_37 ();
 sg13g2_fill_1 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_47 ();
 sg13g2_fill_1 FILLER_71_54 ();
 sg13g2_fill_2 FILLER_71_60 ();
 sg13g2_decap_8 FILLER_71_67 ();
 sg13g2_decap_8 FILLER_71_74 ();
 sg13g2_fill_2 FILLER_71_81 ();
 sg13g2_fill_2 FILLER_71_101 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_4 FILLER_71_119 ();
 sg13g2_fill_2 FILLER_71_133 ();
 sg13g2_fill_2 FILLER_71_145 ();
 sg13g2_fill_1 FILLER_71_155 ();
 sg13g2_decap_8 FILLER_71_160 ();
 sg13g2_decap_8 FILLER_71_167 ();
 sg13g2_decap_8 FILLER_71_174 ();
 sg13g2_decap_8 FILLER_71_181 ();
 sg13g2_decap_8 FILLER_71_188 ();
 sg13g2_decap_8 FILLER_71_195 ();
 sg13g2_decap_8 FILLER_71_202 ();
 sg13g2_decap_8 FILLER_71_209 ();
 sg13g2_decap_8 FILLER_71_216 ();
 sg13g2_decap_8 FILLER_71_223 ();
 sg13g2_decap_8 FILLER_71_230 ();
 sg13g2_decap_8 FILLER_71_237 ();
 sg13g2_decap_8 FILLER_71_244 ();
 sg13g2_decap_8 FILLER_71_251 ();
 sg13g2_decap_8 FILLER_71_258 ();
 sg13g2_fill_2 FILLER_71_269 ();
 sg13g2_fill_1 FILLER_71_271 ();
 sg13g2_decap_8 FILLER_71_285 ();
 sg13g2_decap_8 FILLER_71_292 ();
 sg13g2_decap_8 FILLER_71_299 ();
 sg13g2_decap_8 FILLER_71_306 ();
 sg13g2_decap_8 FILLER_71_313 ();
 sg13g2_fill_1 FILLER_71_320 ();
 sg13g2_fill_1 FILLER_71_326 ();
 sg13g2_decap_8 FILLER_71_334 ();
 sg13g2_decap_4 FILLER_71_341 ();
 sg13g2_decap_8 FILLER_71_353 ();
 sg13g2_decap_8 FILLER_71_360 ();
 sg13g2_decap_8 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_decap_8 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_71_414 ();
 sg13g2_decap_8 FILLER_71_421 ();
 sg13g2_decap_8 FILLER_71_428 ();
 sg13g2_decap_8 FILLER_71_435 ();
 sg13g2_decap_8 FILLER_71_442 ();
 sg13g2_decap_8 FILLER_71_449 ();
 sg13g2_decap_8 FILLER_71_456 ();
 sg13g2_decap_8 FILLER_71_463 ();
 sg13g2_decap_8 FILLER_71_470 ();
 sg13g2_decap_8 FILLER_71_477 ();
 sg13g2_decap_8 FILLER_71_484 ();
 sg13g2_decap_8 FILLER_71_491 ();
 sg13g2_decap_8 FILLER_71_498 ();
 sg13g2_decap_8 FILLER_71_505 ();
 sg13g2_decap_8 FILLER_71_512 ();
 sg13g2_fill_2 FILLER_71_519 ();
 sg13g2_fill_1 FILLER_71_521 ();
 sg13g2_decap_8 FILLER_71_526 ();
 sg13g2_decap_4 FILLER_71_533 ();
 sg13g2_fill_1 FILLER_71_537 ();
 sg13g2_decap_8 FILLER_71_546 ();
 sg13g2_fill_2 FILLER_71_573 ();
 sg13g2_decap_4 FILLER_71_586 ();
 sg13g2_fill_1 FILLER_71_590 ();
 sg13g2_decap_8 FILLER_71_594 ();
 sg13g2_decap_8 FILLER_71_601 ();
 sg13g2_decap_8 FILLER_71_608 ();
 sg13g2_decap_8 FILLER_71_615 ();
 sg13g2_decap_8 FILLER_71_622 ();
 sg13g2_decap_8 FILLER_71_629 ();
 sg13g2_decap_8 FILLER_71_636 ();
 sg13g2_fill_2 FILLER_71_643 ();
 sg13g2_decap_8 FILLER_71_675 ();
 sg13g2_decap_8 FILLER_71_682 ();
 sg13g2_decap_8 FILLER_71_689 ();
 sg13g2_decap_8 FILLER_71_696 ();
 sg13g2_decap_8 FILLER_71_703 ();
 sg13g2_fill_2 FILLER_71_710 ();
 sg13g2_fill_1 FILLER_71_712 ();
 sg13g2_decap_8 FILLER_71_722 ();
 sg13g2_decap_8 FILLER_71_734 ();
 sg13g2_decap_8 FILLER_71_741 ();
 sg13g2_decap_4 FILLER_71_748 ();
 sg13g2_decap_4 FILLER_71_760 ();
 sg13g2_fill_2 FILLER_71_773 ();
 sg13g2_fill_1 FILLER_71_775 ();
 sg13g2_decap_8 FILLER_71_802 ();
 sg13g2_decap_8 FILLER_71_809 ();
 sg13g2_decap_8 FILLER_71_816 ();
 sg13g2_decap_8 FILLER_71_823 ();
 sg13g2_decap_8 FILLER_71_830 ();
 sg13g2_decap_8 FILLER_71_837 ();
 sg13g2_decap_8 FILLER_71_844 ();
 sg13g2_decap_8 FILLER_71_851 ();
 sg13g2_decap_8 FILLER_71_858 ();
 sg13g2_decap_8 FILLER_71_865 ();
 sg13g2_decap_4 FILLER_71_872 ();
 sg13g2_fill_2 FILLER_71_876 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_35 ();
 sg13g2_fill_1 FILLER_72_37 ();
 sg13g2_fill_1 FILLER_72_49 ();
 sg13g2_decap_4 FILLER_72_61 ();
 sg13g2_decap_4 FILLER_72_69 ();
 sg13g2_fill_1 FILLER_72_73 ();
 sg13g2_decap_8 FILLER_72_83 ();
 sg13g2_decap_8 FILLER_72_104 ();
 sg13g2_decap_8 FILLER_72_111 ();
 sg13g2_decap_8 FILLER_72_118 ();
 sg13g2_fill_2 FILLER_72_125 ();
 sg13g2_decap_4 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_164 ();
 sg13g2_decap_8 FILLER_72_171 ();
 sg13g2_decap_8 FILLER_72_178 ();
 sg13g2_decap_8 FILLER_72_185 ();
 sg13g2_decap_4 FILLER_72_192 ();
 sg13g2_decap_8 FILLER_72_200 ();
 sg13g2_fill_2 FILLER_72_207 ();
 sg13g2_decap_8 FILLER_72_235 ();
 sg13g2_decap_8 FILLER_72_242 ();
 sg13g2_decap_8 FILLER_72_249 ();
 sg13g2_decap_8 FILLER_72_291 ();
 sg13g2_decap_8 FILLER_72_298 ();
 sg13g2_decap_4 FILLER_72_305 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_decap_8 FILLER_72_340 ();
 sg13g2_decap_8 FILLER_72_347 ();
 sg13g2_decap_8 FILLER_72_354 ();
 sg13g2_decap_8 FILLER_72_361 ();
 sg13g2_decap_4 FILLER_72_368 ();
 sg13g2_fill_2 FILLER_72_372 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_decap_8 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_413 ();
 sg13g2_decap_8 FILLER_72_440 ();
 sg13g2_decap_8 FILLER_72_447 ();
 sg13g2_decap_8 FILLER_72_454 ();
 sg13g2_decap_8 FILLER_72_461 ();
 sg13g2_decap_8 FILLER_72_468 ();
 sg13g2_decap_8 FILLER_72_475 ();
 sg13g2_decap_8 FILLER_72_482 ();
 sg13g2_decap_8 FILLER_72_489 ();
 sg13g2_decap_4 FILLER_72_496 ();
 sg13g2_decap_8 FILLER_72_526 ();
 sg13g2_fill_2 FILLER_72_537 ();
 sg13g2_fill_1 FILLER_72_539 ();
 sg13g2_decap_8 FILLER_72_543 ();
 sg13g2_decap_8 FILLER_72_550 ();
 sg13g2_fill_2 FILLER_72_557 ();
 sg13g2_decap_8 FILLER_72_567 ();
 sg13g2_decap_8 FILLER_72_574 ();
 sg13g2_fill_1 FILLER_72_581 ();
 sg13g2_fill_1 FILLER_72_591 ();
 sg13g2_fill_2 FILLER_72_595 ();
 sg13g2_fill_1 FILLER_72_597 ();
 sg13g2_fill_1 FILLER_72_602 ();
 sg13g2_decap_8 FILLER_72_611 ();
 sg13g2_decap_8 FILLER_72_618 ();
 sg13g2_decap_8 FILLER_72_625 ();
 sg13g2_decap_8 FILLER_72_632 ();
 sg13g2_decap_8 FILLER_72_639 ();
 sg13g2_fill_2 FILLER_72_646 ();
 sg13g2_decap_4 FILLER_72_656 ();
 sg13g2_fill_1 FILLER_72_660 ();
 sg13g2_decap_8 FILLER_72_675 ();
 sg13g2_decap_8 FILLER_72_682 ();
 sg13g2_decap_8 FILLER_72_689 ();
 sg13g2_decap_8 FILLER_72_696 ();
 sg13g2_decap_8 FILLER_72_703 ();
 sg13g2_decap_8 FILLER_72_710 ();
 sg13g2_decap_8 FILLER_72_717 ();
 sg13g2_decap_8 FILLER_72_724 ();
 sg13g2_decap_8 FILLER_72_731 ();
 sg13g2_decap_8 FILLER_72_738 ();
 sg13g2_fill_1 FILLER_72_745 ();
 sg13g2_decap_8 FILLER_72_761 ();
 sg13g2_decap_8 FILLER_72_768 ();
 sg13g2_decap_8 FILLER_72_775 ();
 sg13g2_decap_8 FILLER_72_786 ();
 sg13g2_decap_8 FILLER_72_793 ();
 sg13g2_decap_8 FILLER_72_800 ();
 sg13g2_decap_8 FILLER_72_807 ();
 sg13g2_decap_8 FILLER_72_814 ();
 sg13g2_decap_8 FILLER_72_821 ();
 sg13g2_decap_8 FILLER_72_828 ();
 sg13g2_decap_8 FILLER_72_835 ();
 sg13g2_decap_8 FILLER_72_842 ();
 sg13g2_decap_8 FILLER_72_849 ();
 sg13g2_decap_8 FILLER_72_856 ();
 sg13g2_decap_8 FILLER_72_863 ();
 sg13g2_decap_8 FILLER_72_870 ();
 sg13g2_fill_1 FILLER_72_877 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_4 FILLER_73_49 ();
 sg13g2_fill_1 FILLER_73_53 ();
 sg13g2_fill_2 FILLER_73_68 ();
 sg13g2_fill_2 FILLER_73_79 ();
 sg13g2_decap_8 FILLER_73_85 ();
 sg13g2_decap_8 FILLER_73_96 ();
 sg13g2_decap_8 FILLER_73_106 ();
 sg13g2_decap_8 FILLER_73_113 ();
 sg13g2_fill_2 FILLER_73_120 ();
 sg13g2_fill_1 FILLER_73_122 ();
 sg13g2_decap_4 FILLER_73_127 ();
 sg13g2_fill_2 FILLER_73_146 ();
 sg13g2_fill_1 FILLER_73_148 ();
 sg13g2_fill_1 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_158 ();
 sg13g2_decap_8 FILLER_73_165 ();
 sg13g2_decap_8 FILLER_73_172 ();
 sg13g2_decap_8 FILLER_73_179 ();
 sg13g2_fill_2 FILLER_73_186 ();
 sg13g2_fill_1 FILLER_73_188 ();
 sg13g2_decap_8 FILLER_73_223 ();
 sg13g2_decap_8 FILLER_73_230 ();
 sg13g2_decap_8 FILLER_73_237 ();
 sg13g2_decap_8 FILLER_73_244 ();
 sg13g2_decap_8 FILLER_73_251 ();
 sg13g2_fill_2 FILLER_73_258 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_decap_4 FILLER_73_287 ();
 sg13g2_fill_2 FILLER_73_291 ();
 sg13g2_decap_8 FILLER_73_302 ();
 sg13g2_fill_1 FILLER_73_309 ();
 sg13g2_fill_2 FILLER_73_332 ();
 sg13g2_fill_2 FILLER_73_338 ();
 sg13g2_decap_8 FILLER_73_352 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_decap_8 FILLER_73_366 ();
 sg13g2_decap_8 FILLER_73_373 ();
 sg13g2_decap_8 FILLER_73_380 ();
 sg13g2_decap_8 FILLER_73_387 ();
 sg13g2_fill_2 FILLER_73_394 ();
 sg13g2_fill_1 FILLER_73_396 ();
 sg13g2_decap_8 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_73_412 ();
 sg13g2_fill_1 FILLER_73_419 ();
 sg13g2_fill_1 FILLER_73_424 ();
 sg13g2_decap_8 FILLER_73_428 ();
 sg13g2_decap_8 FILLER_73_435 ();
 sg13g2_decap_8 FILLER_73_442 ();
 sg13g2_decap_8 FILLER_73_449 ();
 sg13g2_fill_2 FILLER_73_456 ();
 sg13g2_decap_4 FILLER_73_462 ();
 sg13g2_fill_1 FILLER_73_466 ();
 sg13g2_fill_1 FILLER_73_472 ();
 sg13g2_fill_2 FILLER_73_477 ();
 sg13g2_decap_8 FILLER_73_483 ();
 sg13g2_decap_8 FILLER_73_490 ();
 sg13g2_decap_8 FILLER_73_497 ();
 sg13g2_decap_4 FILLER_73_504 ();
 sg13g2_fill_2 FILLER_73_508 ();
 sg13g2_decap_8 FILLER_73_514 ();
 sg13g2_fill_2 FILLER_73_521 ();
 sg13g2_fill_1 FILLER_73_527 ();
 sg13g2_decap_4 FILLER_73_539 ();
 sg13g2_fill_1 FILLER_73_543 ();
 sg13g2_decap_4 FILLER_73_549 ();
 sg13g2_fill_2 FILLER_73_553 ();
 sg13g2_decap_8 FILLER_73_569 ();
 sg13g2_fill_1 FILLER_73_576 ();
 sg13g2_decap_8 FILLER_73_590 ();
 sg13g2_decap_8 FILLER_73_597 ();
 sg13g2_decap_8 FILLER_73_604 ();
 sg13g2_decap_8 FILLER_73_611 ();
 sg13g2_fill_2 FILLER_73_618 ();
 sg13g2_decap_8 FILLER_73_625 ();
 sg13g2_decap_8 FILLER_73_632 ();
 sg13g2_decap_8 FILLER_73_639 ();
 sg13g2_fill_1 FILLER_73_646 ();
 sg13g2_decap_8 FILLER_73_659 ();
 sg13g2_fill_1 FILLER_73_666 ();
 sg13g2_decap_4 FILLER_73_671 ();
 sg13g2_fill_1 FILLER_73_675 ();
 sg13g2_decap_8 FILLER_73_680 ();
 sg13g2_decap_8 FILLER_73_691 ();
 sg13g2_fill_1 FILLER_73_698 ();
 sg13g2_decap_8 FILLER_73_707 ();
 sg13g2_decap_8 FILLER_73_714 ();
 sg13g2_decap_8 FILLER_73_721 ();
 sg13g2_decap_8 FILLER_73_728 ();
 sg13g2_decap_8 FILLER_73_735 ();
 sg13g2_decap_4 FILLER_73_742 ();
 sg13g2_fill_2 FILLER_73_752 ();
 sg13g2_decap_8 FILLER_73_758 ();
 sg13g2_decap_4 FILLER_73_765 ();
 sg13g2_decap_8 FILLER_73_773 ();
 sg13g2_decap_8 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_787 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_8 FILLER_73_857 ();
 sg13g2_decap_8 FILLER_73_864 ();
 sg13g2_decap_8 FILLER_73_871 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_fill_2 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_73 ();
 sg13g2_fill_1 FILLER_74_75 ();
 sg13g2_fill_1 FILLER_74_81 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_fill_2 FILLER_74_124 ();
 sg13g2_fill_1 FILLER_74_160 ();
 sg13g2_decap_4 FILLER_74_170 ();
 sg13g2_fill_1 FILLER_74_174 ();
 sg13g2_decap_8 FILLER_74_201 ();
 sg13g2_decap_4 FILLER_74_208 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_8 FILLER_74_252 ();
 sg13g2_decap_4 FILLER_74_259 ();
 sg13g2_decap_4 FILLER_74_289 ();
 sg13g2_fill_2 FILLER_74_293 ();
 sg13g2_fill_2 FILLER_74_321 ();
 sg13g2_decap_8 FILLER_74_349 ();
 sg13g2_decap_8 FILLER_74_356 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_decap_8 FILLER_74_370 ();
 sg13g2_decap_8 FILLER_74_377 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_fill_1 FILLER_74_406 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_decap_8 FILLER_74_427 ();
 sg13g2_decap_8 FILLER_74_434 ();
 sg13g2_decap_8 FILLER_74_441 ();
 sg13g2_decap_4 FILLER_74_448 ();
 sg13g2_fill_1 FILLER_74_452 ();
 sg13g2_decap_4 FILLER_74_484 ();
 sg13g2_decap_8 FILLER_74_498 ();
 sg13g2_decap_8 FILLER_74_505 ();
 sg13g2_decap_8 FILLER_74_512 ();
 sg13g2_decap_8 FILLER_74_519 ();
 sg13g2_decap_8 FILLER_74_526 ();
 sg13g2_decap_8 FILLER_74_533 ();
 sg13g2_fill_2 FILLER_74_540 ();
 sg13g2_fill_1 FILLER_74_542 ();
 sg13g2_decap_8 FILLER_74_548 ();
 sg13g2_decap_4 FILLER_74_555 ();
 sg13g2_decap_8 FILLER_74_565 ();
 sg13g2_decap_8 FILLER_74_572 ();
 sg13g2_fill_1 FILLER_74_579 ();
 sg13g2_fill_2 FILLER_74_605 ();
 sg13g2_fill_1 FILLER_74_607 ();
 sg13g2_decap_4 FILLER_74_612 ();
 sg13g2_fill_1 FILLER_74_616 ();
 sg13g2_fill_2 FILLER_74_646 ();
 sg13g2_fill_1 FILLER_74_648 ();
 sg13g2_decap_8 FILLER_74_659 ();
 sg13g2_decap_8 FILLER_74_666 ();
 sg13g2_decap_8 FILLER_74_673 ();
 sg13g2_decap_8 FILLER_74_680 ();
 sg13g2_fill_1 FILLER_74_687 ();
 sg13g2_decap_8 FILLER_74_695 ();
 sg13g2_fill_1 FILLER_74_702 ();
 sg13g2_fill_2 FILLER_74_707 ();
 sg13g2_decap_4 FILLER_74_730 ();
 sg13g2_decap_4 FILLER_74_738 ();
 sg13g2_fill_2 FILLER_74_745 ();
 sg13g2_fill_1 FILLER_74_747 ();
 sg13g2_decap_8 FILLER_74_761 ();
 sg13g2_fill_2 FILLER_74_768 ();
 sg13g2_fill_2 FILLER_74_775 ();
 sg13g2_fill_1 FILLER_74_777 ();
 sg13g2_decap_8 FILLER_74_804 ();
 sg13g2_decap_8 FILLER_74_811 ();
 sg13g2_decap_8 FILLER_74_818 ();
 sg13g2_decap_8 FILLER_74_825 ();
 sg13g2_decap_8 FILLER_74_832 ();
 sg13g2_decap_8 FILLER_74_839 ();
 sg13g2_decap_8 FILLER_74_846 ();
 sg13g2_decap_8 FILLER_74_853 ();
 sg13g2_decap_8 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_74_867 ();
 sg13g2_decap_4 FILLER_74_874 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_fill_2 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_52 ();
 sg13g2_fill_2 FILLER_75_56 ();
 sg13g2_fill_2 FILLER_75_66 ();
 sg13g2_decap_4 FILLER_75_71 ();
 sg13g2_fill_2 FILLER_75_75 ();
 sg13g2_decap_8 FILLER_75_81 ();
 sg13g2_decap_8 FILLER_75_88 ();
 sg13g2_decap_8 FILLER_75_95 ();
 sg13g2_decap_8 FILLER_75_102 ();
 sg13g2_decap_8 FILLER_75_109 ();
 sg13g2_decap_8 FILLER_75_116 ();
 sg13g2_fill_2 FILLER_75_123 ();
 sg13g2_fill_1 FILLER_75_125 ();
 sg13g2_decap_8 FILLER_75_144 ();
 sg13g2_decap_4 FILLER_75_151 ();
 sg13g2_decap_8 FILLER_75_159 ();
 sg13g2_decap_8 FILLER_75_166 ();
 sg13g2_decap_8 FILLER_75_173 ();
 sg13g2_fill_2 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_187 ();
 sg13g2_decap_8 FILLER_75_194 ();
 sg13g2_decap_8 FILLER_75_201 ();
 sg13g2_decap_8 FILLER_75_208 ();
 sg13g2_decap_8 FILLER_75_215 ();
 sg13g2_decap_8 FILLER_75_222 ();
 sg13g2_decap_8 FILLER_75_229 ();
 sg13g2_decap_8 FILLER_75_236 ();
 sg13g2_decap_8 FILLER_75_243 ();
 sg13g2_decap_8 FILLER_75_250 ();
 sg13g2_decap_8 FILLER_75_257 ();
 sg13g2_decap_8 FILLER_75_264 ();
 sg13g2_fill_1 FILLER_75_271 ();
 sg13g2_decap_8 FILLER_75_276 ();
 sg13g2_decap_8 FILLER_75_283 ();
 sg13g2_decap_8 FILLER_75_290 ();
 sg13g2_decap_4 FILLER_75_297 ();
 sg13g2_decap_8 FILLER_75_305 ();
 sg13g2_decap_8 FILLER_75_312 ();
 sg13g2_decap_8 FILLER_75_319 ();
 sg13g2_decap_8 FILLER_75_326 ();
 sg13g2_decap_8 FILLER_75_333 ();
 sg13g2_decap_8 FILLER_75_340 ();
 sg13g2_decap_8 FILLER_75_347 ();
 sg13g2_decap_4 FILLER_75_354 ();
 sg13g2_decap_4 FILLER_75_399 ();
 sg13g2_fill_1 FILLER_75_419 ();
 sg13g2_decap_8 FILLER_75_425 ();
 sg13g2_decap_8 FILLER_75_432 ();
 sg13g2_decap_8 FILLER_75_439 ();
 sg13g2_decap_8 FILLER_75_446 ();
 sg13g2_decap_8 FILLER_75_453 ();
 sg13g2_decap_8 FILLER_75_460 ();
 sg13g2_decap_8 FILLER_75_467 ();
 sg13g2_decap_8 FILLER_75_474 ();
 sg13g2_decap_8 FILLER_75_481 ();
 sg13g2_decap_8 FILLER_75_488 ();
 sg13g2_decap_8 FILLER_75_495 ();
 sg13g2_decap_8 FILLER_75_502 ();
 sg13g2_decap_8 FILLER_75_509 ();
 sg13g2_decap_8 FILLER_75_516 ();
 sg13g2_decap_8 FILLER_75_523 ();
 sg13g2_decap_8 FILLER_75_530 ();
 sg13g2_fill_1 FILLER_75_537 ();
 sg13g2_decap_8 FILLER_75_546 ();
 sg13g2_decap_8 FILLER_75_553 ();
 sg13g2_decap_8 FILLER_75_560 ();
 sg13g2_decap_8 FILLER_75_567 ();
 sg13g2_decap_4 FILLER_75_574 ();
 sg13g2_decap_4 FILLER_75_581 ();
 sg13g2_fill_2 FILLER_75_585 ();
 sg13g2_fill_1 FILLER_75_596 ();
 sg13g2_decap_8 FILLER_75_601 ();
 sg13g2_decap_8 FILLER_75_608 ();
 sg13g2_decap_8 FILLER_75_615 ();
 sg13g2_fill_2 FILLER_75_622 ();
 sg13g2_decap_8 FILLER_75_628 ();
 sg13g2_decap_8 FILLER_75_635 ();
 sg13g2_decap_8 FILLER_75_648 ();
 sg13g2_fill_1 FILLER_75_655 ();
 sg13g2_decap_8 FILLER_75_669 ();
 sg13g2_decap_8 FILLER_75_676 ();
 sg13g2_fill_2 FILLER_75_683 ();
 sg13g2_decap_8 FILLER_75_690 ();
 sg13g2_decap_4 FILLER_75_697 ();
 sg13g2_decap_4 FILLER_75_709 ();
 sg13g2_decap_4 FILLER_75_749 ();
 sg13g2_fill_1 FILLER_75_753 ();
 sg13g2_decap_8 FILLER_75_763 ();
 sg13g2_decap_4 FILLER_75_770 ();
 sg13g2_decap_8 FILLER_75_778 ();
 sg13g2_fill_1 FILLER_75_785 ();
 sg13g2_decap_8 FILLER_75_790 ();
 sg13g2_decap_8 FILLER_75_797 ();
 sg13g2_decap_8 FILLER_75_804 ();
 sg13g2_decap_8 FILLER_75_811 ();
 sg13g2_decap_8 FILLER_75_818 ();
 sg13g2_decap_8 FILLER_75_825 ();
 sg13g2_decap_8 FILLER_75_832 ();
 sg13g2_decap_8 FILLER_75_839 ();
 sg13g2_decap_8 FILLER_75_846 ();
 sg13g2_decap_8 FILLER_75_853 ();
 sg13g2_decap_8 FILLER_75_860 ();
 sg13g2_decap_8 FILLER_75_867 ();
 sg13g2_decap_4 FILLER_75_874 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_55 ();
 sg13g2_decap_8 FILLER_76_62 ();
 sg13g2_decap_8 FILLER_76_69 ();
 sg13g2_decap_8 FILLER_76_76 ();
 sg13g2_decap_8 FILLER_76_83 ();
 sg13g2_decap_8 FILLER_76_90 ();
 sg13g2_decap_8 FILLER_76_97 ();
 sg13g2_decap_8 FILLER_76_104 ();
 sg13g2_decap_8 FILLER_76_111 ();
 sg13g2_decap_4 FILLER_76_118 ();
 sg13g2_fill_2 FILLER_76_122 ();
 sg13g2_decap_4 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_141 ();
 sg13g2_decap_8 FILLER_76_148 ();
 sg13g2_decap_8 FILLER_76_155 ();
 sg13g2_decap_8 FILLER_76_162 ();
 sg13g2_decap_8 FILLER_76_169 ();
 sg13g2_decap_8 FILLER_76_176 ();
 sg13g2_decap_8 FILLER_76_183 ();
 sg13g2_decap_8 FILLER_76_190 ();
 sg13g2_decap_8 FILLER_76_197 ();
 sg13g2_decap_8 FILLER_76_204 ();
 sg13g2_decap_8 FILLER_76_211 ();
 sg13g2_decap_8 FILLER_76_218 ();
 sg13g2_decap_8 FILLER_76_225 ();
 sg13g2_decap_8 FILLER_76_232 ();
 sg13g2_decap_8 FILLER_76_239 ();
 sg13g2_decap_8 FILLER_76_246 ();
 sg13g2_decap_8 FILLER_76_253 ();
 sg13g2_decap_8 FILLER_76_260 ();
 sg13g2_decap_8 FILLER_76_267 ();
 sg13g2_decap_8 FILLER_76_274 ();
 sg13g2_decap_8 FILLER_76_281 ();
 sg13g2_decap_8 FILLER_76_288 ();
 sg13g2_decap_8 FILLER_76_295 ();
 sg13g2_decap_8 FILLER_76_302 ();
 sg13g2_decap_8 FILLER_76_309 ();
 sg13g2_decap_8 FILLER_76_316 ();
 sg13g2_decap_8 FILLER_76_323 ();
 sg13g2_decap_8 FILLER_76_330 ();
 sg13g2_decap_8 FILLER_76_337 ();
 sg13g2_fill_1 FILLER_76_344 ();
 sg13g2_decap_8 FILLER_76_348 ();
 sg13g2_decap_8 FILLER_76_355 ();
 sg13g2_fill_2 FILLER_76_362 ();
 sg13g2_decap_8 FILLER_76_368 ();
 sg13g2_decap_8 FILLER_76_375 ();
 sg13g2_decap_8 FILLER_76_382 ();
 sg13g2_decap_8 FILLER_76_389 ();
 sg13g2_decap_4 FILLER_76_396 ();
 sg13g2_fill_1 FILLER_76_400 ();
 sg13g2_fill_2 FILLER_76_409 ();
 sg13g2_fill_1 FILLER_76_411 ();
 sg13g2_decap_8 FILLER_76_442 ();
 sg13g2_decap_8 FILLER_76_449 ();
 sg13g2_decap_8 FILLER_76_456 ();
 sg13g2_decap_8 FILLER_76_463 ();
 sg13g2_decap_8 FILLER_76_470 ();
 sg13g2_decap_8 FILLER_76_477 ();
 sg13g2_decap_8 FILLER_76_484 ();
 sg13g2_decap_8 FILLER_76_491 ();
 sg13g2_decap_8 FILLER_76_498 ();
 sg13g2_decap_8 FILLER_76_505 ();
 sg13g2_decap_8 FILLER_76_512 ();
 sg13g2_decap_8 FILLER_76_519 ();
 sg13g2_decap_8 FILLER_76_526 ();
 sg13g2_fill_2 FILLER_76_533 ();
 sg13g2_decap_8 FILLER_76_561 ();
 sg13g2_decap_8 FILLER_76_568 ();
 sg13g2_decap_4 FILLER_76_583 ();
 sg13g2_fill_1 FILLER_76_594 ();
 sg13g2_decap_8 FILLER_76_600 ();
 sg13g2_decap_8 FILLER_76_607 ();
 sg13g2_decap_8 FILLER_76_614 ();
 sg13g2_decap_8 FILLER_76_621 ();
 sg13g2_decap_8 FILLER_76_628 ();
 sg13g2_decap_8 FILLER_76_635 ();
 sg13g2_decap_8 FILLER_76_647 ();
 sg13g2_decap_4 FILLER_76_654 ();
 sg13g2_fill_1 FILLER_76_658 ();
 sg13g2_decap_4 FILLER_76_682 ();
 sg13g2_fill_1 FILLER_76_686 ();
 sg13g2_fill_1 FILLER_76_690 ();
 sg13g2_decap_8 FILLER_76_701 ();
 sg13g2_decap_8 FILLER_76_708 ();
 sg13g2_fill_2 FILLER_76_734 ();
 sg13g2_fill_1 FILLER_76_736 ();
 sg13g2_fill_1 FILLER_76_742 ();
 sg13g2_decap_8 FILLER_76_746 ();
 sg13g2_decap_8 FILLER_76_753 ();
 sg13g2_decap_8 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_793 ();
 sg13g2_decap_8 FILLER_76_800 ();
 sg13g2_decap_8 FILLER_76_807 ();
 sg13g2_decap_8 FILLER_76_814 ();
 sg13g2_decap_8 FILLER_76_821 ();
 sg13g2_decap_8 FILLER_76_828 ();
 sg13g2_decap_8 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_decap_8 FILLER_76_856 ();
 sg13g2_decap_8 FILLER_76_863 ();
 sg13g2_decap_8 FILLER_76_870 ();
 sg13g2_fill_1 FILLER_76_877 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_4 FILLER_77_126 ();
 sg13g2_fill_2 FILLER_77_130 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_fill_2 FILLER_77_315 ();
 sg13g2_fill_1 FILLER_77_317 ();
 sg13g2_decap_8 FILLER_77_321 ();
 sg13g2_decap_8 FILLER_77_328 ();
 sg13g2_fill_1 FILLER_77_335 ();
 sg13g2_fill_2 FILLER_77_362 ();
 sg13g2_fill_2 FILLER_77_368 ();
 sg13g2_decap_8 FILLER_77_374 ();
 sg13g2_decap_8 FILLER_77_381 ();
 sg13g2_decap_8 FILLER_77_388 ();
 sg13g2_decap_8 FILLER_77_395 ();
 sg13g2_fill_1 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_77_411 ();
 sg13g2_decap_4 FILLER_77_418 ();
 sg13g2_fill_1 FILLER_77_422 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_448 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_8 FILLER_77_462 ();
 sg13g2_fill_2 FILLER_77_469 ();
 sg13g2_decap_8 FILLER_77_481 ();
 sg13g2_decap_8 FILLER_77_488 ();
 sg13g2_decap_8 FILLER_77_495 ();
 sg13g2_decap_8 FILLER_77_502 ();
 sg13g2_decap_8 FILLER_77_509 ();
 sg13g2_decap_8 FILLER_77_516 ();
 sg13g2_decap_8 FILLER_77_523 ();
 sg13g2_decap_4 FILLER_77_530 ();
 sg13g2_decap_4 FILLER_77_568 ();
 sg13g2_fill_1 FILLER_77_572 ();
 sg13g2_decap_8 FILLER_77_577 ();
 sg13g2_decap_4 FILLER_77_584 ();
 sg13g2_decap_8 FILLER_77_596 ();
 sg13g2_decap_8 FILLER_77_603 ();
 sg13g2_fill_2 FILLER_77_610 ();
 sg13g2_fill_1 FILLER_77_612 ();
 sg13g2_decap_8 FILLER_77_617 ();
 sg13g2_decap_8 FILLER_77_624 ();
 sg13g2_decap_8 FILLER_77_631 ();
 sg13g2_decap_8 FILLER_77_646 ();
 sg13g2_decap_8 FILLER_77_653 ();
 sg13g2_fill_1 FILLER_77_660 ();
 sg13g2_decap_4 FILLER_77_664 ();
 sg13g2_decap_8 FILLER_77_676 ();
 sg13g2_decap_8 FILLER_77_683 ();
 sg13g2_decap_8 FILLER_77_690 ();
 sg13g2_decap_8 FILLER_77_697 ();
 sg13g2_decap_8 FILLER_77_704 ();
 sg13g2_decap_8 FILLER_77_711 ();
 sg13g2_decap_8 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_755 ();
 sg13g2_decap_8 FILLER_77_762 ();
 sg13g2_decap_8 FILLER_77_769 ();
 sg13g2_decap_8 FILLER_77_776 ();
 sg13g2_decap_8 FILLER_77_783 ();
 sg13g2_decap_8 FILLER_77_790 ();
 sg13g2_decap_8 FILLER_77_797 ();
 sg13g2_decap_8 FILLER_77_804 ();
 sg13g2_decap_8 FILLER_77_811 ();
 sg13g2_decap_8 FILLER_77_818 ();
 sg13g2_decap_8 FILLER_77_825 ();
 sg13g2_decap_8 FILLER_77_832 ();
 sg13g2_decap_8 FILLER_77_839 ();
 sg13g2_decap_8 FILLER_77_846 ();
 sg13g2_decap_8 FILLER_77_853 ();
 sg13g2_decap_8 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_77_867 ();
 sg13g2_decap_4 FILLER_77_874 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_4 FILLER_78_63 ();
 sg13g2_fill_2 FILLER_78_67 ();
 sg13g2_decap_8 FILLER_78_95 ();
 sg13g2_decap_8 FILLER_78_102 ();
 sg13g2_fill_2 FILLER_78_109 ();
 sg13g2_fill_2 FILLER_78_115 ();
 sg13g2_decap_8 FILLER_78_121 ();
 sg13g2_decap_8 FILLER_78_128 ();
 sg13g2_decap_8 FILLER_78_135 ();
 sg13g2_decap_8 FILLER_78_142 ();
 sg13g2_decap_8 FILLER_78_149 ();
 sg13g2_fill_1 FILLER_78_156 ();
 sg13g2_decap_8 FILLER_78_183 ();
 sg13g2_decap_4 FILLER_78_190 ();
 sg13g2_fill_2 FILLER_78_194 ();
 sg13g2_decap_4 FILLER_78_200 ();
 sg13g2_fill_1 FILLER_78_204 ();
 sg13g2_decap_8 FILLER_78_209 ();
 sg13g2_decap_4 FILLER_78_216 ();
 sg13g2_fill_2 FILLER_78_220 ();
 sg13g2_decap_8 FILLER_78_226 ();
 sg13g2_decap_4 FILLER_78_233 ();
 sg13g2_fill_1 FILLER_78_237 ();
 sg13g2_fill_1 FILLER_78_249 ();
 sg13g2_decap_4 FILLER_78_253 ();
 sg13g2_decap_8 FILLER_78_261 ();
 sg13g2_decap_8 FILLER_78_268 ();
 sg13g2_decap_4 FILLER_78_275 ();
 sg13g2_fill_2 FILLER_78_279 ();
 sg13g2_fill_2 FILLER_78_312 ();
 sg13g2_fill_1 FILLER_78_318 ();
 sg13g2_decap_8 FILLER_78_377 ();
 sg13g2_decap_8 FILLER_78_384 ();
 sg13g2_decap_8 FILLER_78_391 ();
 sg13g2_decap_8 FILLER_78_398 ();
 sg13g2_decap_4 FILLER_78_405 ();
 sg13g2_fill_1 FILLER_78_409 ();
 sg13g2_decap_8 FILLER_78_436 ();
 sg13g2_decap_8 FILLER_78_443 ();
 sg13g2_decap_8 FILLER_78_450 ();
 sg13g2_decap_8 FILLER_78_457 ();
 sg13g2_decap_8 FILLER_78_464 ();
 sg13g2_decap_8 FILLER_78_471 ();
 sg13g2_decap_8 FILLER_78_478 ();
 sg13g2_decap_8 FILLER_78_485 ();
 sg13g2_decap_8 FILLER_78_492 ();
 sg13g2_decap_8 FILLER_78_499 ();
 sg13g2_decap_8 FILLER_78_506 ();
 sg13g2_decap_8 FILLER_78_513 ();
 sg13g2_decap_8 FILLER_78_520 ();
 sg13g2_decap_8 FILLER_78_527 ();
 sg13g2_decap_8 FILLER_78_534 ();
 sg13g2_decap_8 FILLER_78_541 ();
 sg13g2_fill_2 FILLER_78_548 ();
 sg13g2_fill_1 FILLER_78_550 ();
 sg13g2_decap_8 FILLER_78_555 ();
 sg13g2_decap_4 FILLER_78_562 ();
 sg13g2_decap_8 FILLER_78_603 ();
 sg13g2_decap_8 FILLER_78_610 ();
 sg13g2_decap_8 FILLER_78_617 ();
 sg13g2_decap_8 FILLER_78_624 ();
 sg13g2_decap_8 FILLER_78_631 ();
 sg13g2_fill_1 FILLER_78_638 ();
 sg13g2_fill_2 FILLER_78_643 ();
 sg13g2_decap_8 FILLER_78_649 ();
 sg13g2_decap_8 FILLER_78_656 ();
 sg13g2_decap_8 FILLER_78_663 ();
 sg13g2_decap_8 FILLER_78_670 ();
 sg13g2_fill_1 FILLER_78_677 ();
 sg13g2_decap_8 FILLER_78_682 ();
 sg13g2_decap_8 FILLER_78_689 ();
 sg13g2_decap_8 FILLER_78_696 ();
 sg13g2_decap_8 FILLER_78_703 ();
 sg13g2_decap_8 FILLER_78_710 ();
 sg13g2_decap_8 FILLER_78_717 ();
 sg13g2_decap_8 FILLER_78_724 ();
 sg13g2_decap_8 FILLER_78_731 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_decap_8 FILLER_78_745 ();
 sg13g2_decap_8 FILLER_78_752 ();
 sg13g2_decap_8 FILLER_78_759 ();
 sg13g2_decap_8 FILLER_78_766 ();
 sg13g2_decap_8 FILLER_78_773 ();
 sg13g2_decap_8 FILLER_78_780 ();
 sg13g2_decap_8 FILLER_78_787 ();
 sg13g2_decap_8 FILLER_78_794 ();
 sg13g2_decap_8 FILLER_78_801 ();
 sg13g2_decap_8 FILLER_78_808 ();
 sg13g2_decap_8 FILLER_78_815 ();
 sg13g2_decap_8 FILLER_78_822 ();
 sg13g2_decap_8 FILLER_78_829 ();
 sg13g2_decap_8 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_843 ();
 sg13g2_decap_8 FILLER_78_850 ();
 sg13g2_decap_8 FILLER_78_857 ();
 sg13g2_decap_8 FILLER_78_864 ();
 sg13g2_decap_8 FILLER_78_871 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_59 ();
 sg13g2_decap_8 FILLER_79_66 ();
 sg13g2_decap_4 FILLER_79_77 ();
 sg13g2_fill_2 FILLER_79_85 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_fill_1 FILLER_79_98 ();
 sg13g2_fill_2 FILLER_79_103 ();
 sg13g2_fill_1 FILLER_79_105 ();
 sg13g2_fill_2 FILLER_79_136 ();
 sg13g2_decap_8 FILLER_79_142 ();
 sg13g2_decap_8 FILLER_79_149 ();
 sg13g2_fill_2 FILLER_79_186 ();
 sg13g2_fill_1 FILLER_79_188 ();
 sg13g2_fill_2 FILLER_79_241 ();
 sg13g2_fill_1 FILLER_79_243 ();
 sg13g2_decap_8 FILLER_79_276 ();
 sg13g2_decap_4 FILLER_79_283 ();
 sg13g2_fill_1 FILLER_79_287 ();
 sg13g2_decap_4 FILLER_79_292 ();
 sg13g2_decap_8 FILLER_79_300 ();
 sg13g2_decap_8 FILLER_79_307 ();
 sg13g2_decap_8 FILLER_79_314 ();
 sg13g2_decap_4 FILLER_79_321 ();
 sg13g2_fill_1 FILLER_79_325 ();
 sg13g2_fill_1 FILLER_79_356 ();
 sg13g2_decap_8 FILLER_79_361 ();
 sg13g2_decap_8 FILLER_79_368 ();
 sg13g2_decap_8 FILLER_79_375 ();
 sg13g2_decap_8 FILLER_79_382 ();
 sg13g2_decap_8 FILLER_79_389 ();
 sg13g2_fill_2 FILLER_79_396 ();
 sg13g2_fill_1 FILLER_79_398 ();
 sg13g2_decap_8 FILLER_79_403 ();
 sg13g2_decap_4 FILLER_79_410 ();
 sg13g2_decap_8 FILLER_79_418 ();
 sg13g2_decap_8 FILLER_79_425 ();
 sg13g2_decap_8 FILLER_79_432 ();
 sg13g2_decap_8 FILLER_79_439 ();
 sg13g2_decap_8 FILLER_79_446 ();
 sg13g2_decap_8 FILLER_79_453 ();
 sg13g2_decap_8 FILLER_79_460 ();
 sg13g2_decap_8 FILLER_79_467 ();
 sg13g2_decap_8 FILLER_79_474 ();
 sg13g2_decap_8 FILLER_79_481 ();
 sg13g2_decap_8 FILLER_79_488 ();
 sg13g2_decap_8 FILLER_79_495 ();
 sg13g2_decap_8 FILLER_79_502 ();
 sg13g2_decap_8 FILLER_79_509 ();
 sg13g2_decap_8 FILLER_79_516 ();
 sg13g2_decap_8 FILLER_79_523 ();
 sg13g2_decap_8 FILLER_79_530 ();
 sg13g2_fill_2 FILLER_79_537 ();
 sg13g2_decap_8 FILLER_79_569 ();
 sg13g2_decap_8 FILLER_79_576 ();
 sg13g2_decap_8 FILLER_79_583 ();
 sg13g2_decap_8 FILLER_79_616 ();
 sg13g2_decap_8 FILLER_79_623 ();
 sg13g2_decap_8 FILLER_79_630 ();
 sg13g2_fill_2 FILLER_79_637 ();
 sg13g2_decap_4 FILLER_79_665 ();
 sg13g2_fill_2 FILLER_79_669 ();
 sg13g2_decap_8 FILLER_79_697 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_8 FILLER_79_711 ();
 sg13g2_fill_2 FILLER_79_718 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_decap_8 FILLER_79_753 ();
 sg13g2_decap_8 FILLER_79_760 ();
 sg13g2_decap_8 FILLER_79_767 ();
 sg13g2_decap_8 FILLER_79_774 ();
 sg13g2_decap_8 FILLER_79_781 ();
 sg13g2_decap_8 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_8 FILLER_79_858 ();
 sg13g2_decap_8 FILLER_79_865 ();
 sg13g2_decap_4 FILLER_79_872 ();
 sg13g2_fill_2 FILLER_79_876 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_fill_2 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_41 ();
 sg13g2_decap_4 FILLER_80_82 ();
 sg13g2_fill_2 FILLER_80_102 ();
 sg13g2_fill_1 FILLER_80_104 ();
 sg13g2_decap_4 FILLER_80_109 ();
 sg13g2_fill_2 FILLER_80_113 ();
 sg13g2_decap_4 FILLER_80_119 ();
 sg13g2_fill_2 FILLER_80_123 ();
 sg13g2_decap_4 FILLER_80_133 ();
 sg13g2_decap_8 FILLER_80_145 ();
 sg13g2_decap_8 FILLER_80_152 ();
 sg13g2_decap_4 FILLER_80_163 ();
 sg13g2_decap_4 FILLER_80_171 ();
 sg13g2_fill_1 FILLER_80_183 ();
 sg13g2_fill_1 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_201 ();
 sg13g2_decap_4 FILLER_80_209 ();
 sg13g2_decap_4 FILLER_80_217 ();
 sg13g2_fill_1 FILLER_80_225 ();
 sg13g2_fill_1 FILLER_80_230 ();
 sg13g2_decap_4 FILLER_80_235 ();
 sg13g2_fill_2 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_fill_2 FILLER_80_285 ();
 sg13g2_fill_1 FILLER_80_287 ();
 sg13g2_decap_8 FILLER_80_314 ();
 sg13g2_decap_8 FILLER_80_321 ();
 sg13g2_decap_4 FILLER_80_336 ();
 sg13g2_fill_1 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_fill_2 FILLER_80_355 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_decap_8 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_389 ();
 sg13g2_decap_8 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_403 ();
 sg13g2_decap_8 FILLER_80_410 ();
 sg13g2_decap_8 FILLER_80_417 ();
 sg13g2_decap_8 FILLER_80_424 ();
 sg13g2_decap_8 FILLER_80_431 ();
 sg13g2_decap_8 FILLER_80_438 ();
 sg13g2_decap_8 FILLER_80_445 ();
 sg13g2_decap_8 FILLER_80_452 ();
 sg13g2_decap_8 FILLER_80_459 ();
 sg13g2_decap_8 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_473 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_decap_8 FILLER_80_529 ();
 sg13g2_decap_8 FILLER_80_536 ();
 sg13g2_decap_8 FILLER_80_543 ();
 sg13g2_decap_8 FILLER_80_554 ();
 sg13g2_decap_8 FILLER_80_561 ();
 sg13g2_decap_8 FILLER_80_568 ();
 sg13g2_decap_8 FILLER_80_575 ();
 sg13g2_decap_8 FILLER_80_582 ();
 sg13g2_decap_8 FILLER_80_589 ();
 sg13g2_decap_8 FILLER_80_596 ();
 sg13g2_decap_8 FILLER_80_603 ();
 sg13g2_decap_8 FILLER_80_610 ();
 sg13g2_decap_8 FILLER_80_617 ();
 sg13g2_decap_8 FILLER_80_624 ();
 sg13g2_decap_8 FILLER_80_631 ();
 sg13g2_decap_8 FILLER_80_638 ();
 sg13g2_decap_8 FILLER_80_645 ();
 sg13g2_decap_8 FILLER_80_652 ();
 sg13g2_decap_8 FILLER_80_659 ();
 sg13g2_decap_8 FILLER_80_666 ();
 sg13g2_decap_8 FILLER_80_673 ();
 sg13g2_decap_8 FILLER_80_680 ();
 sg13g2_decap_8 FILLER_80_687 ();
 sg13g2_decap_8 FILLER_80_694 ();
 sg13g2_decap_8 FILLER_80_701 ();
 sg13g2_decap_8 FILLER_80_708 ();
 sg13g2_decap_8 FILLER_80_715 ();
 sg13g2_decap_4 FILLER_80_722 ();
 sg13g2_decap_8 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_744 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_8 FILLER_80_856 ();
 sg13g2_decap_8 FILLER_80_863 ();
 sg13g2_decap_8 FILLER_80_870 ();
 sg13g2_fill_1 FILLER_80_877 ();
endmodule
