module tt_um_kianv_bare_metal (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire clknet_leaf_0_clk;
 wire pwm_o;
 wire sclk;
 wire sio0_si_mosi_o;
 wire sio1_so_miso_o;
 wire sio2_o;
 wire sio3_o;
 wire \soc_I.PC[0] ;
 wire \soc_I.PC[10] ;
 wire \soc_I.PC[11] ;
 wire \soc_I.PC[12] ;
 wire \soc_I.PC[13] ;
 wire \soc_I.PC[14] ;
 wire \soc_I.PC[15] ;
 wire \soc_I.PC[16] ;
 wire \soc_I.PC[17] ;
 wire \soc_I.PC[18] ;
 wire \soc_I.PC[19] ;
 wire \soc_I.PC[1] ;
 wire \soc_I.PC[20] ;
 wire \soc_I.PC[21] ;
 wire \soc_I.PC[22] ;
 wire \soc_I.PC[23] ;
 wire \soc_I.PC[24] ;
 wire \soc_I.PC[25] ;
 wire \soc_I.PC[26] ;
 wire \soc_I.PC[27] ;
 wire \soc_I.PC[28] ;
 wire \soc_I.PC[29] ;
 wire \soc_I.PC[2] ;
 wire \soc_I.PC[30] ;
 wire \soc_I.PC[31] ;
 wire \soc_I.PC[3] ;
 wire \soc_I.PC[4] ;
 wire \soc_I.PC[5] ;
 wire \soc_I.PC[6] ;
 wire \soc_I.PC[7] ;
 wire \soc_I.PC[8] ;
 wire \soc_I.PC[9] ;
 wire \soc_I.cpu_mem_addr[0] ;
 wire \soc_I.cpu_mem_addr[1] ;
 wire \soc_I.cpu_mem_wdata[0] ;
 wire \soc_I.cpu_mem_wdata[1] ;
 wire \soc_I.cpu_mem_wdata[2] ;
 wire \soc_I.cpu_mem_wdata[3] ;
 wire \soc_I.cpu_mem_wdata[4] ;
 wire \soc_I.cpu_mem_wdata[5] ;
 wire \soc_I.cpu_mem_wdata[6] ;
 wire \soc_I.cpu_mem_wdata[7] ;
 wire \soc_I.cycle_cnt[0] ;
 wire \soc_I.cycle_cnt[10] ;
 wire \soc_I.cycle_cnt[11] ;
 wire \soc_I.cycle_cnt[12] ;
 wire \soc_I.cycle_cnt[13] ;
 wire \soc_I.cycle_cnt[14] ;
 wire \soc_I.cycle_cnt[15] ;
 wire \soc_I.cycle_cnt[16] ;
 wire \soc_I.cycle_cnt[17] ;
 wire \soc_I.cycle_cnt[18] ;
 wire \soc_I.cycle_cnt[19] ;
 wire \soc_I.cycle_cnt[1] ;
 wire \soc_I.cycle_cnt[20] ;
 wire \soc_I.cycle_cnt[21] ;
 wire \soc_I.cycle_cnt[22] ;
 wire \soc_I.cycle_cnt[23] ;
 wire \soc_I.cycle_cnt[24] ;
 wire \soc_I.cycle_cnt[25] ;
 wire \soc_I.cycle_cnt[26] ;
 wire \soc_I.cycle_cnt[27] ;
 wire \soc_I.cycle_cnt[28] ;
 wire \soc_I.cycle_cnt[29] ;
 wire \soc_I.cycle_cnt[2] ;
 wire \soc_I.cycle_cnt[30] ;
 wire \soc_I.cycle_cnt[31] ;
 wire \soc_I.cycle_cnt[3] ;
 wire \soc_I.cycle_cnt[4] ;
 wire \soc_I.cycle_cnt[5] ;
 wire \soc_I.cycle_cnt[6] ;
 wire \soc_I.cycle_cnt[7] ;
 wire \soc_I.cycle_cnt[8] ;
 wire \soc_I.cycle_cnt[9] ;
 wire \soc_I.cycle_cnt_ready ;
 wire \soc_I.div_ready ;
 wire \soc_I.div_reg[0] ;
 wire \soc_I.div_reg[10] ;
 wire \soc_I.div_reg[11] ;
 wire \soc_I.div_reg[12] ;
 wire \soc_I.div_reg[13] ;
 wire \soc_I.div_reg[14] ;
 wire \soc_I.div_reg[15] ;
 wire \soc_I.div_reg[16] ;
 wire \soc_I.div_reg[17] ;
 wire \soc_I.div_reg[18] ;
 wire \soc_I.div_reg[19] ;
 wire \soc_I.div_reg[1] ;
 wire \soc_I.div_reg[20] ;
 wire \soc_I.div_reg[21] ;
 wire \soc_I.div_reg[22] ;
 wire \soc_I.div_reg[23] ;
 wire \soc_I.div_reg[24] ;
 wire \soc_I.div_reg[25] ;
 wire \soc_I.div_reg[26] ;
 wire \soc_I.div_reg[27] ;
 wire \soc_I.div_reg[28] ;
 wire \soc_I.div_reg[29] ;
 wire \soc_I.div_reg[2] ;
 wire \soc_I.div_reg[30] ;
 wire \soc_I.div_reg[31] ;
 wire \soc_I.div_reg[3] ;
 wire \soc_I.div_reg[4] ;
 wire \soc_I.div_reg[5] ;
 wire \soc_I.div_reg[6] ;
 wire \soc_I.div_reg[7] ;
 wire \soc_I.div_reg[8] ;
 wire \soc_I.div_reg[9] ;
 wire \soc_I.kianv_I.Instr[0] ;
 wire \soc_I.kianv_I.Instr[10] ;
 wire \soc_I.kianv_I.Instr[11] ;
 wire \soc_I.kianv_I.Instr[12] ;
 wire \soc_I.kianv_I.Instr[13] ;
 wire \soc_I.kianv_I.Instr[14] ;
 wire \soc_I.kianv_I.Instr[15] ;
 wire \soc_I.kianv_I.Instr[16] ;
 wire \soc_I.kianv_I.Instr[17] ;
 wire \soc_I.kianv_I.Instr[18] ;
 wire \soc_I.kianv_I.Instr[19] ;
 wire \soc_I.kianv_I.Instr[1] ;
 wire \soc_I.kianv_I.Instr[20] ;
 wire \soc_I.kianv_I.Instr[21] ;
 wire \soc_I.kianv_I.Instr[22] ;
 wire \soc_I.kianv_I.Instr[23] ;
 wire \soc_I.kianv_I.Instr[24] ;
 wire \soc_I.kianv_I.Instr[25] ;
 wire \soc_I.kianv_I.Instr[26] ;
 wire \soc_I.kianv_I.Instr[27] ;
 wire \soc_I.kianv_I.Instr[28] ;
 wire \soc_I.kianv_I.Instr[29] ;
 wire \soc_I.kianv_I.Instr[2] ;
 wire \soc_I.kianv_I.Instr[30] ;
 wire \soc_I.kianv_I.Instr[31] ;
 wire \soc_I.kianv_I.Instr[3] ;
 wire \soc_I.kianv_I.Instr[4] ;
 wire \soc_I.kianv_I.Instr[5] ;
 wire \soc_I.kianv_I.Instr[6] ;
 wire \soc_I.kianv_I.Instr[7] ;
 wire \soc_I.kianv_I.Instr[8] ;
 wire \soc_I.kianv_I.Instr[9] ;
 wire \soc_I.kianv_I.MemWrite ;
 wire \soc_I.kianv_I.control_unit_I.Branch ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.resetn ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[0] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[10] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[11] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[12] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[13] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[1] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[2] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[3] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[4] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[6] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[7] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.ADDR_I.q[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.Addr_I.d0[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_ready ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.alu_I.shift_state ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ;
 wire \soc_I.pwm_I.pcm[0] ;
 wire \soc_I.pwm_I.pcm[1] ;
 wire \soc_I.pwm_I.pcm[2] ;
 wire \soc_I.pwm_I.pcm[3] ;
 wire \soc_I.pwm_I.pcm[4] ;
 wire \soc_I.pwm_I.pcm[5] ;
 wire \soc_I.pwm_I.pcm[6] ;
 wire \soc_I.pwm_I.pcm[7] ;
 wire \soc_I.pwm_I.pwm_accumulator[0] ;
 wire \soc_I.pwm_I.pwm_accumulator[1] ;
 wire \soc_I.pwm_I.pwm_accumulator[2] ;
 wire \soc_I.pwm_I.pwm_accumulator[3] ;
 wire \soc_I.pwm_I.pwm_accumulator[4] ;
 wire \soc_I.pwm_I.pwm_accumulator[5] ;
 wire \soc_I.pwm_I.pwm_accumulator[6] ;
 wire \soc_I.pwm_I.pwm_accumulator[7] ;
 wire \soc_I.pwm_ready ;
 wire \soc_I.qqspi_I.is_quad ;
 wire \soc_I.qqspi_I.rdata[0] ;
 wire \soc_I.qqspi_I.rdata[10] ;
 wire \soc_I.qqspi_I.rdata[11] ;
 wire \soc_I.qqspi_I.rdata[12] ;
 wire \soc_I.qqspi_I.rdata[13] ;
 wire \soc_I.qqspi_I.rdata[14] ;
 wire \soc_I.qqspi_I.rdata[15] ;
 wire \soc_I.qqspi_I.rdata[16] ;
 wire \soc_I.qqspi_I.rdata[17] ;
 wire \soc_I.qqspi_I.rdata[18] ;
 wire \soc_I.qqspi_I.rdata[19] ;
 wire \soc_I.qqspi_I.rdata[1] ;
 wire \soc_I.qqspi_I.rdata[20] ;
 wire \soc_I.qqspi_I.rdata[21] ;
 wire \soc_I.qqspi_I.rdata[22] ;
 wire \soc_I.qqspi_I.rdata[23] ;
 wire \soc_I.qqspi_I.rdata[24] ;
 wire \soc_I.qqspi_I.rdata[25] ;
 wire \soc_I.qqspi_I.rdata[26] ;
 wire \soc_I.qqspi_I.rdata[27] ;
 wire \soc_I.qqspi_I.rdata[28] ;
 wire \soc_I.qqspi_I.rdata[29] ;
 wire \soc_I.qqspi_I.rdata[2] ;
 wire \soc_I.qqspi_I.rdata[30] ;
 wire \soc_I.qqspi_I.rdata[31] ;
 wire \soc_I.qqspi_I.rdata[3] ;
 wire \soc_I.qqspi_I.rdata[4] ;
 wire \soc_I.qqspi_I.rdata[5] ;
 wire \soc_I.qqspi_I.rdata[6] ;
 wire \soc_I.qqspi_I.rdata[7] ;
 wire \soc_I.qqspi_I.rdata[8] ;
 wire \soc_I.qqspi_I.rdata[9] ;
 wire \soc_I.qqspi_I.ready ;
 wire \soc_I.qqspi_I.spi_buf[0] ;
 wire \soc_I.qqspi_I.spi_buf[10] ;
 wire \soc_I.qqspi_I.spi_buf[11] ;
 wire \soc_I.qqspi_I.spi_buf[12] ;
 wire \soc_I.qqspi_I.spi_buf[13] ;
 wire \soc_I.qqspi_I.spi_buf[14] ;
 wire \soc_I.qqspi_I.spi_buf[15] ;
 wire \soc_I.qqspi_I.spi_buf[16] ;
 wire \soc_I.qqspi_I.spi_buf[17] ;
 wire \soc_I.qqspi_I.spi_buf[18] ;
 wire \soc_I.qqspi_I.spi_buf[19] ;
 wire \soc_I.qqspi_I.spi_buf[1] ;
 wire \soc_I.qqspi_I.spi_buf[20] ;
 wire \soc_I.qqspi_I.spi_buf[21] ;
 wire \soc_I.qqspi_I.spi_buf[22] ;
 wire \soc_I.qqspi_I.spi_buf[23] ;
 wire \soc_I.qqspi_I.spi_buf[24] ;
 wire \soc_I.qqspi_I.spi_buf[25] ;
 wire \soc_I.qqspi_I.spi_buf[26] ;
 wire \soc_I.qqspi_I.spi_buf[27] ;
 wire \soc_I.qqspi_I.spi_buf[28] ;
 wire \soc_I.qqspi_I.spi_buf[29] ;
 wire \soc_I.qqspi_I.spi_buf[2] ;
 wire \soc_I.qqspi_I.spi_buf[30] ;
 wire \soc_I.qqspi_I.spi_buf[31] ;
 wire \soc_I.qqspi_I.spi_buf[3] ;
 wire \soc_I.qqspi_I.spi_buf[4] ;
 wire \soc_I.qqspi_I.spi_buf[5] ;
 wire \soc_I.qqspi_I.spi_buf[6] ;
 wire \soc_I.qqspi_I.spi_buf[7] ;
 wire \soc_I.qqspi_I.spi_buf[8] ;
 wire \soc_I.qqspi_I.spi_buf[9] ;
 wire \soc_I.qqspi_I.state[0] ;
 wire \soc_I.qqspi_I.state[1] ;
 wire \soc_I.qqspi_I.state[2] ;
 wire \soc_I.qqspi_I.state[3] ;
 wire \soc_I.qqspi_I.state[4] ;
 wire \soc_I.qqspi_I.state[5] ;
 wire \soc_I.qqspi_I.state[6] ;
 wire \soc_I.qqspi_I.xfer_cycles[0] ;
 wire \soc_I.qqspi_I.xfer_cycles[1] ;
 wire \soc_I.qqspi_I.xfer_cycles[2] ;
 wire \soc_I.qqspi_I.xfer_cycles[3] ;
 wire \soc_I.qqspi_I.xfer_cycles[4] ;
 wire \soc_I.qqspi_I.xfer_cycles[5] ;
 wire \soc_I.rst_cnt[0] ;
 wire \soc_I.rst_cnt[1] ;
 wire \soc_I.rst_cnt[2] ;
 wire \soc_I.rx_uart_i.bit_idx[0] ;
 wire \soc_I.rx_uart_i.bit_idx[1] ;
 wire \soc_I.rx_uart_i.bit_idx[2] ;
 wire \soc_I.rx_uart_i.data_rd ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[0] ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[1] ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[2] ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[3] ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[4] ;
 wire \soc_I.rx_uart_i.fifo_i.din[0] ;
 wire \soc_I.rx_uart_i.fifo_i.din[1] ;
 wire \soc_I.rx_uart_i.fifo_i.din[2] ;
 wire \soc_I.rx_uart_i.fifo_i.din[3] ;
 wire \soc_I.rx_uart_i.fifo_i.din[4] ;
 wire \soc_I.rx_uart_i.fifo_i.din[5] ;
 wire \soc_I.rx_uart_i.fifo_i.din[6] ;
 wire \soc_I.rx_uart_i.fifo_i.din[7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][7] ;
 wire \soc_I.rx_uart_i.fifo_i.rd_ptr[0] ;
 wire \soc_I.rx_uart_i.fifo_i.rd_ptr[1] ;
 wire \soc_I.rx_uart_i.fifo_i.rd_ptr[2] ;
 wire \soc_I.rx_uart_i.fifo_i.rd_ptr[3] ;
 wire \soc_I.rx_uart_i.fifo_i.wr_ptr[0] ;
 wire \soc_I.rx_uart_i.fifo_i.wr_ptr[1] ;
 wire \soc_I.rx_uart_i.fifo_i.wr_ptr[2] ;
 wire \soc_I.rx_uart_i.fifo_i.wr_ptr[3] ;
 wire \soc_I.rx_uart_i.ready ;
 wire \soc_I.rx_uart_i.return_state[0] ;
 wire \soc_I.rx_uart_i.return_state[1] ;
 wire \soc_I.rx_uart_i.rx_in_sync[0] ;
 wire \soc_I.rx_uart_i.rx_in_sync[1] ;
 wire \soc_I.rx_uart_i.rx_in_sync[2] ;
 wire \soc_I.rx_uart_i.state[0] ;
 wire \soc_I.rx_uart_i.state[1] ;
 wire \soc_I.rx_uart_i.state[2] ;
 wire \soc_I.rx_uart_i.wait_states[0] ;
 wire \soc_I.rx_uart_i.wait_states[10] ;
 wire \soc_I.rx_uart_i.wait_states[11] ;
 wire \soc_I.rx_uart_i.wait_states[12] ;
 wire \soc_I.rx_uart_i.wait_states[13] ;
 wire \soc_I.rx_uart_i.wait_states[14] ;
 wire \soc_I.rx_uart_i.wait_states[15] ;
 wire \soc_I.rx_uart_i.wait_states[16] ;
 wire \soc_I.rx_uart_i.wait_states[1] ;
 wire \soc_I.rx_uart_i.wait_states[2] ;
 wire \soc_I.rx_uart_i.wait_states[3] ;
 wire \soc_I.rx_uart_i.wait_states[4] ;
 wire \soc_I.rx_uart_i.wait_states[5] ;
 wire \soc_I.rx_uart_i.wait_states[6] ;
 wire \soc_I.rx_uart_i.wait_states[7] ;
 wire \soc_I.rx_uart_i.wait_states[8] ;
 wire \soc_I.rx_uart_i.wait_states[9] ;
 wire \soc_I.spi0_I.cen ;
 wire \soc_I.spi0_I.div[0] ;
 wire \soc_I.spi0_I.div[10] ;
 wire \soc_I.spi0_I.div[11] ;
 wire \soc_I.spi0_I.div[12] ;
 wire \soc_I.spi0_I.div[13] ;
 wire \soc_I.spi0_I.div[14] ;
 wire \soc_I.spi0_I.div[15] ;
 wire \soc_I.spi0_I.div[1] ;
 wire \soc_I.spi0_I.div[2] ;
 wire \soc_I.spi0_I.div[3] ;
 wire \soc_I.spi0_I.div[4] ;
 wire \soc_I.spi0_I.div[5] ;
 wire \soc_I.spi0_I.div[6] ;
 wire \soc_I.spi0_I.div[7] ;
 wire \soc_I.spi0_I.div[8] ;
 wire \soc_I.spi0_I.div[9] ;
 wire \soc_I.spi0_I.ready_ctrl ;
 wire \soc_I.spi0_I.ready_xfer ;
 wire \soc_I.spi0_I.rx_data[0] ;
 wire \soc_I.spi0_I.rx_data[1] ;
 wire \soc_I.spi0_I.rx_data[2] ;
 wire \soc_I.spi0_I.rx_data[3] ;
 wire \soc_I.spi0_I.rx_data[4] ;
 wire \soc_I.spi0_I.rx_data[5] ;
 wire \soc_I.spi0_I.rx_data[6] ;
 wire \soc_I.spi0_I.rx_data[7] ;
 wire \soc_I.spi0_I.sclk ;
 wire \soc_I.spi0_I.sio0_si_mosi ;
 wire \soc_I.spi0_I.spi_buf[0] ;
 wire \soc_I.spi0_I.spi_buf[1] ;
 wire \soc_I.spi0_I.spi_buf[2] ;
 wire \soc_I.spi0_I.spi_buf[3] ;
 wire \soc_I.spi0_I.spi_buf[4] ;
 wire \soc_I.spi0_I.spi_buf[5] ;
 wire \soc_I.spi0_I.spi_buf[6] ;
 wire \soc_I.spi0_I.spi_buf[7] ;
 wire \soc_I.spi0_I.state ;
 wire \soc_I.spi0_I.tick_cnt[0] ;
 wire \soc_I.spi0_I.tick_cnt[10] ;
 wire \soc_I.spi0_I.tick_cnt[11] ;
 wire \soc_I.spi0_I.tick_cnt[12] ;
 wire \soc_I.spi0_I.tick_cnt[13] ;
 wire \soc_I.spi0_I.tick_cnt[14] ;
 wire \soc_I.spi0_I.tick_cnt[15] ;
 wire \soc_I.spi0_I.tick_cnt[16] ;
 wire \soc_I.spi0_I.tick_cnt[17] ;
 wire \soc_I.spi0_I.tick_cnt[1] ;
 wire \soc_I.spi0_I.tick_cnt[2] ;
 wire \soc_I.spi0_I.tick_cnt[3] ;
 wire \soc_I.spi0_I.tick_cnt[4] ;
 wire \soc_I.spi0_I.tick_cnt[5] ;
 wire \soc_I.spi0_I.tick_cnt[6] ;
 wire \soc_I.spi0_I.tick_cnt[7] ;
 wire \soc_I.spi0_I.tick_cnt[8] ;
 wire \soc_I.spi0_I.tick_cnt[9] ;
 wire \soc_I.spi0_I.xfer_cycles[0] ;
 wire \soc_I.spi0_I.xfer_cycles[1] ;
 wire \soc_I.spi0_I.xfer_cycles[2] ;
 wire \soc_I.spi0_I.xfer_cycles[3] ;
 wire \soc_I.spi0_I.xfer_cycles[4] ;
 wire \soc_I.spi0_I.xfer_cycles[5] ;
 wire \soc_I.spi_div_ready ;
 wire \soc_I.spi_div_reg[16] ;
 wire \soc_I.spi_div_reg[17] ;
 wire \soc_I.spi_div_reg[18] ;
 wire \soc_I.spi_div_reg[19] ;
 wire \soc_I.spi_div_reg[20] ;
 wire \soc_I.spi_div_reg[21] ;
 wire \soc_I.spi_div_reg[22] ;
 wire \soc_I.spi_div_reg[23] ;
 wire \soc_I.spi_div_reg[24] ;
 wire \soc_I.spi_div_reg[25] ;
 wire \soc_I.spi_div_reg[26] ;
 wire \soc_I.spi_div_reg[27] ;
 wire \soc_I.spi_div_reg[28] ;
 wire \soc_I.spi_div_reg[29] ;
 wire \soc_I.spi_div_reg[30] ;
 wire \soc_I.spi_div_reg[31] ;
 wire \soc_I.tx_uart_i.bit_idx[0] ;
 wire \soc_I.tx_uart_i.bit_idx[1] ;
 wire \soc_I.tx_uart_i.bit_idx[2] ;
 wire \soc_I.tx_uart_i.ready ;
 wire \soc_I.tx_uart_i.return_state[0] ;
 wire \soc_I.tx_uart_i.return_state[1] ;
 wire \soc_I.tx_uart_i.state[0] ;
 wire \soc_I.tx_uart_i.state[1] ;
 wire \soc_I.tx_uart_i.tx_data_reg[0] ;
 wire \soc_I.tx_uart_i.tx_data_reg[1] ;
 wire \soc_I.tx_uart_i.tx_data_reg[2] ;
 wire \soc_I.tx_uart_i.tx_data_reg[3] ;
 wire \soc_I.tx_uart_i.tx_data_reg[4] ;
 wire \soc_I.tx_uart_i.tx_data_reg[5] ;
 wire \soc_I.tx_uart_i.tx_data_reg[6] ;
 wire \soc_I.tx_uart_i.tx_data_reg[7] ;
 wire \soc_I.tx_uart_i.tx_out ;
 wire \soc_I.tx_uart_i.wait_states[0] ;
 wire \soc_I.tx_uart_i.wait_states[10] ;
 wire \soc_I.tx_uart_i.wait_states[11] ;
 wire \soc_I.tx_uart_i.wait_states[12] ;
 wire \soc_I.tx_uart_i.wait_states[13] ;
 wire \soc_I.tx_uart_i.wait_states[14] ;
 wire \soc_I.tx_uart_i.wait_states[15] ;
 wire \soc_I.tx_uart_i.wait_states[1] ;
 wire \soc_I.tx_uart_i.wait_states[2] ;
 wire \soc_I.tx_uart_i.wait_states[3] ;
 wire \soc_I.tx_uart_i.wait_states[4] ;
 wire \soc_I.tx_uart_i.wait_states[5] ;
 wire \soc_I.tx_uart_i.wait_states[6] ;
 wire \soc_I.tx_uart_i.wait_states[7] ;
 wire \soc_I.tx_uart_i.wait_states[8] ;
 wire \soc_I.tx_uart_i.wait_states[9] ;
 wire \soc_I.uart_lsr_rdy ;
 wire \soc_I.uart_tx_ready ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _08988_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[11] ),
    .X(_01556_));
 sg13g2_buf_1 _08989_ (.A(\soc_I.kianv_I.MemWrite ),
    .X(_01557_));
 sg13g2_nor2_1 _08990_ (.A(_01556_),
    .B(_01557_),
    .Y(_01558_));
 sg13g2_buf_1 _08991_ (.A(_01558_),
    .X(_01559_));
 sg13g2_buf_1 _08992_ (.A(net530),
    .X(_01560_));
 sg13g2_buf_1 _08993_ (.A(\soc_I.kianv_I.control_unit_I.Branch ),
    .X(_01561_));
 sg13g2_buf_2 _08994_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[4] ),
    .X(_01562_));
 sg13g2_buf_1 _08995_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[12] ),
    .X(_01563_));
 sg13g2_buf_1 _08996_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[6] ),
    .X(_01564_));
 sg13g2_buf_1 _08997_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[1] ),
    .X(_01565_));
 sg13g2_or2_1 _08998_ (.X(_01566_),
    .B(_01565_),
    .A(_01564_));
 sg13g2_buf_1 _08999_ (.A(_01566_),
    .X(_01567_));
 sg13g2_nor4_1 _09000_ (.A(net633),
    .B(_01562_),
    .C(_01563_),
    .D(_01567_),
    .Y(_01568_));
 sg13g2_buf_2 _09001_ (.A(_01568_),
    .X(_01569_));
 sg13g2_buf_8 _09002_ (.A(_01569_),
    .X(_01570_));
 sg13g2_buf_8 _09003_ (.A(net370),
    .X(_01571_));
 sg13g2_buf_1 _09004_ (.A(net343),
    .X(_01572_));
 sg13g2_buf_1 _09005_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[1] ),
    .X(_01573_));
 sg13g2_buf_2 _09006_ (.A(_00032_),
    .X(_01574_));
 sg13g2_inv_1 _09007_ (.Y(_01575_),
    .A(_01574_));
 sg13g2_buf_1 _09008_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[7] ),
    .X(_01576_));
 sg13g2_buf_2 _09009_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[8] ),
    .X(_01577_));
 sg13g2_or2_1 _09010_ (.X(_01578_),
    .B(_01577_),
    .A(net632));
 sg13g2_buf_1 _09011_ (.A(_01578_),
    .X(_01579_));
 sg13g2_nor2_1 _09012_ (.A(_01575_),
    .B(_01579_),
    .Y(_01580_));
 sg13g2_buf_1 _09013_ (.A(_01580_),
    .X(_01581_));
 sg13g2_buf_8 _09014_ (.A(net420),
    .X(_01582_));
 sg13g2_mux2_1 _09015_ (.A0(\soc_I.PC[1] ),
    .A1(_01573_),
    .S(net369),
    .X(_01583_));
 sg13g2_or4_1 _09016_ (.A(net633),
    .B(_01562_),
    .C(_01563_),
    .D(_01567_),
    .X(_01584_));
 sg13g2_buf_1 _09017_ (.A(_01584_),
    .X(_01585_));
 sg13g2_buf_1 _09018_ (.A(net419),
    .X(_01586_));
 sg13g2_and2_1 _09019_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[1] ),
    .B(_01586_),
    .X(_01587_));
 sg13g2_a21o_1 _09020_ (.A2(_01583_),
    .A1(net326),
    .B1(_01587_),
    .X(_01588_));
 sg13g2_buf_1 _09021_ (.A(_01588_),
    .X(_01589_));
 sg13g2_buf_2 _09022_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[3] ),
    .X(_01590_));
 sg13g2_inv_1 _09023_ (.Y(_01591_),
    .A(_01590_));
 sg13g2_nor2_1 _09024_ (.A(_01564_),
    .B(_01565_),
    .Y(_01592_));
 sg13g2_buf_2 _09025_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[10] ),
    .X(_01593_));
 sg13g2_buf_1 _09026_ (.A(_00031_),
    .X(_01594_));
 sg13g2_nand2b_1 _09027_ (.Y(_01595_),
    .B(_01594_),
    .A_N(_01593_));
 sg13g2_nand4_1 _09028_ (.B(net633),
    .C(_01592_),
    .A(_01591_),
    .Y(_01596_),
    .D(_01595_));
 sg13g2_buf_2 _09029_ (.A(_01596_),
    .X(_01597_));
 sg13g2_or2_1 _09030_ (.X(_01598_),
    .B(_01593_),
    .A(_01590_));
 sg13g2_buf_1 _09031_ (.A(_01598_),
    .X(_01599_));
 sg13g2_nor3_1 _09032_ (.A(net633),
    .B(_01592_),
    .C(_01599_),
    .Y(_01600_));
 sg13g2_buf_1 _09033_ (.A(_00028_),
    .X(_01601_));
 sg13g2_nor2_1 _09034_ (.A(\soc_I.kianv_I.Instr[12] ),
    .B(net631),
    .Y(_01602_));
 sg13g2_buf_1 _09035_ (.A(\soc_I.kianv_I.Instr[13] ),
    .X(_01603_));
 sg13g2_inv_1 _09036_ (.Y(_01604_),
    .A(_01603_));
 sg13g2_buf_1 _09037_ (.A(_01604_),
    .X(_01605_));
 sg13g2_nand3b_1 _09038_ (.B(_00027_),
    .C(net529),
    .Y(_01606_),
    .A_N(_01602_));
 sg13g2_buf_1 _09039_ (.A(_01606_),
    .X(_01607_));
 sg13g2_and2_1 _09040_ (.A(_01600_),
    .B(_01607_),
    .X(_01608_));
 sg13g2_buf_1 _09041_ (.A(_01603_),
    .X(_01609_));
 sg13g2_buf_1 _09042_ (.A(\soc_I.kianv_I.Instr[12] ),
    .X(_01610_));
 sg13g2_nand2b_1 _09043_ (.Y(_01611_),
    .B(net630),
    .A_N(net631));
 sg13g2_buf_1 _09044_ (.A(\soc_I.kianv_I.Instr[14] ),
    .X(_01612_));
 sg13g2_buf_1 _09045_ (.A(_01612_),
    .X(_01613_));
 sg13g2_or2_1 _09046_ (.X(_01614_),
    .B(net630),
    .A(net602));
 sg13g2_nand3_1 _09047_ (.B(_01611_),
    .C(_01614_),
    .A(net603),
    .Y(_01615_));
 sg13g2_o21ai_1 _09048_ (.B1(_01615_),
    .Y(_01616_),
    .A1(net603),
    .A2(net631));
 sg13g2_nand2_1 _09049_ (.Y(_01617_),
    .A(net602),
    .B(net529));
 sg13g2_nor2_2 _09050_ (.A(net633),
    .B(_01593_),
    .Y(_01618_));
 sg13g2_nand2_1 _09051_ (.Y(_01619_),
    .A(_01590_),
    .B(_01618_));
 sg13g2_o21ai_1 _09052_ (.B1(_01619_),
    .Y(_01620_),
    .A1(_01617_),
    .A2(_01597_));
 sg13g2_a21o_1 _09053_ (.A2(_01616_),
    .A1(_01608_),
    .B1(_01620_),
    .X(_01621_));
 sg13g2_buf_1 _09054_ (.A(_01621_),
    .X(_01622_));
 sg13g2_buf_8 _09055_ (.A(_01622_),
    .X(_01623_));
 sg13g2_nand3b_1 _09056_ (.B(net631),
    .C(_01612_),
    .Y(_01624_),
    .A_N(_01603_));
 sg13g2_nand2b_1 _09057_ (.Y(_01625_),
    .B(net603),
    .A_N(_01612_));
 sg13g2_and3_1 _09058_ (.X(_01626_),
    .A(net630),
    .B(_01624_),
    .C(_01625_));
 sg13g2_nand3_1 _09059_ (.B(_01600_),
    .C(_01607_),
    .A(_01626_),
    .Y(_01627_));
 sg13g2_buf_2 _09060_ (.A(_01627_),
    .X(_01628_));
 sg13g2_o21ai_1 _09061_ (.B1(_01591_),
    .Y(_01629_),
    .A1(_01625_),
    .A2(_01592_));
 sg13g2_nand2b_1 _09062_ (.Y(_01630_),
    .B(_01593_),
    .A_N(net633));
 sg13g2_nand3b_1 _09063_ (.B(_01594_),
    .C(net633),
    .Y(_01631_),
    .A_N(_01593_));
 sg13g2_or3_1 _09064_ (.A(_01590_),
    .B(_01564_),
    .C(_01565_),
    .X(_01632_));
 sg13g2_a21oi_2 _09065_ (.B1(_01632_),
    .Y(_01633_),
    .A2(_01631_),
    .A1(_01630_));
 sg13g2_a21oi_2 _09066_ (.B1(_01633_),
    .Y(_01634_),
    .A2(_01629_),
    .A1(_01618_));
 sg13g2_nand2_1 _09067_ (.Y(_01635_),
    .A(_01628_),
    .B(_01634_));
 sg13g2_nor2_1 _09068_ (.A(net315),
    .B(_01635_),
    .Y(_01636_));
 sg13g2_a21o_1 _09069_ (.A2(_01636_),
    .A1(_01597_),
    .B1(_01633_),
    .X(_01637_));
 sg13g2_buf_1 _09070_ (.A(_01637_),
    .X(_01638_));
 sg13g2_buf_1 _09071_ (.A(_01638_),
    .X(_01639_));
 sg13g2_buf_1 _09072_ (.A(\soc_I.kianv_I.Instr[4] ),
    .X(_01640_));
 sg13g2_buf_8 _09073_ (.A(_01640_),
    .X(_01641_));
 sg13g2_buf_1 _09074_ (.A(\soc_I.kianv_I.Instr[3] ),
    .X(_01642_));
 sg13g2_nand3b_1 _09075_ (.B(\soc_I.kianv_I.Instr[1] ),
    .C(\soc_I.kianv_I.Instr[0] ),
    .Y(_01643_),
    .A_N(_01642_));
 sg13g2_buf_1 _09076_ (.A(_01643_),
    .X(_01644_));
 sg13g2_buf_1 _09077_ (.A(\soc_I.kianv_I.Instr[6] ),
    .X(_01645_));
 sg13g2_or2_1 _09078_ (.X(_01646_),
    .B(net629),
    .A(\soc_I.kianv_I.Instr[2] ));
 sg13g2_buf_1 _09079_ (.A(_01646_),
    .X(_01647_));
 sg13g2_or3_1 _09080_ (.A(net601),
    .B(net528),
    .C(_01647_),
    .X(_01648_));
 sg13g2_buf_8 _09081_ (.A(\soc_I.kianv_I.Instr[5] ),
    .X(_01649_));
 sg13g2_buf_8 _09082_ (.A(_01649_),
    .X(_01650_));
 sg13g2_nand2_1 _09083_ (.Y(_01651_),
    .A(net600),
    .B(net601));
 sg13g2_buf_8 _09084_ (.A(\soc_I.kianv_I.Instr[2] ),
    .X(_01652_));
 sg13g2_nor2b_1 _09085_ (.A(_01645_),
    .B_N(net628),
    .Y(_01653_));
 sg13g2_buf_1 _09086_ (.A(_00030_),
    .X(_01654_));
 sg13g2_mux2_1 _09087_ (.A0(net600),
    .A1(net601),
    .S(net627),
    .X(_01655_));
 sg13g2_o21ai_1 _09088_ (.B1(_01655_),
    .Y(_01656_),
    .A1(_01651_),
    .A2(_01653_));
 sg13g2_nor2_1 _09089_ (.A(net600),
    .B(_01652_),
    .Y(_01657_));
 sg13g2_nor2_1 _09090_ (.A(net601),
    .B(net629),
    .Y(_01658_));
 sg13g2_and2_1 _09091_ (.A(net601),
    .B(net627),
    .X(_01659_));
 sg13g2_or2_1 _09092_ (.X(_01660_),
    .B(_01659_),
    .A(_01658_));
 sg13g2_nor2b_1 _09093_ (.A(net601),
    .B_N(net600),
    .Y(_01661_));
 sg13g2_nor2b_1 _09094_ (.A(net627),
    .B_N(net628),
    .Y(_01662_));
 sg13g2_a21o_1 _09095_ (.A2(_01662_),
    .A1(_01661_),
    .B1(net528),
    .X(_01663_));
 sg13g2_a221oi_1 _09096_ (.B2(_01660_),
    .C1(_01663_),
    .B1(_01657_),
    .A1(_01648_),
    .Y(_01664_),
    .A2(_01656_));
 sg13g2_buf_2 _09097_ (.A(_01664_),
    .X(_01665_));
 sg13g2_buf_8 _09098_ (.A(_01665_),
    .X(_01666_));
 sg13g2_buf_1 _09099_ (.A(\soc_I.kianv_I.Instr[8] ),
    .X(_01667_));
 sg13g2_nand2b_1 _09100_ (.Y(_01668_),
    .B(_01649_),
    .A_N(_01640_));
 sg13g2_buf_1 _09101_ (.A(_01668_),
    .X(_01669_));
 sg13g2_and2_1 _09102_ (.A(net627),
    .B(net629),
    .X(_01670_));
 sg13g2_nor4_1 _09103_ (.A(net628),
    .B(net528),
    .C(_01669_),
    .D(_01670_),
    .Y(_01671_));
 sg13g2_buf_1 _09104_ (.A(_01671_),
    .X(_01672_));
 sg13g2_or4_1 _09105_ (.A(_01565_),
    .B(_01562_),
    .C(net632),
    .D(_01563_),
    .X(_01673_));
 sg13g2_buf_1 _09106_ (.A(_01673_),
    .X(_01674_));
 sg13g2_nor2_1 _09107_ (.A(_01599_),
    .B(_01674_),
    .Y(_01675_));
 sg13g2_buf_2 _09108_ (.A(_01675_),
    .X(_01676_));
 sg13g2_buf_8 _09109_ (.A(_01676_),
    .X(_01677_));
 sg13g2_a21oi_1 _09110_ (.A1(net626),
    .A2(net418),
    .Y(_01678_),
    .B1(_01677_));
 sg13g2_o21ai_1 _09111_ (.B1(_01678_),
    .Y(_01679_),
    .A1(_00034_),
    .A2(net342));
 sg13g2_buf_1 _09112_ (.A(net367),
    .X(_01680_));
 sg13g2_or2_1 _09113_ (.X(_01681_),
    .B(_01577_),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[0] ));
 sg13g2_buf_2 _09114_ (.A(_01681_),
    .X(_01682_));
 sg13g2_buf_1 _09115_ (.A(_01682_),
    .X(_01683_));
 sg13g2_a21oi_1 _09116_ (.A1(_00033_),
    .A2(_01680_),
    .Y(_01684_),
    .B1(net456));
 sg13g2_nand2_1 _09117_ (.Y(_01685_),
    .A(_01679_),
    .B(_01684_));
 sg13g2_buf_2 _09118_ (.A(_01685_),
    .X(_01686_));
 sg13g2_inv_1 _09119_ (.Y(_01687_),
    .A(_01686_));
 sg13g2_o21ai_1 _09120_ (.B1(_01657_),
    .Y(_01688_),
    .A1(_01658_),
    .A2(_01659_));
 sg13g2_nand2_2 _09121_ (.Y(_01689_),
    .A(_01661_),
    .B(_01662_));
 sg13g2_nand2_1 _09122_ (.Y(_01690_),
    .A(_01688_),
    .B(_01689_));
 sg13g2_buf_1 _09123_ (.A(_00026_),
    .X(_01691_));
 sg13g2_buf_1 _09124_ (.A(net528),
    .X(_01692_));
 sg13g2_or3_1 _09125_ (.A(_00035_),
    .B(net455),
    .C(_01682_),
    .X(_01693_));
 sg13g2_a21oi_1 _09126_ (.A1(_01691_),
    .A2(net341),
    .Y(_01694_),
    .B1(_01693_));
 sg13g2_nor4_1 _09127_ (.A(_01565_),
    .B(_01562_),
    .C(net632),
    .D(_01563_),
    .Y(_01695_));
 sg13g2_buf_2 _09128_ (.A(_01695_),
    .X(_01696_));
 sg13g2_buf_1 _09129_ (.A(_01696_),
    .X(_01697_));
 sg13g2_nor2_1 _09130_ (.A(_01590_),
    .B(_01593_),
    .Y(_01698_));
 sg13g2_buf_2 _09131_ (.A(_01698_),
    .X(_01699_));
 sg13g2_buf_1 _09132_ (.A(_01699_),
    .X(_01700_));
 sg13g2_and2_1 _09133_ (.A(_01691_),
    .B(net453),
    .X(_01701_));
 sg13g2_buf_1 _09134_ (.A(\soc_I.kianv_I.Instr[7] ),
    .X(_01702_));
 sg13g2_inv_1 _09135_ (.Y(_01703_),
    .A(net625));
 sg13g2_or4_1 _09136_ (.A(_01703_),
    .B(net455),
    .C(_01647_),
    .D(_01669_),
    .X(_01704_));
 sg13g2_nand2_1 _09137_ (.Y(_01705_),
    .A(_01699_),
    .B(_01696_));
 sg13g2_buf_2 _09138_ (.A(_01705_),
    .X(_01706_));
 sg13g2_buf_8 _09139_ (.A(_01706_),
    .X(_01707_));
 sg13g2_buf_1 _09140_ (.A(net366),
    .X(_01708_));
 sg13g2_a221oi_1 _09141_ (.B2(net340),
    .C1(net456),
    .B1(_01704_),
    .A1(net454),
    .Y(_01709_),
    .A2(_01701_));
 sg13g2_a21o_1 _09142_ (.A2(_01694_),
    .A1(_01690_),
    .B1(_01709_),
    .X(_01710_));
 sg13g2_buf_2 _09143_ (.A(_01710_),
    .X(_01711_));
 sg13g2_buf_1 _09144_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[0] ),
    .X(_01712_));
 sg13g2_mux2_1 _09145_ (.A0(\soc_I.PC[0] ),
    .A1(_01712_),
    .S(net369),
    .X(_01713_));
 sg13g2_mux2_1 _09146_ (.A0(\soc_I.kianv_I.datapath_unit_I.A1[0] ),
    .A1(_01713_),
    .S(net326),
    .X(_01714_));
 sg13g2_buf_2 _09147_ (.A(_01714_),
    .X(_01715_));
 sg13g2_and2_1 _09148_ (.A(_01711_),
    .B(_01715_),
    .X(_01716_));
 sg13g2_buf_1 _09149_ (.A(_01716_),
    .X(_01717_));
 sg13g2_a21oi_2 _09150_ (.B1(_01709_),
    .Y(_01718_),
    .A2(_01694_),
    .A1(_01690_));
 sg13g2_nor2_1 _09151_ (.A(_01718_),
    .B(_01715_),
    .Y(_01719_));
 sg13g2_and2_1 _09152_ (.A(_01612_),
    .B(net603),
    .X(_01720_));
 sg13g2_buf_2 _09153_ (.A(_01720_),
    .X(_01721_));
 sg13g2_nor2b_1 _09154_ (.A(net602),
    .B_N(net630),
    .Y(_01722_));
 sg13g2_nand2b_1 _09155_ (.Y(_01723_),
    .B(net603),
    .A_N(net631));
 sg13g2_a22oi_1 _09156_ (.Y(_01724_),
    .B1(_01722_),
    .B2(_01723_),
    .A2(_01721_),
    .A1(_01611_));
 sg13g2_buf_1 _09157_ (.A(_01724_),
    .X(_01725_));
 sg13g2_a21oi_1 _09158_ (.A1(net600),
    .A2(_00029_),
    .Y(_01726_),
    .B1(net631));
 sg13g2_nor2_1 _09159_ (.A(net603),
    .B(_01602_),
    .Y(_01727_));
 sg13g2_o21ai_1 _09160_ (.B1(_01727_),
    .Y(_01728_),
    .A1(_00027_),
    .A2(_01726_));
 sg13g2_inv_1 _09161_ (.Y(_01729_),
    .A(\soc_I.kianv_I.Instr[30] ));
 sg13g2_inv_1 _09162_ (.Y(_01730_),
    .A(net600));
 sg13g2_nor2_1 _09163_ (.A(_01729_),
    .B(_01730_),
    .Y(_01731_));
 sg13g2_o21ai_1 _09164_ (.B1(_01600_),
    .Y(_01732_),
    .A1(_01607_),
    .A2(_01731_));
 sg13g2_a221oi_1 _09165_ (.B2(_01628_),
    .C1(_01732_),
    .B1(_01634_),
    .A1(_01725_),
    .Y(_01733_),
    .A2(_01728_));
 sg13g2_buf_1 _09166_ (.A(_01733_),
    .X(_01734_));
 sg13g2_or3_1 _09167_ (.A(_01622_),
    .B(_01633_),
    .C(_01734_),
    .X(_01735_));
 sg13g2_buf_2 _09168_ (.A(_01735_),
    .X(_01736_));
 sg13g2_a21o_1 _09169_ (.A2(_01629_),
    .A1(_01618_),
    .B1(_01633_),
    .X(_01737_));
 sg13g2_buf_1 _09170_ (.A(_01737_),
    .X(_01738_));
 sg13g2_a21oi_1 _09171_ (.A1(net630),
    .A2(_01721_),
    .Y(_01739_),
    .B1(_01597_));
 sg13g2_a21oi_1 _09172_ (.A1(net315),
    .A2(_01738_),
    .Y(_01740_),
    .B1(_01739_));
 sg13g2_buf_2 _09173_ (.A(_01740_),
    .X(_01741_));
 sg13g2_a21oi_1 _09174_ (.A1(_01725_),
    .A2(_01728_),
    .Y(_01742_),
    .B1(_01732_));
 sg13g2_and2_1 _09175_ (.A(_01730_),
    .B(_01725_),
    .X(_01743_));
 sg13g2_o21ai_1 _09176_ (.B1(_01743_),
    .Y(_01744_),
    .A1(_00029_),
    .A2(_01665_));
 sg13g2_a21oi_1 _09177_ (.A1(_01608_),
    .A2(_01616_),
    .Y(_01745_),
    .B1(_01620_));
 sg13g2_buf_1 _09178_ (.A(_01745_),
    .X(_01746_));
 sg13g2_nor2_1 _09179_ (.A(_01590_),
    .B(_01567_),
    .Y(_01747_));
 sg13g2_nand2_1 _09180_ (.Y(_01748_),
    .A(_01630_),
    .B(_01631_));
 sg13g2_a21o_1 _09181_ (.A2(_01626_),
    .A1(net633),
    .B1(_01748_),
    .X(_01749_));
 sg13g2_a21o_1 _09182_ (.A2(_01749_),
    .A1(_01747_),
    .B1(_01739_),
    .X(_01750_));
 sg13g2_a221oi_1 _09183_ (.B2(_01738_),
    .C1(_01750_),
    .B1(_01746_),
    .A1(_01742_),
    .Y(_01751_),
    .A2(_01744_));
 sg13g2_buf_1 _09184_ (.A(_01751_),
    .X(_01752_));
 sg13g2_a21oi_1 _09185_ (.A1(_01736_),
    .A2(_01741_),
    .Y(_01753_),
    .B1(_01752_));
 sg13g2_buf_2 _09186_ (.A(_01753_),
    .X(_01754_));
 sg13g2_buf_8 _09187_ (.A(_01754_),
    .X(_01755_));
 sg13g2_buf_8 _09188_ (.A(net180),
    .X(_01756_));
 sg13g2_buf_8 _09189_ (.A(net171),
    .X(_01757_));
 sg13g2_buf_8 _09190_ (.A(net163),
    .X(_01758_));
 sg13g2_mux2_1 _09191_ (.A0(_01717_),
    .A1(_01719_),
    .S(_01758_),
    .X(_01759_));
 sg13g2_xnor2_1 _09192_ (.Y(_01760_),
    .A(_01687_),
    .B(_01759_));
 sg13g2_and2_1 _09193_ (.A(_01747_),
    .B(_01749_),
    .X(_01761_));
 sg13g2_buf_1 _09194_ (.A(_01761_),
    .X(_01762_));
 sg13g2_a21o_1 _09195_ (.A2(_01744_),
    .A1(_01742_),
    .B1(_01762_),
    .X(_01763_));
 sg13g2_buf_2 _09196_ (.A(_01763_),
    .X(_01764_));
 sg13g2_nor2_1 _09197_ (.A(_01764_),
    .B(_01686_),
    .Y(_01765_));
 sg13g2_inv_1 _09198_ (.Y(_01766_),
    .A(_01628_));
 sg13g2_nand2_1 _09199_ (.Y(_01767_),
    .A(_01766_),
    .B(net325));
 sg13g2_buf_1 _09200_ (.A(_01767_),
    .X(_01768_));
 sg13g2_and4_1 _09201_ (.A(_01628_),
    .B(_01597_),
    .C(_01623_),
    .D(_01634_),
    .X(_01769_));
 sg13g2_buf_1 _09202_ (.A(_01769_),
    .X(_01770_));
 sg13g2_buf_1 _09203_ (.A(_01770_),
    .X(_01771_));
 sg13g2_nor2_1 _09204_ (.A(net213),
    .B(_01765_),
    .Y(_01772_));
 sg13g2_a21oi_1 _09205_ (.A1(_01765_),
    .A2(net310),
    .Y(_01773_),
    .B1(_01772_));
 sg13g2_a21o_1 _09206_ (.A2(_01760_),
    .A1(net187),
    .B1(_01773_),
    .X(_01774_));
 sg13g2_a21oi_2 _09207_ (.B1(_01587_),
    .Y(_01775_),
    .A2(_01583_),
    .A1(_01572_));
 sg13g2_nand2_1 _09208_ (.Y(_01776_),
    .A(_01775_),
    .B(_01639_));
 sg13g2_buf_1 _09209_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[1] ),
    .X(_01777_));
 sg13g2_a21oi_1 _09210_ (.A1(_01742_),
    .A2(_01744_),
    .Y(_01778_),
    .B1(_01762_));
 sg13g2_buf_1 _09211_ (.A(_01778_),
    .X(_01779_));
 sg13g2_a21oi_1 _09212_ (.A1(_01779_),
    .A2(net325),
    .Y(_01780_),
    .B1(_01628_));
 sg13g2_buf_2 _09213_ (.A(_01780_),
    .X(_01781_));
 sg13g2_buf_1 _09214_ (.A(_01781_),
    .X(_01782_));
 sg13g2_nand4_1 _09215_ (.B(_01597_),
    .C(_01623_),
    .A(_01628_),
    .Y(_01783_),
    .D(_01634_));
 sg13g2_buf_1 _09216_ (.A(_01783_),
    .X(_01784_));
 sg13g2_buf_1 _09217_ (.A(_01784_),
    .X(_01785_));
 sg13g2_buf_1 _09218_ (.A(net212),
    .X(_01786_));
 sg13g2_buf_1 _09219_ (.A(_01619_),
    .X(_01787_));
 sg13g2_o21ai_1 _09220_ (.B1(_01787_),
    .Y(_01788_),
    .A1(_01589_),
    .A2(net185));
 sg13g2_a22oi_1 _09221_ (.Y(_01789_),
    .B1(_01687_),
    .B2(_01788_),
    .A2(net186),
    .A1(_01777_));
 sg13g2_o21ai_1 _09222_ (.B1(_01789_),
    .Y(_01790_),
    .A1(_01760_),
    .A2(_01776_));
 sg13g2_a21oi_2 _09223_ (.B1(_01790_),
    .Y(_01791_),
    .A2(_01774_),
    .A1(_01589_));
 sg13g2_buf_2 _09224_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[2] ),
    .X(_01792_));
 sg13g2_buf_1 _09225_ (.A(_01792_),
    .X(_01793_));
 sg13g2_nor2b_1 _09226_ (.A(net599),
    .B_N(\soc_I.kianv_I.datapath_unit_I.ALUOut[1] ),
    .Y(_01794_));
 sg13g2_a21oi_1 _09227_ (.A1(net599),
    .A2(\soc_I.kianv_I.datapath_unit_I.DataLatched[1] ),
    .Y(_01795_),
    .B1(_01794_));
 sg13g2_buf_1 _09228_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[0] ),
    .X(_01796_));
 sg13g2_inv_1 _09229_ (.Y(_01797_),
    .A(net624));
 sg13g2_buf_1 _09230_ (.A(_01797_),
    .X(_01798_));
 sg13g2_mux2_1 _09231_ (.A0(_01791_),
    .A1(_01795_),
    .S(net527),
    .X(_01799_));
 sg13g2_buf_1 _09232_ (.A(_01799_),
    .X(_01800_));
 sg13g2_nand2_1 _09233_ (.Y(_01801_),
    .A(_01573_),
    .B(net457));
 sg13g2_o21ai_1 _09234_ (.B1(_01801_),
    .Y(_01802_),
    .A1(net457),
    .A2(_01800_));
 sg13g2_buf_1 _09235_ (.A(_01802_),
    .X(\soc_I.cpu_mem_addr[1] ));
 sg13g2_buf_8 _09236_ (.A(_01754_),
    .X(_01803_));
 sg13g2_buf_8 _09237_ (.A(net179),
    .X(_01804_));
 sg13g2_nor2_1 _09238_ (.A(_01796_),
    .B(_01577_),
    .Y(_01805_));
 sg13g2_buf_1 _09239_ (.A(_01805_),
    .X(_01806_));
 sg13g2_buf_1 _09240_ (.A(_01806_),
    .X(_01807_));
 sg13g2_buf_1 _09241_ (.A(net451),
    .X(_01808_));
 sg13g2_o21ai_1 _09242_ (.B1(net417),
    .Y(_01809_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[15] ),
    .A2(net340));
 sg13g2_buf_1 _09243_ (.A(_01809_),
    .X(_01810_));
 sg13g2_nand3b_1 _09244_ (.B(_01640_),
    .C(net627),
    .Y(_01811_),
    .A_N(_01649_));
 sg13g2_or2_1 _09245_ (.X(_01812_),
    .B(_01811_),
    .A(net628));
 sg13g2_buf_1 _09246_ (.A(_01812_),
    .X(_01813_));
 sg13g2_nand2b_1 _09247_ (.Y(_01814_),
    .B(_01649_),
    .A_N(_01654_));
 sg13g2_a21o_1 _09248_ (.A2(_01814_),
    .A1(_01647_),
    .B1(net601),
    .X(_01815_));
 sg13g2_buf_1 _09249_ (.A(_01815_),
    .X(_01816_));
 sg13g2_a21o_1 _09250_ (.A2(_01816_),
    .A1(_01813_),
    .B1(net528),
    .X(_01817_));
 sg13g2_buf_1 _09251_ (.A(_01817_),
    .X(_01818_));
 sg13g2_buf_1 _09252_ (.A(\soc_I.kianv_I.Instr[31] ),
    .X(_01819_));
 sg13g2_inv_1 _09253_ (.Y(_01820_),
    .A(net623));
 sg13g2_or2_1 _09254_ (.X(_01821_),
    .B(net528),
    .A(_01820_));
 sg13g2_a21oi_1 _09255_ (.A1(_01813_),
    .A2(_01816_),
    .Y(_01822_),
    .B1(_01821_));
 sg13g2_buf_2 _09256_ (.A(_01822_),
    .X(_01823_));
 sg13g2_a221oi_1 _09257_ (.B2(\soc_I.kianv_I.Instr[15] ),
    .C1(_01823_),
    .B1(net339),
    .A1(net453),
    .Y(_01824_),
    .A2(net454));
 sg13g2_buf_1 _09258_ (.A(_01824_),
    .X(_01825_));
 sg13g2_buf_1 _09259_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[15] ),
    .X(_01826_));
 sg13g2_mux2_1 _09260_ (.A0(\soc_I.PC[15] ),
    .A1(_01826_),
    .S(net420),
    .X(_01827_));
 sg13g2_buf_1 _09261_ (.A(net419),
    .X(_01828_));
 sg13g2_and2_1 _09262_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[15] ),
    .B(net365),
    .X(_01829_));
 sg13g2_a21o_1 _09263_ (.A2(_01827_),
    .A1(net343),
    .B1(_01829_),
    .X(_01830_));
 sg13g2_buf_2 _09264_ (.A(_01830_),
    .X(_01831_));
 sg13g2_o21ai_1 _09265_ (.B1(_01831_),
    .Y(_01832_),
    .A1(_01810_),
    .A2(_01825_));
 sg13g2_buf_2 _09266_ (.A(_01832_),
    .X(_01833_));
 sg13g2_or3_1 _09267_ (.A(_01810_),
    .B(_01825_),
    .C(_01831_),
    .X(_01834_));
 sg13g2_buf_2 _09268_ (.A(_01834_),
    .X(_01835_));
 sg13g2_and2_1 _09269_ (.A(_01833_),
    .B(_01835_),
    .X(_01836_));
 sg13g2_buf_1 _09270_ (.A(_01836_),
    .X(_01837_));
 sg13g2_nor2_1 _09271_ (.A(_01820_),
    .B(net455),
    .Y(_01838_));
 sg13g2_nand2_1 _09272_ (.Y(_01839_),
    .A(_01813_),
    .B(_01816_));
 sg13g2_inv_1 _09273_ (.Y(_01840_),
    .A(net630));
 sg13g2_nor2_2 _09274_ (.A(_01649_),
    .B(net627),
    .Y(_01841_));
 sg13g2_nand2_1 _09275_ (.Y(_01842_),
    .A(_01640_),
    .B(net628));
 sg13g2_and2_1 _09276_ (.A(_01649_),
    .B(net629),
    .X(_01843_));
 sg13g2_buf_1 _09277_ (.A(_01843_),
    .X(_01844_));
 sg13g2_nor4_2 _09278_ (.A(net528),
    .B(_01841_),
    .C(_01842_),
    .Y(_01845_),
    .D(_01844_));
 sg13g2_buf_1 _09279_ (.A(_01845_),
    .X(_01846_));
 sg13g2_nor2_1 _09280_ (.A(_01840_),
    .B(_01846_),
    .Y(_01847_));
 sg13g2_or4_1 _09281_ (.A(net528),
    .B(_01841_),
    .C(_01842_),
    .D(_01844_),
    .X(_01848_));
 sg13g2_buf_2 _09282_ (.A(_01848_),
    .X(_01849_));
 sg13g2_buf_1 _09283_ (.A(_01706_),
    .X(_01850_));
 sg13g2_o21ai_1 _09284_ (.B1(_01850_),
    .Y(_01851_),
    .A1(_00027_),
    .A2(_01849_));
 sg13g2_a221oi_1 _09285_ (.B2(_01847_),
    .C1(_01851_),
    .B1(net339),
    .A1(_01838_),
    .Y(_01852_),
    .A2(_01839_));
 sg13g2_buf_2 _09286_ (.A(_01852_),
    .X(_01853_));
 sg13g2_nand2b_1 _09287_ (.Y(_01854_),
    .B(_01820_),
    .A_N(net455));
 sg13g2_a221oi_1 _09288_ (.B2(_01699_),
    .C1(_01854_),
    .B1(_01696_),
    .A1(_01688_),
    .Y(_01855_),
    .A2(_01689_));
 sg13g2_buf_1 _09289_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[12] ),
    .X(_01856_));
 sg13g2_o21ai_1 _09290_ (.B1(net451),
    .Y(_01857_),
    .A1(_01856_),
    .A2(net364));
 sg13g2_or2_1 _09291_ (.X(_01858_),
    .B(_01857_),
    .A(_01855_));
 sg13g2_buf_1 _09292_ (.A(_01858_),
    .X(_01859_));
 sg13g2_nor2_1 _09293_ (.A(net632),
    .B(_01577_),
    .Y(_01860_));
 sg13g2_buf_8 _09294_ (.A(_01860_),
    .X(_01861_));
 sg13g2_nand2_2 _09295_ (.Y(_01862_),
    .A(_01574_),
    .B(_01861_));
 sg13g2_buf_1 _09296_ (.A(_01575_),
    .X(_01863_));
 sg13g2_buf_1 _09297_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[12] ),
    .X(_01864_));
 sg13g2_inv_1 _09298_ (.Y(_01865_),
    .A(_01864_));
 sg13g2_buf_1 _09299_ (.A(_01579_),
    .X(_01866_));
 sg13g2_nor3_1 _09300_ (.A(net526),
    .B(_01865_),
    .C(net450),
    .Y(_01867_));
 sg13g2_a21oi_1 _09301_ (.A1(\soc_I.PC[12] ),
    .A2(_01862_),
    .Y(_01868_),
    .B1(_01867_));
 sg13g2_nor2_1 _09302_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[12] ),
    .B(net370),
    .Y(_01869_));
 sg13g2_a21oi_1 _09303_ (.A1(net343),
    .A2(_01868_),
    .Y(_01870_),
    .B1(_01869_));
 sg13g2_buf_1 _09304_ (.A(_01870_),
    .X(_01871_));
 sg13g2_o21ai_1 _09305_ (.B1(_01871_),
    .Y(_01872_),
    .A1(_01853_),
    .A2(_01859_));
 sg13g2_buf_2 _09306_ (.A(_01872_),
    .X(_01873_));
 sg13g2_or3_1 _09307_ (.A(_01871_),
    .B(_01853_),
    .C(_01859_),
    .X(_01874_));
 sg13g2_buf_1 _09308_ (.A(_01874_),
    .X(_01875_));
 sg13g2_and2_1 _09309_ (.A(_01873_),
    .B(_01875_),
    .X(_01876_));
 sg13g2_buf_2 _09310_ (.A(_01876_),
    .X(_01877_));
 sg13g2_o21ai_1 _09311_ (.B1(net451),
    .Y(_01878_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[14] ),
    .A2(net364));
 sg13g2_buf_1 _09312_ (.A(_01878_),
    .X(_01879_));
 sg13g2_a221oi_1 _09313_ (.B2(net602),
    .C1(_01823_),
    .B1(_01818_),
    .A1(_01699_),
    .Y(_01880_),
    .A2(_01697_));
 sg13g2_buf_2 _09314_ (.A(_01880_),
    .X(_01881_));
 sg13g2_nand2b_1 _09315_ (.Y(_01882_),
    .B(net419),
    .A_N(\soc_I.kianv_I.datapath_unit_I.A1[14] ));
 sg13g2_buf_1 _09316_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[14] ),
    .X(_01883_));
 sg13g2_nand3_1 _09317_ (.B(_01883_),
    .C(_01861_),
    .A(_01574_),
    .Y(_01884_));
 sg13g2_o21ai_1 _09318_ (.B1(\soc_I.PC[14] ),
    .Y(_01885_),
    .A1(_01575_),
    .A2(net450));
 sg13g2_nand3_1 _09319_ (.B(_01884_),
    .C(_01885_),
    .A(_01569_),
    .Y(_01886_));
 sg13g2_buf_1 _09320_ (.A(_01886_),
    .X(_01887_));
 sg13g2_and2_1 _09321_ (.A(_01882_),
    .B(_01887_),
    .X(_01888_));
 sg13g2_buf_2 _09322_ (.A(_01888_),
    .X(_01889_));
 sg13g2_o21ai_1 _09323_ (.B1(_01889_),
    .Y(_01890_),
    .A1(_01879_),
    .A2(_01881_));
 sg13g2_buf_2 _09324_ (.A(_01890_),
    .X(_01891_));
 sg13g2_nand2_1 _09325_ (.Y(_01892_),
    .A(_01882_),
    .B(_01887_));
 sg13g2_inv_1 _09326_ (.Y(_01893_),
    .A(\soc_I.kianv_I.datapath_unit_I.A2[14] ));
 sg13g2_a21oi_1 _09327_ (.A1(_01893_),
    .A2(net341),
    .Y(_01894_),
    .B1(_01683_));
 sg13g2_nand3b_1 _09328_ (.B(_01892_),
    .C(_01894_),
    .Y(_01895_),
    .A_N(_01881_));
 sg13g2_buf_2 _09329_ (.A(_01895_),
    .X(_01896_));
 sg13g2_o21ai_1 _09330_ (.B1(net451),
    .Y(_01897_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[13] ),
    .A2(net364));
 sg13g2_buf_1 _09331_ (.A(_01897_),
    .X(_01898_));
 sg13g2_a221oi_1 _09332_ (.B2(net603),
    .C1(_01823_),
    .B1(_01818_),
    .A1(net453),
    .Y(_01899_),
    .A2(_01697_));
 sg13g2_buf_2 _09333_ (.A(_01899_),
    .X(_01900_));
 sg13g2_nor2_1 _09334_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[13] ),
    .B(net370),
    .Y(_01901_));
 sg13g2_buf_1 _09335_ (.A(_01574_),
    .X(_01902_));
 sg13g2_buf_1 _09336_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[13] ),
    .X(_01903_));
 sg13g2_buf_1 _09337_ (.A(_01861_),
    .X(_01904_));
 sg13g2_nand3_1 _09338_ (.B(_01903_),
    .C(_01904_),
    .A(net598),
    .Y(_01905_));
 sg13g2_o21ai_1 _09339_ (.B1(\soc_I.PC[13] ),
    .Y(_01906_),
    .A1(net526),
    .A2(net450));
 sg13g2_nand3_1 _09340_ (.B(_01905_),
    .C(_01906_),
    .A(net370),
    .Y(_01907_));
 sg13g2_nor2b_2 _09341_ (.A(_01901_),
    .B_N(_01907_),
    .Y(_01908_));
 sg13g2_o21ai_1 _09342_ (.B1(_01908_),
    .Y(_01909_),
    .A1(_01898_),
    .A2(_01900_));
 sg13g2_buf_2 _09343_ (.A(_01909_),
    .X(_01910_));
 sg13g2_or3_1 _09344_ (.A(_01898_),
    .B(_01900_),
    .C(_01908_),
    .X(_01911_));
 sg13g2_buf_2 _09345_ (.A(_01911_),
    .X(_01912_));
 sg13g2_and4_1 _09346_ (.A(_01891_),
    .B(_01896_),
    .C(_01910_),
    .D(_01912_),
    .X(_01913_));
 sg13g2_buf_1 _09347_ (.A(_01913_),
    .X(_01914_));
 sg13g2_nand4_1 _09348_ (.B(_01837_),
    .C(_01877_),
    .A(net170),
    .Y(_01915_),
    .D(_01914_));
 sg13g2_a21o_1 _09349_ (.A2(_01741_),
    .A1(_01736_),
    .B1(_01752_),
    .X(_01916_));
 sg13g2_buf_8 _09350_ (.A(_01916_),
    .X(_01917_));
 sg13g2_buf_8 _09351_ (.A(_01917_),
    .X(_01918_));
 sg13g2_buf_8 _09352_ (.A(net178),
    .X(_01919_));
 sg13g2_buf_8 _09353_ (.A(net169),
    .X(_01920_));
 sg13g2_nand2_1 _09354_ (.Y(_01921_),
    .A(_01833_),
    .B(_01835_));
 sg13g2_nand2_1 _09355_ (.Y(_01922_),
    .A(_01873_),
    .B(_01875_));
 sg13g2_a22oi_1 _09356_ (.Y(_01923_),
    .B1(_01910_),
    .B2(_01912_),
    .A2(_01896_),
    .A1(_01891_));
 sg13g2_nand4_1 _09357_ (.B(_01921_),
    .C(_01922_),
    .A(net162),
    .Y(_01924_),
    .D(_01923_));
 sg13g2_nand2_1 _09358_ (.Y(_01925_),
    .A(_01915_),
    .B(_01924_));
 sg13g2_buf_8 _09359_ (.A(net162),
    .X(_01926_));
 sg13g2_buf_1 _09360_ (.A(net417),
    .X(_01927_));
 sg13g2_nand2b_1 _09361_ (.Y(_01928_),
    .B(net365),
    .A_N(\soc_I.kianv_I.datapath_unit_I.A1[8] ));
 sg13g2_buf_2 _09362_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[8] ),
    .X(_01929_));
 sg13g2_and3_1 _09363_ (.X(_01930_),
    .A(_01574_),
    .B(_01929_),
    .C(_01861_));
 sg13g2_inv_1 _09364_ (.Y(_01931_),
    .A(\soc_I.PC[8] ));
 sg13g2_a21oi_1 _09365_ (.A1(_01574_),
    .A2(_01861_),
    .Y(_01932_),
    .B1(_01931_));
 sg13g2_or3_1 _09366_ (.A(net419),
    .B(_01930_),
    .C(_01932_),
    .X(_01933_));
 sg13g2_buf_1 _09367_ (.A(\soc_I.kianv_I.Instr[28] ),
    .X(_01934_));
 sg13g2_o21ai_1 _09368_ (.B1(_01934_),
    .Y(_01935_),
    .A1(_01599_),
    .A2(_01674_));
 sg13g2_buf_1 _09369_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[8] ),
    .X(_01936_));
 sg13g2_nand3_1 _09370_ (.B(_01699_),
    .C(_01696_),
    .A(_01936_),
    .Y(_01937_));
 sg13g2_o21ai_1 _09371_ (.B1(_01937_),
    .Y(_01938_),
    .A1(_01845_),
    .A2(_01935_));
 sg13g2_nand3_1 _09372_ (.B(_01933_),
    .C(_01938_),
    .A(_01928_),
    .Y(_01939_));
 sg13g2_buf_1 _09373_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[9] ),
    .X(_01940_));
 sg13g2_buf_8 _09374_ (.A(net368),
    .X(_01941_));
 sg13g2_nand2b_1 _09375_ (.Y(_01942_),
    .B(net338),
    .A_N(_01940_));
 sg13g2_buf_2 _09376_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[9] ),
    .X(_01943_));
 sg13g2_and3_1 _09377_ (.X(_01944_),
    .A(_01574_),
    .B(_01943_),
    .C(_01861_));
 sg13g2_buf_1 _09378_ (.A(_01944_),
    .X(_01945_));
 sg13g2_inv_1 _09379_ (.Y(_01946_),
    .A(\soc_I.PC[9] ));
 sg13g2_a21oi_1 _09380_ (.A1(net598),
    .A2(net449),
    .Y(_01947_),
    .B1(_01946_));
 sg13g2_or3_1 _09381_ (.A(_01586_),
    .B(_01945_),
    .C(_01947_),
    .X(_01948_));
 sg13g2_buf_1 _09382_ (.A(_01948_),
    .X(_01949_));
 sg13g2_buf_1 _09383_ (.A(\soc_I.kianv_I.Instr[29] ),
    .X(_01950_));
 sg13g2_o21ai_1 _09384_ (.B1(_01950_),
    .Y(_01951_),
    .A1(_01599_),
    .A2(_01674_));
 sg13g2_buf_2 _09385_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[9] ),
    .X(_01952_));
 sg13g2_nand3_1 _09386_ (.B(_01699_),
    .C(_01696_),
    .A(_01952_),
    .Y(_01953_));
 sg13g2_o21ai_1 _09387_ (.B1(_01953_),
    .Y(_01954_),
    .A1(_01845_),
    .A2(_01951_));
 sg13g2_buf_2 _09388_ (.A(_01954_),
    .X(_01955_));
 sg13g2_a21oi_1 _09389_ (.A1(_01942_),
    .A2(_01949_),
    .Y(_01956_),
    .B1(_01955_));
 sg13g2_nand3_1 _09390_ (.B(_01949_),
    .C(_01955_),
    .A(_01942_),
    .Y(_01957_));
 sg13g2_o21ai_1 _09391_ (.B1(_01957_),
    .Y(_01958_),
    .A1(_01939_),
    .A2(_01956_));
 sg13g2_buf_1 _09392_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[10] ),
    .X(_01959_));
 sg13g2_mux2_1 _09393_ (.A0(\soc_I.PC[10] ),
    .A1(_01959_),
    .S(net420),
    .X(_01960_));
 sg13g2_and2_1 _09394_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[10] ),
    .B(net365),
    .X(_01961_));
 sg13g2_a21o_1 _09395_ (.A2(_01960_),
    .A1(net326),
    .B1(_01961_),
    .X(_01962_));
 sg13g2_buf_1 _09396_ (.A(_01962_),
    .X(_01963_));
 sg13g2_or2_1 _09397_ (.X(_01964_),
    .B(_01656_),
    .A(_01692_));
 sg13g2_nor3_2 _09398_ (.A(_01641_),
    .B(_01644_),
    .C(_01647_),
    .Y(_01965_));
 sg13g2_nor2_1 _09399_ (.A(_00035_),
    .B(_01965_),
    .Y(_01966_));
 sg13g2_nor3_1 _09400_ (.A(net628),
    .B(net455),
    .C(_01669_),
    .Y(_01967_));
 sg13g2_nand2b_1 _09401_ (.Y(_01968_),
    .B(net625),
    .A_N(_01654_));
 sg13g2_nand2b_1 _09402_ (.Y(_01969_),
    .B(net623),
    .A_N(net629));
 sg13g2_o21ai_1 _09403_ (.B1(_01969_),
    .Y(_01970_),
    .A1(_01658_),
    .A2(_01968_));
 sg13g2_a21o_1 _09404_ (.A2(_01970_),
    .A1(_01967_),
    .B1(_01677_),
    .X(_01971_));
 sg13g2_a221oi_1 _09405_ (.B2(_01966_),
    .C1(_01971_),
    .B1(_01964_),
    .A1(_01690_),
    .Y(_01972_),
    .A2(_01838_));
 sg13g2_buf_2 _09406_ (.A(_01972_),
    .X(_01973_));
 sg13g2_o21ai_1 _09407_ (.B1(net451),
    .Y(_01974_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[11] ),
    .A2(net366));
 sg13g2_or2_1 _09408_ (.X(_01975_),
    .B(_01974_),
    .A(_01855_));
 sg13g2_buf_2 _09409_ (.A(_01975_),
    .X(_01976_));
 sg13g2_buf_8 _09410_ (.A(net370),
    .X(_01977_));
 sg13g2_buf_8 _09411_ (.A(net337),
    .X(_01978_));
 sg13g2_buf_1 _09412_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[11] ),
    .X(_01979_));
 sg13g2_and3_1 _09413_ (.X(_01980_),
    .A(net598),
    .B(_01979_),
    .C(net449));
 sg13g2_a21oi_1 _09414_ (.A1(\soc_I.PC[11] ),
    .A2(_01862_),
    .Y(_01981_),
    .B1(_01980_));
 sg13g2_nor2_1 _09415_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[11] ),
    .B(net337),
    .Y(_01982_));
 sg13g2_a21o_1 _09416_ (.A2(_01981_),
    .A1(_01978_),
    .B1(_01982_),
    .X(_01983_));
 sg13g2_buf_2 _09417_ (.A(_01983_),
    .X(_01984_));
 sg13g2_o21ai_1 _09418_ (.B1(_01984_),
    .Y(_01985_),
    .A1(_01973_),
    .A2(_01976_));
 sg13g2_buf_1 _09419_ (.A(_01985_),
    .X(_01986_));
 sg13g2_nand4_1 _09420_ (.B(_01958_),
    .C(_01963_),
    .A(_01927_),
    .Y(_01987_),
    .D(_01986_));
 sg13g2_nor2_1 _09421_ (.A(_00046_),
    .B(net364),
    .Y(_01988_));
 sg13g2_and3_1 _09422_ (.X(_01989_),
    .A(\soc_I.kianv_I.Instr[30] ),
    .B(net364),
    .C(net418));
 sg13g2_o21ai_1 _09423_ (.B1(net417),
    .Y(_01990_),
    .A1(_01988_),
    .A2(_01989_));
 sg13g2_buf_2 _09424_ (.A(_01990_),
    .X(_01991_));
 sg13g2_a21oi_1 _09425_ (.A1(_00046_),
    .A2(net367),
    .Y(_01992_),
    .B1(_00029_));
 sg13g2_nand3b_1 _09426_ (.B(net417),
    .C(_01992_),
    .Y(_01993_),
    .A_N(net342));
 sg13g2_buf_2 _09427_ (.A(_01993_),
    .X(_01994_));
 sg13g2_nand2_2 _09428_ (.Y(_01995_),
    .A(_01991_),
    .B(_01994_));
 sg13g2_nand4_1 _09429_ (.B(_01958_),
    .C(_01995_),
    .A(net363),
    .Y(_01996_),
    .D(_01986_));
 sg13g2_a21oi_1 _09430_ (.A1(_01571_),
    .A2(_01960_),
    .Y(_01997_),
    .B1(_01961_));
 sg13g2_buf_2 _09431_ (.A(_01997_),
    .X(_01998_));
 sg13g2_a21oi_1 _09432_ (.A1(_01991_),
    .A2(_01994_),
    .Y(_01999_),
    .B1(_01998_));
 sg13g2_nor3_2 _09433_ (.A(_01984_),
    .B(_01973_),
    .C(_01976_),
    .Y(_02000_));
 sg13g2_a21oi_1 _09434_ (.A1(_01986_),
    .A2(_01999_),
    .Y(_02001_),
    .B1(_02000_));
 sg13g2_and3_1 _09435_ (.X(_02002_),
    .A(_01987_),
    .B(_01996_),
    .C(_02001_));
 sg13g2_nor2_1 _09436_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[8] ),
    .B(_01940_),
    .Y(_02003_));
 sg13g2_a21oi_1 _09437_ (.A1(net338),
    .A2(_02003_),
    .Y(_02004_),
    .B1(_01808_));
 sg13g2_nor3_1 _09438_ (.A(_01929_),
    .B(_01943_),
    .C(_01862_),
    .Y(_02005_));
 sg13g2_nor3_1 _09439_ (.A(\soc_I.PC[8] ),
    .B(\soc_I.PC[9] ),
    .C(net369),
    .Y(_02006_));
 sg13g2_buf_8 _09440_ (.A(net324),
    .X(_02007_));
 sg13g2_o21ai_1 _09441_ (.B1(net314),
    .Y(_02008_),
    .A1(_02005_),
    .A2(_02006_));
 sg13g2_nor2_1 _09442_ (.A(_01940_),
    .B(net370),
    .Y(_02009_));
 sg13g2_nor3_1 _09443_ (.A(net419),
    .B(_01945_),
    .C(_01947_),
    .Y(_02010_));
 sg13g2_o21ai_1 _09444_ (.B1(_01955_),
    .Y(_02011_),
    .A1(_02009_),
    .A2(_02010_));
 sg13g2_nand2_1 _09445_ (.Y(_02012_),
    .A(\soc_I.kianv_I.datapath_unit_I.A1[8] ),
    .B(net365));
 sg13g2_o21ai_1 _09446_ (.B1(_01569_),
    .Y(_02013_),
    .A1(_01930_),
    .A2(_01932_));
 sg13g2_buf_1 _09447_ (.A(_02013_),
    .X(_02014_));
 sg13g2_a21oi_1 _09448_ (.A1(_02012_),
    .A2(_02014_),
    .Y(_02015_),
    .B1(_01938_));
 sg13g2_nor3_1 _09449_ (.A(_02009_),
    .B(_02010_),
    .C(_01955_),
    .Y(_02016_));
 sg13g2_a221oi_1 _09450_ (.B2(_02015_),
    .C1(_02016_),
    .B1(_02011_),
    .A1(_02004_),
    .Y(_02017_),
    .A2(_02008_));
 sg13g2_buf_1 _09451_ (.A(_02017_),
    .X(_02018_));
 sg13g2_a21oi_1 _09452_ (.A1(_01995_),
    .A2(_02018_),
    .Y(_02019_),
    .B1(_01998_));
 sg13g2_nor2_1 _09453_ (.A(_01995_),
    .B(_02018_),
    .Y(_02020_));
 sg13g2_a21oi_1 _09454_ (.A1(_01978_),
    .A2(_01981_),
    .Y(_02021_),
    .B1(_01982_));
 sg13g2_or3_1 _09455_ (.A(_02021_),
    .B(_01973_),
    .C(_01976_),
    .X(_02022_));
 sg13g2_buf_1 _09456_ (.A(_02022_),
    .X(_02023_));
 sg13g2_o21ai_1 _09457_ (.B1(_02023_),
    .Y(_02024_),
    .A1(_02019_),
    .A2(_02020_));
 sg13g2_o21ai_1 _09458_ (.B1(_02021_),
    .Y(_02025_),
    .A1(_01973_),
    .A2(_01976_));
 sg13g2_buf_2 _09459_ (.A(_02025_),
    .X(_02026_));
 sg13g2_and2_1 _09460_ (.A(net163),
    .B(_02026_),
    .X(_02027_));
 sg13g2_a22oi_1 _09461_ (.Y(_02028_),
    .B1(_02024_),
    .B2(_02027_),
    .A2(_02002_),
    .A1(net157));
 sg13g2_buf_1 _09462_ (.A(_02028_),
    .X(_02029_));
 sg13g2_buf_8 _09463_ (.A(net178),
    .X(_02030_));
 sg13g2_buf_2 _09464_ (.A(\soc_I.kianv_I.Instr[21] ),
    .X(_02031_));
 sg13g2_nand2_1 _09465_ (.Y(_02032_),
    .A(_02031_),
    .B(net416));
 sg13g2_a21oi_1 _09466_ (.A1(net623),
    .A2(_01849_),
    .Y(_02033_),
    .B1(_01676_));
 sg13g2_buf_1 _09467_ (.A(_02033_),
    .X(_02034_));
 sg13g2_buf_1 _09468_ (.A(_01806_),
    .X(_02035_));
 sg13g2_o21ai_1 _09469_ (.B1(net448),
    .Y(_02036_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[21] ),
    .A2(net366));
 sg13g2_a21oi_1 _09470_ (.A1(_02032_),
    .A2(_02034_),
    .Y(_02037_),
    .B1(_02036_));
 sg13g2_buf_2 _09471_ (.A(_02037_),
    .X(_02038_));
 sg13g2_buf_1 _09472_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[21] ),
    .X(_02039_));
 sg13g2_mux2_1 _09473_ (.A0(\soc_I.PC[21] ),
    .A1(_02039_),
    .S(net420),
    .X(_02040_));
 sg13g2_mux2_1 _09474_ (.A0(\soc_I.kianv_I.datapath_unit_I.A1[21] ),
    .A1(_02040_),
    .S(net337),
    .X(_02041_));
 sg13g2_buf_2 _09475_ (.A(_02041_),
    .X(_02042_));
 sg13g2_xnor2_1 _09476_ (.Y(_02043_),
    .A(_02038_),
    .B(_02042_));
 sg13g2_buf_1 _09477_ (.A(_02043_),
    .X(_02044_));
 sg13g2_nand2_1 _09478_ (.Y(_02045_),
    .A(\soc_I.kianv_I.Instr[20] ),
    .B(net416));
 sg13g2_o21ai_1 _09479_ (.B1(net448),
    .Y(_02046_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[20] ),
    .A2(net366));
 sg13g2_a21o_1 _09480_ (.A2(_02045_),
    .A1(_02034_),
    .B1(_02046_),
    .X(_02047_));
 sg13g2_buf_2 _09481_ (.A(_02047_),
    .X(_02048_));
 sg13g2_buf_2 _09482_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[20] ),
    .X(_02049_));
 sg13g2_and3_1 _09483_ (.X(_02050_),
    .A(net598),
    .B(_02049_),
    .C(net449));
 sg13g2_a21oi_1 _09484_ (.A1(\soc_I.PC[20] ),
    .A2(_01862_),
    .Y(_02051_),
    .B1(_02050_));
 sg13g2_nor2_1 _09485_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[20] ),
    .B(net370),
    .Y(_02052_));
 sg13g2_a21o_1 _09486_ (.A2(_02051_),
    .A1(net337),
    .B1(_02052_),
    .X(_02053_));
 sg13g2_buf_2 _09487_ (.A(_02053_),
    .X(_02054_));
 sg13g2_xnor2_1 _09488_ (.Y(_02055_),
    .A(_02048_),
    .B(_02054_));
 sg13g2_buf_2 _09489_ (.A(_02055_),
    .X(_02056_));
 sg13g2_nor2_1 _09490_ (.A(net272),
    .B(_02056_),
    .Y(_02057_));
 sg13g2_buf_1 _09491_ (.A(\soc_I.kianv_I.Instr[22] ),
    .X(_02058_));
 sg13g2_nand2_1 _09492_ (.Y(_02059_),
    .A(net622),
    .B(net416));
 sg13g2_o21ai_1 _09493_ (.B1(net448),
    .Y(_02060_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[22] ),
    .A2(net366));
 sg13g2_a21oi_1 _09494_ (.A1(_02034_),
    .A2(_02059_),
    .Y(_02061_),
    .B1(_02060_));
 sg13g2_buf_2 _09495_ (.A(_02061_),
    .X(_02062_));
 sg13g2_o21ai_1 _09496_ (.B1(\soc_I.PC[22] ),
    .Y(_02063_),
    .A1(net526),
    .A2(net450));
 sg13g2_buf_2 _09497_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[22] ),
    .X(_02064_));
 sg13g2_nand3_1 _09498_ (.B(_02064_),
    .C(net449),
    .A(net598),
    .Y(_02065_));
 sg13g2_nand3_1 _09499_ (.B(_02063_),
    .C(_02065_),
    .A(net337),
    .Y(_02066_));
 sg13g2_buf_1 _09500_ (.A(_02066_),
    .X(_02067_));
 sg13g2_nand2b_1 _09501_ (.Y(_02068_),
    .B(net368),
    .A_N(\soc_I.kianv_I.datapath_unit_I.A1[22] ));
 sg13g2_and2_1 _09502_ (.A(_02067_),
    .B(_02068_),
    .X(_02069_));
 sg13g2_buf_2 _09503_ (.A(_02069_),
    .X(_02070_));
 sg13g2_xnor2_1 _09504_ (.Y(_02071_),
    .A(_02062_),
    .B(_02070_));
 sg13g2_buf_2 _09505_ (.A(_02071_),
    .X(_02072_));
 sg13g2_o21ai_1 _09506_ (.B1(\soc_I.PC[23] ),
    .Y(_02073_),
    .A1(net526),
    .A2(net450));
 sg13g2_buf_1 _09507_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[23] ),
    .X(_02074_));
 sg13g2_nand3_1 _09508_ (.B(_02074_),
    .C(net449),
    .A(net598),
    .Y(_02075_));
 sg13g2_nand3_1 _09509_ (.B(_02073_),
    .C(_02075_),
    .A(_01977_),
    .Y(_02076_));
 sg13g2_nand2b_1 _09510_ (.Y(_02077_),
    .B(net368),
    .A_N(\soc_I.kianv_I.datapath_unit_I.A1[23] ));
 sg13g2_and2_1 _09511_ (.A(_02076_),
    .B(_02077_),
    .X(_02078_));
 sg13g2_buf_1 _09512_ (.A(_02078_),
    .X(_02079_));
 sg13g2_buf_8 _09513_ (.A(_02034_),
    .X(_02080_));
 sg13g2_buf_2 _09514_ (.A(\soc_I.kianv_I.Instr[23] ),
    .X(_02081_));
 sg13g2_nand2_1 _09515_ (.Y(_02082_),
    .A(_02081_),
    .B(net416));
 sg13g2_o21ai_1 _09516_ (.B1(net448),
    .Y(_02083_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[23] ),
    .A2(net366));
 sg13g2_a21oi_1 _09517_ (.A1(net323),
    .A2(_02082_),
    .Y(_02084_),
    .B1(_02083_));
 sg13g2_buf_1 _09518_ (.A(_02084_),
    .X(_02085_));
 sg13g2_xnor2_1 _09519_ (.Y(_02086_),
    .A(_02079_),
    .B(net309));
 sg13g2_buf_2 _09520_ (.A(_02086_),
    .X(_02087_));
 sg13g2_nor2_1 _09521_ (.A(_02072_),
    .B(_02087_),
    .Y(_02088_));
 sg13g2_nand3_1 _09522_ (.B(_02057_),
    .C(_02088_),
    .A(net168),
    .Y(_02089_));
 sg13g2_nand2_1 _09523_ (.Y(_02090_),
    .A(_02067_),
    .B(_02068_));
 sg13g2_xnor2_1 _09524_ (.Y(_02091_),
    .A(_02062_),
    .B(_02090_));
 sg13g2_nand2_2 _09525_ (.Y(_02092_),
    .A(_02076_),
    .B(_02077_));
 sg13g2_xnor2_1 _09526_ (.Y(_02093_),
    .A(_02092_),
    .B(_02085_));
 sg13g2_nor2_1 _09527_ (.A(_02091_),
    .B(_02093_),
    .Y(_02094_));
 sg13g2_buf_2 _09528_ (.A(_02094_),
    .X(_02095_));
 sg13g2_and2_1 _09529_ (.A(net272),
    .B(_02056_),
    .X(_02096_));
 sg13g2_buf_1 _09530_ (.A(_02096_),
    .X(_02097_));
 sg13g2_nand3_1 _09531_ (.B(_02095_),
    .C(_02097_),
    .A(net171),
    .Y(_02098_));
 sg13g2_buf_1 _09532_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[19] ),
    .X(_02099_));
 sg13g2_mux2_1 _09533_ (.A0(\soc_I.PC[19] ),
    .A1(_02099_),
    .S(_01580_),
    .X(_02100_));
 sg13g2_mux2_1 _09534_ (.A0(\soc_I.kianv_I.datapath_unit_I.A1[19] ),
    .A1(_02100_),
    .S(net370),
    .X(_02101_));
 sg13g2_buf_1 _09535_ (.A(_02101_),
    .X(_02102_));
 sg13g2_a221oi_1 _09536_ (.B2(\soc_I.kianv_I.Instr[19] ),
    .C1(_01823_),
    .B1(net339),
    .A1(net453),
    .Y(_02103_),
    .A2(net454));
 sg13g2_buf_2 _09537_ (.A(_02103_),
    .X(_02104_));
 sg13g2_o21ai_1 _09538_ (.B1(net451),
    .Y(_02105_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[19] ),
    .A2(net364));
 sg13g2_buf_1 _09539_ (.A(_02105_),
    .X(_02106_));
 sg13g2_or3_1 _09540_ (.A(_02102_),
    .B(_02104_),
    .C(_02106_),
    .X(_02107_));
 sg13g2_buf_2 _09541_ (.A(_02107_),
    .X(_02108_));
 sg13g2_o21ai_1 _09542_ (.B1(_02102_),
    .Y(_02109_),
    .A1(_02104_),
    .A2(_02106_));
 sg13g2_buf_1 _09543_ (.A(_02109_),
    .X(_02110_));
 sg13g2_nand2_1 _09544_ (.Y(_02111_),
    .A(_02108_),
    .B(net271));
 sg13g2_o21ai_1 _09545_ (.B1(net417),
    .Y(_02112_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[18] ),
    .A2(net340));
 sg13g2_buf_1 _09546_ (.A(_02112_),
    .X(_02113_));
 sg13g2_buf_1 _09547_ (.A(\soc_I.kianv_I.Instr[18] ),
    .X(_02114_));
 sg13g2_a221oi_1 _09548_ (.B2(net621),
    .C1(_01823_),
    .B1(net339),
    .A1(net453),
    .Y(_02115_),
    .A2(net454));
 sg13g2_buf_1 _09549_ (.A(_02115_),
    .X(_02116_));
 sg13g2_buf_1 _09550_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[18] ),
    .X(_02117_));
 sg13g2_mux2_1 _09551_ (.A0(\soc_I.PC[18] ),
    .A1(_02117_),
    .S(net420),
    .X(_02118_));
 sg13g2_and2_1 _09552_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[18] ),
    .B(net365),
    .X(_02119_));
 sg13g2_a21o_1 _09553_ (.A2(_02118_),
    .A1(net324),
    .B1(_02119_),
    .X(_02120_));
 sg13g2_o21ai_1 _09554_ (.B1(_02120_),
    .Y(_02121_),
    .A1(_02113_),
    .A2(_02116_));
 sg13g2_buf_2 _09555_ (.A(_02121_),
    .X(_02122_));
 sg13g2_a21oi_1 _09556_ (.A1(_01571_),
    .A2(_02118_),
    .Y(_02123_),
    .B1(_02119_));
 sg13g2_buf_2 _09557_ (.A(_02123_),
    .X(_02124_));
 sg13g2_inv_1 _09558_ (.Y(_02125_),
    .A(\soc_I.kianv_I.datapath_unit_I.A2[18] ));
 sg13g2_a21oi_1 _09559_ (.A1(_02125_),
    .A2(net341),
    .Y(_02126_),
    .B1(net456));
 sg13g2_nand3b_1 _09560_ (.B(_02124_),
    .C(_02126_),
    .Y(_02127_),
    .A_N(_02116_));
 sg13g2_buf_2 _09561_ (.A(_02127_),
    .X(_02128_));
 sg13g2_o21ai_1 _09562_ (.B1(_01807_),
    .Y(_02129_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[17] ),
    .A2(net364));
 sg13g2_buf_2 _09563_ (.A(_02129_),
    .X(_02130_));
 sg13g2_buf_2 _09564_ (.A(\soc_I.kianv_I.Instr[17] ),
    .X(_02131_));
 sg13g2_a221oi_1 _09565_ (.B2(net620),
    .C1(_01823_),
    .B1(net339),
    .A1(net453),
    .Y(_02132_),
    .A2(net454));
 sg13g2_buf_2 _09566_ (.A(_02132_),
    .X(_02133_));
 sg13g2_buf_1 _09567_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[17] ),
    .X(_02134_));
 sg13g2_mux2_1 _09568_ (.A0(\soc_I.PC[17] ),
    .A1(_02134_),
    .S(net420),
    .X(_02135_));
 sg13g2_and2_1 _09569_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[17] ),
    .B(net419),
    .X(_02136_));
 sg13g2_a21o_1 _09570_ (.A2(_02135_),
    .A1(net337),
    .B1(_02136_),
    .X(_02137_));
 sg13g2_buf_1 _09571_ (.A(_02137_),
    .X(_02138_));
 sg13g2_o21ai_1 _09572_ (.B1(_02138_),
    .Y(_02139_),
    .A1(_02130_),
    .A2(_02133_));
 sg13g2_buf_1 _09573_ (.A(_02139_),
    .X(_02140_));
 sg13g2_or3_1 _09574_ (.A(_02138_),
    .B(_02130_),
    .C(_02133_),
    .X(_02141_));
 sg13g2_buf_2 _09575_ (.A(_02141_),
    .X(_02142_));
 sg13g2_nand4_1 _09576_ (.B(_02128_),
    .C(net270),
    .A(_02122_),
    .Y(_02143_),
    .D(_02142_));
 sg13g2_buf_1 _09577_ (.A(_02143_),
    .X(_02144_));
 sg13g2_o21ai_1 _09578_ (.B1(net417),
    .Y(_02145_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[16] ),
    .A2(net364));
 sg13g2_buf_1 _09579_ (.A(_02145_),
    .X(_02146_));
 sg13g2_buf_2 _09580_ (.A(\soc_I.kianv_I.Instr[16] ),
    .X(_02147_));
 sg13g2_a221oi_1 _09581_ (.B2(_02147_),
    .C1(_01823_),
    .B1(net339),
    .A1(net453),
    .Y(_02148_),
    .A2(net454));
 sg13g2_buf_2 _09582_ (.A(_02148_),
    .X(_02149_));
 sg13g2_buf_2 _09583_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[16] ),
    .X(_02150_));
 sg13g2_mux2_1 _09584_ (.A0(\soc_I.PC[16] ),
    .A1(_02150_),
    .S(net420),
    .X(_02151_));
 sg13g2_and2_1 _09585_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[16] ),
    .B(net365),
    .X(_02152_));
 sg13g2_a21o_1 _09586_ (.A2(_02151_),
    .A1(net343),
    .B1(_02152_),
    .X(_02153_));
 sg13g2_buf_1 _09587_ (.A(_02153_),
    .X(_02154_));
 sg13g2_o21ai_1 _09588_ (.B1(_02154_),
    .Y(_02155_),
    .A1(_02146_),
    .A2(_02149_));
 sg13g2_buf_1 _09589_ (.A(_02155_),
    .X(_02156_));
 sg13g2_or3_1 _09590_ (.A(_02154_),
    .B(_02146_),
    .C(_02149_),
    .X(_02157_));
 sg13g2_buf_2 _09591_ (.A(_02157_),
    .X(_02158_));
 sg13g2_nand2_2 _09592_ (.Y(_02159_),
    .A(net269),
    .B(_02158_));
 sg13g2_or4_1 _09593_ (.A(net169),
    .B(_02111_),
    .C(_02144_),
    .D(_02159_),
    .X(_02160_));
 sg13g2_a22oi_1 _09594_ (.Y(_02161_),
    .B1(net270),
    .B2(_02142_),
    .A2(_02128_),
    .A1(_02122_));
 sg13g2_buf_2 _09595_ (.A(_02161_),
    .X(_02162_));
 sg13g2_nand4_1 _09596_ (.B(_02111_),
    .C(_02159_),
    .A(net168),
    .Y(_02163_),
    .D(_02162_));
 sg13g2_a22oi_1 _09597_ (.Y(_02164_),
    .B1(_02160_),
    .B2(_02163_),
    .A2(_02098_),
    .A1(_02089_));
 sg13g2_buf_2 _09598_ (.A(_02164_),
    .X(_02165_));
 sg13g2_nand3_1 _09599_ (.B(_02029_),
    .C(_02165_),
    .A(_01925_),
    .Y(_02166_));
 sg13g2_and2_1 _09600_ (.A(_01891_),
    .B(_01896_),
    .X(_02167_));
 sg13g2_buf_1 _09601_ (.A(_02167_),
    .X(_02168_));
 sg13g2_nor2_1 _09602_ (.A(_01898_),
    .B(_01900_),
    .Y(_02169_));
 sg13g2_buf_2 _09603_ (.A(_02169_),
    .X(_02170_));
 sg13g2_nand2_1 _09604_ (.Y(_02171_),
    .A(_02170_),
    .B(_01873_));
 sg13g2_nand2b_1 _09605_ (.Y(_02172_),
    .B(_01907_),
    .A_N(_01901_));
 sg13g2_buf_2 _09606_ (.A(_02172_),
    .X(_02173_));
 sg13g2_o21ai_1 _09607_ (.B1(_02173_),
    .Y(_02174_),
    .A1(_02170_),
    .A2(_01873_));
 sg13g2_nand4_1 _09608_ (.B(_01837_),
    .C(_02171_),
    .A(_02168_),
    .Y(_02175_),
    .D(_02174_));
 sg13g2_buf_8 _09609_ (.A(net162),
    .X(_02176_));
 sg13g2_nor3_1 _09610_ (.A(_01810_),
    .B(_01825_),
    .C(_01831_),
    .Y(_02177_));
 sg13g2_a21oi_1 _09611_ (.A1(_01891_),
    .A2(_01833_),
    .Y(_02178_),
    .B1(_02177_));
 sg13g2_nor2_1 _09612_ (.A(_02176_),
    .B(_02178_),
    .Y(_02179_));
 sg13g2_buf_8 _09613_ (.A(net170),
    .X(_02180_));
 sg13g2_nor2_1 _09614_ (.A(_01810_),
    .B(_01825_),
    .Y(_02181_));
 sg13g2_buf_1 _09615_ (.A(_02181_),
    .X(_02182_));
 sg13g2_nand3_1 _09616_ (.B(_01882_),
    .C(_01887_),
    .A(_01894_),
    .Y(_02183_));
 sg13g2_buf_1 _09617_ (.A(_02183_),
    .X(_02184_));
 sg13g2_a21oi_2 _09618_ (.B1(_01829_),
    .Y(_02185_),
    .A2(_01827_),
    .A1(net314));
 sg13g2_o21ai_1 _09619_ (.B1(_02185_),
    .Y(_02186_),
    .A1(_01881_),
    .A2(_02184_));
 sg13g2_nor3_1 _09620_ (.A(_01881_),
    .B(_02185_),
    .C(_02184_),
    .Y(_02187_));
 sg13g2_a21o_1 _09621_ (.A2(_02186_),
    .A1(_02182_),
    .B1(_02187_),
    .X(_02188_));
 sg13g2_nor2_1 _09622_ (.A(net161),
    .B(_02188_),
    .Y(_02189_));
 sg13g2_nor3_2 _09623_ (.A(_01898_),
    .B(_01900_),
    .C(_02173_),
    .Y(_02190_));
 sg13g2_nor2_1 _09624_ (.A(_01853_),
    .B(_01859_),
    .Y(_02191_));
 sg13g2_buf_2 _09625_ (.A(_02191_),
    .X(_02192_));
 sg13g2_o21ai_1 _09626_ (.B1(_02173_),
    .Y(_02193_),
    .A1(_01898_),
    .A2(_01900_));
 sg13g2_and3_1 _09627_ (.X(_02194_),
    .A(_01871_),
    .B(_02192_),
    .C(_02193_));
 sg13g2_a22oi_1 _09628_ (.Y(_02195_),
    .B1(_01833_),
    .B2(_01835_),
    .A2(_01896_),
    .A1(_01891_));
 sg13g2_buf_1 _09629_ (.A(_02195_),
    .X(_02196_));
 sg13g2_o21ai_1 _09630_ (.B1(_02196_),
    .Y(_02197_),
    .A1(_02190_),
    .A2(_02194_));
 sg13g2_a22oi_1 _09631_ (.Y(_02198_),
    .B1(_02189_),
    .B2(_02197_),
    .A2(_02179_),
    .A1(_02175_));
 sg13g2_buf_1 _09632_ (.A(_02198_),
    .X(_02199_));
 sg13g2_and2_1 _09633_ (.A(_02108_),
    .B(_02110_),
    .X(_02200_));
 sg13g2_buf_2 _09634_ (.A(_02200_),
    .X(_02201_));
 sg13g2_and2_1 _09635_ (.A(_02122_),
    .B(_02128_),
    .X(_02202_));
 sg13g2_buf_1 _09636_ (.A(_02202_),
    .X(_02203_));
 sg13g2_a21oi_1 _09637_ (.A1(_01572_),
    .A2(_02135_),
    .Y(_02204_),
    .B1(_02136_));
 sg13g2_buf_2 _09638_ (.A(_02204_),
    .X(_02205_));
 sg13g2_nor2_2 _09639_ (.A(_02130_),
    .B(_02133_),
    .Y(_02206_));
 sg13g2_o21ai_1 _09640_ (.B1(_02206_),
    .Y(_02207_),
    .A1(_02205_),
    .A2(net269));
 sg13g2_nand2_1 _09641_ (.Y(_02208_),
    .A(_02205_),
    .B(net269));
 sg13g2_nand4_1 _09642_ (.B(_02203_),
    .C(_02207_),
    .A(_02201_),
    .Y(_02209_),
    .D(_02208_));
 sg13g2_nor3_1 _09643_ (.A(_02102_),
    .B(_02104_),
    .C(_02106_),
    .Y(_02210_));
 sg13g2_a21oi_1 _09644_ (.A1(net271),
    .A2(_02122_),
    .Y(_02211_),
    .B1(_02210_));
 sg13g2_nor2_1 _09645_ (.A(_02176_),
    .B(_02211_),
    .Y(_02212_));
 sg13g2_buf_1 _09646_ (.A(_01779_),
    .X(_02213_));
 sg13g2_a21oi_1 _09647_ (.A1(net325),
    .A2(_01738_),
    .Y(_02214_),
    .B1(_01739_));
 sg13g2_nand2_1 _09648_ (.Y(_02215_),
    .A(net268),
    .B(_02214_));
 sg13g2_nand2_1 _09649_ (.Y(_02216_),
    .A(_01736_),
    .B(_01741_));
 sg13g2_a21oi_2 _09650_ (.B1(_02152_),
    .Y(_02217_),
    .A2(_02151_),
    .A1(net314));
 sg13g2_nor3_1 _09651_ (.A(_02217_),
    .B(_02146_),
    .C(_02149_),
    .Y(_02218_));
 sg13g2_o21ai_1 _09652_ (.B1(_02205_),
    .Y(_02219_),
    .A1(_02130_),
    .A2(_02133_));
 sg13g2_nor3_1 _09653_ (.A(_02205_),
    .B(_02130_),
    .C(_02133_),
    .Y(_02220_));
 sg13g2_a21o_1 _09654_ (.A2(_02219_),
    .A1(_02218_),
    .B1(_02220_),
    .X(_02221_));
 sg13g2_a22oi_1 _09655_ (.Y(_02222_),
    .B1(_02122_),
    .B2(_02128_),
    .A2(net271),
    .A1(_02108_));
 sg13g2_nor3_1 _09656_ (.A(_02113_),
    .B(_02116_),
    .C(_02124_),
    .Y(_02223_));
 sg13g2_nand2b_1 _09657_ (.Y(_02224_),
    .B(net368),
    .A_N(\soc_I.kianv_I.datapath_unit_I.A1[19] ));
 sg13g2_o21ai_1 _09658_ (.B1(_02224_),
    .Y(_02225_),
    .A1(net368),
    .A2(_02100_));
 sg13g2_buf_1 _09659_ (.A(_02225_),
    .X(_02226_));
 sg13g2_o21ai_1 _09660_ (.B1(_02226_),
    .Y(_02227_),
    .A1(_02104_),
    .A2(_02106_));
 sg13g2_nor3_1 _09661_ (.A(_02226_),
    .B(_02104_),
    .C(_02106_),
    .Y(_02228_));
 sg13g2_a21o_1 _09662_ (.A2(_02227_),
    .A1(_02223_),
    .B1(_02228_),
    .X(_02229_));
 sg13g2_a221oi_1 _09663_ (.B2(_02222_),
    .C1(_02229_),
    .B1(_02221_),
    .A1(_02215_),
    .Y(_02230_),
    .A2(_02216_));
 sg13g2_a221oi_1 _09664_ (.B2(_02212_),
    .C1(_02230_),
    .B1(_02209_),
    .A1(_02089_),
    .Y(_02231_),
    .A2(_02098_));
 sg13g2_a21oi_2 _09665_ (.B1(_02231_),
    .Y(_02232_),
    .A2(_02165_),
    .A1(_02199_));
 sg13g2_and2_1 _09666_ (.A(_02166_),
    .B(_02232_),
    .X(_02233_));
 sg13g2_buf_2 _09667_ (.A(_02233_),
    .X(_02234_));
 sg13g2_inv_1 _09668_ (.Y(_02235_),
    .A(_02038_));
 sg13g2_a21oi_1 _09669_ (.A1(net323),
    .A2(_02045_),
    .Y(_02236_),
    .B1(_02046_));
 sg13g2_buf_1 _09670_ (.A(_02236_),
    .X(_02237_));
 sg13g2_a21oi_1 _09671_ (.A1(net343),
    .A2(_02051_),
    .Y(_02238_),
    .B1(_02052_));
 sg13g2_buf_2 _09672_ (.A(_02238_),
    .X(_02239_));
 sg13g2_nand3_1 _09673_ (.B(_02237_),
    .C(_02239_),
    .A(_02042_),
    .Y(_02240_));
 sg13g2_a21oi_1 _09674_ (.A1(_02237_),
    .A2(_02239_),
    .Y(_02241_),
    .B1(_02042_));
 sg13g2_a21oi_1 _09675_ (.A1(_02235_),
    .A2(_02240_),
    .Y(_02242_),
    .B1(_02241_));
 sg13g2_buf_1 _09676_ (.A(_02079_),
    .X(_02243_));
 sg13g2_nor2_1 _09677_ (.A(net267),
    .B(net309),
    .Y(_02244_));
 sg13g2_nand2_1 _09678_ (.Y(_02245_),
    .A(_02062_),
    .B(_02070_));
 sg13g2_nor2_1 _09679_ (.A(_02244_),
    .B(_02245_),
    .Y(_02246_));
 sg13g2_nor2_1 _09680_ (.A(_02062_),
    .B(_02070_),
    .Y(_02247_));
 sg13g2_nor2_1 _09681_ (.A(_02244_),
    .B(_02247_),
    .Y(_02248_));
 sg13g2_o21ai_1 _09682_ (.B1(_02248_),
    .Y(_02249_),
    .A1(_02242_),
    .A2(_02246_));
 sg13g2_nand2_1 _09683_ (.Y(_02250_),
    .A(net267),
    .B(net309));
 sg13g2_and2_1 _09684_ (.A(net156),
    .B(_02250_),
    .X(_02251_));
 sg13g2_nand2_1 _09685_ (.Y(_02252_),
    .A(_02249_),
    .B(_02251_));
 sg13g2_nand2b_1 _09686_ (.Y(_02253_),
    .B(net338),
    .A_N(\soc_I.kianv_I.datapath_unit_I.A1[21] ));
 sg13g2_o21ai_1 _09687_ (.B1(_02253_),
    .Y(_02254_),
    .A1(net338),
    .A2(_02040_));
 sg13g2_buf_1 _09688_ (.A(_02254_),
    .X(_02255_));
 sg13g2_nand2_1 _09689_ (.Y(_02256_),
    .A(_02048_),
    .B(_02239_));
 sg13g2_o21ai_1 _09690_ (.B1(_02038_),
    .Y(_02257_),
    .A1(_02255_),
    .A2(_02256_));
 sg13g2_nand2_1 _09691_ (.Y(_02258_),
    .A(_02255_),
    .B(_02256_));
 sg13g2_nand3_1 _09692_ (.B(_02257_),
    .C(_02258_),
    .A(_02095_),
    .Y(_02259_));
 sg13g2_nand2b_1 _09693_ (.Y(_02260_),
    .B(_02070_),
    .A_N(_02062_));
 sg13g2_a21o_1 _09694_ (.A2(_02082_),
    .A1(net323),
    .B1(_02083_),
    .X(_02261_));
 sg13g2_buf_1 _09695_ (.A(_02261_),
    .X(_02262_));
 sg13g2_nor2_1 _09696_ (.A(net267),
    .B(_02262_),
    .Y(_02263_));
 sg13g2_nand2_1 _09697_ (.Y(_02264_),
    .A(net267),
    .B(_02262_));
 sg13g2_o21ai_1 _09698_ (.B1(_02264_),
    .Y(_02265_),
    .A1(_02260_),
    .A2(_02263_));
 sg13g2_nor2_1 _09699_ (.A(net157),
    .B(_02265_),
    .Y(_02266_));
 sg13g2_nand2_1 _09700_ (.Y(_02267_),
    .A(_02259_),
    .B(_02266_));
 sg13g2_buf_1 _09701_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[2] ),
    .X(_02268_));
 sg13g2_mux2_1 _09702_ (.A0(\soc_I.PC[2] ),
    .A1(_02268_),
    .S(net369),
    .X(_02269_));
 sg13g2_and2_1 _09703_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[2] ),
    .B(net365),
    .X(_02270_));
 sg13g2_a21o_1 _09704_ (.A2(_02269_),
    .A1(net324),
    .B1(_02270_),
    .X(_02271_));
 sg13g2_buf_1 _09705_ (.A(_02271_),
    .X(_02272_));
 sg13g2_buf_2 _09706_ (.A(\soc_I.kianv_I.Instr[9] ),
    .X(_02273_));
 sg13g2_a221oi_1 _09707_ (.B2(_02273_),
    .C1(_01682_),
    .B1(_01672_),
    .A1(_01700_),
    .Y(_02274_),
    .A2(net454));
 sg13g2_nor3_1 _09708_ (.A(net622),
    .B(net367),
    .C(_01683_),
    .Y(_02275_));
 sg13g2_nand2_1 _09709_ (.Y(_02276_),
    .A(_02273_),
    .B(net418));
 sg13g2_buf_1 _09710_ (.A(\soc_I.cpu_mem_wdata[2] ),
    .X(_02277_));
 sg13g2_nor3_1 _09711_ (.A(net619),
    .B(_01850_),
    .C(net456),
    .Y(_02278_));
 sg13g2_a221oi_1 _09712_ (.B2(_02276_),
    .C1(_02278_),
    .B1(_02275_),
    .A1(net342),
    .Y(_02279_),
    .A2(_02274_));
 sg13g2_buf_2 _09713_ (.A(_02279_),
    .X(_02280_));
 sg13g2_buf_1 _09714_ (.A(_02280_),
    .X(_02281_));
 sg13g2_buf_1 _09715_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[3] ),
    .X(_02282_));
 sg13g2_mux2_1 _09716_ (.A0(\soc_I.PC[3] ),
    .A1(_02282_),
    .S(net369),
    .X(_02283_));
 sg13g2_mux2_1 _09717_ (.A0(\soc_I.kianv_I.datapath_unit_I.A1[3] ),
    .A1(_02283_),
    .S(net324),
    .X(_02284_));
 sg13g2_buf_2 _09718_ (.A(_02284_),
    .X(_02285_));
 sg13g2_buf_2 _09719_ (.A(_02285_),
    .X(_02286_));
 sg13g2_a21o_1 _09720_ (.A2(_01676_),
    .A1(_00036_),
    .B1(_01682_),
    .X(_02287_));
 sg13g2_buf_1 _09721_ (.A(_02287_),
    .X(_02288_));
 sg13g2_buf_2 _09722_ (.A(\soc_I.kianv_I.Instr[10] ),
    .X(_02289_));
 sg13g2_a21oi_1 _09723_ (.A1(_02289_),
    .A2(net418),
    .Y(_02290_),
    .B1(_01676_));
 sg13g2_or2_1 _09724_ (.X(_02291_),
    .B(_02290_),
    .A(_02288_));
 sg13g2_buf_1 _09725_ (.A(_02291_),
    .X(_02292_));
 sg13g2_or3_1 _09726_ (.A(_00037_),
    .B(_01665_),
    .C(_02288_),
    .X(_02293_));
 sg13g2_buf_1 _09727_ (.A(_02293_),
    .X(_02294_));
 sg13g2_nand2_1 _09728_ (.Y(_02295_),
    .A(_02292_),
    .B(_02294_));
 sg13g2_buf_2 _09729_ (.A(_02295_),
    .X(_02296_));
 sg13g2_a22oi_1 _09730_ (.Y(_02297_),
    .B1(net266),
    .B2(_02296_),
    .A2(net308),
    .A1(_02272_));
 sg13g2_a21oi_1 _09731_ (.A1(net324),
    .A2(_02269_),
    .Y(_02298_),
    .B1(_02270_));
 sg13g2_buf_2 _09732_ (.A(_02298_),
    .X(_02299_));
 sg13g2_or2_1 _09733_ (.X(_02300_),
    .B(_02280_),
    .A(_02299_));
 sg13g2_buf_1 _09734_ (.A(_02300_),
    .X(_02301_));
 sg13g2_nand3_1 _09735_ (.B(_02292_),
    .C(_02294_),
    .A(_02285_),
    .Y(_02302_));
 sg13g2_and2_1 _09736_ (.A(_02301_),
    .B(_02302_),
    .X(_02303_));
 sg13g2_mux2_1 _09737_ (.A0(_02297_),
    .A1(_02303_),
    .S(net180),
    .X(_02304_));
 sg13g2_buf_1 _09738_ (.A(_02304_),
    .X(_02305_));
 sg13g2_and3_1 _09739_ (.X(_02306_),
    .A(_01679_),
    .B(_01684_),
    .C(_01775_));
 sg13g2_buf_1 _09740_ (.A(_02306_),
    .X(_02307_));
 sg13g2_a21o_1 _09741_ (.A2(_01684_),
    .A1(_01679_),
    .B1(_01775_),
    .X(_02308_));
 sg13g2_o21ai_1 _09742_ (.B1(_02308_),
    .Y(_02309_),
    .A1(_01719_),
    .A2(_02307_));
 sg13g2_nand2_1 _09743_ (.Y(_02310_),
    .A(_02272_),
    .B(_02280_));
 sg13g2_buf_2 _09744_ (.A(_02310_),
    .X(_02311_));
 sg13g2_nand2b_1 _09745_ (.Y(_02312_),
    .B(_02299_),
    .A_N(_02280_));
 sg13g2_buf_1 _09746_ (.A(_02312_),
    .X(_02313_));
 sg13g2_nand2_1 _09747_ (.Y(_02314_),
    .A(_02311_),
    .B(_02313_));
 sg13g2_nand3_1 _09748_ (.B(_02309_),
    .C(_02314_),
    .A(net171),
    .Y(_02315_));
 sg13g2_a21oi_1 _09749_ (.A1(_01711_),
    .A2(_01715_),
    .Y(_02316_),
    .B1(_01589_));
 sg13g2_nand3_1 _09750_ (.B(_01711_),
    .C(_01715_),
    .A(_01589_),
    .Y(_02317_));
 sg13g2_o21ai_1 _09751_ (.B1(_02317_),
    .Y(_02318_),
    .A1(_01686_),
    .A2(_02316_));
 sg13g2_nand4_1 _09752_ (.B(_02311_),
    .C(_02313_),
    .A(_02030_),
    .Y(_02319_),
    .D(_02318_));
 sg13g2_nand3_1 _09753_ (.B(_02315_),
    .C(_02319_),
    .A(_02305_),
    .Y(_02320_));
 sg13g2_buf_2 _09754_ (.A(_02320_),
    .X(_02321_));
 sg13g2_buf_1 _09755_ (.A(\soc_I.kianv_I.Instr[27] ),
    .X(_02322_));
 sg13g2_nand4_1 _09756_ (.B(_01706_),
    .C(net418),
    .A(_02322_),
    .Y(_02323_),
    .D(net448));
 sg13g2_nand3b_1 _09757_ (.B(net367),
    .C(net448),
    .Y(_02324_),
    .A_N(_00044_));
 sg13g2_nand2_2 _09758_ (.Y(_02325_),
    .A(_02323_),
    .B(_02324_));
 sg13g2_and3_1 _09759_ (.X(_02326_),
    .A(_00044_),
    .B(_01699_),
    .C(_01696_));
 sg13g2_nor3_1 _09760_ (.A(_00045_),
    .B(_01682_),
    .C(_02326_),
    .Y(_02327_));
 sg13g2_nor2b_1 _09761_ (.A(_01666_),
    .B_N(_02327_),
    .Y(_02328_));
 sg13g2_buf_2 _09762_ (.A(_02328_),
    .X(_02329_));
 sg13g2_buf_1 _09763_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[7] ),
    .X(_02330_));
 sg13g2_mux2_1 _09764_ (.A0(\soc_I.PC[7] ),
    .A1(_02330_),
    .S(_01581_),
    .X(_02331_));
 sg13g2_and2_1 _09765_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[7] ),
    .B(net419),
    .X(_02332_));
 sg13g2_a21o_1 _09766_ (.A2(_02331_),
    .A1(net337),
    .B1(_02332_),
    .X(_02333_));
 sg13g2_buf_2 _09767_ (.A(_02333_),
    .X(_02334_));
 sg13g2_nor3_2 _09768_ (.A(_02325_),
    .B(_02329_),
    .C(_02334_),
    .Y(_02335_));
 sg13g2_nor2_1 _09769_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[6] ),
    .B(_01570_),
    .Y(_02336_));
 sg13g2_buf_1 _09770_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[6] ),
    .X(_02337_));
 sg13g2_nand3_1 _09771_ (.B(_02337_),
    .C(_01861_),
    .A(_01574_),
    .Y(_02338_));
 sg13g2_o21ai_1 _09772_ (.B1(\soc_I.PC[6] ),
    .Y(_02339_),
    .A1(net526),
    .A2(net450));
 sg13g2_and3_1 _09773_ (.X(_02340_),
    .A(_01569_),
    .B(_02338_),
    .C(_02339_));
 sg13g2_buf_1 _09774_ (.A(_02340_),
    .X(_02341_));
 sg13g2_nor2_1 _09775_ (.A(_02336_),
    .B(_02341_),
    .Y(_02342_));
 sg13g2_buf_2 _09776_ (.A(_02342_),
    .X(_02343_));
 sg13g2_a21oi_1 _09777_ (.A1(\soc_I.kianv_I.Instr[26] ),
    .A2(net418),
    .Y(_02344_),
    .B1(_01676_));
 sg13g2_a21o_1 _09778_ (.A2(_01676_),
    .A1(_00042_),
    .B1(_01682_),
    .X(_02345_));
 sg13g2_buf_2 _09779_ (.A(_02345_),
    .X(_02346_));
 sg13g2_nor2_2 _09780_ (.A(_02344_),
    .B(_02346_),
    .Y(_02347_));
 sg13g2_nor3_2 _09781_ (.A(_00043_),
    .B(net342),
    .C(_02346_),
    .Y(_02348_));
 sg13g2_nor3_1 _09782_ (.A(_02343_),
    .B(_02347_),
    .C(_02348_),
    .Y(_02349_));
 sg13g2_o21ai_1 _09783_ (.B1(_02334_),
    .Y(_02350_),
    .A1(_02325_),
    .A2(_02329_));
 sg13g2_buf_2 _09784_ (.A(_02350_),
    .X(_02351_));
 sg13g2_o21ai_1 _09785_ (.B1(_02351_),
    .Y(_02352_),
    .A1(_02335_),
    .A2(_02349_));
 sg13g2_nand2_1 _09786_ (.Y(_02353_),
    .A(_02023_),
    .B(_02026_));
 sg13g2_a21o_1 _09787_ (.A2(_01994_),
    .A1(_01991_),
    .B1(_01998_),
    .X(_02354_));
 sg13g2_buf_8 _09788_ (.A(_02354_),
    .X(_02355_));
 sg13g2_nand4_1 _09789_ (.B(_01706_),
    .C(_01806_),
    .A(_01934_),
    .Y(_02356_),
    .D(_01849_));
 sg13g2_buf_1 _09790_ (.A(_02356_),
    .X(_02357_));
 sg13g2_nand3_1 _09791_ (.B(_01676_),
    .C(_01806_),
    .A(_01936_),
    .Y(_02358_));
 sg13g2_buf_1 _09792_ (.A(_02358_),
    .X(_02359_));
 sg13g2_nand4_1 _09793_ (.B(_01933_),
    .C(_02357_),
    .A(_01928_),
    .Y(_02360_),
    .D(_02359_));
 sg13g2_buf_1 _09794_ (.A(_02360_),
    .X(_02361_));
 sg13g2_nand4_1 _09795_ (.B(_02012_),
    .C(_02014_),
    .A(_01807_),
    .Y(_02362_),
    .D(_01938_));
 sg13g2_buf_2 _09796_ (.A(_02362_),
    .X(_02363_));
 sg13g2_and4_1 _09797_ (.A(_01950_),
    .B(_01707_),
    .C(net448),
    .D(_01849_),
    .X(_02364_));
 sg13g2_and3_1 _09798_ (.X(_02365_),
    .A(_01952_),
    .B(net367),
    .C(net448));
 sg13g2_or4_1 _09799_ (.A(_02009_),
    .B(_02010_),
    .C(_02364_),
    .D(_02365_),
    .X(_02366_));
 sg13g2_buf_2 _09800_ (.A(_02366_),
    .X(_02367_));
 sg13g2_nand2_1 _09801_ (.Y(_02368_),
    .A(_01940_),
    .B(_01828_));
 sg13g2_o21ai_1 _09802_ (.B1(_01977_),
    .Y(_02369_),
    .A1(_01945_),
    .A2(_01947_));
 sg13g2_nand4_1 _09803_ (.B(_02368_),
    .C(_02369_),
    .A(_01808_),
    .Y(_02370_),
    .D(_01955_));
 sg13g2_buf_1 _09804_ (.A(_02370_),
    .X(_02371_));
 sg13g2_a22oi_1 _09805_ (.Y(_02372_),
    .B1(_02367_),
    .B2(_02371_),
    .A2(_02363_),
    .A1(_02361_));
 sg13g2_buf_1 _09806_ (.A(_02372_),
    .X(_02373_));
 sg13g2_nand3_1 _09807_ (.B(_01994_),
    .C(_01998_),
    .A(_01991_),
    .Y(_02374_));
 sg13g2_buf_2 _09808_ (.A(_02374_),
    .X(_02375_));
 sg13g2_and3_1 _09809_ (.X(_02376_),
    .A(_02355_),
    .B(_02373_),
    .C(_02375_));
 sg13g2_nand4_1 _09810_ (.B(_02352_),
    .C(_02353_),
    .A(net162),
    .Y(_02377_),
    .D(_02376_));
 sg13g2_and2_1 _09811_ (.A(_02023_),
    .B(_02026_),
    .X(_02378_));
 sg13g2_buf_2 _09812_ (.A(_02378_),
    .X(_02379_));
 sg13g2_and2_1 _09813_ (.A(_02323_),
    .B(_02324_),
    .X(_02380_));
 sg13g2_buf_1 _09814_ (.A(_02380_),
    .X(_02381_));
 sg13g2_nand2b_1 _09815_ (.Y(_02382_),
    .B(_02327_),
    .A_N(net342));
 sg13g2_buf_1 _09816_ (.A(_02382_),
    .X(_02383_));
 sg13g2_a21oi_1 _09817_ (.A1(_02381_),
    .A2(_02383_),
    .Y(_02384_),
    .B1(_02334_));
 sg13g2_or2_1 _09818_ (.X(_02385_),
    .B(_02346_),
    .A(_02344_));
 sg13g2_buf_2 _09819_ (.A(_02385_),
    .X(_02386_));
 sg13g2_or3_1 _09820_ (.A(_00043_),
    .B(_01665_),
    .C(_02346_),
    .X(_02387_));
 sg13g2_buf_2 _09821_ (.A(_02387_),
    .X(_02388_));
 sg13g2_a21oi_1 _09822_ (.A1(_02386_),
    .A2(_02388_),
    .Y(_02389_),
    .B1(_02343_));
 sg13g2_nand3_1 _09823_ (.B(_02383_),
    .C(_02334_),
    .A(_02381_),
    .Y(_02390_));
 sg13g2_buf_1 _09824_ (.A(_02390_),
    .X(_02391_));
 sg13g2_o21ai_1 _09825_ (.B1(_02391_),
    .Y(_02392_),
    .A1(_02384_),
    .A2(_02389_));
 sg13g2_nand4_1 _09826_ (.B(_02363_),
    .C(_02367_),
    .A(_02361_),
    .Y(_02393_),
    .D(_02371_));
 sg13g2_buf_1 _09827_ (.A(_02393_),
    .X(_02394_));
 sg13g2_a21oi_1 _09828_ (.A1(_02355_),
    .A2(_02375_),
    .Y(_02395_),
    .B1(_02394_));
 sg13g2_nand4_1 _09829_ (.B(_02379_),
    .C(_02392_),
    .A(net171),
    .Y(_02396_),
    .D(_02395_));
 sg13g2_buf_1 _09830_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[4] ),
    .X(_02397_));
 sg13g2_mux2_1 _09831_ (.A0(\soc_I.PC[4] ),
    .A1(_02397_),
    .S(_01581_),
    .X(_02398_));
 sg13g2_and2_1 _09832_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[4] ),
    .B(_01585_),
    .X(_02399_));
 sg13g2_a21oi_1 _09833_ (.A1(net324),
    .A2(_02398_),
    .Y(_02400_),
    .B1(_02399_));
 sg13g2_buf_2 _09834_ (.A(_02400_),
    .X(_02401_));
 sg13g2_nand4_1 _09835_ (.B(net366),
    .C(net418),
    .A(\soc_I.kianv_I.Instr[11] ),
    .Y(_02402_),
    .D(_02035_));
 sg13g2_nand3b_1 _09836_ (.B(net367),
    .C(_02035_),
    .Y(_02403_),
    .A_N(_00038_));
 sg13g2_nand2_2 _09837_ (.Y(_02404_),
    .A(_02402_),
    .B(_02403_));
 sg13g2_and3_1 _09838_ (.X(_02405_),
    .A(_00038_),
    .B(_01699_),
    .C(_01696_));
 sg13g2_nor3_1 _09839_ (.A(_00039_),
    .B(_01682_),
    .C(_02405_),
    .Y(_02406_));
 sg13g2_nor2b_2 _09840_ (.A(net342),
    .B_N(_02406_),
    .Y(_02407_));
 sg13g2_nor3_2 _09841_ (.A(_02401_),
    .B(_02404_),
    .C(_02407_),
    .Y(_02408_));
 sg13g2_and2_1 _09842_ (.A(_02402_),
    .B(_02403_),
    .X(_02409_));
 sg13g2_buf_2 _09843_ (.A(_02409_),
    .X(_02410_));
 sg13g2_nand2b_1 _09844_ (.Y(_02411_),
    .B(_02406_),
    .A_N(net342));
 sg13g2_buf_1 _09845_ (.A(_02411_),
    .X(_02412_));
 sg13g2_a21o_1 _09846_ (.A2(_02398_),
    .A1(net343),
    .B1(_02399_),
    .X(_02413_));
 sg13g2_buf_1 _09847_ (.A(_02413_),
    .X(_02414_));
 sg13g2_a21oi_2 _09848_ (.B1(_02414_),
    .Y(_02415_),
    .A2(_02412_),
    .A1(_02410_));
 sg13g2_a21oi_1 _09849_ (.A1(_02292_),
    .A2(_02294_),
    .Y(_02416_),
    .B1(net266));
 sg13g2_nor3_2 _09850_ (.A(_02408_),
    .B(_02415_),
    .C(_02416_),
    .Y(_02417_));
 sg13g2_a21oi_1 _09851_ (.A1(_00040_),
    .A2(net367),
    .Y(_02418_),
    .B1(_01682_));
 sg13g2_buf_2 _09852_ (.A(_02418_),
    .X(_02419_));
 sg13g2_buf_1 _09853_ (.A(_00041_),
    .X(_02420_));
 sg13g2_a21oi_1 _09854_ (.A1(\soc_I.kianv_I.Instr[25] ),
    .A2(net418),
    .Y(_02421_),
    .B1(_01676_));
 sg13g2_o21ai_1 _09855_ (.B1(_02421_),
    .Y(_02422_),
    .A1(_02420_),
    .A2(_01665_));
 sg13g2_buf_2 _09856_ (.A(_02422_),
    .X(_02423_));
 sg13g2_nor2_2 _09857_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[5] ),
    .B(_01570_),
    .Y(_02424_));
 sg13g2_buf_1 _09858_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[5] ),
    .X(_02425_));
 sg13g2_inv_1 _09859_ (.Y(_02426_),
    .A(_02425_));
 sg13g2_nor3_1 _09860_ (.A(_01863_),
    .B(_02426_),
    .C(_01866_),
    .Y(_02427_));
 sg13g2_inv_1 _09861_ (.Y(_02428_),
    .A(\soc_I.PC[5] ));
 sg13g2_a21oi_1 _09862_ (.A1(_01902_),
    .A2(_01861_),
    .Y(_02429_),
    .B1(_02428_));
 sg13g2_or3_1 _09863_ (.A(net419),
    .B(_02427_),
    .C(_02429_),
    .X(_02430_));
 sg13g2_nand2b_1 _09864_ (.Y(_02431_),
    .B(_02430_),
    .A_N(_02424_));
 sg13g2_buf_2 _09865_ (.A(_02431_),
    .X(_02432_));
 sg13g2_a21oi_2 _09866_ (.B1(_02432_),
    .Y(_02433_),
    .A2(_02423_),
    .A1(_02419_));
 sg13g2_and3_1 _09867_ (.X(_02434_),
    .A(_02432_),
    .B(_02419_),
    .C(_02423_));
 sg13g2_buf_2 _09868_ (.A(_02434_),
    .X(_02435_));
 sg13g2_nor2_1 _09869_ (.A(_02433_),
    .B(_02435_),
    .Y(_02436_));
 sg13g2_buf_1 _09870_ (.A(_02436_),
    .X(_02437_));
 sg13g2_nand3_1 _09871_ (.B(_02417_),
    .C(_02437_),
    .A(net170),
    .Y(_02438_));
 sg13g2_buf_8 _09872_ (.A(net168),
    .X(_02439_));
 sg13g2_a21o_1 _09873_ (.A2(_02423_),
    .A1(_02419_),
    .B1(_02432_),
    .X(_02440_));
 sg13g2_buf_1 _09874_ (.A(_02440_),
    .X(_02441_));
 sg13g2_nand3_1 _09875_ (.B(_02419_),
    .C(_02423_),
    .A(_02432_),
    .Y(_02442_));
 sg13g2_buf_1 _09876_ (.A(_02442_),
    .X(_02443_));
 sg13g2_o21ai_1 _09877_ (.B1(_02401_),
    .Y(_02444_),
    .A1(_02404_),
    .A2(_02407_));
 sg13g2_nand3_1 _09878_ (.B(_02410_),
    .C(_02412_),
    .A(_02414_),
    .Y(_02445_));
 sg13g2_buf_1 _09879_ (.A(_02445_),
    .X(_02446_));
 sg13g2_nor2_1 _09880_ (.A(_02288_),
    .B(_02290_),
    .Y(_02447_));
 sg13g2_nor3_1 _09881_ (.A(_00037_),
    .B(net342),
    .C(_02288_),
    .Y(_02448_));
 sg13g2_nor3_1 _09882_ (.A(net266),
    .B(_02447_),
    .C(_02448_),
    .Y(_02449_));
 sg13g2_a221oi_1 _09883_ (.B2(_02446_),
    .C1(_02449_),
    .B1(_02444_),
    .A1(_02441_),
    .Y(_02450_),
    .A2(_02443_));
 sg13g2_buf_1 _09884_ (.A(_02450_),
    .X(_02451_));
 sg13g2_nand2_1 _09885_ (.Y(_02452_),
    .A(net160),
    .B(_02451_));
 sg13g2_a22oi_1 _09886_ (.Y(_02453_),
    .B1(_02438_),
    .B2(_02452_),
    .A2(_02396_),
    .A1(_02377_));
 sg13g2_o21ai_1 _09887_ (.B1(_02441_),
    .Y(_02454_),
    .A1(_02446_),
    .A2(_02435_));
 sg13g2_buf_2 _09888_ (.A(_02454_),
    .X(_02455_));
 sg13g2_nand3_1 _09889_ (.B(_02386_),
    .C(_02388_),
    .A(_02343_),
    .Y(_02456_));
 sg13g2_buf_2 _09890_ (.A(_02456_),
    .X(_02457_));
 sg13g2_a21oi_1 _09891_ (.A1(_02391_),
    .A2(_02457_),
    .Y(_02458_),
    .B1(_02384_));
 sg13g2_nor2_1 _09892_ (.A(_02455_),
    .B(_02458_),
    .Y(_02459_));
 sg13g2_a21oi_1 _09893_ (.A1(_02410_),
    .A2(_02412_),
    .Y(_02460_),
    .B1(_02401_));
 sg13g2_nor3_1 _09894_ (.A(_01828_),
    .B(_02427_),
    .C(_02429_),
    .Y(_02461_));
 sg13g2_nor2_1 _09895_ (.A(_02424_),
    .B(_02461_),
    .Y(_02462_));
 sg13g2_a21o_1 _09896_ (.A2(_02423_),
    .A1(_02419_),
    .B1(_02462_),
    .X(_02463_));
 sg13g2_buf_1 _09897_ (.A(_02463_),
    .X(_02464_));
 sg13g2_nand3b_1 _09898_ (.B(_02430_),
    .C(_02419_),
    .Y(_02465_),
    .A_N(_02424_));
 sg13g2_nor2b_1 _09899_ (.A(_02465_),
    .B_N(_02423_),
    .Y(_02466_));
 sg13g2_a21o_1 _09900_ (.A2(_02464_),
    .A1(_02460_),
    .B1(_02466_),
    .X(_02467_));
 sg13g2_buf_2 _09901_ (.A(_02467_),
    .X(_02468_));
 sg13g2_o21ai_1 _09902_ (.B1(_02343_),
    .Y(_02469_),
    .A1(_02347_),
    .A2(_02348_));
 sg13g2_buf_2 _09903_ (.A(_02469_),
    .X(_02470_));
 sg13g2_o21ai_1 _09904_ (.B1(_02351_),
    .Y(_02471_),
    .A1(_02335_),
    .A2(_02470_));
 sg13g2_buf_1 _09905_ (.A(_02471_),
    .X(_02472_));
 sg13g2_nor3_1 _09906_ (.A(_01757_),
    .B(_02468_),
    .C(_02472_),
    .Y(_02473_));
 sg13g2_a221oi_1 _09907_ (.B2(_02180_),
    .C1(_02473_),
    .B1(_02459_),
    .A1(_02377_),
    .Y(_02474_),
    .A2(_02396_));
 sg13g2_a21o_1 _09908_ (.A2(_02453_),
    .A1(_02321_),
    .B1(_02474_),
    .X(_02475_));
 sg13g2_buf_1 _09909_ (.A(_02475_),
    .X(_02476_));
 sg13g2_and2_1 _09910_ (.A(_01925_),
    .B(_02165_),
    .X(_02477_));
 sg13g2_buf_1 _09911_ (.A(_02477_),
    .X(_02478_));
 sg13g2_buf_1 _09912_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[25] ),
    .X(_02479_));
 sg13g2_mux2_1 _09913_ (.A0(\soc_I.PC[25] ),
    .A1(_02479_),
    .S(net369),
    .X(_02480_));
 sg13g2_and2_1 _09914_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[25] ),
    .B(net365),
    .X(_02481_));
 sg13g2_a21o_1 _09915_ (.A2(_02480_),
    .A1(net324),
    .B1(_02481_),
    .X(_02482_));
 sg13g2_buf_1 _09916_ (.A(_02482_),
    .X(_02483_));
 sg13g2_nand2_1 _09917_ (.Y(_02484_),
    .A(\soc_I.kianv_I.Instr[25] ),
    .B(net416));
 sg13g2_o21ai_1 _09918_ (.B1(net451),
    .Y(_02485_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[25] ),
    .A2(_01707_));
 sg13g2_a21oi_1 _09919_ (.A1(_02080_),
    .A2(_02484_),
    .Y(_02486_),
    .B1(_02485_));
 sg13g2_buf_1 _09920_ (.A(_02486_),
    .X(_02487_));
 sg13g2_nor2_1 _09921_ (.A(_02483_),
    .B(net307),
    .Y(_02488_));
 sg13g2_buf_1 _09922_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[24] ),
    .X(_02489_));
 sg13g2_mux2_1 _09923_ (.A0(\soc_I.PC[24] ),
    .A1(_02489_),
    .S(net420),
    .X(_02490_));
 sg13g2_mux2_1 _09924_ (.A0(\soc_I.kianv_I.datapath_unit_I.A1[24] ),
    .A1(_02490_),
    .S(net343),
    .X(_02491_));
 sg13g2_buf_1 _09925_ (.A(_02491_),
    .X(_02492_));
 sg13g2_buf_1 _09926_ (.A(_02492_),
    .X(_02493_));
 sg13g2_nand2_1 _09927_ (.Y(_02494_),
    .A(\soc_I.kianv_I.Instr[24] ),
    .B(net416));
 sg13g2_o21ai_1 _09928_ (.B1(net451),
    .Y(_02495_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[24] ),
    .A2(net366));
 sg13g2_a21oi_1 _09929_ (.A1(net323),
    .A2(_02494_),
    .Y(_02496_),
    .B1(_02495_));
 sg13g2_buf_2 _09930_ (.A(_02496_),
    .X(_02497_));
 sg13g2_nand2_1 _09931_ (.Y(_02498_),
    .A(net306),
    .B(_02497_));
 sg13g2_or2_1 _09932_ (.X(_02499_),
    .B(_02498_),
    .A(_02488_));
 sg13g2_a21o_1 _09933_ (.A2(_02494_),
    .A1(net323),
    .B1(_02495_),
    .X(_02500_));
 sg13g2_buf_2 _09934_ (.A(_02500_),
    .X(_02501_));
 sg13g2_nand2_1 _09935_ (.Y(_02502_),
    .A(net306),
    .B(_02501_));
 sg13g2_a21oi_2 _09936_ (.B1(_02481_),
    .Y(_02503_),
    .A2(_02480_),
    .A1(net343));
 sg13g2_nand2_1 _09937_ (.Y(_02504_),
    .A(_02503_),
    .B(net307));
 sg13g2_nand2b_1 _09938_ (.Y(_02505_),
    .B(_02504_),
    .A_N(_02502_));
 sg13g2_mux2_1 _09939_ (.A0(_02499_),
    .A1(_02505_),
    .S(_01754_),
    .X(_02506_));
 sg13g2_buf_1 _09940_ (.A(_02506_),
    .X(_02507_));
 sg13g2_or2_1 _09941_ (.X(_02508_),
    .B(net307),
    .A(_02503_));
 sg13g2_buf_1 _09942_ (.A(_02508_),
    .X(_02509_));
 sg13g2_nand2_1 _09943_ (.Y(_02510_),
    .A(_02483_),
    .B(net307));
 sg13g2_mux2_1 _09944_ (.A0(_02509_),
    .A1(_02510_),
    .S(_01917_),
    .X(_02511_));
 sg13g2_buf_1 _09945_ (.A(_02511_),
    .X(_02512_));
 sg13g2_nand2_1 _09946_ (.Y(_02513_),
    .A(_02507_),
    .B(_02512_));
 sg13g2_buf_1 _09947_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[28] ),
    .X(_02514_));
 sg13g2_mux2_1 _09948_ (.A0(\soc_I.PC[28] ),
    .A1(_02514_),
    .S(_01582_),
    .X(_02515_));
 sg13g2_and2_1 _09949_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[28] ),
    .B(net338),
    .X(_02516_));
 sg13g2_a21oi_2 _09950_ (.B1(_02516_),
    .Y(_02517_),
    .A2(_02515_),
    .A1(net314));
 sg13g2_nand2_1 _09951_ (.Y(_02518_),
    .A(_01934_),
    .B(net416));
 sg13g2_o21ai_1 _09952_ (.B1(net417),
    .Y(_02519_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[28] ),
    .A2(_01708_));
 sg13g2_a21oi_1 _09953_ (.A1(_02080_),
    .A2(_02518_),
    .Y(_02520_),
    .B1(_02519_));
 sg13g2_buf_2 _09954_ (.A(_02520_),
    .X(_02521_));
 sg13g2_xnor2_1 _09955_ (.Y(_02522_),
    .A(_02517_),
    .B(_02521_));
 sg13g2_buf_2 _09956_ (.A(_02522_),
    .X(_02523_));
 sg13g2_nand2_1 _09957_ (.Y(_02524_),
    .A(_01950_),
    .B(net416));
 sg13g2_o21ai_1 _09958_ (.B1(net417),
    .Y(_02525_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[29] ),
    .A2(net340));
 sg13g2_a21oi_2 _09959_ (.B1(_02525_),
    .Y(_02526_),
    .A2(_02524_),
    .A1(net323));
 sg13g2_buf_1 _09960_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[29] ),
    .X(_02527_));
 sg13g2_mux2_1 _09961_ (.A0(\soc_I.PC[29] ),
    .A1(_02527_),
    .S(net369),
    .X(_02528_));
 sg13g2_and2_1 _09962_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[29] ),
    .B(net368),
    .X(_02529_));
 sg13g2_a21oi_1 _09963_ (.A1(net314),
    .A2(_02528_),
    .Y(_02530_),
    .B1(_02529_));
 sg13g2_buf_2 _09964_ (.A(_02530_),
    .X(_02531_));
 sg13g2_xnor2_1 _09965_ (.Y(_02532_),
    .A(_02526_),
    .B(_02531_));
 sg13g2_buf_2 _09966_ (.A(_02532_),
    .X(_02533_));
 sg13g2_inv_1 _09967_ (.Y(_02534_),
    .A(_02322_));
 sg13g2_nor3_1 _09968_ (.A(_02534_),
    .B(_01841_),
    .C(_01844_),
    .Y(_02535_));
 sg13g2_nor2_1 _09969_ (.A(net455),
    .B(_01842_),
    .Y(_02536_));
 sg13g2_a221oi_1 _09970_ (.B2(_02536_),
    .C1(net341),
    .B1(_02535_),
    .A1(net623),
    .Y(_02537_),
    .A2(_01849_));
 sg13g2_buf_1 _09971_ (.A(_02537_),
    .X(_02538_));
 sg13g2_inv_1 _09972_ (.Y(_02539_),
    .A(\soc_I.kianv_I.datapath_unit_I.A2[27] ));
 sg13g2_a21oi_1 _09973_ (.A1(_02539_),
    .A2(net341),
    .Y(_02540_),
    .B1(net456));
 sg13g2_nand2b_1 _09974_ (.Y(_02541_),
    .B(_02540_),
    .A_N(_02538_));
 sg13g2_buf_2 _09975_ (.A(_02541_),
    .X(_02542_));
 sg13g2_nor2_1 _09976_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[27] ),
    .B(net326),
    .Y(_02543_));
 sg13g2_buf_1 _09977_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[27] ),
    .X(_02544_));
 sg13g2_nand3_1 _09978_ (.B(_02544_),
    .C(_01904_),
    .A(net598),
    .Y(_02545_));
 sg13g2_o21ai_1 _09979_ (.B1(\soc_I.PC[27] ),
    .Y(_02546_),
    .A1(net526),
    .A2(net450));
 sg13g2_nand3_1 _09980_ (.B(_02545_),
    .C(_02546_),
    .A(net324),
    .Y(_02547_));
 sg13g2_nand2b_1 _09981_ (.Y(_02548_),
    .B(_02547_),
    .A_N(_02543_));
 sg13g2_buf_1 _09982_ (.A(_02548_),
    .X(_02549_));
 sg13g2_nor2_1 _09983_ (.A(_02542_),
    .B(_02549_),
    .Y(_02550_));
 sg13g2_buf_1 _09984_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[26] ),
    .X(_02551_));
 sg13g2_mux2_1 _09985_ (.A0(\soc_I.PC[26] ),
    .A1(_02551_),
    .S(net369),
    .X(_02552_));
 sg13g2_and2_1 _09986_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[26] ),
    .B(net368),
    .X(_02553_));
 sg13g2_a21o_1 _09987_ (.A2(_02552_),
    .A1(net326),
    .B1(_02553_),
    .X(_02554_));
 sg13g2_buf_2 _09988_ (.A(_02554_),
    .X(_02555_));
 sg13g2_inv_1 _09989_ (.Y(_02556_),
    .A(\soc_I.kianv_I.Instr[26] ));
 sg13g2_nor3_1 _09990_ (.A(_02556_),
    .B(_01841_),
    .C(_01844_),
    .Y(_02557_));
 sg13g2_a221oi_1 _09991_ (.B2(_02536_),
    .C1(net367),
    .B1(_02557_),
    .A1(net623),
    .Y(_02558_),
    .A2(_01849_));
 sg13g2_buf_1 _09992_ (.A(_02558_),
    .X(_02559_));
 sg13g2_nor2_1 _09993_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ),
    .B(net340),
    .Y(_02560_));
 sg13g2_nor2_1 _09994_ (.A(_02559_),
    .B(_02560_),
    .Y(_02561_));
 sg13g2_xnor2_1 _09995_ (.Y(_02562_),
    .A(_02555_),
    .B(_02561_));
 sg13g2_or2_1 _09996_ (.X(_02563_),
    .B(_02560_),
    .A(_02559_));
 sg13g2_buf_1 _09997_ (.A(_02563_),
    .X(_02564_));
 sg13g2_nor3_1 _09998_ (.A(net456),
    .B(_02559_),
    .C(_02560_),
    .Y(_02565_));
 sg13g2_buf_2 _09999_ (.A(_02565_),
    .X(_02566_));
 sg13g2_mux2_1 _10000_ (.A0(_02564_),
    .A1(_02566_),
    .S(_02555_),
    .X(_02567_));
 sg13g2_a21oi_1 _10001_ (.A1(_02539_),
    .A2(net341),
    .Y(_02568_),
    .B1(_02538_));
 sg13g2_nor2b_1 _10002_ (.A(_02543_),
    .B_N(_02547_),
    .Y(_02569_));
 sg13g2_buf_2 _10003_ (.A(_02569_),
    .X(_02570_));
 sg13g2_nor2_1 _10004_ (.A(_02568_),
    .B(_02570_),
    .Y(_02571_));
 sg13g2_nor3_1 _10005_ (.A(net363),
    .B(_02570_),
    .C(_02555_),
    .Y(_02572_));
 sg13g2_a221oi_1 _10006_ (.B2(_02571_),
    .C1(_02572_),
    .B1(_02567_),
    .A1(_02550_),
    .Y(_02573_),
    .A2(_02562_));
 sg13g2_buf_1 _10007_ (.A(_02573_),
    .X(_02574_));
 sg13g2_nor4_1 _10008_ (.A(net168),
    .B(_02523_),
    .C(_02533_),
    .D(_02574_),
    .Y(_02575_));
 sg13g2_nand2_2 _10009_ (.Y(_02576_),
    .A(_02523_),
    .B(_02533_));
 sg13g2_a21oi_1 _10010_ (.A1(net326),
    .A2(_02552_),
    .Y(_02577_),
    .B1(_02553_));
 sg13g2_buf_2 _10011_ (.A(_02577_),
    .X(_02578_));
 sg13g2_mux2_1 _10012_ (.A0(_02564_),
    .A1(_02566_),
    .S(_02578_),
    .X(_02579_));
 sg13g2_nor2_1 _10013_ (.A(_02568_),
    .B(_02549_),
    .Y(_02580_));
 sg13g2_nor2_2 _10014_ (.A(_02542_),
    .B(_02570_),
    .Y(_02581_));
 sg13g2_xnor2_1 _10015_ (.Y(_02582_),
    .A(_02578_),
    .B(_02561_));
 sg13g2_nor3_1 _10016_ (.A(net363),
    .B(_02549_),
    .C(_02578_),
    .Y(_02583_));
 sg13g2_a221oi_1 _10017_ (.B2(_02582_),
    .C1(_02583_),
    .B1(_02581_),
    .A1(_02579_),
    .Y(_02584_),
    .A2(_02580_));
 sg13g2_buf_1 _10018_ (.A(_02584_),
    .X(_02585_));
 sg13g2_nor3_1 _10019_ (.A(net171),
    .B(_02576_),
    .C(_02585_),
    .Y(_02586_));
 sg13g2_or2_1 _10020_ (.X(_02587_),
    .B(_02586_),
    .A(_02575_));
 sg13g2_nor2b_1 _10021_ (.A(_02538_),
    .B_N(_02540_),
    .Y(_02588_));
 sg13g2_buf_1 _10022_ (.A(_02588_),
    .X(_02589_));
 sg13g2_nand2_1 _10023_ (.Y(_02590_),
    .A(_02589_),
    .B(_02570_));
 sg13g2_buf_1 _10024_ (.A(_02549_),
    .X(_02591_));
 sg13g2_nand2_1 _10025_ (.Y(_02592_),
    .A(_02542_),
    .B(net211));
 sg13g2_nand3_1 _10026_ (.B(_02566_),
    .C(_02592_),
    .A(_02555_),
    .Y(_02593_));
 sg13g2_a21o_1 _10027_ (.A2(_02593_),
    .A1(_02590_),
    .B1(_02576_),
    .X(_02594_));
 sg13g2_a21o_1 _10028_ (.A2(_02515_),
    .A1(net314),
    .B1(_02516_),
    .X(_02595_));
 sg13g2_buf_1 _10029_ (.A(_02595_),
    .X(_02596_));
 sg13g2_nand2_1 _10030_ (.Y(_02597_),
    .A(_02596_),
    .B(_02521_));
 sg13g2_nor2_1 _10031_ (.A(_02531_),
    .B(_02597_),
    .Y(_02598_));
 sg13g2_a21o_1 _10032_ (.A2(_02524_),
    .A1(net323),
    .B1(_02525_),
    .X(_02599_));
 sg13g2_buf_1 _10033_ (.A(_02599_),
    .X(_02600_));
 sg13g2_a21oi_1 _10034_ (.A1(_02531_),
    .A2(_02597_),
    .Y(_02601_),
    .B1(_02600_));
 sg13g2_nor3_1 _10035_ (.A(net179),
    .B(_02598_),
    .C(_02601_),
    .Y(_02602_));
 sg13g2_o21ai_1 _10036_ (.B1(net211),
    .Y(_02603_),
    .A1(_02578_),
    .A2(_02566_));
 sg13g2_buf_1 _10037_ (.A(_02578_),
    .X(_02604_));
 sg13g2_nor2_1 _10038_ (.A(net211),
    .B(net265),
    .Y(_02605_));
 sg13g2_nand2_1 _10039_ (.Y(_02606_),
    .A(net363),
    .B(_02561_));
 sg13g2_a22oi_1 _10040_ (.Y(_02607_),
    .B1(_02605_),
    .B2(_02606_),
    .A2(_02603_),
    .A1(_02542_));
 sg13g2_nor2_2 _10041_ (.A(_02523_),
    .B(_02533_),
    .Y(_02608_));
 sg13g2_nand2b_1 _10042_ (.Y(_02609_),
    .B(_02608_),
    .A_N(_02607_));
 sg13g2_nor2_1 _10043_ (.A(_02517_),
    .B(_02521_),
    .Y(_02610_));
 sg13g2_a21o_1 _10044_ (.A2(_02528_),
    .A1(net314),
    .B1(_02529_),
    .X(_02611_));
 sg13g2_buf_1 _10045_ (.A(_02611_),
    .X(_02612_));
 sg13g2_nand2_1 _10046_ (.Y(_02613_),
    .A(_02610_),
    .B(_02612_));
 sg13g2_o21ai_1 _10047_ (.B1(_02600_),
    .Y(_02614_),
    .A1(_02610_),
    .A2(_02612_));
 sg13g2_and3_1 _10048_ (.X(_02615_),
    .A(net171),
    .B(_02613_),
    .C(_02614_));
 sg13g2_a22oi_1 _10049_ (.Y(_02616_),
    .B1(_02609_),
    .B2(_02615_),
    .A2(_02602_),
    .A1(_02594_));
 sg13g2_a21o_1 _10050_ (.A2(_02587_),
    .A1(_02513_),
    .B1(_02616_),
    .X(_02617_));
 sg13g2_a221oi_1 _10051_ (.B2(_02478_),
    .C1(_02617_),
    .B1(_02476_),
    .A1(_02252_),
    .Y(_02618_),
    .A2(_02267_));
 sg13g2_buf_1 _10052_ (.A(_02618_),
    .X(_02619_));
 sg13g2_nand2_1 _10053_ (.Y(_02620_),
    .A(_02234_),
    .B(_02619_));
 sg13g2_buf_1 _10054_ (.A(net268),
    .X(_02621_));
 sg13g2_buf_1 _10055_ (.A(net210),
    .X(_02622_));
 sg13g2_buf_1 _10056_ (.A(net184),
    .X(_02623_));
 sg13g2_o21ai_1 _10057_ (.B1(_01721_),
    .Y(_02624_),
    .A1(net177),
    .A2(_01635_));
 sg13g2_buf_1 _10058_ (.A(_02566_),
    .X(_02625_));
 sg13g2_nand2_1 _10059_ (.Y(_02626_),
    .A(net264),
    .B(_02592_));
 sg13g2_or2_1 _10060_ (.X(_02627_),
    .B(_02581_),
    .A(net264));
 sg13g2_mux2_1 _10061_ (.A0(_02626_),
    .A1(_02627_),
    .S(net163),
    .X(_02628_));
 sg13g2_nand2_1 _10062_ (.Y(_02629_),
    .A(_02570_),
    .B(_02555_));
 sg13g2_a22oi_1 _10063_ (.Y(_02630_),
    .B1(_02628_),
    .B2(_02629_),
    .A2(_02512_),
    .A1(_02507_));
 sg13g2_nand2_1 _10064_ (.Y(_02631_),
    .A(net156),
    .B(_02589_));
 sg13g2_nand2_1 _10065_ (.Y(_02632_),
    .A(net161),
    .B(_02542_));
 sg13g2_a221oi_1 _10066_ (.B2(_02632_),
    .C1(net265),
    .B1(_02631_),
    .A1(_02507_),
    .Y(_02633_),
    .A2(_02512_));
 sg13g2_nor2_1 _10067_ (.A(net265),
    .B(_02628_),
    .Y(_02634_));
 sg13g2_a21oi_1 _10068_ (.A1(_02631_),
    .A2(_02632_),
    .Y(_02635_),
    .B1(net211));
 sg13g2_or4_1 _10069_ (.A(_02630_),
    .B(_02633_),
    .C(_02634_),
    .D(_02635_),
    .X(_02636_));
 sg13g2_buf_1 _10070_ (.A(_02636_),
    .X(_02637_));
 sg13g2_xnor2_1 _10071_ (.Y(_02638_),
    .A(_02503_),
    .B(_02487_));
 sg13g2_buf_1 _10072_ (.A(_02638_),
    .X(_02639_));
 sg13g2_xnor2_1 _10073_ (.Y(_02640_),
    .A(_02492_),
    .B(_02501_));
 sg13g2_buf_1 _10074_ (.A(_02640_),
    .X(_02641_));
 sg13g2_and2_1 _10075_ (.A(net209),
    .B(_02641_),
    .X(_02642_));
 sg13g2_buf_1 _10076_ (.A(_02642_),
    .X(_02643_));
 sg13g2_nand2_1 _10077_ (.Y(_02644_),
    .A(net162),
    .B(_02643_));
 sg13g2_nor2_1 _10078_ (.A(net209),
    .B(_02641_),
    .Y(_02645_));
 sg13g2_nand3b_1 _10079_ (.B(_02645_),
    .C(net170),
    .Y(_02646_),
    .A_N(_02574_));
 sg13g2_o21ai_1 _10080_ (.B1(_02646_),
    .Y(_02647_),
    .A1(_02585_),
    .A2(_02644_));
 sg13g2_buf_2 _10081_ (.A(_02647_),
    .X(_02648_));
 sg13g2_or2_1 _10082_ (.X(_02649_),
    .B(_02615_),
    .A(_02602_));
 sg13g2_nand2b_1 _10083_ (.Y(_02650_),
    .B(_02649_),
    .A_N(_02648_));
 sg13g2_buf_8 _10084_ (.A(net158),
    .X(_02651_));
 sg13g2_buf_1 _10085_ (.A(net153),
    .X(_02652_));
 sg13g2_nor2_1 _10086_ (.A(net153),
    .B(_02576_),
    .Y(_02653_));
 sg13g2_a21oi_1 _10087_ (.A1(net148),
    .A2(_02608_),
    .Y(_02654_),
    .B1(_02653_));
 sg13g2_nand2_1 _10088_ (.Y(_02655_),
    .A(\soc_I.kianv_I.datapath_unit_I.A2[31] ),
    .B(net341));
 sg13g2_nand2_1 _10089_ (.Y(_02656_),
    .A(net623),
    .B(net340));
 sg13g2_a21oi_1 _10090_ (.A1(_02655_),
    .A2(_02656_),
    .Y(_02657_),
    .B1(net456));
 sg13g2_buf_1 _10091_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[31] ),
    .X(_02658_));
 sg13g2_nand2_1 _10092_ (.Y(_02659_),
    .A(_02658_),
    .B(_01582_));
 sg13g2_nand2_1 _10093_ (.Y(_02660_),
    .A(\soc_I.PC[31] ),
    .B(_01862_));
 sg13g2_a21oi_1 _10094_ (.A1(_02659_),
    .A2(_02660_),
    .Y(_02661_),
    .B1(net338));
 sg13g2_a21oi_2 _10095_ (.B1(_02661_),
    .Y(_02662_),
    .A2(_01941_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[31] ));
 sg13g2_xnor2_1 _10096_ (.Y(_02663_),
    .A(_02657_),
    .B(_02662_));
 sg13g2_nor2_1 _10097_ (.A(\soc_I.kianv_I.datapath_unit_I.A1[30] ),
    .B(net314),
    .Y(_02664_));
 sg13g2_buf_1 _10098_ (.A(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[30] ),
    .X(_02665_));
 sg13g2_nand3_1 _10099_ (.B(_02665_),
    .C(net449),
    .A(_01902_),
    .Y(_02666_));
 sg13g2_o21ai_1 _10100_ (.B1(\soc_I.PC[30] ),
    .Y(_02667_),
    .A1(net526),
    .A2(net450));
 sg13g2_nand3_1 _10101_ (.B(_02666_),
    .C(_02667_),
    .A(_02007_),
    .Y(_02668_));
 sg13g2_nand2b_1 _10102_ (.Y(_02669_),
    .B(_02668_),
    .A_N(_02664_));
 sg13g2_buf_1 _10103_ (.A(_02669_),
    .X(_02670_));
 sg13g2_nand3_1 _10104_ (.B(net340),
    .C(_01849_),
    .A(net623),
    .Y(_02671_));
 sg13g2_buf_1 _10105_ (.A(_02671_),
    .X(_02672_));
 sg13g2_a21oi_1 _10106_ (.A1(net453),
    .A2(net454),
    .Y(_02673_),
    .B1(_01729_));
 sg13g2_a22oi_1 _10107_ (.Y(_02674_),
    .B1(_01846_),
    .B2(_02673_),
    .A2(net341),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[30] ));
 sg13g2_buf_1 _10108_ (.A(_02674_),
    .X(_02675_));
 sg13g2_a21oi_1 _10109_ (.A1(_02672_),
    .A2(_02675_),
    .Y(_02676_),
    .B1(net456));
 sg13g2_buf_2 _10110_ (.A(_02676_),
    .X(_02677_));
 sg13g2_or2_1 _10111_ (.X(_02678_),
    .B(_02677_),
    .A(_02670_));
 sg13g2_buf_1 _10112_ (.A(_02678_),
    .X(_02679_));
 sg13g2_nand2_1 _10113_ (.Y(_02680_),
    .A(net208),
    .B(_02677_));
 sg13g2_and2_1 _10114_ (.A(_02679_),
    .B(_02680_),
    .X(_02681_));
 sg13g2_buf_1 _10115_ (.A(_02681_),
    .X(_02682_));
 sg13g2_nor2b_1 _10116_ (.A(_02663_),
    .B_N(_02682_),
    .Y(_02683_));
 sg13g2_buf_8 _10117_ (.A(net161),
    .X(_02684_));
 sg13g2_buf_8 _10118_ (.A(net155),
    .X(_02685_));
 sg13g2_nor2_1 _10119_ (.A(net152),
    .B(_02682_),
    .Y(_02686_));
 sg13g2_a22oi_1 _10120_ (.Y(_02687_),
    .B1(_02686_),
    .B2(_02663_),
    .A2(_02683_),
    .A1(net148));
 sg13g2_a21oi_1 _10121_ (.A1(_02649_),
    .A2(_02654_),
    .Y(_02688_),
    .B1(_02687_));
 sg13g2_o21ai_1 _10122_ (.B1(_02688_),
    .Y(_02689_),
    .A1(_02637_),
    .A2(_02650_));
 sg13g2_nor2_1 _10123_ (.A(_02624_),
    .B(_02689_),
    .Y(_02690_));
 sg13g2_nand2_1 _10124_ (.Y(_02691_),
    .A(_02620_),
    .B(_02690_));
 sg13g2_inv_1 _10125_ (.Y(_02692_),
    .A(_02624_));
 sg13g2_buf_1 _10126_ (.A(_02657_),
    .X(_02693_));
 sg13g2_a21oi_1 _10127_ (.A1(net305),
    .A2(_02662_),
    .Y(_02694_),
    .B1(_02677_));
 sg13g2_a21o_1 _10128_ (.A2(_01941_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[31] ),
    .B1(_02661_),
    .X(_02695_));
 sg13g2_buf_2 _10129_ (.A(_02695_),
    .X(_02696_));
 sg13g2_o21ai_1 _10130_ (.B1(_02677_),
    .Y(_02697_),
    .A1(net305),
    .A2(_02696_));
 sg13g2_nor2_1 _10131_ (.A(net152),
    .B(_02697_),
    .Y(_02698_));
 sg13g2_a21oi_1 _10132_ (.A1(_02652_),
    .A2(_02694_),
    .Y(_02699_),
    .B1(_02698_));
 sg13g2_buf_8 _10133_ (.A(net156),
    .X(_02700_));
 sg13g2_buf_8 _10134_ (.A(net151),
    .X(_02701_));
 sg13g2_xnor2_1 _10135_ (.Y(_02702_),
    .A(net147),
    .B(net305));
 sg13g2_nand2_1 _10136_ (.Y(_02703_),
    .A(_02696_),
    .B(_02702_));
 sg13g2_o21ai_1 _10137_ (.B1(_02703_),
    .Y(_02704_),
    .A1(net208),
    .A2(_02699_));
 sg13g2_buf_1 _10138_ (.A(_02704_),
    .X(_02705_));
 sg13g2_a21oi_1 _10139_ (.A1(_02692_),
    .A2(_02705_),
    .Y(_02706_),
    .B1(_01597_));
 sg13g2_nand2_1 _10140_ (.Y(_02707_),
    .A(net602),
    .B(net603));
 sg13g2_a21o_1 _10141_ (.A2(_02619_),
    .A1(_02234_),
    .B1(_02689_),
    .X(_02708_));
 sg13g2_nor2_1 _10142_ (.A(_02707_),
    .B(_02705_),
    .Y(_02709_));
 sg13g2_a22oi_1 _10143_ (.Y(_02710_),
    .B1(_02708_),
    .B2(_02709_),
    .A2(net325),
    .A1(_02707_));
 sg13g2_nand3_1 _10144_ (.B(_02706_),
    .C(_02710_),
    .A(_02691_),
    .Y(_02711_));
 sg13g2_buf_1 _10145_ (.A(net177),
    .X(_02712_));
 sg13g2_nor3_2 _10146_ (.A(_01721_),
    .B(net167),
    .C(_01597_),
    .Y(_02713_));
 sg13g2_nand2_1 _10147_ (.Y(_02714_),
    .A(_02517_),
    .B(_02521_));
 sg13g2_nor2_1 _10148_ (.A(_02589_),
    .B(net211),
    .Y(_02715_));
 sg13g2_a21oi_1 _10149_ (.A1(_02714_),
    .A2(_02715_),
    .Y(_02716_),
    .B1(_02610_));
 sg13g2_nor2_1 _10150_ (.A(_02596_),
    .B(_02521_),
    .Y(_02717_));
 sg13g2_a21o_1 _10151_ (.A2(_02597_),
    .A1(_02590_),
    .B1(_02717_),
    .X(_02718_));
 sg13g2_mux2_1 _10152_ (.A0(_02716_),
    .A1(_02718_),
    .S(net169),
    .X(_02719_));
 sg13g2_buf_2 _10153_ (.A(_02719_),
    .X(_02720_));
 sg13g2_nor2b_1 _10154_ (.A(_02664_),
    .B_N(_02668_),
    .Y(_02721_));
 sg13g2_buf_2 _10155_ (.A(_02721_),
    .X(_02722_));
 sg13g2_xnor2_1 _10156_ (.Y(_02723_),
    .A(net160),
    .B(_02677_));
 sg13g2_o21ai_1 _10157_ (.B1(_02723_),
    .Y(_02724_),
    .A1(_02722_),
    .A2(_02612_));
 sg13g2_a21o_1 _10158_ (.A2(_02720_),
    .A1(net208),
    .B1(_02724_),
    .X(_02725_));
 sg13g2_o21ai_1 _10159_ (.B1(_02526_),
    .Y(_02726_),
    .A1(_02722_),
    .A2(_02677_));
 sg13g2_nand2b_1 _10160_ (.Y(_02727_),
    .B(net160),
    .A_N(_02726_));
 sg13g2_nand3_1 _10161_ (.B(_02600_),
    .C(_02680_),
    .A(net163),
    .Y(_02728_));
 sg13g2_a22oi_1 _10162_ (.Y(_02729_),
    .B1(_02720_),
    .B2(_02531_),
    .A2(_02728_),
    .A1(_02727_));
 sg13g2_nor3_1 _10163_ (.A(net208),
    .B(_02531_),
    .C(_02720_),
    .Y(_02730_));
 sg13g2_nor2_1 _10164_ (.A(_02729_),
    .B(_02730_),
    .Y(_02731_));
 sg13g2_nor2_1 _10165_ (.A(_02048_),
    .B(_02239_),
    .Y(_02732_));
 sg13g2_o21ai_1 _10166_ (.B1(_02256_),
    .Y(_02733_),
    .A1(_02732_),
    .A2(net271));
 sg13g2_nand3_1 _10167_ (.B(_02072_),
    .C(_02733_),
    .A(net272),
    .Y(_02734_));
 sg13g2_a221oi_1 _10168_ (.B2(_02068_),
    .C1(_02060_),
    .B1(_02067_),
    .A1(net323),
    .Y(_02735_),
    .A2(_02059_));
 sg13g2_or3_1 _10169_ (.A(_02038_),
    .B(_02255_),
    .C(_02735_),
    .X(_02736_));
 sg13g2_and3_1 _10170_ (.X(_02737_),
    .A(net179),
    .B(_02260_),
    .C(_02736_));
 sg13g2_nor2_1 _10171_ (.A(net272),
    .B(_02072_),
    .Y(_02738_));
 sg13g2_nand2_1 _10172_ (.Y(_02739_),
    .A(_02048_),
    .B(_02054_));
 sg13g2_nor2_1 _10173_ (.A(_02048_),
    .B(_02054_),
    .Y(_02740_));
 sg13g2_a21o_1 _10174_ (.A2(_02739_),
    .A1(_02228_),
    .B1(_02740_),
    .X(_02741_));
 sg13g2_buf_1 _10175_ (.A(_02741_),
    .X(_02742_));
 sg13g2_a22oi_1 _10176_ (.Y(_02743_),
    .B1(_02062_),
    .B2(_02070_),
    .A2(_02042_),
    .A1(_02038_));
 sg13g2_nor2_1 _10177_ (.A(_02247_),
    .B(_02743_),
    .Y(_02744_));
 sg13g2_a21oi_1 _10178_ (.A1(_02738_),
    .A2(_02742_),
    .Y(_02745_),
    .B1(_02744_));
 sg13g2_a22oi_1 _10179_ (.Y(_02746_),
    .B1(_02745_),
    .B2(net162),
    .A2(_02737_),
    .A1(_02734_));
 sg13g2_buf_1 _10180_ (.A(_02746_),
    .X(_02747_));
 sg13g2_o21ai_1 _10181_ (.B1(_02217_),
    .Y(_02748_),
    .A1(_02146_),
    .A2(_02149_));
 sg13g2_and3_1 _10182_ (.X(_02749_),
    .A(_02182_),
    .B(_01831_),
    .C(_02748_));
 sg13g2_o21ai_1 _10183_ (.B1(_02162_),
    .Y(_02750_),
    .A1(_02218_),
    .A2(_02749_));
 sg13g2_or3_1 _10184_ (.A(_02205_),
    .B(_02130_),
    .C(_02133_),
    .X(_02751_));
 sg13g2_and2_1 _10185_ (.A(net621),
    .B(net339),
    .X(_02752_));
 sg13g2_inv_1 _10186_ (.Y(_02753_),
    .A(_02134_));
 sg13g2_inv_1 _10187_ (.Y(_02754_),
    .A(_02117_));
 sg13g2_nor4_1 _10188_ (.A(net526),
    .B(_02753_),
    .C(_02754_),
    .D(_01866_),
    .Y(_02755_));
 sg13g2_nand2_1 _10189_ (.Y(_02756_),
    .A(\soc_I.PC[17] ),
    .B(\soc_I.PC[18] ));
 sg13g2_a21oi_1 _10190_ (.A1(net598),
    .A2(net449),
    .Y(_02757_),
    .B1(_02756_));
 sg13g2_o21ai_1 _10191_ (.B1(net326),
    .Y(_02758_),
    .A1(_02755_),
    .A2(_02757_));
 sg13g2_nand3_1 _10192_ (.B(\soc_I.kianv_I.datapath_unit_I.A1[18] ),
    .C(net368),
    .A(\soc_I.kianv_I.datapath_unit_I.A1[17] ),
    .Y(_02759_));
 sg13g2_a21oi_1 _10193_ (.A1(_02758_),
    .A2(_02759_),
    .Y(_02760_),
    .B1(_02130_));
 sg13g2_and2_1 _10194_ (.A(net620),
    .B(net339),
    .X(_02761_));
 sg13g2_a22oi_1 _10195_ (.Y(_02762_),
    .B1(_02760_),
    .B2(_02761_),
    .A2(_02752_),
    .A1(_02126_));
 sg13g2_or2_1 _10196_ (.X(_02763_),
    .B(_01823_),
    .A(_01680_));
 sg13g2_o21ai_1 _10197_ (.B1(_02763_),
    .Y(_02764_),
    .A1(_02126_),
    .A2(_02760_));
 sg13g2_a22oi_1 _10198_ (.Y(_02765_),
    .B1(_02762_),
    .B2(_02764_),
    .A2(_02124_),
    .A1(_02751_));
 sg13g2_buf_1 _10199_ (.A(_02765_),
    .X(_02766_));
 sg13g2_nor2_1 _10200_ (.A(net180),
    .B(_02766_),
    .Y(_02767_));
 sg13g2_nand4_1 _10201_ (.B(_02072_),
    .C(_02097_),
    .A(net179),
    .Y(_02768_),
    .D(_02201_));
 sg13g2_nand2_1 _10202_ (.Y(_02769_),
    .A(_02237_),
    .B(_02054_));
 sg13g2_a221oi_1 _10203_ (.B2(net271),
    .C1(net272),
    .B1(_02108_),
    .A1(_02256_),
    .Y(_02770_),
    .A2(_02769_));
 sg13g2_buf_1 _10204_ (.A(_02770_),
    .X(_02771_));
 sg13g2_nand3_1 _10205_ (.B(_02091_),
    .C(_02771_),
    .A(net169),
    .Y(_02772_));
 sg13g2_and4_1 _10206_ (.A(_02122_),
    .B(_02128_),
    .C(net270),
    .D(_02142_),
    .X(_02773_));
 sg13g2_nor3_1 _10207_ (.A(_02154_),
    .B(_02146_),
    .C(_02149_),
    .Y(_02774_));
 sg13g2_a21oi_1 _10208_ (.A1(_02156_),
    .A2(_01833_),
    .Y(_02775_),
    .B1(_02774_));
 sg13g2_nor2_2 _10209_ (.A(_02113_),
    .B(_02116_),
    .Y(_02776_));
 sg13g2_nand2_1 _10210_ (.Y(_02777_),
    .A(_02758_),
    .B(_02759_));
 sg13g2_o21ai_1 _10211_ (.B1(_02777_),
    .Y(_02778_),
    .A1(_02130_),
    .A2(_02133_));
 sg13g2_nand2_1 _10212_ (.Y(_02779_),
    .A(_02776_),
    .B(_02778_));
 sg13g2_nand2_1 _10213_ (.Y(_02780_),
    .A(_02124_),
    .B(net270));
 sg13g2_a221oi_1 _10214_ (.B2(_02780_),
    .C1(net178),
    .B1(_02779_),
    .A1(_02773_),
    .Y(_02781_),
    .A2(_02775_));
 sg13g2_buf_1 _10215_ (.A(_02781_),
    .X(_02782_));
 sg13g2_a221oi_1 _10216_ (.B2(_02772_),
    .C1(_02782_),
    .B1(_02768_),
    .A1(_02750_),
    .Y(_02783_),
    .A2(_02767_));
 sg13g2_buf_1 _10217_ (.A(_02783_),
    .X(_02784_));
 sg13g2_nand2_2 _10218_ (.Y(_02785_),
    .A(_02672_),
    .B(_02675_));
 sg13g2_xnor2_1 _10219_ (.Y(_02786_),
    .A(_02722_),
    .B(_02785_));
 sg13g2_o21ai_1 _10220_ (.B1(net363),
    .Y(_02787_),
    .A1(_02785_),
    .A2(_02568_));
 sg13g2_nor2_1 _10221_ (.A(_02722_),
    .B(_02570_),
    .Y(_02788_));
 sg13g2_mux2_1 _10222_ (.A0(_02322_),
    .A1(net623),
    .S(_01849_),
    .X(_02789_));
 sg13g2_nor2_1 _10223_ (.A(_02539_),
    .B(_01708_),
    .Y(_02790_));
 sg13g2_a221oi_1 _10224_ (.B2(net340),
    .C1(_02790_),
    .B1(_02789_),
    .A1(_02672_),
    .Y(_02791_),
    .A2(_02675_));
 sg13g2_and4_1 _10225_ (.A(net363),
    .B(_02722_),
    .C(net211),
    .D(_02791_),
    .X(_02792_));
 sg13g2_a221oi_1 _10226_ (.B2(_02788_),
    .C1(_02792_),
    .B1(_02787_),
    .A1(_02550_),
    .Y(_02793_),
    .A2(_02786_));
 sg13g2_nand3b_1 _10227_ (.B(_02608_),
    .C(net170),
    .Y(_02794_),
    .A_N(_02793_));
 sg13g2_xnor2_1 _10228_ (.Y(_02795_),
    .A(net208),
    .B(_02785_));
 sg13g2_nor2_1 _10229_ (.A(net208),
    .B(net211),
    .Y(_02796_));
 sg13g2_and4_1 _10230_ (.A(net363),
    .B(net208),
    .C(_02570_),
    .D(_02791_),
    .X(_02797_));
 sg13g2_a221oi_1 _10231_ (.B2(_02796_),
    .C1(_02797_),
    .B1(_02787_),
    .A1(_02581_),
    .Y(_02798_),
    .A2(_02795_));
 sg13g2_or3_1 _10232_ (.A(net170),
    .B(_02576_),
    .C(_02798_),
    .X(_02799_));
 sg13g2_xnor2_1 _10233_ (.Y(_02800_),
    .A(_02492_),
    .B(_02497_));
 sg13g2_xnor2_1 _10234_ (.Y(_02801_),
    .A(_02578_),
    .B(_02566_));
 sg13g2_nor2_1 _10235_ (.A(net209),
    .B(_02801_),
    .Y(_02802_));
 sg13g2_nand4_1 _10236_ (.B(_02087_),
    .C(_02800_),
    .A(net170),
    .Y(_02803_),
    .D(_02802_));
 sg13g2_and2_1 _10237_ (.A(net209),
    .B(_02801_),
    .X(_02804_));
 sg13g2_nor2_1 _10238_ (.A(_02087_),
    .B(_02800_),
    .Y(_02805_));
 sg13g2_nand3_1 _10239_ (.B(_02804_),
    .C(_02805_),
    .A(net162),
    .Y(_02806_));
 sg13g2_a22oi_1 _10240_ (.Y(_02807_),
    .B1(_02803_),
    .B2(_02806_),
    .A2(_02799_),
    .A1(_02794_));
 sg13g2_o21ai_1 _10241_ (.B1(_02807_),
    .Y(_02808_),
    .A1(_02747_),
    .A2(_02784_));
 sg13g2_nand2_1 _10242_ (.Y(_02809_),
    .A(_02794_),
    .B(_02799_));
 sg13g2_nor2_1 _10243_ (.A(net171),
    .B(net264),
    .Y(_02810_));
 sg13g2_nand3_1 _10244_ (.B(net309),
    .C(_02497_),
    .A(net267),
    .Y(_02811_));
 sg13g2_nand3_1 _10245_ (.B(net309),
    .C(net306),
    .A(net267),
    .Y(_02812_));
 sg13g2_nand4_1 _10246_ (.B(_02510_),
    .C(_02811_),
    .A(_02498_),
    .Y(_02813_),
    .D(_02812_));
 sg13g2_nor2_1 _10247_ (.A(net265),
    .B(_02488_),
    .Y(_02814_));
 sg13g2_nand2_1 _10248_ (.Y(_02815_),
    .A(_02813_),
    .B(_02814_));
 sg13g2_nor2_1 _10249_ (.A(net170),
    .B(_02555_),
    .Y(_02816_));
 sg13g2_nand2b_1 _10250_ (.Y(_02817_),
    .B(_02813_),
    .A_N(_02488_));
 sg13g2_nand3_1 _10251_ (.B(_02262_),
    .C(net306),
    .A(net267),
    .Y(_02818_));
 sg13g2_nand3_1 _10252_ (.B(_02262_),
    .C(_02501_),
    .A(net267),
    .Y(_02819_));
 sg13g2_nand3_1 _10253_ (.B(_02818_),
    .C(_02819_),
    .A(_02502_),
    .Y(_02820_));
 sg13g2_o21ai_1 _10254_ (.B1(net265),
    .Y(_02821_),
    .A1(net264),
    .A2(_02509_));
 sg13g2_nand2_1 _10255_ (.Y(_02822_),
    .A(net264),
    .B(_02509_));
 sg13g2_a221oi_1 _10256_ (.B2(_02822_),
    .C1(net162),
    .B1(_02821_),
    .A1(_02802_),
    .Y(_02823_),
    .A2(_02820_));
 sg13g2_a221oi_1 _10257_ (.B2(_02817_),
    .C1(_02823_),
    .B1(_02816_),
    .A1(_02810_),
    .Y(_02824_),
    .A2(_02815_));
 sg13g2_nand2_1 _10258_ (.Y(_02825_),
    .A(_02809_),
    .B(_02824_));
 sg13g2_nand4_1 _10259_ (.B(_02731_),
    .C(_02808_),
    .A(_02725_),
    .Y(_02826_),
    .D(_02825_));
 sg13g2_buf_1 _10260_ (.A(_02826_),
    .X(_02827_));
 sg13g2_nor3_1 _10261_ (.A(_01871_),
    .B(_01853_),
    .C(_01859_),
    .Y(_02828_));
 sg13g2_o21ai_1 _10262_ (.B1(_01873_),
    .Y(_02829_),
    .A1(_02828_),
    .A2(_02026_));
 sg13g2_nor3_1 _10263_ (.A(_01879_),
    .B(_01881_),
    .C(_01889_),
    .Y(_02830_));
 sg13g2_o21ai_1 _10264_ (.B1(_01891_),
    .Y(_02831_),
    .A1(_02830_),
    .A2(_01910_));
 sg13g2_a21o_1 _10265_ (.A2(_02829_),
    .A1(_01914_),
    .B1(_02831_),
    .X(_02832_));
 sg13g2_buf_2 _10266_ (.A(_02832_),
    .X(_02833_));
 sg13g2_nor2_2 _10267_ (.A(_01879_),
    .B(_01881_),
    .Y(_02834_));
 sg13g2_o21ai_1 _10268_ (.B1(_02834_),
    .Y(_02835_),
    .A1(_01889_),
    .A2(_02190_));
 sg13g2_a21o_1 _10269_ (.A2(_01868_),
    .A1(net326),
    .B1(_01869_),
    .X(_02836_));
 sg13g2_buf_2 _10270_ (.A(_02836_),
    .X(_02837_));
 sg13g2_o21ai_1 _10271_ (.B1(_02837_),
    .Y(_02838_),
    .A1(_01853_),
    .A2(_01859_));
 sg13g2_nor3_1 _10272_ (.A(_02837_),
    .B(_01853_),
    .C(_01859_),
    .Y(_02839_));
 sg13g2_a221oi_1 _10273_ (.B2(_02838_),
    .C1(_02839_),
    .B1(_02000_),
    .A1(_01889_),
    .Y(_02840_),
    .A2(_02190_));
 sg13g2_nand2_1 _10274_ (.Y(_02841_),
    .A(_01889_),
    .B(_02193_));
 sg13g2_o21ai_1 _10275_ (.B1(_02834_),
    .Y(_02842_),
    .A1(_01889_),
    .A2(_02193_));
 sg13g2_a221oi_1 _10276_ (.B2(_02842_),
    .C1(_01803_),
    .B1(_02841_),
    .A1(_02835_),
    .Y(_02843_),
    .A2(_02840_));
 sg13g2_a21oi_2 _10277_ (.B1(_02843_),
    .Y(_02844_),
    .A2(_02833_),
    .A1(net161));
 sg13g2_nand4_1 _10278_ (.B(_01877_),
    .C(_01914_),
    .A(_01803_),
    .Y(_02845_),
    .D(_02379_));
 sg13g2_buf_2 _10279_ (.A(_02845_),
    .X(_02846_));
 sg13g2_a22oi_1 _10280_ (.Y(_02847_),
    .B1(_02023_),
    .B2(_02026_),
    .A2(_01875_),
    .A1(_01873_));
 sg13g2_buf_1 _10281_ (.A(_02847_),
    .X(_02848_));
 sg13g2_nand3_1 _10282_ (.B(_01923_),
    .C(_02848_),
    .A(_01919_),
    .Y(_02849_));
 sg13g2_buf_2 _10283_ (.A(_02849_),
    .X(_02850_));
 sg13g2_and2_1 _10284_ (.A(_02846_),
    .B(_02850_),
    .X(_02851_));
 sg13g2_buf_1 _10285_ (.A(_02851_),
    .X(_02852_));
 sg13g2_nor2_2 _10286_ (.A(_02404_),
    .B(_02407_),
    .Y(_02853_));
 sg13g2_xnor2_1 _10287_ (.Y(_02854_),
    .A(net178),
    .B(_02853_));
 sg13g2_nand2b_1 _10288_ (.Y(_02855_),
    .B(net338),
    .A_N(\soc_I.kianv_I.datapath_unit_I.A1[3] ));
 sg13g2_or2_1 _10289_ (.X(_02856_),
    .B(_02283_),
    .A(net338));
 sg13g2_and3_1 _10290_ (.X(_02857_),
    .A(_02272_),
    .B(net308),
    .C(_02296_));
 sg13g2_or4_1 _10291_ (.A(_02299_),
    .B(_02280_),
    .C(_02447_),
    .D(_02448_),
    .X(_02858_));
 sg13g2_a221oi_1 _10292_ (.B2(_01741_),
    .C1(_02858_),
    .B1(_01736_),
    .A1(_01779_),
    .Y(_02859_),
    .A2(_02214_));
 sg13g2_a221oi_1 _10293_ (.B2(net178),
    .C1(_02859_),
    .B1(_02857_),
    .A1(_02855_),
    .Y(_02860_),
    .A2(_02856_));
 sg13g2_o21ai_1 _10294_ (.B1(_02860_),
    .Y(_02861_),
    .A1(_02401_),
    .A2(_02854_));
 sg13g2_a21oi_1 _10295_ (.A1(net337),
    .A2(_02331_),
    .Y(_02862_),
    .B1(_02332_));
 sg13g2_buf_2 _10296_ (.A(_02862_),
    .X(_02863_));
 sg13g2_nand3_1 _10297_ (.B(_02383_),
    .C(_02863_),
    .A(_02381_),
    .Y(_02864_));
 sg13g2_buf_1 _10298_ (.A(_02864_),
    .X(_02865_));
 sg13g2_or2_1 _10299_ (.X(_02866_),
    .B(_02341_),
    .A(_02336_));
 sg13g2_buf_2 _10300_ (.A(_02866_),
    .X(_02867_));
 sg13g2_nand3_1 _10301_ (.B(_02386_),
    .C(_02388_),
    .A(_02867_),
    .Y(_02868_));
 sg13g2_buf_2 _10302_ (.A(_02868_),
    .X(_02869_));
 sg13g2_a22oi_1 _10303_ (.Y(_02870_),
    .B1(_02869_),
    .B2(_02470_),
    .A2(_02865_),
    .A1(_02351_));
 sg13g2_buf_1 _10304_ (.A(_02870_),
    .X(_02871_));
 sg13g2_nand2_1 _10305_ (.Y(_02872_),
    .A(_02361_),
    .B(_02363_));
 sg13g2_buf_2 _10306_ (.A(_02872_),
    .X(_02873_));
 sg13g2_nor3_1 _10307_ (.A(_02873_),
    .B(_02433_),
    .C(_02435_),
    .Y(_02874_));
 sg13g2_nand2_1 _10308_ (.Y(_02875_),
    .A(_02367_),
    .B(_02371_));
 sg13g2_buf_2 _10309_ (.A(_02875_),
    .X(_02876_));
 sg13g2_a21oi_1 _10310_ (.A1(_02355_),
    .A2(_02375_),
    .Y(_02877_),
    .B1(_02876_));
 sg13g2_nand4_1 _10311_ (.B(_02871_),
    .C(_02874_),
    .A(net180),
    .Y(_02878_),
    .D(_02877_));
 sg13g2_o21ai_1 _10312_ (.B1(_02867_),
    .Y(_02879_),
    .A1(_02347_),
    .A2(_02348_));
 sg13g2_a22oi_1 _10313_ (.Y(_02880_),
    .B1(_02457_),
    .B2(_02879_),
    .A2(_02443_),
    .A1(_02441_));
 sg13g2_buf_1 _10314_ (.A(_02880_),
    .X(_02881_));
 sg13g2_a21oi_1 _10315_ (.A1(_02381_),
    .A2(_02383_),
    .Y(_02882_),
    .B1(_02863_));
 sg13g2_and2_1 _10316_ (.A(_02361_),
    .B(_02363_),
    .X(_02883_));
 sg13g2_buf_1 _10317_ (.A(_02883_),
    .X(_02884_));
 sg13g2_nor3_1 _10318_ (.A(_02882_),
    .B(_02335_),
    .C(_02884_),
    .Y(_02885_));
 sg13g2_and3_1 _10319_ (.X(_02886_),
    .A(_02355_),
    .B(_02876_),
    .C(_02375_));
 sg13g2_nand4_1 _10320_ (.B(_02881_),
    .C(_02885_),
    .A(net178),
    .Y(_02887_),
    .D(_02886_));
 sg13g2_a21oi_1 _10321_ (.A1(_02296_),
    .A2(_02301_),
    .Y(_02888_),
    .B1(_02415_));
 sg13g2_nor2_1 _10322_ (.A(_02408_),
    .B(_02888_),
    .Y(_02889_));
 sg13g2_nor2_1 _10323_ (.A(_02447_),
    .B(_02448_),
    .Y(_02890_));
 sg13g2_buf_2 _10324_ (.A(_02890_),
    .X(_02891_));
 sg13g2_a22oi_1 _10325_ (.Y(_02892_),
    .B1(_02311_),
    .B2(_02891_),
    .A2(_02853_),
    .A1(_02401_));
 sg13g2_nor3_1 _10326_ (.A(_01754_),
    .B(_02460_),
    .C(_02892_),
    .Y(_02893_));
 sg13g2_a221oi_1 _10327_ (.B2(net179),
    .C1(_02893_),
    .B1(_02889_),
    .A1(_02878_),
    .Y(_02894_),
    .A2(_02887_));
 sg13g2_nand2_2 _10328_ (.Y(_02895_),
    .A(_02446_),
    .B(_02444_));
 sg13g2_xnor2_1 _10329_ (.Y(_02896_),
    .A(_02285_),
    .B(_02891_));
 sg13g2_buf_2 _10330_ (.A(_02896_),
    .X(_02897_));
 sg13g2_nand4_1 _10331_ (.B(_02313_),
    .C(_02895_),
    .A(net178),
    .Y(_02898_),
    .D(_02897_));
 sg13g2_buf_1 _10332_ (.A(_02898_),
    .X(_02899_));
 sg13g2_nand2_1 _10333_ (.Y(_02900_),
    .A(_02299_),
    .B(net308));
 sg13g2_nor2_1 _10334_ (.A(_02408_),
    .B(_02415_),
    .Y(_02901_));
 sg13g2_xnor2_1 _10335_ (.Y(_02902_),
    .A(_02285_),
    .B(_02296_));
 sg13g2_buf_1 _10336_ (.A(_02902_),
    .X(_02903_));
 sg13g2_nand4_1 _10337_ (.B(_02900_),
    .C(_02901_),
    .A(net180),
    .Y(_02904_),
    .D(net183));
 sg13g2_buf_1 _10338_ (.A(_02904_),
    .X(_02905_));
 sg13g2_a22oi_1 _10339_ (.Y(_02906_),
    .B1(_02899_),
    .B2(_02905_),
    .A2(_02887_),
    .A1(_02878_));
 sg13g2_a221oi_1 _10340_ (.B2(_01741_),
    .C1(_01686_),
    .B1(_01736_),
    .A1(_01779_),
    .Y(_02907_),
    .A2(_02214_));
 sg13g2_o21ai_1 _10341_ (.B1(_01719_),
    .Y(_02908_),
    .A1(_01775_),
    .A2(_02907_));
 sg13g2_nand3_1 _10342_ (.B(_01917_),
    .C(_02317_),
    .A(_01686_),
    .Y(_02909_));
 sg13g2_o21ai_1 _10343_ (.B1(_02307_),
    .Y(_02910_),
    .A1(_01718_),
    .A2(_01754_));
 sg13g2_and3_1 _10344_ (.X(_02911_),
    .A(_02908_),
    .B(_02909_),
    .C(_02910_));
 sg13g2_buf_2 _10345_ (.A(_02911_),
    .X(_02912_));
 sg13g2_a22oi_1 _10346_ (.Y(_02913_),
    .B1(_02906_),
    .B2(_02912_),
    .A2(_02894_),
    .A1(_02861_));
 sg13g2_buf_2 _10347_ (.A(_02913_),
    .X(_02914_));
 sg13g2_a21o_1 _10348_ (.A2(_02833_),
    .A1(_01804_),
    .B1(_02843_),
    .X(_02915_));
 sg13g2_nor2_2 _10349_ (.A(_02347_),
    .B(_02348_),
    .Y(_02916_));
 sg13g2_o21ai_1 _10350_ (.B1(_02916_),
    .Y(_02917_),
    .A1(_02343_),
    .A2(_02433_));
 sg13g2_nand2_1 _10351_ (.Y(_02918_),
    .A(_02419_),
    .B(_02423_));
 sg13g2_nor4_2 _10352_ (.A(_02336_),
    .B(_02341_),
    .C(_02424_),
    .Y(_02919_),
    .D(_02461_));
 sg13g2_nor2_2 _10353_ (.A(_02325_),
    .B(_02329_),
    .Y(_02920_));
 sg13g2_a221oi_1 _10354_ (.B2(_02919_),
    .C1(_02920_),
    .B1(_02918_),
    .A1(_02357_),
    .Y(_02921_),
    .A2(_02359_));
 sg13g2_nand2_2 _10355_ (.Y(_02922_),
    .A(_02357_),
    .B(_02359_));
 sg13g2_nor2_1 _10356_ (.A(_02863_),
    .B(_02922_),
    .Y(_02923_));
 sg13g2_nand2_1 _10357_ (.Y(_02924_),
    .A(_02863_),
    .B(_02922_));
 sg13g2_nand2_2 _10358_ (.Y(_02925_),
    .A(_02012_),
    .B(_02014_));
 sg13g2_a22oi_1 _10359_ (.Y(_02926_),
    .B1(_02924_),
    .B2(_02925_),
    .A2(_02923_),
    .A1(_02920_));
 sg13g2_a21o_1 _10360_ (.A2(_02921_),
    .A1(_02917_),
    .B1(_02926_),
    .X(_02927_));
 sg13g2_a21oi_1 _10361_ (.A1(_02920_),
    .A2(_02363_),
    .Y(_02928_),
    .B1(_02923_));
 sg13g2_nor3_1 _10362_ (.A(_02867_),
    .B(_02347_),
    .C(_02348_),
    .Y(_02929_));
 sg13g2_a221oi_1 _10363_ (.B2(_02918_),
    .C1(_02929_),
    .B1(_02919_),
    .A1(_02916_),
    .Y(_02930_),
    .A2(_02433_));
 sg13g2_buf_1 _10364_ (.A(_02930_),
    .X(_02931_));
 sg13g2_or2_1 _10365_ (.X(_02932_),
    .B(_02931_),
    .A(_02928_));
 sg13g2_nand2_1 _10366_ (.Y(_02933_),
    .A(net171),
    .B(_02877_));
 sg13g2_a21oi_1 _10367_ (.A1(_02927_),
    .A2(_02932_),
    .Y(_02934_),
    .B1(_02933_));
 sg13g2_nand2_1 _10368_ (.Y(_02935_),
    .A(_01942_),
    .B(_01949_));
 sg13g2_and2_1 _10369_ (.A(_01927_),
    .B(_01955_),
    .X(_02936_));
 sg13g2_nor2b_1 _10370_ (.A(_02935_),
    .B_N(_02936_),
    .Y(_02937_));
 sg13g2_a21oi_1 _10371_ (.A1(_02375_),
    .A2(_02937_),
    .Y(_02938_),
    .B1(_01999_));
 sg13g2_a21oi_1 _10372_ (.A1(_01991_),
    .A2(_01994_),
    .Y(_02939_),
    .B1(_01963_));
 sg13g2_nand3_1 _10373_ (.B(_01994_),
    .C(_01963_),
    .A(_01991_),
    .Y(_02940_));
 sg13g2_buf_1 _10374_ (.A(_02940_),
    .X(_02941_));
 sg13g2_o21ai_1 _10375_ (.B1(_02941_),
    .Y(_02942_),
    .A1(_02939_),
    .A2(_02367_));
 sg13g2_nand2_1 _10376_ (.Y(_02943_),
    .A(_01756_),
    .B(_02942_));
 sg13g2_o21ai_1 _10377_ (.B1(_02943_),
    .Y(_02944_),
    .A1(_01804_),
    .A2(_02938_));
 sg13g2_and2_1 _10378_ (.A(_02367_),
    .B(_02371_),
    .X(_02945_));
 sg13g2_buf_1 _10379_ (.A(_02945_),
    .X(_02946_));
 sg13g2_nand2_1 _10380_ (.Y(_02947_),
    .A(_02355_),
    .B(_02375_));
 sg13g2_nand2_1 _10381_ (.Y(_02948_),
    .A(_02381_),
    .B(_02383_));
 sg13g2_a21oi_1 _10382_ (.A1(_02386_),
    .A2(_02388_),
    .Y(_02949_),
    .B1(_02867_));
 sg13g2_and3_1 _10383_ (.X(_02950_),
    .A(_02419_),
    .B(_02423_),
    .C(_02919_));
 sg13g2_or2_1 _10384_ (.X(_02951_),
    .B(_01666_),
    .A(_02420_));
 sg13g2_a221oi_1 _10385_ (.B2(_02951_),
    .C1(_02465_),
    .B1(_02421_),
    .A1(_02386_),
    .Y(_02952_),
    .A2(_02388_));
 sg13g2_or4_1 _10386_ (.A(_02948_),
    .B(_02949_),
    .C(_02950_),
    .D(_02952_),
    .X(_02953_));
 sg13g2_nor2_1 _10387_ (.A(_02925_),
    .B(_02922_),
    .Y(_02954_));
 sg13g2_nor2_1 _10388_ (.A(_02863_),
    .B(_02954_),
    .Y(_02955_));
 sg13g2_nor2_1 _10389_ (.A(_02920_),
    .B(_02954_),
    .Y(_02956_));
 sg13g2_or3_1 _10390_ (.A(_02949_),
    .B(_02950_),
    .C(_02952_),
    .X(_02957_));
 sg13g2_buf_1 _10391_ (.A(_02957_),
    .X(_02958_));
 sg13g2_and2_1 _10392_ (.A(_02925_),
    .B(_02922_),
    .X(_02959_));
 sg13g2_buf_1 _10393_ (.A(_02959_),
    .X(_02960_));
 sg13g2_a221oi_1 _10394_ (.B2(_02958_),
    .C1(_02960_),
    .B1(_02956_),
    .A1(_02953_),
    .Y(_02961_),
    .A2(_02955_));
 sg13g2_buf_1 _10395_ (.A(_02961_),
    .X(_02962_));
 sg13g2_nor4_1 _10396_ (.A(_01756_),
    .B(_02946_),
    .C(_02947_),
    .D(_02962_),
    .Y(_02963_));
 sg13g2_nor4_1 _10397_ (.A(_02915_),
    .B(_02934_),
    .C(_02944_),
    .D(_02963_),
    .Y(_02964_));
 sg13g2_a22oi_1 _10398_ (.Y(_02965_),
    .B1(_01833_),
    .B2(_01835_),
    .A2(_02158_),
    .A1(net269));
 sg13g2_buf_1 _10399_ (.A(_02965_),
    .X(_02966_));
 sg13g2_and3_1 _10400_ (.X(_02967_),
    .A(net169),
    .B(_02162_),
    .C(_02966_));
 sg13g2_nand4_1 _10401_ (.B(_02158_),
    .C(_01833_),
    .A(net269),
    .Y(_02968_),
    .D(_01835_));
 sg13g2_buf_2 _10402_ (.A(_02968_),
    .X(_02969_));
 sg13g2_nor3_1 _10403_ (.A(net169),
    .B(_02144_),
    .C(_02969_),
    .Y(_02970_));
 sg13g2_or2_1 _10404_ (.X(_02971_),
    .B(_02970_),
    .A(_02967_));
 sg13g2_buf_2 _10405_ (.A(_02971_),
    .X(_02972_));
 sg13g2_nand2_1 _10406_ (.Y(_02973_),
    .A(net179),
    .B(_02802_));
 sg13g2_nand2_1 _10407_ (.Y(_02974_),
    .A(net169),
    .B(_02804_));
 sg13g2_nand4_1 _10408_ (.B(_02091_),
    .C(_02771_),
    .A(net178),
    .Y(_02975_),
    .D(_02805_));
 sg13g2_buf_1 _10409_ (.A(_02975_),
    .X(_02976_));
 sg13g2_and3_1 _10410_ (.X(_02977_),
    .A(_02056_),
    .B(_02108_),
    .C(net271));
 sg13g2_buf_1 _10411_ (.A(_02977_),
    .X(_02978_));
 sg13g2_and2_1 _10412_ (.A(net272),
    .B(_02800_),
    .X(_02979_));
 sg13g2_nand4_1 _10413_ (.B(_02095_),
    .C(_02978_),
    .A(net180),
    .Y(_02980_),
    .D(_02979_));
 sg13g2_buf_1 _10414_ (.A(_02980_),
    .X(_02981_));
 sg13g2_a22oi_1 _10415_ (.Y(_02982_),
    .B1(_02976_),
    .B2(_02981_),
    .A2(_02974_),
    .A1(_02973_));
 sg13g2_buf_1 _10416_ (.A(_02982_),
    .X(_02983_));
 sg13g2_nand3_1 _10417_ (.B(_02972_),
    .C(_02983_),
    .A(_02809_),
    .Y(_02984_));
 sg13g2_a221oi_1 _10418_ (.B2(_02964_),
    .C1(_02984_),
    .B1(net146),
    .A1(_02844_),
    .Y(_02985_),
    .A2(_02852_));
 sg13g2_buf_1 _10419_ (.A(_02985_),
    .X(_02986_));
 sg13g2_nor2_1 _10420_ (.A(_02827_),
    .B(_02986_),
    .Y(_02987_));
 sg13g2_xnor2_1 _10421_ (.Y(_02988_),
    .A(_02652_),
    .B(_02663_));
 sg13g2_xor2_1 _10422_ (.B(_02988_),
    .A(_02987_),
    .X(_02989_));
 sg13g2_and2_1 _10423_ (.A(net167),
    .B(_02706_),
    .X(_02990_));
 sg13g2_a22oi_1 _10424_ (.Y(_02991_),
    .B1(_02990_),
    .B2(_02691_),
    .A2(_02989_),
    .A1(_02713_));
 sg13g2_a21o_1 _10425_ (.A2(_02991_),
    .A1(_02711_),
    .B1(net315),
    .X(_02992_));
 sg13g2_nand2b_1 _10426_ (.Y(_02993_),
    .B(_02706_),
    .A_N(_02713_));
 sg13g2_a21oi_1 _10427_ (.A1(_02620_),
    .A2(_02690_),
    .Y(_02994_),
    .B1(_02993_));
 sg13g2_o21ai_1 _10428_ (.B1(_02994_),
    .Y(_02995_),
    .A1(net167),
    .A2(_02710_));
 sg13g2_o21ai_1 _10429_ (.B1(_02713_),
    .Y(_02996_),
    .A1(_02712_),
    .A2(_02710_));
 sg13g2_a21oi_2 _10430_ (.B1(_02689_),
    .Y(_02997_),
    .A2(_02619_),
    .A1(_02234_));
 sg13g2_nor2_1 _10431_ (.A(net305),
    .B(_02705_),
    .Y(_02998_));
 sg13g2_nor2b_1 _10432_ (.A(_02997_),
    .B_N(_02998_),
    .Y(_02999_));
 sg13g2_buf_1 _10433_ (.A(net152),
    .X(_03000_));
 sg13g2_o21ai_1 _10434_ (.B1(net145),
    .Y(_03001_),
    .A1(_02679_),
    .A2(_02662_));
 sg13g2_o21ai_1 _10435_ (.B1(net305),
    .Y(_03002_),
    .A1(_02997_),
    .A2(_03001_));
 sg13g2_o21ai_1 _10436_ (.B1(_03002_),
    .Y(_03003_),
    .A1(_02696_),
    .A2(_02999_));
 sg13g2_mux2_1 _10437_ (.A0(_02995_),
    .A1(_02996_),
    .S(_03003_),
    .X(_03004_));
 sg13g2_buf_1 _10438_ (.A(_01764_),
    .X(_03005_));
 sg13g2_nor3_1 _10439_ (.A(_01721_),
    .B(net263),
    .C(net315),
    .Y(_03006_));
 sg13g2_buf_1 _10440_ (.A(net147),
    .X(_03007_));
 sg13g2_a21oi_2 _10441_ (.B1(_02474_),
    .Y(_03008_),
    .A2(_02453_),
    .A1(_02321_));
 sg13g2_nor2_1 _10442_ (.A(_02199_),
    .B(_02029_),
    .Y(_03009_));
 sg13g2_nor2_1 _10443_ (.A(_02199_),
    .B(_01925_),
    .Y(_03010_));
 sg13g2_a21oi_1 _10444_ (.A1(_03008_),
    .A2(_03009_),
    .Y(_03011_),
    .B1(_03010_));
 sg13g2_xnor2_1 _10445_ (.Y(_03012_),
    .A(_02159_),
    .B(_03011_));
 sg13g2_buf_8 _10446_ (.A(net160),
    .X(_03013_));
 sg13g2_buf_8 _10447_ (.A(net154),
    .X(_03014_));
 sg13g2_nand2_1 _10448_ (.Y(_03015_),
    .A(_02927_),
    .B(_02932_));
 sg13g2_nand2_1 _10449_ (.Y(_03016_),
    .A(net150),
    .B(_02962_));
 sg13g2_o21ai_1 _10450_ (.B1(_03016_),
    .Y(_03017_),
    .A1(net150),
    .A2(_03015_));
 sg13g2_buf_1 _10451_ (.A(_03017_),
    .X(_03018_));
 sg13g2_nand3_1 _10452_ (.B(_02871_),
    .C(_02874_),
    .A(_01757_),
    .Y(_03019_));
 sg13g2_nand3_1 _10453_ (.B(_02881_),
    .C(_02885_),
    .A(_02439_),
    .Y(_03020_));
 sg13g2_a221oi_1 _10454_ (.B2(_03020_),
    .C1(_02893_),
    .B1(_03019_),
    .A1(net158),
    .Y(_03021_),
    .A2(_02889_));
 sg13g2_a22oi_1 _10455_ (.Y(_03022_),
    .B1(_03019_),
    .B2(_03020_),
    .A2(_02905_),
    .A1(_02899_));
 sg13g2_a22oi_1 _10456_ (.Y(_03023_),
    .B1(_03022_),
    .B2(_02912_),
    .A2(_03021_),
    .A1(_02861_));
 sg13g2_buf_2 _10457_ (.A(_03023_),
    .X(_03024_));
 sg13g2_nand2_1 _10458_ (.Y(_03025_),
    .A(_03018_),
    .B(_03024_));
 sg13g2_xnor2_1 _10459_ (.Y(_03026_),
    .A(_02876_),
    .B(_03025_));
 sg13g2_a22oi_1 _10460_ (.Y(_03027_),
    .B1(_02259_),
    .B2(_02266_),
    .A2(_02251_),
    .A1(_02249_));
 sg13g2_buf_1 _10461_ (.A(_03027_),
    .X(_03028_));
 sg13g2_nor2_1 _10462_ (.A(_03028_),
    .B(_02641_),
    .Y(_03029_));
 sg13g2_nand3b_1 _10463_ (.B(_02232_),
    .C(_03029_),
    .Y(_03030_),
    .A_N(_02478_));
 sg13g2_nand4_1 _10464_ (.B(_02232_),
    .C(_03008_),
    .A(_02166_),
    .Y(_03031_),
    .D(_03029_));
 sg13g2_a21o_1 _10465_ (.A2(_02232_),
    .A1(_02166_),
    .B1(_02800_),
    .X(_03032_));
 sg13g2_and3_1 _10466_ (.X(_03033_),
    .A(_01925_),
    .B(_02165_),
    .C(_02641_));
 sg13g2_a22oi_1 _10467_ (.Y(_03034_),
    .B1(_03033_),
    .B2(_02476_),
    .A2(_02641_),
    .A1(_03028_));
 sg13g2_nand4_1 _10468_ (.B(_03031_),
    .C(_03032_),
    .A(_03030_),
    .Y(_03035_),
    .D(_03034_));
 sg13g2_buf_2 _10469_ (.A(_03035_),
    .X(_03036_));
 sg13g2_nor4_1 _10470_ (.A(net142),
    .B(_03012_),
    .C(_03026_),
    .D(_03036_),
    .Y(_03037_));
 sg13g2_and4_1 _10471_ (.A(net142),
    .B(_03012_),
    .C(_03026_),
    .D(_03036_),
    .X(_03038_));
 sg13g2_nand2_1 _10472_ (.Y(_03039_),
    .A(_02140_),
    .B(_02142_));
 sg13g2_nand4_1 _10473_ (.B(_01896_),
    .C(_01833_),
    .A(_01891_),
    .Y(_03040_),
    .D(_01835_));
 sg13g2_or3_1 _10474_ (.A(_01919_),
    .B(_02159_),
    .C(_03040_),
    .X(_03041_));
 sg13g2_a22oi_1 _10475_ (.Y(_03042_),
    .B1(_02158_),
    .B2(net269),
    .A2(_02142_),
    .A1(net270));
 sg13g2_nand3_1 _10476_ (.B(_02196_),
    .C(_03042_),
    .A(_01920_),
    .Y(_03043_));
 sg13g2_o21ai_1 _10477_ (.B1(_03043_),
    .Y(_03044_),
    .A1(_03039_),
    .A2(_03041_));
 sg13g2_buf_1 _10478_ (.A(_03044_),
    .X(_03045_));
 sg13g2_a21o_1 _10479_ (.A2(_01999_),
    .A1(_01986_),
    .B1(_02000_),
    .X(_03046_));
 sg13g2_a22oi_1 _10480_ (.Y(_03047_),
    .B1(_01912_),
    .B2(_01910_),
    .A2(_01875_),
    .A1(_01873_));
 sg13g2_a221oi_1 _10481_ (.B2(_03047_),
    .C1(_02194_),
    .B1(_03046_),
    .A1(_02170_),
    .Y(_03048_),
    .A2(_01908_));
 sg13g2_and2_1 _10482_ (.A(_01910_),
    .B(_01912_),
    .X(_03049_));
 sg13g2_buf_1 _10483_ (.A(_03049_),
    .X(_03050_));
 sg13g2_nor2_2 _10484_ (.A(_01973_),
    .B(_01976_),
    .Y(_03051_));
 sg13g2_nand2_1 _10485_ (.Y(_03052_),
    .A(_03051_),
    .B(_02941_));
 sg13g2_o21ai_1 _10486_ (.B1(_01984_),
    .Y(_03053_),
    .A1(_03051_),
    .A2(_02941_));
 sg13g2_nand4_1 _10487_ (.B(_03050_),
    .C(_03052_),
    .A(_01877_),
    .Y(_03054_),
    .D(_03053_));
 sg13g2_a21oi_1 _10488_ (.A1(_02171_),
    .A2(_02174_),
    .Y(_03055_),
    .B1(net168));
 sg13g2_a22oi_1 _10489_ (.Y(_03056_),
    .B1(_03054_),
    .B2(_03055_),
    .A2(_03048_),
    .A1(_01920_));
 sg13g2_a21oi_1 _10490_ (.A1(_02188_),
    .A2(_03042_),
    .Y(_03057_),
    .B1(_02221_));
 sg13g2_and4_1 _10491_ (.A(net269),
    .B(net270),
    .C(_02142_),
    .D(_02158_),
    .X(_03058_));
 sg13g2_a221oi_1 _10492_ (.B2(_03058_),
    .C1(net168),
    .B1(_02178_),
    .A1(_02207_),
    .Y(_03059_),
    .A2(_02208_));
 sg13g2_a21oi_1 _10493_ (.A1(net160),
    .A2(_03057_),
    .Y(_03060_),
    .B1(_03059_));
 sg13g2_a21o_1 _10494_ (.A2(_03056_),
    .A1(_03045_),
    .B1(_03060_),
    .X(_03061_));
 sg13g2_buf_1 _10495_ (.A(_03061_),
    .X(_03062_));
 sg13g2_nand3_1 _10496_ (.B(_02909_),
    .C(_02910_),
    .A(_02908_),
    .Y(_03063_));
 sg13g2_buf_2 _10497_ (.A(_03063_),
    .X(_03064_));
 sg13g2_nand2_1 _10498_ (.Y(_03065_),
    .A(_01918_),
    .B(_02895_));
 sg13g2_nand2_1 _10499_ (.Y(_03066_),
    .A(_02441_),
    .B(_02443_));
 sg13g2_o21ai_1 _10500_ (.B1(_02863_),
    .Y(_03067_),
    .A1(_02325_),
    .A2(_02329_));
 sg13g2_a22oi_1 _10501_ (.Y(_03068_),
    .B1(_02879_),
    .B2(_02457_),
    .A2(_03067_),
    .A1(_02391_));
 sg13g2_nor3_1 _10502_ (.A(_02272_),
    .B(_02280_),
    .C(net266),
    .Y(_03069_));
 sg13g2_o21ai_1 _10503_ (.B1(net266),
    .Y(_03070_),
    .A1(_02272_),
    .A2(net308));
 sg13g2_o21ai_1 _10504_ (.B1(_03070_),
    .Y(_03071_),
    .A1(_02891_),
    .A2(_03069_));
 sg13g2_nand4_1 _10505_ (.B(_03066_),
    .C(_03068_),
    .A(_02373_),
    .Y(_03072_),
    .D(_03071_));
 sg13g2_or2_1 _10506_ (.X(_03073_),
    .B(_03072_),
    .A(_03065_));
 sg13g2_a221oi_1 _10507_ (.B2(_02470_),
    .C1(_02394_),
    .B1(_02869_),
    .A1(_02351_),
    .Y(_03074_),
    .A2(_02865_));
 sg13g2_and2_1 _10508_ (.A(_02299_),
    .B(_02280_),
    .X(_03075_));
 sg13g2_nand2_1 _10509_ (.Y(_03076_),
    .A(_02302_),
    .B(_03075_));
 sg13g2_nand3b_1 _10510_ (.B(_03074_),
    .C(_03076_),
    .Y(_03077_),
    .A_N(_02438_));
 sg13g2_nor3_1 _10511_ (.A(net156),
    .B(_01922_),
    .C(_02353_),
    .Y(_03078_));
 sg13g2_nand2_1 _10512_ (.Y(_03079_),
    .A(_01910_),
    .B(_01912_));
 sg13g2_and2_1 _10513_ (.A(_02355_),
    .B(_02375_),
    .X(_03080_));
 sg13g2_buf_2 _10514_ (.A(_03080_),
    .X(_03081_));
 sg13g2_nand4_1 _10515_ (.B(net270),
    .C(_02142_),
    .A(net269),
    .Y(_03082_),
    .D(_02158_));
 sg13g2_nor4_1 _10516_ (.A(_03040_),
    .B(_03079_),
    .C(_03081_),
    .D(_03082_),
    .Y(_03083_));
 sg13g2_nor4_1 _10517_ (.A(_01877_),
    .B(_03050_),
    .C(_02379_),
    .D(_02947_),
    .Y(_03084_));
 sg13g2_and3_1 _10518_ (.X(_03085_),
    .A(net154),
    .B(_02196_),
    .C(_03042_));
 sg13g2_a22oi_1 _10519_ (.Y(_03086_),
    .B1(_03084_),
    .B2(_03085_),
    .A2(_03083_),
    .A1(_03078_));
 sg13g2_a221oi_1 _10520_ (.B2(_03077_),
    .C1(_03086_),
    .B1(_03073_),
    .A1(_02305_),
    .Y(_03087_),
    .A2(_03064_));
 sg13g2_buf_1 _10521_ (.A(_03087_),
    .X(_03088_));
 sg13g2_and2_1 _10522_ (.A(net180),
    .B(_02018_),
    .X(_03089_));
 sg13g2_nor2_1 _10523_ (.A(_02873_),
    .B(_02876_),
    .Y(_03090_));
 sg13g2_a22oi_1 _10524_ (.Y(_03091_),
    .B1(_03074_),
    .B2(_02455_),
    .A2(_02458_),
    .A1(_03090_));
 sg13g2_nor2_2 _10525_ (.A(_02882_),
    .B(_02335_),
    .Y(_03092_));
 sg13g2_nor2_1 _10526_ (.A(_02349_),
    .B(_02949_),
    .Y(_03093_));
 sg13g2_nand4_1 _10527_ (.B(_02468_),
    .C(_03092_),
    .A(_02373_),
    .Y(_03094_),
    .D(_03093_));
 sg13g2_a221oi_1 _10528_ (.B2(_02472_),
    .C1(net180),
    .B1(_02373_),
    .A1(net363),
    .Y(_03095_),
    .A2(_01958_));
 sg13g2_a22oi_1 _10529_ (.Y(_03096_),
    .B1(_03094_),
    .B2(_03095_),
    .A2(_03091_),
    .A1(_03089_));
 sg13g2_buf_2 _10530_ (.A(_03096_),
    .X(_03097_));
 sg13g2_nor2b_1 _10531_ (.A(_03086_),
    .B_N(_03097_),
    .Y(_03098_));
 sg13g2_xnor2_1 _10532_ (.Y(_03099_),
    .A(_02555_),
    .B(_02625_));
 sg13g2_nand3_1 _10533_ (.B(_02265_),
    .C(_02645_),
    .A(net179),
    .Y(_03100_));
 sg13g2_o21ai_1 _10534_ (.B1(_02250_),
    .Y(_03101_),
    .A1(_02244_),
    .A2(_02245_));
 sg13g2_nand3_1 _10535_ (.B(_02643_),
    .C(_03101_),
    .A(net169),
    .Y(_03102_));
 sg13g2_nand4_1 _10536_ (.B(_02512_),
    .C(_03100_),
    .A(_02507_),
    .Y(_03103_),
    .D(_03102_));
 sg13g2_buf_1 _10537_ (.A(_03103_),
    .X(_03104_));
 sg13g2_a21oi_1 _10538_ (.A1(_02057_),
    .A2(_02229_),
    .Y(_03105_),
    .B1(_02242_));
 sg13g2_nand3_1 _10539_ (.B(_02088_),
    .C(_02643_),
    .A(net157),
    .Y(_03106_));
 sg13g2_nand3_1 _10540_ (.B(_02095_),
    .C(_02645_),
    .A(net158),
    .Y(_03107_));
 sg13g2_a221oi_1 _10541_ (.B2(_02258_),
    .C1(net168),
    .B1(_02257_),
    .A1(_02097_),
    .Y(_03108_),
    .A2(_02211_));
 sg13g2_a221oi_1 _10542_ (.B2(_03107_),
    .C1(_03108_),
    .B1(_03106_),
    .A1(net151),
    .Y(_03109_),
    .A2(_03105_));
 sg13g2_buf_1 _10543_ (.A(_03109_),
    .X(_03110_));
 sg13g2_or3_1 _10544_ (.A(_03099_),
    .B(_03104_),
    .C(_03110_),
    .X(_03111_));
 sg13g2_or4_1 _10545_ (.A(_03062_),
    .B(_03088_),
    .C(_03098_),
    .D(_03111_),
    .X(_03112_));
 sg13g2_or2_1 _10546_ (.X(_03113_),
    .B(_03110_),
    .A(_03104_));
 sg13g2_nand3_1 _10547_ (.B(_02057_),
    .C(_02222_),
    .A(net168),
    .Y(_03114_));
 sg13g2_nand4_1 _10548_ (.B(_02097_),
    .C(_02201_),
    .A(net179),
    .Y(_03115_),
    .D(_02203_));
 sg13g2_a22oi_1 _10549_ (.Y(_03116_),
    .B1(_03114_),
    .B2(_03115_),
    .A2(_03107_),
    .A1(_03106_));
 sg13g2_and2_1 _10550_ (.A(_03099_),
    .B(_03116_),
    .X(_03117_));
 sg13g2_nor4_1 _10551_ (.A(_03099_),
    .B(_03104_),
    .C(_03110_),
    .D(_03116_),
    .Y(_03118_));
 sg13g2_a221oi_1 _10552_ (.B2(_03117_),
    .C1(_03118_),
    .B1(_03062_),
    .A1(_03099_),
    .Y(_03119_),
    .A2(_03113_));
 sg13g2_o21ai_1 _10553_ (.B1(_03117_),
    .Y(_03120_),
    .A1(_03088_),
    .A2(_03098_));
 sg13g2_and3_1 _10554_ (.X(_03121_),
    .A(_03112_),
    .B(_03119_),
    .C(_03120_));
 sg13g2_mux2_1 _10555_ (.A0(_03037_),
    .A1(_03038_),
    .S(_03121_),
    .X(_03122_));
 sg13g2_xnor2_1 _10556_ (.Y(_03123_),
    .A(net145),
    .B(_02168_));
 sg13g2_nand2_1 _10557_ (.Y(_03124_),
    .A(_03114_),
    .B(_03115_));
 sg13g2_a21oi_1 _10558_ (.A1(net156),
    .A2(_03105_),
    .Y(_03125_),
    .B1(_03108_));
 sg13g2_a21oi_1 _10559_ (.A1(_03124_),
    .A2(_03060_),
    .Y(_03126_),
    .B1(_03125_));
 sg13g2_buf_1 _10560_ (.A(_03126_),
    .X(_03127_));
 sg13g2_nand2_1 _10561_ (.Y(_03128_),
    .A(_03124_),
    .B(_03045_));
 sg13g2_xnor2_1 _10562_ (.Y(_03129_),
    .A(net142),
    .B(_02072_));
 sg13g2_a21o_1 _10563_ (.A2(_03128_),
    .A1(net141),
    .B1(_03129_),
    .X(_03130_));
 sg13g2_nand3_1 _10564_ (.B(_03129_),
    .C(_03128_),
    .A(net141),
    .Y(_03131_));
 sg13g2_nand2_1 _10565_ (.Y(_03132_),
    .A(_02305_),
    .B(_03064_));
 sg13g2_nor3_1 _10566_ (.A(_02394_),
    .B(_02433_),
    .C(_02435_),
    .Y(_03133_));
 sg13g2_a221oi_1 _10567_ (.B2(_03075_),
    .C1(_01752_),
    .B1(_02302_),
    .A1(_01736_),
    .Y(_03134_),
    .A2(_01741_));
 sg13g2_nand4_1 _10568_ (.B(_02871_),
    .C(_03133_),
    .A(_02417_),
    .Y(_03135_),
    .D(_03134_));
 sg13g2_o21ai_1 _10569_ (.B1(_03135_),
    .Y(_03136_),
    .A1(_03065_),
    .A2(_03072_));
 sg13g2_buf_1 _10570_ (.A(_03136_),
    .X(_03137_));
 sg13g2_xnor2_1 _10571_ (.Y(_03138_),
    .A(_01755_),
    .B(_02170_));
 sg13g2_nand3_1 _10572_ (.B(_02379_),
    .C(_02947_),
    .A(_01755_),
    .Y(_03139_));
 sg13g2_nand3_1 _10573_ (.B(_02353_),
    .C(_03081_),
    .A(_01918_),
    .Y(_03140_));
 sg13g2_or2_1 _10574_ (.X(_03141_),
    .B(_02838_),
    .A(_02190_));
 sg13g2_a221oi_1 _10575_ (.B2(_02828_),
    .C1(_01752_),
    .B1(_01910_),
    .A1(_01736_),
    .Y(_03142_),
    .A2(_01741_));
 sg13g2_a21oi_1 _10576_ (.A1(_02030_),
    .A2(_03141_),
    .Y(_03143_),
    .B1(_03142_));
 sg13g2_a221oi_1 _10577_ (.B2(_03140_),
    .C1(_03143_),
    .B1(_03139_),
    .A1(_02173_),
    .Y(_03144_),
    .A2(_03138_));
 sg13g2_and2_1 _10578_ (.A(_03137_),
    .B(_03144_),
    .X(_03145_));
 sg13g2_a21o_1 _10579_ (.A2(_03144_),
    .A1(_03097_),
    .B1(_03056_),
    .X(_03146_));
 sg13g2_a21oi_1 _10580_ (.A1(_03132_),
    .A2(_03145_),
    .Y(_03147_),
    .B1(_03146_));
 sg13g2_a21oi_1 _10581_ (.A1(_03130_),
    .A2(_03131_),
    .Y(_03148_),
    .B1(_03147_));
 sg13g2_a21o_1 _10582_ (.A2(_03145_),
    .A1(_03132_),
    .B1(_03146_),
    .X(_03149_));
 sg13g2_buf_8 _10583_ (.A(_03149_),
    .X(_03150_));
 sg13g2_xnor2_1 _10584_ (.Y(_03151_),
    .A(net152),
    .B(_02072_));
 sg13g2_xnor2_1 _10585_ (.Y(_03152_),
    .A(net141),
    .B(_03151_));
 sg13g2_nor3_1 _10586_ (.A(_03150_),
    .B(_03123_),
    .C(_03152_),
    .Y(_03153_));
 sg13g2_a21o_1 _10587_ (.A2(_03148_),
    .A1(_03123_),
    .B1(_03153_),
    .X(_03154_));
 sg13g2_a21oi_1 _10588_ (.A1(_02192_),
    .A2(_02000_),
    .Y(_03155_),
    .B1(_01871_));
 sg13g2_nor2_1 _10589_ (.A(_02192_),
    .B(_02000_),
    .Y(_03156_));
 sg13g2_or3_1 _10590_ (.A(net163),
    .B(_03155_),
    .C(_03156_),
    .X(_03157_));
 sg13g2_o21ai_1 _10591_ (.B1(_02837_),
    .Y(_03158_),
    .A1(_02192_),
    .A2(_02026_));
 sg13g2_nand2_1 _10592_ (.Y(_03159_),
    .A(_02192_),
    .B(_02026_));
 sg13g2_nand3_1 _10593_ (.B(_03158_),
    .C(_03159_),
    .A(net163),
    .Y(_03160_));
 sg13g2_nand4_1 _10594_ (.B(_01877_),
    .C(_02379_),
    .A(_02180_),
    .Y(_03161_),
    .D(_02942_));
 sg13g2_nand3b_1 _10595_ (.B(net156),
    .C(_02848_),
    .Y(_03162_),
    .A_N(_02938_));
 sg13g2_nand4_1 _10596_ (.B(_03160_),
    .C(_03161_),
    .A(_03157_),
    .Y(_03163_),
    .D(_03162_));
 sg13g2_nand4_1 _10597_ (.B(_02159_),
    .C(_02196_),
    .A(_01926_),
    .Y(_03164_),
    .D(_03079_));
 sg13g2_o21ai_1 _10598_ (.B1(_03164_),
    .Y(_03165_),
    .A1(_03079_),
    .A2(_03041_));
 sg13g2_nor2b_1 _10599_ (.A(_02969_),
    .B_N(_02831_),
    .Y(_03166_));
 sg13g2_or3_1 _10600_ (.A(net154),
    .B(_02775_),
    .C(_03166_),
    .X(_03167_));
 sg13g2_nor2_1 _10601_ (.A(_02146_),
    .B(_02149_),
    .Y(_03168_));
 sg13g2_nand2_1 _10602_ (.Y(_03169_),
    .A(_02154_),
    .B(_03168_));
 sg13g2_o21ai_1 _10603_ (.B1(_01892_),
    .Y(_03170_),
    .A1(_01879_),
    .A2(_01881_));
 sg13g2_nor2_1 _10604_ (.A(_01881_),
    .B(_02184_),
    .Y(_03171_));
 sg13g2_a21oi_1 _10605_ (.A1(_02190_),
    .A2(_03170_),
    .Y(_03172_),
    .B1(_03171_));
 sg13g2_nand3b_1 _10606_ (.B(_02748_),
    .C(_01831_),
    .Y(_03173_),
    .A_N(_03172_));
 sg13g2_nand2_1 _10607_ (.Y(_03174_),
    .A(_02182_),
    .B(_02748_));
 sg13g2_a21o_1 _10608_ (.A2(_03172_),
    .A1(_02185_),
    .B1(_03174_),
    .X(_03175_));
 sg13g2_nand4_1 _10609_ (.B(_03169_),
    .C(_03173_),
    .A(net151),
    .Y(_03176_),
    .D(_03175_));
 sg13g2_a22oi_1 _10610_ (.Y(_03177_),
    .B1(_03167_),
    .B2(_03176_),
    .A2(_03165_),
    .A1(_03163_));
 sg13g2_buf_2 _10611_ (.A(_03177_),
    .X(_03178_));
 sg13g2_xnor2_1 _10612_ (.Y(_03179_),
    .A(net154),
    .B(net209));
 sg13g2_buf_1 _10613_ (.A(_03179_),
    .X(_03180_));
 sg13g2_nand4_1 _10614_ (.B(_02264_),
    .C(_02502_),
    .A(_02260_),
    .Y(_03181_),
    .D(_02736_));
 sg13g2_nor2_1 _10615_ (.A(net306),
    .B(_02501_),
    .Y(_03182_));
 sg13g2_a21oi_1 _10616_ (.A1(_02263_),
    .A2(_02502_),
    .Y(_03183_),
    .B1(_03182_));
 sg13g2_nand3_1 _10617_ (.B(_03181_),
    .C(_03183_),
    .A(net155),
    .Y(_03184_));
 sg13g2_a22oi_1 _10618_ (.Y(_03185_),
    .B1(net306),
    .B2(_02497_),
    .A2(net309),
    .A1(_02243_));
 sg13g2_o21ai_1 _10619_ (.B1(_03185_),
    .Y(_03186_),
    .A1(_02247_),
    .A2(_02743_));
 sg13g2_nor2_1 _10620_ (.A(net306),
    .B(_02497_),
    .Y(_03187_));
 sg13g2_a21oi_1 _10621_ (.A1(_02244_),
    .A2(_02498_),
    .Y(_03188_),
    .B1(_03187_));
 sg13g2_nand3_1 _10622_ (.B(_03186_),
    .C(_03188_),
    .A(net151),
    .Y(_03189_));
 sg13g2_nand2_1 _10623_ (.Y(_03190_),
    .A(_03184_),
    .B(_03189_));
 sg13g2_nand3_1 _10624_ (.B(_02095_),
    .C(_02979_),
    .A(net163),
    .Y(_03191_));
 sg13g2_nand3_1 _10625_ (.B(_02738_),
    .C(_02805_),
    .A(net160),
    .Y(_03192_));
 sg13g2_a22oi_1 _10626_ (.Y(_03193_),
    .B1(_02778_),
    .B2(_02776_),
    .A2(net270),
    .A1(_02124_));
 sg13g2_nand2_1 _10627_ (.Y(_03194_),
    .A(_03193_),
    .B(_02978_));
 sg13g2_nor2_1 _10628_ (.A(net156),
    .B(_02733_),
    .Y(_03195_));
 sg13g2_a21oi_1 _10629_ (.A1(_02108_),
    .A2(net271),
    .Y(_03196_),
    .B1(_02056_));
 sg13g2_a221oi_1 _10630_ (.B2(_03196_),
    .C1(_02742_),
    .B1(_02766_),
    .A1(_02215_),
    .Y(_03197_),
    .A2(_02216_));
 sg13g2_a221oi_1 _10631_ (.B2(_03195_),
    .C1(_03197_),
    .B1(_03194_),
    .A1(_03191_),
    .Y(_03198_),
    .A2(_03192_));
 sg13g2_buf_1 _10632_ (.A(_03198_),
    .X(_03199_));
 sg13g2_nor3_1 _10633_ (.A(_03180_),
    .B(_03190_),
    .C(_03199_),
    .Y(_03200_));
 sg13g2_nand4_1 _10634_ (.B(_03024_),
    .C(_03178_),
    .A(_03018_),
    .Y(_03201_),
    .D(_03200_));
 sg13g2_or2_1 _10635_ (.X(_03202_),
    .B(_03199_),
    .A(_03190_));
 sg13g2_nand3_1 _10636_ (.B(_02966_),
    .C(_02886_),
    .A(_03013_),
    .Y(_03203_));
 sg13g2_or4_1 _10637_ (.A(_01926_),
    .B(_02876_),
    .C(_03081_),
    .D(_02969_),
    .X(_03204_));
 sg13g2_a22oi_1 _10638_ (.Y(_03205_),
    .B1(_03203_),
    .B2(_03204_),
    .A2(_02850_),
    .A1(_02846_));
 sg13g2_nor4_1 _10639_ (.A(_03180_),
    .B(_03190_),
    .C(_03199_),
    .D(_03205_),
    .Y(_03206_));
 sg13g2_nand2_1 _10640_ (.Y(_03207_),
    .A(net155),
    .B(_02773_));
 sg13g2_nand2_1 _10641_ (.Y(_03208_),
    .A(net151),
    .B(_02162_));
 sg13g2_a22oi_1 _10642_ (.Y(_03209_),
    .B1(_02976_),
    .B2(_02981_),
    .A2(_03208_),
    .A1(_03207_));
 sg13g2_nor4_1 _10643_ (.A(_03180_),
    .B(_03190_),
    .C(_03199_),
    .D(_03209_),
    .Y(_03210_));
 sg13g2_a221oi_1 _10644_ (.B2(_03206_),
    .C1(_03210_),
    .B1(_03178_),
    .A1(_03180_),
    .Y(_03211_),
    .A2(_03202_));
 sg13g2_nand3b_1 _10645_ (.B(_03209_),
    .C(_03180_),
    .Y(_03212_),
    .A_N(_03178_));
 sg13g2_nand3_1 _10646_ (.B(_03209_),
    .C(_03205_),
    .A(_03180_),
    .Y(_03213_));
 sg13g2_a21o_1 _10647_ (.A2(_03024_),
    .A1(_03018_),
    .B1(_03213_),
    .X(_03214_));
 sg13g2_and4_1 _10648_ (.A(_03201_),
    .B(_03211_),
    .C(_03212_),
    .D(_03214_),
    .X(_03215_));
 sg13g2_buf_1 _10649_ (.A(_03215_),
    .X(_03216_));
 sg13g2_buf_8 _10650_ (.A(net150),
    .X(_03217_));
 sg13g2_nor2_1 _10651_ (.A(_02581_),
    .B(_02715_),
    .Y(_03218_));
 sg13g2_xnor2_1 _10652_ (.Y(_03219_),
    .A(net144),
    .B(_03218_));
 sg13g2_nand2_1 _10653_ (.Y(_03220_),
    .A(_02803_),
    .B(_02806_));
 sg13g2_a21o_1 _10654_ (.A2(_03220_),
    .A1(_02747_),
    .B1(_02824_),
    .X(_03221_));
 sg13g2_buf_1 _10655_ (.A(_03221_),
    .X(_03222_));
 sg13g2_a22oi_1 _10656_ (.Y(_03223_),
    .B1(_02841_),
    .B2(_02842_),
    .A2(_02840_),
    .A1(_02835_));
 sg13g2_nor3_1 _10657_ (.A(net154),
    .B(_02144_),
    .C(_02969_),
    .Y(_03224_));
 sg13g2_a22oi_1 _10658_ (.Y(_03225_),
    .B1(_03224_),
    .B2(_02833_),
    .A2(_03223_),
    .A1(_02967_));
 sg13g2_a21o_1 _10659_ (.A2(_02767_),
    .A1(_02750_),
    .B1(_02782_),
    .X(_03226_));
 sg13g2_buf_1 _10660_ (.A(_03226_),
    .X(_03227_));
 sg13g2_and2_1 _10661_ (.A(_02976_),
    .B(_02981_),
    .X(_03228_));
 sg13g2_a221oi_1 _10662_ (.B2(_03227_),
    .C1(_03228_),
    .B1(_03225_),
    .A1(_02973_),
    .Y(_03229_),
    .A2(_02974_));
 sg13g2_buf_1 _10663_ (.A(_03229_),
    .X(_03230_));
 sg13g2_buf_1 _10664_ (.A(net146),
    .X(_03231_));
 sg13g2_nor3_1 _10665_ (.A(_02934_),
    .B(_02944_),
    .C(_02963_),
    .Y(_03232_));
 sg13g2_buf_2 _10666_ (.A(_03232_),
    .X(_03233_));
 sg13g2_buf_8 _10667_ (.A(_03233_),
    .X(_03234_));
 sg13g2_nand2_1 _10668_ (.Y(_03235_),
    .A(_02846_),
    .B(_02850_));
 sg13g2_nand3_1 _10669_ (.B(_02983_),
    .C(_03235_),
    .A(_02972_),
    .Y(_03236_));
 sg13g2_a21oi_1 _10670_ (.A1(net140),
    .A2(net139),
    .Y(_03237_),
    .B1(_03236_));
 sg13g2_nor4_1 _10671_ (.A(_03219_),
    .B(_03222_),
    .C(_03230_),
    .D(_03237_),
    .Y(_03238_));
 sg13g2_xnor2_1 _10672_ (.Y(_03239_),
    .A(_02439_),
    .B(_01837_));
 sg13g2_nand2b_1 _10673_ (.Y(_03240_),
    .B(_03235_),
    .A_N(_03239_));
 sg13g2_nor2_1 _10674_ (.A(net146),
    .B(_03240_),
    .Y(_03241_));
 sg13g2_and4_1 _10675_ (.A(_02844_),
    .B(net146),
    .C(_03233_),
    .D(_03239_),
    .X(_03242_));
 sg13g2_nand3_1 _10676_ (.B(_02850_),
    .C(_03239_),
    .A(_02846_),
    .Y(_03243_));
 sg13g2_mux2_1 _10677_ (.A0(_03239_),
    .A1(_03243_),
    .S(_02844_),
    .X(_03244_));
 sg13g2_o21ai_1 _10678_ (.B1(_03244_),
    .Y(_03245_),
    .A1(_03233_),
    .A2(_03240_));
 sg13g2_nor3_1 _10679_ (.A(_03241_),
    .B(_03242_),
    .C(_03245_),
    .Y(_03246_));
 sg13g2_nor3_1 _10680_ (.A(_03216_),
    .B(_03238_),
    .C(_03246_),
    .Y(_03247_));
 sg13g2_nand2_1 _10681_ (.Y(_03248_),
    .A(_03157_),
    .B(_03160_));
 sg13g2_buf_2 _10682_ (.A(_03248_),
    .X(_03249_));
 sg13g2_nor2_1 _10683_ (.A(net157),
    .B(_02144_),
    .Y(_03250_));
 sg13g2_or2_1 _10684_ (.X(_03251_),
    .B(_03166_),
    .A(_02775_));
 sg13g2_nand3_1 _10685_ (.B(_03173_),
    .C(_03175_),
    .A(_03169_),
    .Y(_03252_));
 sg13g2_and2_1 _10686_ (.A(net156),
    .B(_02162_),
    .X(_03253_));
 sg13g2_o21ai_1 _10687_ (.B1(net161),
    .Y(_03254_),
    .A1(_02733_),
    .A2(_03193_));
 sg13g2_o21ai_1 _10688_ (.B1(net160),
    .Y(_03255_),
    .A1(_02742_),
    .A2(_02766_));
 sg13g2_nand2_1 _10689_ (.Y(_03256_),
    .A(_03254_),
    .B(_03255_));
 sg13g2_a221oi_1 _10690_ (.B2(_03253_),
    .C1(_03256_),
    .B1(_03252_),
    .A1(_03250_),
    .Y(_03257_),
    .A2(_03251_));
 sg13g2_buf_2 _10691_ (.A(_03257_),
    .X(_03258_));
 sg13g2_a21oi_1 _10692_ (.A1(_02239_),
    .A2(_02227_),
    .Y(_03259_),
    .B1(_02237_));
 sg13g2_nor2_1 _10693_ (.A(_02239_),
    .B(_02227_),
    .Y(_03260_));
 sg13g2_nor2_1 _10694_ (.A(_03259_),
    .B(_03260_),
    .Y(_03261_));
 sg13g2_a21oi_1 _10695_ (.A1(_02239_),
    .A2(_02108_),
    .Y(_03262_),
    .B1(_02048_));
 sg13g2_a21oi_1 _10696_ (.A1(_02054_),
    .A2(_02210_),
    .Y(_03263_),
    .B1(_03262_));
 sg13g2_and2_1 _10697_ (.A(net158),
    .B(_03263_),
    .X(_03264_));
 sg13g2_a21oi_2 _10698_ (.B1(_03264_),
    .Y(_03265_),
    .A2(_03261_),
    .A1(net150));
 sg13g2_nor2_1 _10699_ (.A(_03258_),
    .B(_03265_),
    .Y(_03266_));
 sg13g2_nand3_1 _10700_ (.B(_03186_),
    .C(_03188_),
    .A(net209),
    .Y(_03267_));
 sg13g2_nand4_1 _10701_ (.B(_02639_),
    .C(_03186_),
    .A(_02625_),
    .Y(_03268_),
    .D(_03188_));
 sg13g2_nor2_1 _10702_ (.A(net157),
    .B(_02606_),
    .Y(_03269_));
 sg13g2_a221oi_1 _10703_ (.B2(net265),
    .C1(_03269_),
    .B1(_03268_),
    .A1(_02810_),
    .Y(_03270_),
    .A2(_03267_));
 sg13g2_nor2_1 _10704_ (.A(_02503_),
    .B(net307),
    .Y(_03271_));
 sg13g2_nand2_1 _10705_ (.Y(_03272_),
    .A(net265),
    .B(net264));
 sg13g2_nand3_1 _10706_ (.B(_03271_),
    .C(_03272_),
    .A(net161),
    .Y(_03273_));
 sg13g2_nand2_1 _10707_ (.Y(_03274_),
    .A(net265),
    .B(_02564_));
 sg13g2_nand4_1 _10708_ (.B(_02483_),
    .C(net307),
    .A(net157),
    .Y(_03275_),
    .D(_03274_));
 sg13g2_and2_1 _10709_ (.A(_02504_),
    .B(_03272_),
    .X(_03276_));
 sg13g2_nand4_1 _10710_ (.B(_03181_),
    .C(_03183_),
    .A(net161),
    .Y(_03277_),
    .D(_03276_));
 sg13g2_nand4_1 _10711_ (.B(_03273_),
    .C(_03275_),
    .A(_02720_),
    .Y(_03278_),
    .D(_03277_));
 sg13g2_inv_1 _10712_ (.Y(_03279_),
    .A(_02523_));
 sg13g2_nand3_1 _10713_ (.B(_03279_),
    .C(_03218_),
    .A(net158),
    .Y(_03280_));
 sg13g2_or2_1 _10714_ (.X(_03281_),
    .B(_02715_),
    .A(_02581_));
 sg13g2_nand3_1 _10715_ (.B(_02523_),
    .C(_03281_),
    .A(net154),
    .Y(_03282_));
 sg13g2_nand3_1 _10716_ (.B(_03280_),
    .C(_03282_),
    .A(_02720_),
    .Y(_03283_));
 sg13g2_o21ai_1 _10717_ (.B1(_03283_),
    .Y(_03284_),
    .A1(_03270_),
    .A2(_03278_));
 sg13g2_xnor2_1 _10718_ (.Y(_03285_),
    .A(net147),
    .B(_02533_));
 sg13g2_nand2_1 _10719_ (.Y(_03286_),
    .A(_03284_),
    .B(_03285_));
 sg13g2_a21oi_2 _10720_ (.B1(_03078_),
    .Y(_03287_),
    .A2(_02848_),
    .A1(net150));
 sg13g2_a21oi_1 _10721_ (.A1(net146),
    .A2(_03233_),
    .Y(_03288_),
    .B1(_03287_));
 sg13g2_or4_1 _10722_ (.A(_03249_),
    .B(_03266_),
    .C(_03286_),
    .D(_03288_),
    .X(_03289_));
 sg13g2_and4_1 _10723_ (.A(net157),
    .B(_02162_),
    .C(_01923_),
    .D(_02966_),
    .X(_03290_));
 sg13g2_and2_1 _10724_ (.A(_01914_),
    .B(_02978_),
    .X(_03291_));
 sg13g2_a22oi_1 _10725_ (.Y(_03292_),
    .B1(_03291_),
    .B2(_02970_),
    .A2(_03290_),
    .A1(_03196_));
 sg13g2_buf_1 _10726_ (.A(_03292_),
    .X(_03293_));
 sg13g2_xnor2_1 _10727_ (.Y(_03294_),
    .A(net155),
    .B(_02533_));
 sg13g2_or4_1 _10728_ (.A(net160),
    .B(_02523_),
    .C(_02574_),
    .D(net209),
    .X(_03295_));
 sg13g2_nand2_1 _10729_ (.Y(_03296_),
    .A(_02523_),
    .B(net209));
 sg13g2_or3_1 _10730_ (.A(net163),
    .B(_02585_),
    .C(_03296_),
    .X(_03297_));
 sg13g2_a22oi_1 _10731_ (.Y(_03298_),
    .B1(_03295_),
    .B2(_03297_),
    .A2(_03192_),
    .A1(_03191_));
 sg13g2_buf_1 _10732_ (.A(_03298_),
    .X(_03299_));
 sg13g2_nand2_1 _10733_ (.Y(_03300_),
    .A(_03294_),
    .B(_03299_));
 sg13g2_nor2_1 _10734_ (.A(_03293_),
    .B(_03300_),
    .Y(_03301_));
 sg13g2_o21ai_1 _10735_ (.B1(_03301_),
    .Y(_03302_),
    .A1(_03249_),
    .A2(_03288_));
 sg13g2_nor2_1 _10736_ (.A(_03270_),
    .B(_03278_),
    .Y(_03303_));
 sg13g2_nor2b_1 _10737_ (.A(_03303_),
    .B_N(_03283_),
    .Y(_03304_));
 sg13g2_inv_1 _10738_ (.Y(_03305_),
    .A(_03300_));
 sg13g2_a22oi_1 _10739_ (.Y(_03306_),
    .B1(_03305_),
    .B2(_03266_),
    .A2(_03294_),
    .A1(_03304_));
 sg13g2_and2_1 _10740_ (.A(_03285_),
    .B(_03293_),
    .X(_03307_));
 sg13g2_o21ai_1 _10741_ (.B1(_03307_),
    .Y(_03308_),
    .A1(_03258_),
    .A2(_03265_));
 sg13g2_inv_1 _10742_ (.Y(_03309_),
    .A(_03299_));
 sg13g2_nand2_1 _10743_ (.Y(_03310_),
    .A(_03285_),
    .B(_03309_));
 sg13g2_a21o_1 _10744_ (.A2(_03310_),
    .A1(_03308_),
    .B1(_03304_),
    .X(_03311_));
 sg13g2_and4_1 _10745_ (.A(_03289_),
    .B(_03302_),
    .C(_03306_),
    .D(_03311_),
    .X(_03312_));
 sg13g2_and2_1 _10746_ (.A(_03163_),
    .B(_03165_),
    .X(_03313_));
 sg13g2_a21o_1 _10747_ (.A2(_03176_),
    .A1(_03167_),
    .B1(_03313_),
    .X(_03314_));
 sg13g2_a21o_1 _10748_ (.A2(_03204_),
    .A1(_03203_),
    .B1(_02852_),
    .X(_03315_));
 sg13g2_a21oi_1 _10749_ (.A1(_03018_),
    .A2(_03024_),
    .Y(_03316_),
    .B1(_03315_));
 sg13g2_xnor2_1 _10750_ (.Y(_03317_),
    .A(net145),
    .B(_03039_));
 sg13g2_nor3_1 _10751_ (.A(_03314_),
    .B(_03316_),
    .C(_03317_),
    .Y(_03318_));
 sg13g2_a21o_1 _10752_ (.A2(_03024_),
    .A1(_03018_),
    .B1(_03315_),
    .X(_03319_));
 sg13g2_xnor2_1 _10753_ (.Y(_03320_),
    .A(net142),
    .B(_03039_));
 sg13g2_a21oi_1 _10754_ (.A1(_03178_),
    .A2(_03319_),
    .Y(_03321_),
    .B1(_03320_));
 sg13g2_or3_1 _10755_ (.A(net150),
    .B(_02093_),
    .C(_02833_),
    .X(_03322_));
 sg13g2_nand2_1 _10756_ (.Y(_03323_),
    .A(net154),
    .B(_02093_));
 sg13g2_or2_1 _10757_ (.X(_03324_),
    .B(_03223_),
    .A(_03323_));
 sg13g2_a21o_1 _10758_ (.A2(_03324_),
    .A1(_03322_),
    .B1(_02747_),
    .X(_03325_));
 sg13g2_buf_1 _10759_ (.A(_03325_),
    .X(_03326_));
 sg13g2_xnor2_1 _10760_ (.Y(_03327_),
    .A(net153),
    .B(_02201_));
 sg13g2_buf_2 _10761_ (.A(_03327_),
    .X(_03328_));
 sg13g2_nand3_1 _10762_ (.B(_03225_),
    .C(_03328_),
    .A(_03227_),
    .Y(_03329_));
 sg13g2_a21oi_1 _10763_ (.A1(_03326_),
    .A2(_03329_),
    .Y(_03330_),
    .B1(_02784_));
 sg13g2_nand2_1 _10764_ (.Y(_03331_),
    .A(_02983_),
    .B(_03218_));
 sg13g2_and4_1 _10765_ (.A(_02091_),
    .B(_02162_),
    .C(_02771_),
    .D(_02966_),
    .X(_03332_));
 sg13g2_nor2_1 _10766_ (.A(net158),
    .B(_02093_),
    .Y(_03333_));
 sg13g2_nand4_1 _10767_ (.B(_02056_),
    .C(_02108_),
    .A(net272),
    .Y(_03334_),
    .D(net271));
 sg13g2_nor4_1 _10768_ (.A(_02091_),
    .B(_02144_),
    .C(_03334_),
    .D(_02969_),
    .Y(_03335_));
 sg13g2_nor2_1 _10769_ (.A(net151),
    .B(_02087_),
    .Y(_03336_));
 sg13g2_a22oi_1 _10770_ (.Y(_03337_),
    .B1(_03335_),
    .B2(_03336_),
    .A2(_03333_),
    .A1(_03332_));
 sg13g2_buf_1 _10771_ (.A(_03337_),
    .X(_03338_));
 sg13g2_and3_1 _10772_ (.X(_03339_),
    .A(net142),
    .B(_02111_),
    .C(_03338_));
 sg13g2_and3_1 _10773_ (.X(_03340_),
    .A(net145),
    .B(_02201_),
    .C(_03338_));
 sg13g2_nand2_1 _10774_ (.Y(_03341_),
    .A(_02983_),
    .B(_03281_));
 sg13g2_inv_1 _10775_ (.Y(_03342_),
    .A(_02972_));
 sg13g2_a221oi_1 _10776_ (.B2(_03341_),
    .C1(_03342_),
    .B1(_03340_),
    .A1(_03331_),
    .Y(_03343_),
    .A2(_03339_));
 sg13g2_a21oi_1 _10777_ (.A1(net140),
    .A2(net139),
    .Y(_03344_),
    .B1(_02852_));
 sg13g2_mux2_1 _10778_ (.A0(_03330_),
    .A1(_03343_),
    .S(_03344_),
    .X(_03345_));
 sg13g2_nor3_1 _10779_ (.A(_03318_),
    .B(_03321_),
    .C(_03345_),
    .Y(_03346_));
 sg13g2_and4_1 _10780_ (.A(_03154_),
    .B(_03247_),
    .C(_03312_),
    .D(_03346_),
    .X(_03347_));
 sg13g2_a21oi_1 _10781_ (.A1(_02209_),
    .A2(_02212_),
    .Y(_03348_),
    .B1(_02230_));
 sg13g2_a21oi_1 _10782_ (.A1(_03052_),
    .A2(_03053_),
    .Y(_03349_),
    .B1(net144));
 sg13g2_a221oi_1 _10783_ (.B2(_01924_),
    .C1(_03349_),
    .B1(_01915_),
    .A1(net144),
    .Y(_03350_),
    .A2(_02001_));
 sg13g2_nand2_1 _10784_ (.Y(_03351_),
    .A(_02160_),
    .B(_02163_));
 sg13g2_o21ai_1 _10785_ (.B1(_03351_),
    .Y(_03352_),
    .A1(_02199_),
    .A2(_03350_));
 sg13g2_nand2b_1 _10786_ (.Y(_03353_),
    .B(_03352_),
    .A_N(_03348_));
 sg13g2_inv_1 _10787_ (.Y(_03354_),
    .A(_03097_));
 sg13g2_and2_1 _10788_ (.A(net158),
    .B(_02303_),
    .X(_03355_));
 sg13g2_a21oi_1 _10789_ (.A1(_02700_),
    .A2(_02297_),
    .Y(_03356_),
    .B1(_03355_));
 sg13g2_o21ai_1 _10790_ (.B1(_03137_),
    .Y(_03357_),
    .A1(_03356_),
    .A2(_02912_));
 sg13g2_nand2_1 _10791_ (.Y(_03358_),
    .A(_03351_),
    .B(_01925_));
 sg13g2_a221oi_1 _10792_ (.B2(_03140_),
    .C1(_03358_),
    .B1(_03139_),
    .A1(_03354_),
    .Y(_03359_),
    .A2(_03357_));
 sg13g2_buf_1 _10793_ (.A(_03359_),
    .X(_03360_));
 sg13g2_nor2_1 _10794_ (.A(_03353_),
    .B(_03360_),
    .Y(_03361_));
 sg13g2_xnor2_1 _10795_ (.Y(_03362_),
    .A(net145),
    .B(_02056_));
 sg13g2_xor2_1 _10796_ (.B(_03362_),
    .A(_03361_),
    .X(_03363_));
 sg13g2_xnor2_1 _10797_ (.Y(_03364_),
    .A(net151),
    .B(_03050_));
 sg13g2_xnor2_1 _10798_ (.Y(_03365_),
    .A(net152),
    .B(net272));
 sg13g2_nor2_1 _10799_ (.A(_03293_),
    .B(_03365_),
    .Y(_03366_));
 sg13g2_nor2_1 _10800_ (.A(_03364_),
    .B(_03366_),
    .Y(_03367_));
 sg13g2_o21ai_1 _10801_ (.B1(_03365_),
    .Y(_03368_),
    .A1(_03258_),
    .A2(_03265_));
 sg13g2_and2_1 _10802_ (.A(_03364_),
    .B(_03368_),
    .X(_03369_));
 sg13g2_nor2_1 _10803_ (.A(_03249_),
    .B(_03288_),
    .Y(_03370_));
 sg13g2_mux2_1 _10804_ (.A0(_03367_),
    .A1(_03369_),
    .S(_03370_),
    .X(_03371_));
 sg13g2_nor3_1 _10805_ (.A(_03062_),
    .B(_03088_),
    .C(_03098_),
    .Y(_03372_));
 sg13g2_xnor2_1 _10806_ (.Y(_03373_),
    .A(net145),
    .B(_02203_));
 sg13g2_xnor2_1 _10807_ (.Y(_03374_),
    .A(_03372_),
    .B(_03373_));
 sg13g2_nor2_1 _10808_ (.A(net153),
    .B(_01877_),
    .Y(_03375_));
 sg13g2_and4_1 _10809_ (.A(net155),
    .B(_01877_),
    .C(_02024_),
    .D(_02026_),
    .X(_03376_));
 sg13g2_a21oi_1 _10810_ (.A1(_02002_),
    .A2(_03375_),
    .Y(_03377_),
    .B1(_03376_));
 sg13g2_nor2_1 _10811_ (.A(_02476_),
    .B(_03377_),
    .Y(_03378_));
 sg13g2_nand2b_1 _10812_ (.Y(_03379_),
    .B(_03008_),
    .A_N(_02029_));
 sg13g2_xnor2_1 _10813_ (.Y(_03380_),
    .A(net151),
    .B(_01877_));
 sg13g2_a21oi_1 _10814_ (.A1(net155),
    .A2(_02889_),
    .Y(_03381_),
    .B1(_02893_));
 sg13g2_nand2_1 _10815_ (.Y(_03382_),
    .A(_02899_),
    .B(_02905_));
 sg13g2_a22oi_1 _10816_ (.Y(_03383_),
    .B1(_02912_),
    .B2(_03382_),
    .A2(_03381_),
    .A1(_02861_));
 sg13g2_buf_2 _10817_ (.A(_03383_),
    .X(_03384_));
 sg13g2_xnor2_1 _10818_ (.Y(_03385_),
    .A(net148),
    .B(_02437_));
 sg13g2_xnor2_1 _10819_ (.Y(_03386_),
    .A(_03384_),
    .B(_03385_));
 sg13g2_a21o_1 _10820_ (.A2(_03380_),
    .A1(_03379_),
    .B1(_03386_),
    .X(_03387_));
 sg13g2_xnor2_1 _10821_ (.Y(_03388_),
    .A(net155),
    .B(_02379_));
 sg13g2_buf_2 _10822_ (.A(_03388_),
    .X(_03389_));
 sg13g2_nand3_1 _10823_ (.B(net139),
    .C(_03389_),
    .A(net140),
    .Y(_03390_));
 sg13g2_o21ai_1 _10824_ (.B1(_03390_),
    .Y(_03391_),
    .A1(net139),
    .A2(_03389_));
 sg13g2_nor4_1 _10825_ (.A(_03374_),
    .B(_03378_),
    .C(_03387_),
    .D(_03391_),
    .Y(_03392_));
 sg13g2_nand3_1 _10826_ (.B(_02044_),
    .C(_03261_),
    .A(net142),
    .Y(_03393_));
 sg13g2_nand3b_1 _10827_ (.B(_03263_),
    .C(net148),
    .Y(_03394_),
    .A_N(_02044_));
 sg13g2_a21o_1 _10828_ (.A2(_03394_),
    .A1(_03393_),
    .B1(_03258_),
    .X(_03395_));
 sg13g2_buf_1 _10829_ (.A(_03395_),
    .X(_03396_));
 sg13g2_and2_1 _10830_ (.A(_03293_),
    .B(_03365_),
    .X(_03397_));
 sg13g2_o21ai_1 _10831_ (.B1(_03397_),
    .Y(_03398_),
    .A1(_03258_),
    .A2(_03265_));
 sg13g2_nand2_1 _10832_ (.Y(_03399_),
    .A(_03396_),
    .B(_03398_));
 sg13g2_or2_1 _10833_ (.X(_03400_),
    .B(_03336_),
    .A(_03333_));
 sg13g2_nand3b_1 _10834_ (.B(_02087_),
    .C(net152),
    .Y(_03401_),
    .A_N(_03335_));
 sg13g2_o21ai_1 _10835_ (.B1(_03401_),
    .Y(_03402_),
    .A1(_03323_),
    .A2(_03332_));
 sg13g2_nor2_1 _10836_ (.A(_02747_),
    .B(_02784_),
    .Y(_03403_));
 sg13g2_mux2_1 _10837_ (.A0(_03400_),
    .A1(_03402_),
    .S(_03403_),
    .X(_03404_));
 sg13g2_nand2_1 _10838_ (.Y(_03405_),
    .A(_03227_),
    .B(_03225_));
 sg13g2_a21oi_1 _10839_ (.A1(_02750_),
    .A2(_02767_),
    .Y(_03406_),
    .B1(_02782_));
 sg13g2_nor2_1 _10840_ (.A(_03406_),
    .B(_02972_),
    .Y(_03407_));
 sg13g2_mux2_1 _10841_ (.A0(_03405_),
    .A1(_03407_),
    .S(_03328_),
    .X(_03408_));
 sg13g2_nand2_2 _10842_ (.Y(_03409_),
    .A(_02869_),
    .B(_02470_));
 sg13g2_nor3_1 _10843_ (.A(net155),
    .B(_02468_),
    .C(_03409_),
    .Y(_03410_));
 sg13g2_nor3_1 _10844_ (.A(_02700_),
    .B(_02455_),
    .C(_03093_),
    .Y(_03411_));
 sg13g2_or2_1 _10845_ (.X(_03412_),
    .B(_03411_),
    .A(_03410_));
 sg13g2_nand2_1 _10846_ (.Y(_03413_),
    .A(net148),
    .B(_02901_));
 sg13g2_nand3b_1 _10847_ (.B(_03413_),
    .C(_03065_),
    .Y(_03414_),
    .A_N(_03412_));
 sg13g2_nand2_1 _10848_ (.Y(_03415_),
    .A(_02417_),
    .B(_02437_));
 sg13g2_nand2_1 _10849_ (.Y(_03416_),
    .A(_02684_),
    .B(_03093_));
 sg13g2_nand3_1 _10850_ (.B(_02451_),
    .C(_03409_),
    .A(net150),
    .Y(_03417_));
 sg13g2_o21ai_1 _10851_ (.B1(_03417_),
    .Y(_03418_),
    .A1(_03415_),
    .A2(_03416_));
 sg13g2_xnor2_1 _10852_ (.Y(_03419_),
    .A(_02684_),
    .B(_02895_));
 sg13g2_nand2b_1 _10853_ (.Y(_03420_),
    .B(_02296_),
    .A_N(_02286_));
 sg13g2_nand2b_1 _10854_ (.Y(_03421_),
    .B(_02891_),
    .A_N(_02286_));
 sg13g2_mux2_1 _10855_ (.A0(_03420_),
    .A1(_03421_),
    .S(_03013_),
    .X(_03422_));
 sg13g2_buf_1 _10856_ (.A(_03422_),
    .X(_03423_));
 sg13g2_xor2_1 _10857_ (.B(_03423_),
    .A(_03419_),
    .X(_03424_));
 sg13g2_nand2b_1 _10858_ (.Y(_03425_),
    .B(_03424_),
    .A_N(_03418_));
 sg13g2_mux2_1 _10859_ (.A0(_03414_),
    .A1(_03425_),
    .S(_02321_),
    .X(_03426_));
 sg13g2_nor2_1 _10860_ (.A(_01711_),
    .B(_01715_),
    .Y(_03427_));
 sg13g2_a21oi_1 _10861_ (.A1(net152),
    .A2(_01717_),
    .Y(_03428_),
    .B1(_03427_));
 sg13g2_nor2b_1 _10862_ (.A(_02307_),
    .B_N(_02308_),
    .Y(_03429_));
 sg13g2_and2_1 _10863_ (.A(_03428_),
    .B(_03429_),
    .X(_03430_));
 sg13g2_a21oi_1 _10864_ (.A1(net144),
    .A2(_01717_),
    .Y(_03431_),
    .B1(_03429_));
 sg13g2_nor2_1 _10865_ (.A(_02844_),
    .B(_03338_),
    .Y(_03432_));
 sg13g2_nor3_1 _10866_ (.A(_02468_),
    .B(_02451_),
    .C(_03409_),
    .Y(_03433_));
 sg13g2_a221oi_1 _10867_ (.B2(_03409_),
    .C1(_03433_),
    .B1(_02468_),
    .A1(_02215_),
    .Y(_03434_),
    .A2(_02216_));
 sg13g2_a221oi_1 _10868_ (.B2(_02437_),
    .C1(_02455_),
    .B1(_02417_),
    .A1(_02869_),
    .Y(_03435_),
    .A2(_02470_));
 sg13g2_and2_1 _10869_ (.A(_02455_),
    .B(_03093_),
    .X(_03436_));
 sg13g2_nor3_1 _10870_ (.A(net147),
    .B(_03435_),
    .C(_03436_),
    .Y(_03437_));
 sg13g2_nor2_1 _10871_ (.A(_03434_),
    .B(_03437_),
    .Y(_03438_));
 sg13g2_or4_1 _10872_ (.A(_03430_),
    .B(_03431_),
    .C(_03432_),
    .D(_03438_),
    .X(_03439_));
 sg13g2_or4_1 _10873_ (.A(_03404_),
    .B(_03408_),
    .C(_03426_),
    .D(_03439_),
    .X(_03440_));
 sg13g2_or2_1 _10874_ (.X(_03441_),
    .B(_02458_),
    .A(_02455_));
 sg13g2_nor2_1 _10875_ (.A(_02884_),
    .B(_03441_),
    .Y(_03442_));
 sg13g2_nor3_1 _10876_ (.A(_02873_),
    .B(_02468_),
    .C(_02472_),
    .Y(_03443_));
 sg13g2_and2_1 _10877_ (.A(_02884_),
    .B(_02392_),
    .X(_03444_));
 sg13g2_nor2b_1 _10878_ (.A(_03415_),
    .B_N(_03444_),
    .Y(_03445_));
 sg13g2_and2_1 _10879_ (.A(_02352_),
    .B(_02873_),
    .X(_03446_));
 sg13g2_and2_1 _10880_ (.A(_02451_),
    .B(_03446_),
    .X(_03447_));
 sg13g2_mux4_1 _10881_ (.S0(net144),
    .A0(_03442_),
    .A1(_03443_),
    .A2(_03445_),
    .A3(_03447_),
    .S1(_02321_),
    .X(_03448_));
 sg13g2_or2_1 _10882_ (.X(_03449_),
    .B(_02472_),
    .A(_02468_));
 sg13g2_nand3_1 _10883_ (.B(_03066_),
    .C(_03421_),
    .A(_02895_),
    .Y(_03450_));
 sg13g2_o21ai_1 _10884_ (.B1(net147),
    .Y(_03451_),
    .A1(_02352_),
    .A2(_02873_));
 sg13g2_a221oi_1 _10885_ (.B2(_03450_),
    .C1(_03451_),
    .B1(_03443_),
    .A1(_03449_),
    .Y(_03452_),
    .A2(_03446_));
 sg13g2_nand2_1 _10886_ (.Y(_03453_),
    .A(_02391_),
    .B(_02457_));
 sg13g2_a221oi_1 _10887_ (.B2(_02437_),
    .C1(_02455_),
    .B1(_02417_),
    .A1(_03067_),
    .Y(_03454_),
    .A2(_03453_));
 sg13g2_o21ai_1 _10888_ (.B1(net153),
    .Y(_03455_),
    .A1(_02884_),
    .A2(_02392_));
 sg13g2_a221oi_1 _10889_ (.B2(_02873_),
    .C1(_03455_),
    .B1(_03454_),
    .A1(_03441_),
    .Y(_03456_),
    .A2(_03444_));
 sg13g2_nor2_1 _10890_ (.A(_03452_),
    .B(_03456_),
    .Y(_03457_));
 sg13g2_nor2_1 _10891_ (.A(_03448_),
    .B(_03457_),
    .Y(_03458_));
 sg13g2_xnor2_1 _10892_ (.Y(_03459_),
    .A(net158),
    .B(_02682_));
 sg13g2_a21oi_1 _10893_ (.A1(_02587_),
    .A2(_03104_),
    .Y(_03460_),
    .B1(_02616_));
 sg13g2_buf_2 _10894_ (.A(_03460_),
    .X(_03461_));
 sg13g2_or2_1 _10895_ (.X(_03462_),
    .B(_03461_),
    .A(_03459_));
 sg13g2_nor3_1 _10896_ (.A(_03007_),
    .B(_02900_),
    .C(net183),
    .Y(_03463_));
 sg13g2_nor3_1 _10897_ (.A(net145),
    .B(_02311_),
    .C(net183),
    .Y(_03464_));
 sg13g2_o21ai_1 _10898_ (.B1(_03064_),
    .Y(_03465_),
    .A1(_03463_),
    .A2(_03464_));
 sg13g2_nor3_1 _10899_ (.A(net148),
    .B(_02313_),
    .C(_02897_),
    .Y(_03466_));
 sg13g2_nor3_1 _10900_ (.A(net144),
    .B(_02301_),
    .C(_02897_),
    .Y(_03467_));
 sg13g2_o21ai_1 _10901_ (.B1(_03064_),
    .Y(_03468_),
    .A1(_03466_),
    .A2(_03467_));
 sg13g2_nor3_1 _10902_ (.A(net148),
    .B(_02900_),
    .C(net183),
    .Y(_03469_));
 sg13g2_nor3_1 _10903_ (.A(net148),
    .B(_02301_),
    .C(net183),
    .Y(_03470_));
 sg13g2_o21ai_1 _10904_ (.B1(_02912_),
    .Y(_03471_),
    .A1(_03469_),
    .A2(_03470_));
 sg13g2_nor3_1 _10905_ (.A(net144),
    .B(_02311_),
    .C(_02897_),
    .Y(_03472_));
 sg13g2_nor3_1 _10906_ (.A(net144),
    .B(_02313_),
    .C(_02897_),
    .Y(_03473_));
 sg13g2_o21ai_1 _10907_ (.B1(_02912_),
    .Y(_03474_),
    .A1(_03472_),
    .A2(_03473_));
 sg13g2_nand4_1 _10908_ (.B(_03468_),
    .C(_03471_),
    .A(_03465_),
    .Y(_03475_),
    .D(_03474_));
 sg13g2_nand3b_1 _10909_ (.B(_03462_),
    .C(_03475_),
    .Y(_03476_),
    .A_N(_03458_));
 sg13g2_inv_1 _10910_ (.Y(_03477_),
    .A(_02931_));
 sg13g2_nand2_2 _10911_ (.Y(_03478_),
    .A(_02386_),
    .B(_02388_));
 sg13g2_a21o_1 _10912_ (.A2(_02464_),
    .A1(_03478_),
    .B1(_02343_),
    .X(_03479_));
 sg13g2_o21ai_1 _10913_ (.B1(_03479_),
    .Y(_03480_),
    .A1(_03478_),
    .A2(_02464_));
 sg13g2_o21ai_1 _10914_ (.B1(_02867_),
    .Y(_03481_),
    .A1(_03478_),
    .A2(_02435_));
 sg13g2_o21ai_1 _10915_ (.B1(_03481_),
    .Y(_03482_),
    .A1(_02916_),
    .A2(_02443_));
 sg13g2_nand2_1 _10916_ (.Y(_03483_),
    .A(_02351_),
    .B(_02865_));
 sg13g2_mux4_1 _10917_ (.S0(_03014_),
    .A0(_03477_),
    .A1(_03480_),
    .A2(_03482_),
    .A3(_02958_),
    .S1(_03483_),
    .X(_03484_));
 sg13g2_nand3_1 _10918_ (.B(_03483_),
    .C(_02881_),
    .A(net147),
    .Y(_03485_));
 sg13g2_nand4_1 _10919_ (.B(_02437_),
    .C(_03092_),
    .A(net153),
    .Y(_03486_),
    .D(_03409_));
 sg13g2_and2_1 _10920_ (.A(_03485_),
    .B(_03486_),
    .X(_03487_));
 sg13g2_nor2b_1 _10921_ (.A(_03484_),
    .B_N(_03487_),
    .Y(_03488_));
 sg13g2_nor2_1 _10922_ (.A(_02701_),
    .B(_03092_),
    .Y(_03489_));
 sg13g2_nor2_1 _10923_ (.A(net153),
    .B(_02958_),
    .Y(_03490_));
 sg13g2_a22oi_1 _10924_ (.Y(_03491_),
    .B1(_03490_),
    .B2(_03092_),
    .A2(_03489_),
    .A1(_02931_));
 sg13g2_nor2b_1 _10925_ (.A(_03484_),
    .B_N(_03491_),
    .Y(_03492_));
 sg13g2_mux2_1 _10926_ (.A0(_03488_),
    .A1(_03492_),
    .S(_03384_),
    .X(_03493_));
 sg13g2_o21ai_1 _10927_ (.B1(_03219_),
    .Y(_03494_),
    .A1(_03222_),
    .A2(_03230_));
 sg13g2_or2_1 _10928_ (.X(_03495_),
    .B(_03389_),
    .A(net140));
 sg13g2_xnor2_1 _10929_ (.Y(_03496_),
    .A(net153),
    .B(_03081_));
 sg13g2_nor2_1 _10930_ (.A(_03097_),
    .B(_03496_),
    .Y(_03497_));
 sg13g2_and2_1 _10931_ (.A(_03137_),
    .B(_03496_),
    .X(_03498_));
 sg13g2_and2_1 _10932_ (.A(_03097_),
    .B(_03496_),
    .X(_03499_));
 sg13g2_a221oi_1 _10933_ (.B2(_03132_),
    .C1(_03499_),
    .B1(_03498_),
    .A1(_03357_),
    .Y(_03500_),
    .A2(_03497_));
 sg13g2_nand4_1 _10934_ (.B(_03494_),
    .C(_03495_),
    .A(_03493_),
    .Y(_03501_),
    .D(_03500_));
 sg13g2_nor4_1 _10935_ (.A(_03399_),
    .B(_03440_),
    .C(_03476_),
    .D(_03501_),
    .Y(_03502_));
 sg13g2_and4_1 _10936_ (.A(_03363_),
    .B(_03371_),
    .C(_03392_),
    .D(_03502_),
    .X(_03503_));
 sg13g2_nand2_1 _10937_ (.Y(_03504_),
    .A(net157),
    .B(_02088_));
 sg13g2_nand3_1 _10938_ (.B(_02095_),
    .C(_02608_),
    .A(net161),
    .Y(_03505_));
 sg13g2_o21ai_1 _10939_ (.B1(_03505_),
    .Y(_03506_),
    .A1(_03504_),
    .A2(_02576_));
 sg13g2_nand2_1 _10940_ (.Y(_03507_),
    .A(_02648_),
    .B(_03506_));
 sg13g2_inv_1 _10941_ (.Y(_03508_),
    .A(_03507_));
 sg13g2_o21ai_1 _10942_ (.B1(net141),
    .Y(_03509_),
    .A1(_03147_),
    .A2(_03128_));
 sg13g2_nand2_1 _10943_ (.Y(_03510_),
    .A(_03459_),
    .B(_03461_));
 sg13g2_a21oi_1 _10944_ (.A1(_03508_),
    .A2(_03509_),
    .Y(_03511_),
    .B1(_03510_));
 sg13g2_xnor2_1 _10945_ (.Y(_03512_),
    .A(net154),
    .B(_02682_));
 sg13g2_and3_1 _10946_ (.X(_03513_),
    .A(_03508_),
    .B(_03509_),
    .C(_03512_));
 sg13g2_a21oi_1 _10947_ (.A1(_02478_),
    .A2(_02476_),
    .Y(_03514_),
    .B1(_03028_));
 sg13g2_o21ai_1 _10948_ (.B1(_02648_),
    .Y(_03515_),
    .A1(_02231_),
    .A2(_03028_));
 sg13g2_xnor2_1 _10949_ (.Y(_03516_),
    .A(net147),
    .B(_03279_));
 sg13g2_nand3b_1 _10950_ (.B(_03515_),
    .C(_03516_),
    .Y(_03517_),
    .A_N(_02637_));
 sg13g2_inv_1 _10951_ (.Y(_03518_),
    .A(_03516_));
 sg13g2_nand2_1 _10952_ (.Y(_03519_),
    .A(_02637_),
    .B(_03518_));
 sg13g2_nand4_1 _10953_ (.B(_03514_),
    .C(_03517_),
    .A(_02234_),
    .Y(_03520_),
    .D(_03519_));
 sg13g2_buf_1 _10954_ (.A(_03520_),
    .X(_03521_));
 sg13g2_and3_1 _10955_ (.X(_03522_),
    .A(_02165_),
    .B(_02648_),
    .C(_03516_));
 sg13g2_o21ai_1 _10956_ (.B1(_03518_),
    .Y(_03523_),
    .A1(_02637_),
    .A2(_02648_));
 sg13g2_a22oi_1 _10957_ (.Y(_03524_),
    .B1(_03523_),
    .B2(_03517_),
    .A2(_03522_),
    .A1(_03011_));
 sg13g2_nand2_1 _10958_ (.Y(_03525_),
    .A(_03521_),
    .B(_03524_));
 sg13g2_nor4_1 _10959_ (.A(_02989_),
    .B(_03511_),
    .C(_03513_),
    .D(_03525_),
    .Y(_03526_));
 sg13g2_nand4_1 _10960_ (.B(_03347_),
    .C(_03503_),
    .A(_03122_),
    .Y(_03527_),
    .D(_03526_));
 sg13g2_a22oi_1 _10961_ (.Y(_03528_),
    .B1(_03006_),
    .B2(_03527_),
    .A2(_03004_),
    .A1(_02992_));
 sg13g2_buf_1 _10962_ (.A(_03528_),
    .X(_03529_));
 sg13g2_nand2_1 _10963_ (.Y(_03530_),
    .A(net325),
    .B(_02713_));
 sg13g2_inv_1 _10964_ (.Y(_03531_),
    .A(_03530_));
 sg13g2_nor3_1 _10965_ (.A(_03511_),
    .B(_03513_),
    .C(_03525_),
    .Y(_03532_));
 sg13g2_nand4_1 _10966_ (.B(_03347_),
    .C(_03503_),
    .A(_03122_),
    .Y(_03533_),
    .D(_03532_));
 sg13g2_nor2_1 _10967_ (.A(net527),
    .B(_01558_),
    .Y(_03534_));
 sg13g2_buf_1 _10968_ (.A(net186),
    .X(_03535_));
 sg13g2_buf_2 _10969_ (.A(net176),
    .X(_03536_));
 sg13g2_buf_1 _10970_ (.A(net452),
    .X(_03537_));
 sg13g2_buf_1 _10971_ (.A(net415),
    .X(_03538_));
 sg13g2_nor2_1 _10972_ (.A(_01628_),
    .B(net315),
    .Y(_03539_));
 sg13g2_buf_1 _10973_ (.A(_03539_),
    .X(_03540_));
 sg13g2_buf_1 _10974_ (.A(net262),
    .X(_03541_));
 sg13g2_nand3_1 _10975_ (.B(_03541_),
    .C(_01715_),
    .A(net167),
    .Y(_03542_));
 sg13g2_nand2_1 _10976_ (.Y(_03543_),
    .A(net362),
    .B(_03542_));
 sg13g2_buf_1 _10977_ (.A(net187),
    .X(_03544_));
 sg13g2_buf_1 _10978_ (.A(net175),
    .X(_03545_));
 sg13g2_buf_1 _10979_ (.A(net165),
    .X(_03546_));
 sg13g2_nand2b_1 _10980_ (.Y(_03547_),
    .B(net159),
    .A_N(_01717_));
 sg13g2_buf_1 _10981_ (.A(net212),
    .X(_03548_));
 sg13g2_buf_1 _10982_ (.A(net182),
    .X(_03549_));
 sg13g2_a221oi_1 _10983_ (.B2(net174),
    .C1(_03427_),
    .B1(_03547_),
    .A1(net167),
    .Y(_03550_),
    .A2(_01717_));
 sg13g2_a221oi_1 _10984_ (.B2(_03543_),
    .C1(_03550_),
    .B1(_01711_),
    .A1(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[0] ),
    .Y(_03551_),
    .A2(net166));
 sg13g2_nand2b_1 _10985_ (.Y(_03552_),
    .B(net315),
    .A_N(_02705_));
 sg13g2_o21ai_1 _10986_ (.B1(net263),
    .Y(_03553_),
    .A1(_02997_),
    .A2(_03552_));
 sg13g2_nand2_1 _10987_ (.Y(_03554_),
    .A(_02712_),
    .B(net315));
 sg13g2_nand4_1 _10988_ (.B(net305),
    .C(_02679_),
    .A(_03000_),
    .Y(_03555_),
    .D(_02696_));
 sg13g2_nor2b_1 _10989_ (.A(_02998_),
    .B_N(_03555_),
    .Y(_03556_));
 sg13g2_inv_1 _10990_ (.Y(_03557_),
    .A(net305));
 sg13g2_a21oi_1 _10991_ (.A1(_03557_),
    .A2(_02696_),
    .Y(_03558_),
    .B1(net263));
 sg13g2_o21ai_1 _10992_ (.B1(_03558_),
    .Y(_03559_),
    .A1(_02997_),
    .A2(_03556_));
 sg13g2_nand4_1 _10993_ (.B(_03553_),
    .C(_03554_),
    .A(_01738_),
    .Y(_03560_),
    .D(_03559_));
 sg13g2_nand3_1 _10994_ (.B(_03551_),
    .C(_03560_),
    .A(_03534_),
    .Y(_03561_));
 sg13g2_a21o_1 _10995_ (.A2(_03533_),
    .A1(_03531_),
    .B1(_03561_),
    .X(_03562_));
 sg13g2_buf_1 _10996_ (.A(net624),
    .X(_03563_));
 sg13g2_buf_1 _10997_ (.A(net597),
    .X(_03564_));
 sg13g2_buf_1 _10998_ (.A(net525),
    .X(_03565_));
 sg13g2_buf_1 _10999_ (.A(net599),
    .X(_03566_));
 sg13g2_buf_1 _11000_ (.A(net524),
    .X(_03567_));
 sg13g2_mux2_1 _11001_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[0] ),
    .S(net446),
    .X(_03568_));
 sg13g2_nor2_1 _11002_ (.A(net447),
    .B(_03568_),
    .Y(_03569_));
 sg13g2_nand2_1 _11003_ (.Y(_03570_),
    .A(_01712_),
    .B(net457));
 sg13g2_o21ai_1 _11004_ (.B1(_03570_),
    .Y(_03571_),
    .A1(net457),
    .A2(_03569_));
 sg13g2_o21ai_1 _11005_ (.B1(_03571_),
    .Y(_03572_),
    .A1(_03529_),
    .A2(_03562_));
 sg13g2_buf_1 _11006_ (.A(_03572_),
    .X(_03573_));
 sg13g2_buf_2 _11007_ (.A(_03573_),
    .X(_03574_));
 sg13g2_inv_2 _11008_ (.Y(\soc_I.cpu_mem_addr[0] ),
    .A(net76));
 sg13g2_inv_1 _11009_ (.Y(_03575_),
    .A(net629));
 sg13g2_buf_1 _11010_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.resetn ),
    .X(_03576_));
 sg13g2_buf_1 _11011_ (.A(_03576_),
    .X(_03577_));
 sg13g2_buf_1 _11012_ (.A(_03577_),
    .X(_03578_));
 sg13g2_nand4_1 _11013_ (.B(_03575_),
    .C(net632),
    .A(net600),
    .Y(_03579_),
    .D(net523));
 sg13g2_nand3_1 _11014_ (.B(_02007_),
    .C(net449),
    .A(_01700_),
    .Y(_03580_));
 sg13g2_inv_1 _11015_ (.Y(_03581_),
    .A(_01556_));
 sg13g2_inv_1 _11016_ (.Y(_03582_),
    .A(_01557_));
 sg13g2_nand2_1 _11017_ (.Y(_03583_),
    .A(_03581_),
    .B(_03582_));
 sg13g2_buf_1 _11018_ (.A(_03583_),
    .X(_03584_));
 sg13g2_nand2_1 _11019_ (.Y(_03585_),
    .A(net187),
    .B(_03294_));
 sg13g2_nand3_1 _11020_ (.B(_03284_),
    .C(_03285_),
    .A(net175),
    .Y(_03586_));
 sg13g2_nor2_1 _11021_ (.A(_03293_),
    .B(_03309_),
    .Y(_03587_));
 sg13g2_inv_1 _11022_ (.Y(_03588_),
    .A(_03249_));
 sg13g2_o21ai_1 _11023_ (.B1(_03588_),
    .Y(_03589_),
    .A1(_03233_),
    .A2(_03287_));
 sg13g2_nor4_1 _11024_ (.A(net146),
    .B(_03293_),
    .C(_03287_),
    .D(_03309_),
    .Y(_03590_));
 sg13g2_a221oi_1 _11025_ (.B2(_03589_),
    .C1(_03590_),
    .B1(_03587_),
    .A1(_03266_),
    .Y(_03591_),
    .A2(_03299_));
 sg13g2_mux2_1 _11026_ (.A0(_03585_),
    .A1(_03586_),
    .S(_03591_),
    .X(_03592_));
 sg13g2_nand2_1 _11027_ (.Y(_03593_),
    .A(net210),
    .B(_02526_));
 sg13g2_mux2_1 _11028_ (.A0(net310),
    .A1(net182),
    .S(_03593_),
    .X(_03594_));
 sg13g2_buf_1 _11029_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[29] ),
    .X(_03595_));
 sg13g2_o21ai_1 _11030_ (.B1(net452),
    .Y(_03596_),
    .A1(net185),
    .A2(_02612_));
 sg13g2_a22oi_1 _11031_ (.Y(_03597_),
    .B1(_02526_),
    .B2(_03596_),
    .A2(net186),
    .A1(_03595_));
 sg13g2_o21ai_1 _11032_ (.B1(_03597_),
    .Y(_03598_),
    .A1(_02531_),
    .A2(_03594_));
 sg13g2_nor2_1 _11033_ (.A(_03284_),
    .B(_03585_),
    .Y(_03599_));
 sg13g2_nor2_1 _11034_ (.A(_03598_),
    .B(_03599_),
    .Y(_03600_));
 sg13g2_and2_1 _11035_ (.A(net597),
    .B(_03600_),
    .X(_03601_));
 sg13g2_buf_1 _11036_ (.A(net597),
    .X(_03602_));
 sg13g2_buf_1 _11037_ (.A(_01792_),
    .X(_03603_));
 sg13g2_mux2_1 _11038_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[29] ),
    .S(net595),
    .X(_03604_));
 sg13g2_nor2_1 _11039_ (.A(_03602_),
    .B(_03604_),
    .Y(_03605_));
 sg13g2_a21o_1 _11040_ (.A2(_03601_),
    .A1(_03592_),
    .B1(_03605_),
    .X(_03606_));
 sg13g2_buf_1 _11041_ (.A(_03606_),
    .X(_03607_));
 sg13g2_o21ai_1 _11042_ (.B1(_01597_),
    .Y(_03608_),
    .A1(_01762_),
    .A2(_01636_));
 sg13g2_buf_1 _11043_ (.A(_03608_),
    .X(_03609_));
 sg13g2_buf_1 _11044_ (.A(_03609_),
    .X(_03610_));
 sg13g2_nor2_1 _11045_ (.A(_01797_),
    .B(net181),
    .Y(_03611_));
 sg13g2_buf_1 _11046_ (.A(_03611_),
    .X(_03612_));
 sg13g2_nand3_1 _11047_ (.B(net262),
    .C(_02693_),
    .A(net184),
    .Y(_03613_));
 sg13g2_o21ai_1 _11048_ (.B1(_03613_),
    .Y(_03614_),
    .A1(net182),
    .A2(_02693_));
 sg13g2_and2_1 _11049_ (.A(_01590_),
    .B(_01618_),
    .X(_03615_));
 sg13g2_buf_1 _11050_ (.A(_03615_),
    .X(_03616_));
 sg13g2_a21oi_1 _11051_ (.A1(net210),
    .A2(_02696_),
    .Y(_03617_),
    .B1(_01786_));
 sg13g2_o21ai_1 _11052_ (.B1(net305),
    .Y(_03618_),
    .A1(_03616_),
    .A2(_03617_));
 sg13g2_inv_1 _11053_ (.Y(_03619_),
    .A(_03618_));
 sg13g2_a221oi_1 _11054_ (.B2(_03614_),
    .C1(_03619_),
    .B1(_02696_),
    .A1(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[31] ),
    .Y(_03620_),
    .A2(_03535_));
 sg13g2_mux2_1 _11055_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[31] ),
    .S(_01792_),
    .X(_03621_));
 sg13g2_nand2_1 _11056_ (.Y(_03622_),
    .A(net527),
    .B(_03621_));
 sg13g2_o21ai_1 _11057_ (.B1(_03622_),
    .Y(_03623_),
    .A1(net527),
    .A2(_03620_));
 sg13g2_a21oi_1 _11058_ (.A1(_02989_),
    .A2(_03612_),
    .Y(_03624_),
    .B1(_03623_));
 sg13g2_buf_8 _11059_ (.A(_03624_),
    .X(_03625_));
 sg13g2_o21ai_1 _11060_ (.B1(_03461_),
    .Y(_03626_),
    .A1(_03127_),
    .A2(_03507_));
 sg13g2_nand3_1 _11061_ (.B(_03512_),
    .C(_03626_),
    .A(net175),
    .Y(_03627_));
 sg13g2_and3_1 _11062_ (.X(_03628_),
    .A(net187),
    .B(_03507_),
    .C(_03459_));
 sg13g2_nand2_1 _11063_ (.Y(_03629_),
    .A(net268),
    .B(_02677_));
 sg13g2_mux2_1 _11064_ (.A0(_01767_),
    .A1(_01784_),
    .S(_03629_),
    .X(_03630_));
 sg13g2_buf_1 _11065_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[30] ),
    .X(_03631_));
 sg13g2_o21ai_1 _11066_ (.B1(net452),
    .Y(_03632_),
    .A1(_01784_),
    .A2(_02722_));
 sg13g2_a22oi_1 _11067_ (.Y(_03633_),
    .B1(_02677_),
    .B2(_03632_),
    .A2(_01781_),
    .A1(_03631_));
 sg13g2_o21ai_1 _11068_ (.B1(_03633_),
    .Y(_03634_),
    .A1(_02670_),
    .A2(_03630_));
 sg13g2_a21oi_1 _11069_ (.A1(_03461_),
    .A2(_03628_),
    .Y(_03635_),
    .B1(_03634_));
 sg13g2_and2_1 _11070_ (.A(_03124_),
    .B(_03045_),
    .X(_03636_));
 sg13g2_buf_1 _11071_ (.A(_03636_),
    .X(_03637_));
 sg13g2_nand2b_1 _11072_ (.Y(_03638_),
    .B(_03609_),
    .A_N(_03634_));
 sg13g2_nand4_1 _11073_ (.B(_03459_),
    .C(_03461_),
    .A(net141),
    .Y(_03639_),
    .D(_03638_));
 sg13g2_a21o_1 _11074_ (.A2(_03637_),
    .A1(_03150_),
    .B1(_03639_),
    .X(_03640_));
 sg13g2_o21ai_1 _11075_ (.B1(_03512_),
    .Y(_03641_),
    .A1(_01638_),
    .A2(_03634_));
 sg13g2_a21oi_1 _11076_ (.A1(_03507_),
    .A2(_03461_),
    .Y(_03642_),
    .B1(_03641_));
 sg13g2_nand3_1 _11077_ (.B(_03637_),
    .C(_03642_),
    .A(_03150_),
    .Y(_03643_));
 sg13g2_nand4_1 _11078_ (.B(_03635_),
    .C(_03640_),
    .A(_03627_),
    .Y(_03644_),
    .D(_03643_));
 sg13g2_buf_1 _11079_ (.A(_03644_),
    .X(_03645_));
 sg13g2_nand2_1 _11080_ (.Y(_03646_),
    .A(net595),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[30] ));
 sg13g2_nand2b_1 _11081_ (.Y(_03647_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[30] ),
    .A_N(net595));
 sg13g2_a21oi_1 _11082_ (.A1(_03646_),
    .A2(_03647_),
    .Y(_03648_),
    .B1(net522));
 sg13g2_a21oi_1 _11083_ (.A1(net525),
    .A2(_03645_),
    .Y(_03649_),
    .B1(_03648_));
 sg13g2_buf_8 _11084_ (.A(_03649_),
    .X(_03650_));
 sg13g2_nand4_1 _11085_ (.B(_03607_),
    .C(_03625_),
    .A(net445),
    .Y(_03651_),
    .D(net113));
 sg13g2_buf_1 _11086_ (.A(_03651_),
    .X(_03652_));
 sg13g2_or4_1 _11087_ (.A(_02527_),
    .B(_02665_),
    .C(_02658_),
    .D(net445),
    .X(_03653_));
 sg13g2_buf_1 _11088_ (.A(_03653_),
    .X(_03654_));
 sg13g2_nand2_1 _11089_ (.Y(_03655_),
    .A(_03652_),
    .B(_03654_));
 sg13g2_nand2_1 _11090_ (.Y(_03656_),
    .A(_03216_),
    .B(_03612_));
 sg13g2_buf_1 _11091_ (.A(net527),
    .X(_03657_));
 sg13g2_buf_1 _11092_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[25] ),
    .X(_03658_));
 sg13g2_nand2_1 _11093_ (.Y(_03659_),
    .A(net177),
    .B(net307));
 sg13g2_mux2_1 _11094_ (.A0(net207),
    .A1(net213),
    .S(_03659_),
    .X(_03660_));
 sg13g2_o21ai_1 _11095_ (.B1(net362),
    .Y(_03661_),
    .A1(net174),
    .A2(_02483_));
 sg13g2_and2_1 _11096_ (.A(net307),
    .B(_03661_),
    .X(_03662_));
 sg13g2_a221oi_1 _11097_ (.B2(_03660_),
    .C1(_03662_),
    .B1(_02483_),
    .A1(_03658_),
    .Y(_03663_),
    .A2(net166));
 sg13g2_mux2_1 _11098_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[25] ),
    .S(net524),
    .X(_03664_));
 sg13g2_nand2_1 _11099_ (.Y(_03665_),
    .A(net444),
    .B(_03664_));
 sg13g2_o21ai_1 _11100_ (.B1(_03665_),
    .Y(_03666_),
    .A1(net444),
    .A2(_03663_));
 sg13g2_inv_1 _11101_ (.Y(_03667_),
    .A(_03666_));
 sg13g2_nand3_1 _11102_ (.B(_03656_),
    .C(_03667_),
    .A(net445),
    .Y(_03668_));
 sg13g2_buf_1 _11103_ (.A(_03668_),
    .X(_03669_));
 sg13g2_nand2b_1 _11104_ (.Y(_03670_),
    .B(net530),
    .A_N(_02479_));
 sg13g2_nand2_1 _11105_ (.Y(_03671_),
    .A(_03669_),
    .B(_03670_));
 sg13g2_nand2_1 _11106_ (.Y(_03672_),
    .A(_03655_),
    .B(_03671_));
 sg13g2_and2_1 _11107_ (.A(_03669_),
    .B(_03670_),
    .X(_03673_));
 sg13g2_buf_1 _11108_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[18] ),
    .X(_03674_));
 sg13g2_o21ai_1 _11109_ (.B1(_03538_),
    .Y(_03675_),
    .A1(_03549_),
    .A2(_02120_));
 sg13g2_nand3_1 _11110_ (.B(net207),
    .C(_02776_),
    .A(net177),
    .Y(_03676_));
 sg13g2_a21o_1 _11111_ (.A2(_02776_),
    .A1(net177),
    .B1(_03549_),
    .X(_03677_));
 sg13g2_a21oi_1 _11112_ (.A1(_03676_),
    .A2(_03677_),
    .Y(_03678_),
    .B1(_02124_));
 sg13g2_a221oi_1 _11113_ (.B2(_03675_),
    .C1(_03678_),
    .B1(_02776_),
    .A1(_03674_),
    .Y(_03679_),
    .A2(net166));
 sg13g2_inv_1 _11114_ (.Y(_03680_),
    .A(_03679_));
 sg13g2_a21oi_2 _11115_ (.B1(_03680_),
    .Y(_03681_),
    .A2(_03374_),
    .A1(net159));
 sg13g2_nand2_1 _11116_ (.Y(_03682_),
    .A(net165),
    .B(net142));
 sg13g2_nand2_1 _11117_ (.Y(_03683_),
    .A(net165),
    .B(net145));
 sg13g2_mux2_1 _11118_ (.A0(_03682_),
    .A1(_03683_),
    .S(_03012_),
    .X(_03684_));
 sg13g2_nand2_1 _11119_ (.Y(_03685_),
    .A(net167),
    .B(_03168_));
 sg13g2_mux2_1 _11120_ (.A0(net310),
    .A1(net174),
    .S(_03685_),
    .X(_03686_));
 sg13g2_buf_1 _11121_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[16] ),
    .X(_03687_));
 sg13g2_o21ai_1 _11122_ (.B1(net362),
    .Y(_03688_),
    .A1(net174),
    .A2(_02154_));
 sg13g2_a22oi_1 _11123_ (.Y(_03689_),
    .B1(_03168_),
    .B2(_03688_),
    .A2(net166),
    .A1(_03687_));
 sg13g2_o21ai_1 _11124_ (.B1(_03689_),
    .Y(_03690_),
    .A1(_02217_),
    .A2(_03686_));
 sg13g2_inv_1 _11125_ (.Y(_03691_),
    .A(_03690_));
 sg13g2_and4_1 _11126_ (.A(_03564_),
    .B(_03681_),
    .C(_03684_),
    .D(_03691_),
    .X(_03692_));
 sg13g2_nor2_1 _11127_ (.A(\soc_I.kianv_I.datapath_unit_I.DataLatched[16] ),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[18] ),
    .Y(_03693_));
 sg13g2_nor3_1 _11128_ (.A(_03567_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[16] ),
    .C(\soc_I.kianv_I.datapath_unit_I.ALUOut[18] ),
    .Y(_03694_));
 sg13g2_a21oi_1 _11129_ (.A1(net446),
    .A2(_03693_),
    .Y(_03695_),
    .B1(_03694_));
 sg13g2_nor2_1 _11130_ (.A(net447),
    .B(_03695_),
    .Y(_03696_));
 sg13g2_a221oi_1 _11131_ (.B2(_02964_),
    .C1(_03338_),
    .B1(net146),
    .A1(_02844_),
    .Y(_03697_),
    .A2(_02852_));
 sg13g2_o21ai_1 _11132_ (.B1(net165),
    .Y(_03698_),
    .A1(_03404_),
    .A2(_03697_));
 sg13g2_nand2b_1 _11133_ (.Y(_03699_),
    .B(net175),
    .A_N(_02784_));
 sg13g2_buf_1 _11134_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[23] ),
    .X(_03700_));
 sg13g2_o21ai_1 _11135_ (.B1(net452),
    .Y(_03701_),
    .A1(net212),
    .A2(_02243_));
 sg13g2_nand3_1 _11136_ (.B(net262),
    .C(net309),
    .A(net268),
    .Y(_03702_));
 sg13g2_o21ai_1 _11137_ (.B1(_01770_),
    .Y(_03703_),
    .A1(_01764_),
    .A2(_02262_));
 sg13g2_a21oi_1 _11138_ (.A1(_03702_),
    .A2(_03703_),
    .Y(_03704_),
    .B1(_02092_));
 sg13g2_a221oi_1 _11139_ (.B2(_03701_),
    .C1(_03704_),
    .B1(net309),
    .A1(_03700_),
    .Y(_03705_),
    .A2(_01781_));
 sg13g2_buf_1 _11140_ (.A(_03705_),
    .X(_03706_));
 sg13g2_o21ai_1 _11141_ (.B1(_03706_),
    .Y(_03707_),
    .A1(_03326_),
    .A2(_03699_));
 sg13g2_nand2_1 _11142_ (.Y(_03708_),
    .A(_03235_),
    .B(_03706_));
 sg13g2_a21o_1 _11143_ (.A2(net139),
    .A1(net140),
    .B1(_03708_),
    .X(_03709_));
 sg13g2_a21oi_1 _11144_ (.A1(_03707_),
    .A2(_03709_),
    .Y(_03710_),
    .B1(_01798_));
 sg13g2_mux2_1 _11145_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[23] ),
    .S(net595),
    .X(_03711_));
 sg13g2_nor2_1 _11146_ (.A(net522),
    .B(_03711_),
    .Y(_03712_));
 sg13g2_a21o_1 _11147_ (.A2(_03710_),
    .A1(_03698_),
    .B1(_03712_),
    .X(_03713_));
 sg13g2_buf_2 _11148_ (.A(_03713_),
    .X(_03714_));
 sg13g2_buf_1 _11149_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[17] ),
    .X(_03715_));
 sg13g2_o21ai_1 _11150_ (.B1(net415),
    .Y(_03716_),
    .A1(net182),
    .A2(_02138_));
 sg13g2_nand3_1 _11151_ (.B(net262),
    .C(_02206_),
    .A(net210),
    .Y(_03717_));
 sg13g2_a21o_1 _11152_ (.A2(_02206_),
    .A1(net210),
    .B1(net212),
    .X(_03718_));
 sg13g2_a21oi_1 _11153_ (.A1(_03717_),
    .A2(_03718_),
    .Y(_03719_),
    .B1(_02205_));
 sg13g2_a221oi_1 _11154_ (.B2(_03716_),
    .C1(_03719_),
    .B1(_02206_),
    .A1(_03715_),
    .Y(_03720_),
    .A2(net186));
 sg13g2_buf_1 _11155_ (.A(_03720_),
    .X(_03721_));
 sg13g2_mux2_1 _11156_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[17] ),
    .S(_01792_),
    .X(_03722_));
 sg13g2_nand2_1 _11157_ (.Y(_03723_),
    .A(net527),
    .B(_03722_));
 sg13g2_o21ai_1 _11158_ (.B1(_03723_),
    .Y(_03724_),
    .A1(net527),
    .A2(_03721_));
 sg13g2_nand2_1 _11159_ (.Y(_03725_),
    .A(_03317_),
    .B(net164));
 sg13g2_a21oi_1 _11160_ (.A1(_03178_),
    .A2(_03319_),
    .Y(_03726_),
    .B1(_03725_));
 sg13g2_nand2_2 _11161_ (.Y(_03727_),
    .A(net624),
    .B(_03544_));
 sg13g2_nor4_1 _11162_ (.A(_03314_),
    .B(_03316_),
    .C(_03317_),
    .D(_03727_),
    .Y(_03728_));
 sg13g2_nor3_1 _11163_ (.A(_03724_),
    .B(_03726_),
    .C(_03728_),
    .Y(_03729_));
 sg13g2_buf_1 _11164_ (.A(_03729_),
    .X(_03730_));
 sg13g2_o21ai_1 _11165_ (.B1(_03328_),
    .Y(_03731_),
    .A1(_03406_),
    .A2(_02972_));
 sg13g2_a221oi_1 _11166_ (.B2(_03233_),
    .C1(_03731_),
    .B1(net146),
    .A1(_02846_),
    .Y(_03732_),
    .A2(_02850_));
 sg13g2_xor2_1 _11167_ (.B(_03328_),
    .A(_03405_),
    .X(_03733_));
 sg13g2_nand3b_1 _11168_ (.B(_03733_),
    .C(net165),
    .Y(_03734_),
    .A_N(_03732_));
 sg13g2_nand2_1 _11169_ (.Y(_03735_),
    .A(_03231_),
    .B(_03234_));
 sg13g2_nor4_2 _11170_ (.A(net181),
    .B(_03342_),
    .C(_02852_),
    .Y(_03736_),
    .D(_03328_));
 sg13g2_buf_1 _11171_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[19] ),
    .X(_03737_));
 sg13g2_nor2_1 _11172_ (.A(_02104_),
    .B(_02106_),
    .Y(_03738_));
 sg13g2_o21ai_1 _11173_ (.B1(net415),
    .Y(_03739_),
    .A1(net182),
    .A2(_02102_));
 sg13g2_nand2_1 _11174_ (.Y(_03740_),
    .A(net210),
    .B(_03738_));
 sg13g2_mux2_1 _11175_ (.A0(net310),
    .A1(net185),
    .S(_03740_),
    .X(_03741_));
 sg13g2_nor2_1 _11176_ (.A(_02226_),
    .B(_03741_),
    .Y(_03742_));
 sg13g2_a221oi_1 _11177_ (.B2(_03739_),
    .C1(_03742_),
    .B1(_03738_),
    .A1(_03737_),
    .Y(_03743_),
    .A2(net186));
 sg13g2_nand2_1 _11178_ (.Y(_03744_),
    .A(net597),
    .B(_03743_));
 sg13g2_a21oi_1 _11179_ (.A1(_03735_),
    .A2(_03736_),
    .Y(_03745_),
    .B1(_03744_));
 sg13g2_mux2_1 _11180_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[19] ),
    .S(net595),
    .X(_03746_));
 sg13g2_nor2_1 _11181_ (.A(net522),
    .B(_03746_),
    .Y(_03747_));
 sg13g2_a21o_1 _11182_ (.A2(_03745_),
    .A1(_03734_),
    .B1(_03747_),
    .X(_03748_));
 sg13g2_buf_2 _11183_ (.A(_03748_),
    .X(_03749_));
 sg13g2_and3_1 _11184_ (.X(_03750_),
    .A(net122),
    .B(_03730_),
    .C(_03749_));
 sg13g2_o21ai_1 _11185_ (.B1(_03750_),
    .Y(_03751_),
    .A1(_03692_),
    .A2(_03696_));
 sg13g2_buf_1 _11186_ (.A(_03584_),
    .X(_03752_));
 sg13g2_a21oi_1 _11187_ (.A1(_03521_),
    .A2(_03524_),
    .Y(_03753_),
    .B1(_03727_));
 sg13g2_mux2_1 _11188_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[28] ),
    .S(_03566_),
    .X(_03754_));
 sg13g2_buf_1 _11189_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[28] ),
    .X(_03755_));
 sg13g2_nand2_1 _11190_ (.Y(_03756_),
    .A(net177),
    .B(_02521_));
 sg13g2_mux2_1 _11191_ (.A0(net207),
    .A1(net213),
    .S(_03756_),
    .X(_03757_));
 sg13g2_o21ai_1 _11192_ (.B1(net362),
    .Y(_03758_),
    .A1(net174),
    .A2(_02596_));
 sg13g2_and2_1 _11193_ (.A(_02521_),
    .B(_03758_),
    .X(_03759_));
 sg13g2_a221oi_1 _11194_ (.B2(_03757_),
    .C1(_03759_),
    .B1(_02596_),
    .A1(_03755_),
    .Y(_03760_),
    .A2(net166));
 sg13g2_buf_1 _11195_ (.A(_03760_),
    .X(_03761_));
 sg13g2_nand2_1 _11196_ (.Y(_03762_),
    .A(_03564_),
    .B(_03761_));
 sg13g2_o21ai_1 _11197_ (.B1(_03762_),
    .Y(_03763_),
    .A1(net525),
    .A2(_03754_));
 sg13g2_nand2b_1 _11198_ (.Y(_03764_),
    .B(_03763_),
    .A_N(_03753_));
 sg13g2_buf_1 _11199_ (.A(_03582_),
    .X(_03765_));
 sg13g2_or3_1 _11200_ (.A(_03249_),
    .B(_03288_),
    .C(_03368_),
    .X(_03766_));
 sg13g2_nor2b_1 _11201_ (.A(_03249_),
    .B_N(_03287_),
    .Y(_03767_));
 sg13g2_nand3_1 _11202_ (.B(net139),
    .C(_03588_),
    .A(net140),
    .Y(_03768_));
 sg13g2_nand3b_1 _11203_ (.B(_03366_),
    .C(_03768_),
    .Y(_03769_),
    .A_N(_03767_));
 sg13g2_nand4_1 _11204_ (.B(_03398_),
    .C(_03766_),
    .A(_03396_),
    .Y(_03770_),
    .D(_03769_));
 sg13g2_buf_1 _11205_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[21] ),
    .X(_03771_));
 sg13g2_buf_1 _11206_ (.A(net185),
    .X(_03772_));
 sg13g2_o21ai_1 _11207_ (.B1(net362),
    .Y(_03773_),
    .A1(net173),
    .A2(_02042_));
 sg13g2_nand3_1 _11208_ (.B(net262),
    .C(_02038_),
    .A(net177),
    .Y(_03774_));
 sg13g2_o21ai_1 _11209_ (.B1(net213),
    .Y(_03775_),
    .A1(net263),
    .A2(_02235_));
 sg13g2_a21oi_1 _11210_ (.A1(_03774_),
    .A2(_03775_),
    .Y(_03776_),
    .B1(_02255_));
 sg13g2_a221oi_1 _11211_ (.B2(_03773_),
    .C1(_03776_),
    .B1(_02038_),
    .A1(_03771_),
    .Y(_03777_),
    .A2(net176));
 sg13g2_buf_1 _11212_ (.A(_03777_),
    .X(_03778_));
 sg13g2_mux2_1 _11213_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[21] ),
    .S(net524),
    .X(_03779_));
 sg13g2_nand2_1 _11214_ (.Y(_03780_),
    .A(net444),
    .B(_03779_));
 sg13g2_o21ai_1 _11215_ (.B1(_03780_),
    .Y(_03781_),
    .A1(net444),
    .A2(_03778_));
 sg13g2_a221oi_1 _11216_ (.B2(_03770_),
    .C1(_03781_),
    .B1(net164),
    .A1(_03581_),
    .Y(_03782_),
    .A2(net521));
 sg13g2_inv_1 _11217_ (.Y(_03783_),
    .A(_02514_));
 sg13g2_or4_1 _11218_ (.A(_02099_),
    .B(_02039_),
    .C(_02074_),
    .D(_03783_),
    .X(_03784_));
 sg13g2_nor4_1 _11219_ (.A(_02150_),
    .B(_02134_),
    .C(_02117_),
    .D(_03784_),
    .Y(_03785_));
 sg13g2_a22oi_1 _11220_ (.Y(_03786_),
    .B1(_03785_),
    .B2(net457),
    .A2(_03782_),
    .A1(_03764_));
 sg13g2_a221oi_1 _11221_ (.B2(_03752_),
    .C1(_03786_),
    .B1(_03751_),
    .A1(_03652_),
    .Y(_03787_),
    .A2(_03654_));
 sg13g2_buf_2 _11222_ (.A(_03787_),
    .X(_03788_));
 sg13g2_mux2_1 _11223_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[4] ),
    .S(net524),
    .X(_03789_));
 sg13g2_a21oi_1 _11224_ (.A1(_02321_),
    .A2(_03423_),
    .Y(_03790_),
    .B1(_03419_));
 sg13g2_and3_1 _11225_ (.X(_03791_),
    .A(_01639_),
    .B(_03419_),
    .C(_03423_));
 sg13g2_buf_1 _11226_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[4] ),
    .X(_03792_));
 sg13g2_nand2_1 _11227_ (.Y(_03793_),
    .A(_02410_),
    .B(_02412_));
 sg13g2_o21ai_1 _11228_ (.B1(_03537_),
    .Y(_03794_),
    .A1(net185),
    .A2(_02414_));
 sg13g2_nand3_1 _11229_ (.B(net262),
    .C(_03793_),
    .A(net210),
    .Y(_03795_));
 sg13g2_o21ai_1 _11230_ (.B1(_01771_),
    .Y(_03796_),
    .A1(_01764_),
    .A2(_02853_));
 sg13g2_a21oi_1 _11231_ (.A1(_03795_),
    .A2(_03796_),
    .Y(_03797_),
    .B1(_02401_));
 sg13g2_a221oi_1 _11232_ (.B2(_03794_),
    .C1(_03797_),
    .B1(_03793_),
    .A1(_03792_),
    .Y(_03798_),
    .A2(_01782_));
 sg13g2_inv_1 _11233_ (.Y(_03799_),
    .A(_03798_));
 sg13g2_a221oi_1 _11234_ (.B2(_02321_),
    .C1(_03799_),
    .B1(_03791_),
    .A1(_03544_),
    .Y(_03800_),
    .A2(_03790_));
 sg13g2_buf_1 _11235_ (.A(_03800_),
    .X(_03801_));
 sg13g2_nor2_1 _11236_ (.A(net444),
    .B(_03801_),
    .Y(_03802_));
 sg13g2_a21oi_1 _11237_ (.A1(net444),
    .A2(_03789_),
    .Y(_03803_),
    .B1(_03802_));
 sg13g2_buf_1 _11238_ (.A(_03803_),
    .X(_03804_));
 sg13g2_nand2_1 _11239_ (.Y(_03805_),
    .A(_02397_),
    .B(net530));
 sg13g2_o21ai_1 _11240_ (.B1(_03805_),
    .Y(_03806_),
    .A1(net530),
    .A2(net119));
 sg13g2_buf_1 _11241_ (.A(_03806_),
    .X(_03807_));
 sg13g2_nor2_1 _11242_ (.A(_01573_),
    .B(_02282_),
    .Y(_03808_));
 sg13g2_nand3_1 _11243_ (.B(_02311_),
    .C(_02897_),
    .A(net147),
    .Y(_03809_));
 sg13g2_nand3_1 _11244_ (.B(_02301_),
    .C(net183),
    .A(_02651_),
    .Y(_03810_));
 sg13g2_nand3_1 _11245_ (.B(_03809_),
    .C(_03810_),
    .A(_03064_),
    .Y(_03811_));
 sg13g2_nand3_1 _11246_ (.B(_02900_),
    .C(_02897_),
    .A(_02651_),
    .Y(_03812_));
 sg13g2_nand3_1 _11247_ (.B(_02313_),
    .C(_02903_),
    .A(_03014_),
    .Y(_03813_));
 sg13g2_nand3_1 _11248_ (.B(_03812_),
    .C(_03813_),
    .A(_02912_),
    .Y(_03814_));
 sg13g2_xnor2_1 _11249_ (.Y(_03815_),
    .A(_01758_),
    .B(_02299_));
 sg13g2_nor3_1 _11250_ (.A(net308),
    .B(net183),
    .C(_03815_),
    .Y(_03816_));
 sg13g2_nand3_1 _11251_ (.B(net183),
    .C(_03815_),
    .A(net308),
    .Y(_03817_));
 sg13g2_nand2b_1 _11252_ (.Y(_03818_),
    .B(_03817_),
    .A_N(_03816_));
 sg13g2_a21oi_1 _11253_ (.A1(_03811_),
    .A2(_03814_),
    .Y(_03819_),
    .B1(_03818_));
 sg13g2_nor3_1 _11254_ (.A(_01764_),
    .B(_01768_),
    .C(_02891_),
    .Y(_03820_));
 sg13g2_a21oi_1 _11255_ (.A1(_02621_),
    .A2(_02296_),
    .Y(_03821_),
    .B1(_01786_));
 sg13g2_o21ai_1 _11256_ (.B1(net266),
    .Y(_03822_),
    .A1(_03820_),
    .A2(_03821_));
 sg13g2_buf_1 _11257_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[3] ),
    .X(_03823_));
 sg13g2_o21ai_1 _11258_ (.B1(net452),
    .Y(_03824_),
    .A1(net185),
    .A2(net266));
 sg13g2_a22oi_1 _11259_ (.Y(_03825_),
    .B1(_02296_),
    .B2(_03824_),
    .A2(net186),
    .A1(_03823_));
 sg13g2_and2_1 _11260_ (.A(_03822_),
    .B(_03825_),
    .X(_03826_));
 sg13g2_o21ai_1 _11261_ (.B1(_03826_),
    .Y(_03827_),
    .A1(net181),
    .A2(_03819_));
 sg13g2_nand2_1 _11262_ (.Y(_03828_),
    .A(net595),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[3] ));
 sg13g2_nand2b_1 _11263_ (.Y(_03829_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[3] ),
    .A_N(net599));
 sg13g2_a21oi_1 _11264_ (.A1(_03828_),
    .A2(_03829_),
    .Y(_03830_),
    .B1(net597));
 sg13g2_a21oi_1 _11265_ (.A1(_03602_),
    .A2(_03827_),
    .Y(_03831_),
    .B1(_03830_));
 sg13g2_buf_1 _11266_ (.A(_03831_),
    .X(_03832_));
 sg13g2_and2_1 _11267_ (.A(net445),
    .B(_01800_),
    .X(_03833_));
 sg13g2_a22oi_1 _11268_ (.Y(_03834_),
    .B1(net118),
    .B2(_03833_),
    .A2(_03808_),
    .A1(net530));
 sg13g2_buf_1 _11269_ (.A(_03834_),
    .X(_03835_));
 sg13g2_nand2_1 _11270_ (.Y(_03836_),
    .A(_02622_),
    .B(net308));
 sg13g2_mux2_1 _11271_ (.A0(_01768_),
    .A1(net173),
    .S(_03836_),
    .X(_03837_));
 sg13g2_buf_1 _11272_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[2] ),
    .X(_03838_));
 sg13g2_o21ai_1 _11273_ (.B1(net415),
    .Y(_03839_),
    .A1(_03548_),
    .A2(_02272_));
 sg13g2_a22oi_1 _11274_ (.Y(_03840_),
    .B1(net308),
    .B2(_03839_),
    .A2(net186),
    .A1(_03838_));
 sg13g2_o21ai_1 _11275_ (.B1(_03840_),
    .Y(_03841_),
    .A1(_02299_),
    .A2(_03837_));
 sg13g2_xnor2_1 _11276_ (.Y(_03842_),
    .A(_03217_),
    .B(_02314_));
 sg13g2_nand3_1 _11277_ (.B(_02315_),
    .C(_02319_),
    .A(net187),
    .Y(_03843_));
 sg13g2_a21oi_1 _11278_ (.A1(_03064_),
    .A2(_03842_),
    .Y(_03844_),
    .B1(_03843_));
 sg13g2_nor2_1 _11279_ (.A(_03841_),
    .B(_03844_),
    .Y(_03845_));
 sg13g2_inv_1 _11280_ (.Y(_03846_),
    .A(\soc_I.kianv_I.datapath_unit_I.ALUOut[2] ));
 sg13g2_nand2_1 _11281_ (.Y(_03847_),
    .A(net599),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[2] ));
 sg13g2_o21ai_1 _11282_ (.B1(_03847_),
    .Y(_03848_),
    .A1(_03603_),
    .A2(_03846_));
 sg13g2_nand2_1 _11283_ (.Y(_03849_),
    .A(_01798_),
    .B(_03848_));
 sg13g2_o21ai_1 _11284_ (.B1(_03849_),
    .Y(_03850_),
    .A1(net527),
    .A2(_03845_));
 sg13g2_buf_1 _11285_ (.A(_03850_),
    .X(_03851_));
 sg13g2_and2_1 _11286_ (.A(_02268_),
    .B(net530),
    .X(_03852_));
 sg13g2_a21oi_1 _11287_ (.A1(net445),
    .A2(_03851_),
    .Y(_03853_),
    .B1(_03852_));
 sg13g2_buf_2 _11288_ (.A(_03853_),
    .X(_03854_));
 sg13g2_nand2b_1 _11289_ (.Y(_03855_),
    .B(_03854_),
    .A_N(_03835_));
 sg13g2_and2_1 _11290_ (.A(_02881_),
    .B(_02885_),
    .X(_03856_));
 sg13g2_buf_1 _11291_ (.A(_03856_),
    .X(_03857_));
 sg13g2_nor2_1 _11292_ (.A(net152),
    .B(_02876_),
    .Y(_03858_));
 sg13g2_and2_1 _11293_ (.A(_02871_),
    .B(_02874_),
    .X(_03859_));
 sg13g2_and3_1 _11294_ (.X(_03860_),
    .A(_02685_),
    .B(_02876_),
    .C(_03859_));
 sg13g2_a21oi_1 _11295_ (.A1(_03857_),
    .A2(_03858_),
    .Y(_03861_),
    .B1(_03860_));
 sg13g2_nor2_1 _11296_ (.A(_02685_),
    .B(_02946_),
    .Y(_03862_));
 sg13g2_a21oi_1 _11297_ (.A1(_02917_),
    .A2(_02921_),
    .Y(_03863_),
    .B1(_02926_));
 sg13g2_nor2_1 _11298_ (.A(_02928_),
    .B(_02931_),
    .Y(_03864_));
 sg13g2_nor4_1 _11299_ (.A(_02701_),
    .B(_02876_),
    .C(_03863_),
    .D(_03864_),
    .Y(_03865_));
 sg13g2_a21oi_1 _11300_ (.A1(_03862_),
    .A2(_02962_),
    .Y(_03866_),
    .B1(_03865_));
 sg13g2_mux2_1 _11301_ (.A0(_03861_),
    .A1(_03866_),
    .S(_03384_),
    .X(_03867_));
 sg13g2_a21oi_1 _11302_ (.A1(net268),
    .A2(_02937_),
    .Y(_03868_),
    .B1(net212));
 sg13g2_or2_1 _11303_ (.X(_03869_),
    .B(_03868_),
    .A(_03616_));
 sg13g2_inv_1 _11304_ (.Y(_03870_),
    .A(_02936_));
 sg13g2_o21ai_1 _11305_ (.B1(_03870_),
    .Y(_03871_),
    .A1(net212),
    .A2(_02935_));
 sg13g2_buf_1 _11306_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[9] ),
    .X(_03872_));
 sg13g2_nand2_1 _11307_ (.Y(_03873_),
    .A(_02213_),
    .B(net325));
 sg13g2_mux2_1 _11308_ (.A0(_02937_),
    .A1(_03872_),
    .S(_03873_),
    .X(_03874_));
 sg13g2_a22oi_1 _11309_ (.Y(_03875_),
    .B1(_03874_),
    .B2(_01766_),
    .A2(_03871_),
    .A1(_03869_));
 sg13g2_inv_1 _11310_ (.Y(_03876_),
    .A(_03875_));
 sg13g2_nor2b_1 _11311_ (.A(_03857_),
    .B_N(_02962_),
    .Y(_03877_));
 sg13g2_nor3_1 _11312_ (.A(_03859_),
    .B(_03863_),
    .C(_03864_),
    .Y(_03878_));
 sg13g2_nand2_1 _11313_ (.Y(_03879_),
    .A(_02958_),
    .B(_02956_));
 sg13g2_a21oi_1 _11314_ (.A1(_02953_),
    .A2(_02955_),
    .Y(_03880_),
    .B1(_02960_));
 sg13g2_nand2_1 _11315_ (.Y(_03881_),
    .A(_03879_),
    .B(_03880_));
 sg13g2_mux4_1 _11316_ (.S0(_03217_),
    .A0(_03015_),
    .A1(_03877_),
    .A2(_03878_),
    .A3(_03881_),
    .S1(_02946_),
    .X(_03882_));
 sg13g2_nor3_1 _11317_ (.A(_01797_),
    .B(_03876_),
    .C(_03882_),
    .Y(_03883_));
 sg13g2_mux2_1 _11318_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[9] ),
    .S(_01792_),
    .X(_03884_));
 sg13g2_nand3_1 _11319_ (.B(net181),
    .C(_03875_),
    .A(net624),
    .Y(_03885_));
 sg13g2_o21ai_1 _11320_ (.B1(_03885_),
    .Y(_03886_),
    .A1(net624),
    .A2(_03884_));
 sg13g2_a21oi_1 _11321_ (.A1(_03867_),
    .A2(_03883_),
    .Y(_03887_),
    .B1(_03886_));
 sg13g2_buf_1 _11322_ (.A(_03887_),
    .X(_03888_));
 sg13g2_mux2_1 _11323_ (.A0(_03412_),
    .A1(_03418_),
    .S(_02321_),
    .X(_03889_));
 sg13g2_buf_1 _11324_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[6] ),
    .X(_03890_));
 sg13g2_o21ai_1 _11325_ (.B1(net452),
    .Y(_03891_),
    .A1(net212),
    .A2(_02343_));
 sg13g2_nand3_1 _11326_ (.B(net262),
    .C(_03478_),
    .A(_02621_),
    .Y(_03892_));
 sg13g2_o21ai_1 _11327_ (.B1(_01770_),
    .Y(_03893_),
    .A1(_01764_),
    .A2(_02916_));
 sg13g2_a21oi_1 _11328_ (.A1(_03892_),
    .A2(_03893_),
    .Y(_03894_),
    .B1(_02867_));
 sg13g2_a221oi_1 _11329_ (.B2(_03891_),
    .C1(_03894_),
    .B1(_03478_),
    .A1(_03890_),
    .Y(_03895_),
    .A2(_01782_));
 sg13g2_o21ai_1 _11330_ (.B1(_03895_),
    .Y(_03896_),
    .A1(_03434_),
    .A2(_03437_));
 sg13g2_nand2_1 _11331_ (.Y(_03897_),
    .A(_03610_),
    .B(_03895_));
 sg13g2_o21ai_1 _11332_ (.B1(_03897_),
    .Y(_03898_),
    .A1(_03889_),
    .A2(_03896_));
 sg13g2_buf_1 _11333_ (.A(_03898_),
    .X(_03899_));
 sg13g2_mux2_1 _11334_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[6] ),
    .S(net599),
    .X(_03900_));
 sg13g2_nor2_1 _11335_ (.A(net597),
    .B(_03900_),
    .Y(_03901_));
 sg13g2_a21oi_1 _11336_ (.A1(net525),
    .A2(_03899_),
    .Y(_03902_),
    .B1(_03901_));
 sg13g2_nor2_1 _11337_ (.A(net128),
    .B(_03902_),
    .Y(_03903_));
 sg13g2_nand2_1 _11338_ (.Y(_03904_),
    .A(net268),
    .B(_02192_));
 sg13g2_mux2_1 _11339_ (.A0(net310),
    .A1(net212),
    .S(_03904_),
    .X(_03905_));
 sg13g2_buf_1 _11340_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[12] ),
    .X(_03906_));
 sg13g2_o21ai_1 _11341_ (.B1(net452),
    .Y(_03907_),
    .A1(_01784_),
    .A2(_01871_));
 sg13g2_a22oi_1 _11342_ (.Y(_03908_),
    .B1(_02192_),
    .B2(_03907_),
    .A2(_01781_),
    .A1(_03906_));
 sg13g2_o21ai_1 _11343_ (.B1(_03908_),
    .Y(_03909_),
    .A1(_02837_),
    .A2(_03905_));
 sg13g2_nor2_1 _11344_ (.A(_02029_),
    .B(_03909_),
    .Y(_03910_));
 sg13g2_a21oi_1 _11345_ (.A1(_01638_),
    .A2(_03380_),
    .Y(_03911_),
    .B1(_03909_));
 sg13g2_a21oi_1 _11346_ (.A1(_03008_),
    .A2(_03910_),
    .Y(_03912_),
    .B1(_03911_));
 sg13g2_nand2_1 _11347_ (.Y(_03913_),
    .A(_01792_),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[12] ));
 sg13g2_nand2b_1 _11348_ (.Y(_03914_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[12] ),
    .A_N(_01792_));
 sg13g2_a21oi_1 _11349_ (.A1(_03913_),
    .A2(_03914_),
    .Y(_03915_),
    .B1(_01796_));
 sg13g2_a221oi_1 _11350_ (.B2(_03563_),
    .C1(_03915_),
    .B1(_03912_),
    .A1(_03378_),
    .Y(_03916_),
    .A2(net164));
 sg13g2_buf_8 _11351_ (.A(_03916_),
    .X(_03917_));
 sg13g2_and2_1 _11352_ (.A(_03583_),
    .B(net131),
    .X(_03918_));
 sg13g2_nor4_1 _11353_ (.A(_02337_),
    .B(_01943_),
    .C(_01864_),
    .D(net445),
    .Y(_03919_));
 sg13g2_a21o_1 _11354_ (.A2(_03918_),
    .A1(_03903_),
    .B1(_03919_),
    .X(_03920_));
 sg13g2_buf_1 _11355_ (.A(_03920_),
    .X(_03921_));
 sg13g2_buf_1 _11356_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[15] ),
    .X(_03922_));
 sg13g2_o21ai_1 _11357_ (.B1(net415),
    .Y(_03923_),
    .A1(net182),
    .A2(_01831_));
 sg13g2_nand3_1 _11358_ (.B(net262),
    .C(_02182_),
    .A(net184),
    .Y(_03924_));
 sg13g2_a21o_1 _11359_ (.A2(_02182_),
    .A1(net184),
    .B1(net185),
    .X(_03925_));
 sg13g2_a21oi_1 _11360_ (.A1(_03924_),
    .A2(_03925_),
    .Y(_03926_),
    .B1(_02185_));
 sg13g2_a221oi_1 _11361_ (.B2(_03923_),
    .C1(_03926_),
    .B1(_02182_),
    .A1(_03922_),
    .Y(_03927_),
    .A2(net176));
 sg13g2_inv_1 _11362_ (.Y(_03928_),
    .A(_03927_));
 sg13g2_nand2_1 _11363_ (.Y(_03929_),
    .A(net599),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[15] ));
 sg13g2_nand2b_1 _11364_ (.Y(_03930_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[15] ),
    .A_N(net599));
 sg13g2_a21oi_1 _11365_ (.A1(_03929_),
    .A2(_03930_),
    .Y(_03931_),
    .B1(net597));
 sg13g2_a221oi_1 _11366_ (.B2(_03563_),
    .C1(_03931_),
    .B1(_03928_),
    .A1(_03246_),
    .Y(_03932_),
    .A2(net164));
 sg13g2_buf_1 _11367_ (.A(_03932_),
    .X(_03933_));
 sg13g2_buf_1 _11368_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[7] ),
    .X(_03934_));
 sg13g2_o21ai_1 _11369_ (.B1(net452),
    .Y(_03935_),
    .A1(_01785_),
    .A2(_02334_));
 sg13g2_nand3_1 _11370_ (.B(_03540_),
    .C(_02948_),
    .A(_02213_),
    .Y(_03936_));
 sg13g2_o21ai_1 _11371_ (.B1(_01770_),
    .Y(_03937_),
    .A1(_01764_),
    .A2(_02920_));
 sg13g2_a21oi_1 _11372_ (.A1(_03936_),
    .A2(_03937_),
    .Y(_03938_),
    .B1(_02863_));
 sg13g2_a221oi_1 _11373_ (.B2(_03935_),
    .C1(_03938_),
    .B1(_02948_),
    .A1(_03934_),
    .Y(_03939_),
    .A2(_01781_));
 sg13g2_buf_1 _11374_ (.A(_03939_),
    .X(_03940_));
 sg13g2_nand3b_1 _11375_ (.B(_03487_),
    .C(_03940_),
    .Y(_03941_),
    .A_N(_03484_));
 sg13g2_nand3b_1 _11376_ (.B(_03491_),
    .C(_03940_),
    .Y(_03942_),
    .A_N(_03484_));
 sg13g2_mux2_1 _11377_ (.A0(_03941_),
    .A1(_03942_),
    .S(_03384_),
    .X(_03943_));
 sg13g2_buf_1 _11378_ (.A(_03610_),
    .X(_03944_));
 sg13g2_nand2_1 _11379_ (.Y(_03945_),
    .A(net172),
    .B(_03940_));
 sg13g2_nor2_1 _11380_ (.A(_03005_),
    .B(_02918_),
    .Y(_03946_));
 sg13g2_nor2_1 _11381_ (.A(net173),
    .B(_03946_),
    .Y(_03947_));
 sg13g2_a21oi_1 _11382_ (.A1(net207),
    .A2(_03946_),
    .Y(_03948_),
    .B1(_03947_));
 sg13g2_buf_1 _11383_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[5] ),
    .X(_03949_));
 sg13g2_inv_1 _11384_ (.Y(_03950_),
    .A(_02918_));
 sg13g2_o21ai_1 _11385_ (.B1(_03537_),
    .Y(_03951_),
    .A1(_03772_),
    .A2(_02462_));
 sg13g2_a22oi_1 _11386_ (.Y(_03952_),
    .B1(_03950_),
    .B2(_03951_),
    .A2(_03535_),
    .A1(_03949_));
 sg13g2_o21ai_1 _11387_ (.B1(_03952_),
    .Y(_03953_),
    .A1(_02432_),
    .A2(_03948_));
 sg13g2_a221oi_1 _11388_ (.B2(_03945_),
    .C1(_03953_),
    .B1(_03943_),
    .A1(_03545_),
    .Y(_03954_),
    .A2(_03386_));
 sg13g2_nor2_1 _11389_ (.A(\soc_I.kianv_I.datapath_unit_I.DataLatched[5] ),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[7] ),
    .Y(_03955_));
 sg13g2_nor3_1 _11390_ (.A(_03603_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[5] ),
    .C(\soc_I.kianv_I.datapath_unit_I.ALUOut[7] ),
    .Y(_03956_));
 sg13g2_a21oi_1 _11391_ (.A1(net524),
    .A2(_03955_),
    .Y(_03957_),
    .B1(_03956_));
 sg13g2_nor3_1 _11392_ (.A(net522),
    .B(_01559_),
    .C(_03957_),
    .Y(_03958_));
 sg13g2_a21o_1 _11393_ (.A2(_03954_),
    .A1(_03534_),
    .B1(_03958_),
    .X(_03959_));
 sg13g2_nor4_1 _11394_ (.A(_02425_),
    .B(_02330_),
    .C(_01826_),
    .D(net445),
    .Y(_03960_));
 sg13g2_a21o_1 _11395_ (.A2(_03959_),
    .A1(_03933_),
    .B1(_03960_),
    .X(_03961_));
 sg13g2_buf_1 _11396_ (.A(_03961_),
    .X(_03962_));
 sg13g2_buf_1 _11397_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[13] ),
    .X(_03963_));
 sg13g2_o21ai_1 _11398_ (.B1(net362),
    .Y(_03964_),
    .A1(net174),
    .A2(_01908_));
 sg13g2_nand3_1 _11399_ (.B(_03541_),
    .C(_02170_),
    .A(_02623_),
    .Y(_03965_));
 sg13g2_a21o_1 _11400_ (.A2(_02170_),
    .A1(_02622_),
    .B1(net173),
    .X(_03966_));
 sg13g2_a21oi_1 _11401_ (.A1(_03965_),
    .A2(_03966_),
    .Y(_03967_),
    .B1(_02173_));
 sg13g2_a221oi_1 _11402_ (.B2(_03964_),
    .C1(_03967_),
    .B1(_02170_),
    .A1(_03963_),
    .Y(_03968_),
    .A2(net176));
 sg13g2_nor2_1 _11403_ (.A(net181),
    .B(_03364_),
    .Y(_03969_));
 sg13g2_nand4_1 _11404_ (.B(net139),
    .C(_03588_),
    .A(net140),
    .Y(_03970_),
    .D(_03969_));
 sg13g2_and2_1 _11405_ (.A(net187),
    .B(_03364_),
    .X(_03971_));
 sg13g2_a22oi_1 _11406_ (.Y(_03972_),
    .B1(_03971_),
    .B2(_03249_),
    .A2(_03969_),
    .A1(_03767_));
 sg13g2_nand2b_1 _11407_ (.Y(_03973_),
    .B(_03971_),
    .A_N(_03287_));
 sg13g2_a21o_1 _11408_ (.A2(net139),
    .A1(net140),
    .B1(_03973_),
    .X(_03974_));
 sg13g2_nand4_1 _11409_ (.B(_03970_),
    .C(_03972_),
    .A(_03968_),
    .Y(_03975_),
    .D(_03974_));
 sg13g2_buf_1 _11410_ (.A(_03975_),
    .X(_03976_));
 sg13g2_nand2_1 _11411_ (.Y(_03977_),
    .A(net175),
    .B(_03123_));
 sg13g2_xnor2_1 _11412_ (.Y(_03978_),
    .A(_03007_),
    .B(_02168_));
 sg13g2_nand2_1 _11413_ (.Y(_03979_),
    .A(net175),
    .B(_03978_));
 sg13g2_mux2_1 _11414_ (.A0(_03977_),
    .A1(_03979_),
    .S(_03150_),
    .X(_03980_));
 sg13g2_buf_1 _11415_ (.A(_03980_),
    .X(_03981_));
 sg13g2_buf_1 _11416_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[14] ),
    .X(_03982_));
 sg13g2_o21ai_1 _11417_ (.B1(_03538_),
    .Y(_03983_),
    .A1(net173),
    .A2(_01889_));
 sg13g2_nand3_1 _11418_ (.B(net207),
    .C(_02834_),
    .A(_02623_),
    .Y(_03984_));
 sg13g2_a21o_1 _11419_ (.A2(_02834_),
    .A1(net184),
    .B1(net173),
    .X(_03985_));
 sg13g2_a21oi_1 _11420_ (.A1(_03984_),
    .A2(_03985_),
    .Y(_03986_),
    .B1(_01892_));
 sg13g2_a221oi_1 _11421_ (.B2(_03983_),
    .C1(_03986_),
    .B1(_02834_),
    .A1(_03982_),
    .Y(_03987_),
    .A2(net176));
 sg13g2_buf_1 _11422_ (.A(_03987_),
    .X(_03988_));
 sg13g2_and2_1 _11423_ (.A(net525),
    .B(_03988_),
    .X(_03989_));
 sg13g2_nand3b_1 _11424_ (.B(_03981_),
    .C(_03989_),
    .Y(_03990_),
    .A_N(_03976_));
 sg13g2_nor2_1 _11425_ (.A(\soc_I.kianv_I.datapath_unit_I.DataLatched[13] ),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[14] ),
    .Y(_03991_));
 sg13g2_nor3_1 _11426_ (.A(net524),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[13] ),
    .C(\soc_I.kianv_I.datapath_unit_I.ALUOut[14] ),
    .Y(_03992_));
 sg13g2_a21o_1 _11427_ (.A2(_03991_),
    .A1(_03566_),
    .B1(_03992_),
    .X(_03993_));
 sg13g2_a21oi_1 _11428_ (.A1(_03657_),
    .A2(_03993_),
    .Y(_03994_),
    .B1(net530));
 sg13g2_inv_1 _11429_ (.Y(_03995_),
    .A(_01883_));
 sg13g2_nor4_1 _11430_ (.A(_01929_),
    .B(_01959_),
    .C(_01979_),
    .D(_01903_),
    .Y(_03996_));
 sg13g2_nand3_1 _11431_ (.B(net530),
    .C(_03996_),
    .A(_03995_),
    .Y(_03997_));
 sg13g2_mux2_1 _11432_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[11] ),
    .S(_01792_),
    .X(_03998_));
 sg13g2_nor2_1 _11433_ (.A(net624),
    .B(_03998_),
    .Y(_03999_));
 sg13g2_buf_1 _11434_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[11] ),
    .X(_04000_));
 sg13g2_o21ai_1 _11435_ (.B1(_01787_),
    .Y(_04001_),
    .A1(_01785_),
    .A2(_02021_));
 sg13g2_nand3_1 _11436_ (.B(_03540_),
    .C(_03051_),
    .A(net268),
    .Y(_04002_));
 sg13g2_a21o_1 _11437_ (.A2(_03051_),
    .A1(net268),
    .B1(_01784_),
    .X(_04003_));
 sg13g2_a21oi_1 _11438_ (.A1(_04002_),
    .A2(_04003_),
    .Y(_04004_),
    .B1(_01984_));
 sg13g2_a221oi_1 _11439_ (.B2(_04001_),
    .C1(_04004_),
    .B1(_03051_),
    .A1(_04000_),
    .Y(_04005_),
    .A2(_01781_));
 sg13g2_buf_1 _11440_ (.A(_04005_),
    .X(_04006_));
 sg13g2_nor2_1 _11441_ (.A(_01797_),
    .B(_03389_),
    .Y(_04007_));
 sg13g2_and4_1 _11442_ (.A(_02914_),
    .B(_03233_),
    .C(_04006_),
    .D(_04007_),
    .X(_04008_));
 sg13g2_nand3_1 _11443_ (.B(_03389_),
    .C(_04006_),
    .A(net624),
    .Y(_04009_));
 sg13g2_nor2_1 _11444_ (.A(_03231_),
    .B(_04009_),
    .Y(_04010_));
 sg13g2_nand3_1 _11445_ (.B(net181),
    .C(_04006_),
    .A(net624),
    .Y(_04011_));
 sg13g2_o21ai_1 _11446_ (.B1(_04011_),
    .Y(_04012_),
    .A1(_03234_),
    .A2(_04009_));
 sg13g2_nor4_1 _11447_ (.A(_03999_),
    .B(_04008_),
    .C(_04010_),
    .D(_04012_),
    .Y(_04013_));
 sg13g2_buf_2 _11448_ (.A(_04013_),
    .X(_04014_));
 sg13g2_xnor2_1 _11449_ (.Y(_04015_),
    .A(net150),
    .B(_03081_));
 sg13g2_nand2_1 _11450_ (.Y(_04016_),
    .A(net187),
    .B(_04015_));
 sg13g2_nor4_2 _11451_ (.A(_03356_),
    .B(_02912_),
    .C(_03097_),
    .Y(_04017_),
    .D(_04016_));
 sg13g2_nor3_1 _11452_ (.A(_03097_),
    .B(_03137_),
    .C(_04016_),
    .Y(_04018_));
 sg13g2_nand2_1 _11453_ (.Y(_04019_),
    .A(net187),
    .B(_03496_));
 sg13g2_a221oi_1 _11454_ (.B2(_03077_),
    .C1(_04019_),
    .B1(_03073_),
    .A1(_02305_),
    .Y(_04020_),
    .A2(_03064_));
 sg13g2_nor2_1 _11455_ (.A(net181),
    .B(_04015_),
    .Y(_04021_));
 sg13g2_nand2_1 _11456_ (.Y(_04022_),
    .A(net210),
    .B(_01995_));
 sg13g2_mux2_1 _11457_ (.A0(net310),
    .A1(_03548_),
    .S(_04022_),
    .X(_04023_));
 sg13g2_buf_1 _11458_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[10] ),
    .X(_04024_));
 sg13g2_o21ai_1 _11459_ (.B1(net415),
    .Y(_04025_),
    .A1(net185),
    .A2(_01963_));
 sg13g2_a22oi_1 _11460_ (.Y(_04026_),
    .B1(_01995_),
    .B2(_04025_),
    .A2(net186),
    .A1(_04024_));
 sg13g2_o21ai_1 _11461_ (.B1(_04026_),
    .Y(_04027_),
    .A1(_01998_),
    .A2(_04023_));
 sg13g2_a21o_1 _11462_ (.A2(_04021_),
    .A1(_03097_),
    .B1(_04027_),
    .X(_04028_));
 sg13g2_or4_1 _11463_ (.A(_04017_),
    .B(_04018_),
    .C(_04020_),
    .D(_04028_),
    .X(_04029_));
 sg13g2_o21ai_1 _11464_ (.B1(net165),
    .Y(_04030_),
    .A1(_03452_),
    .A2(_03456_));
 sg13g2_a21oi_1 _11465_ (.A1(net184),
    .A2(_02960_),
    .Y(_04031_),
    .B1(_03772_));
 sg13g2_a21o_1 _11466_ (.A2(_02925_),
    .A1(_01771_),
    .B1(_02922_),
    .X(_04032_));
 sg13g2_o21ai_1 _11467_ (.B1(_04032_),
    .Y(_04033_),
    .A1(_03616_),
    .A2(_04031_));
 sg13g2_buf_1 _11468_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[8] ),
    .X(_04034_));
 sg13g2_mux2_1 _11469_ (.A0(_02960_),
    .A1(_04034_),
    .S(_03873_),
    .X(_04035_));
 sg13g2_nand2_1 _11470_ (.Y(_04036_),
    .A(_01766_),
    .B(_04035_));
 sg13g2_and3_1 _11471_ (.X(_04037_),
    .A(net597),
    .B(_04033_),
    .C(_04036_));
 sg13g2_o21ai_1 _11472_ (.B1(_04037_),
    .Y(_04038_),
    .A1(_03448_),
    .A2(_04030_));
 sg13g2_mux2_1 _11473_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[10] ),
    .S(_01793_),
    .X(_04039_));
 sg13g2_mux2_1 _11474_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[8] ),
    .S(_01793_),
    .X(_04040_));
 sg13g2_or3_1 _11475_ (.A(net522),
    .B(_04039_),
    .C(_04040_),
    .X(_04041_));
 sg13g2_o21ai_1 _11476_ (.B1(_04041_),
    .Y(_04042_),
    .A1(_04029_),
    .A2(_04038_));
 sg13g2_nand3b_1 _11477_ (.B(_04042_),
    .C(_03584_),
    .Y(_04043_),
    .A_N(_04014_));
 sg13g2_a22oi_1 _11478_ (.Y(_04044_),
    .B1(_03997_),
    .B2(_04043_),
    .A2(_03994_),
    .A1(_03990_));
 sg13g2_nand3_1 _11479_ (.B(_03962_),
    .C(_04044_),
    .A(_03921_),
    .Y(_04045_));
 sg13g2_nor3_1 _11480_ (.A(_03807_),
    .B(_03855_),
    .C(_04045_),
    .Y(_04046_));
 sg13g2_xnor2_1 _11481_ (.Y(_04047_),
    .A(_03000_),
    .B(_03036_));
 sg13g2_mux2_1 _11482_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[24] ),
    .S(net595),
    .X(_04048_));
 sg13g2_buf_1 _11483_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[24] ),
    .X(_04049_));
 sg13g2_o21ai_1 _11484_ (.B1(net415),
    .Y(_04050_),
    .A1(net182),
    .A2(net306));
 sg13g2_a22oi_1 _11485_ (.Y(_04051_),
    .B1(_02497_),
    .B2(_04050_),
    .A2(net176),
    .A1(_04049_));
 sg13g2_nor3_1 _11486_ (.A(net263),
    .B(net310),
    .C(_02501_),
    .Y(_04052_));
 sg13g2_a21oi_1 _11487_ (.A1(net184),
    .A2(_02497_),
    .Y(_04053_),
    .B1(net182));
 sg13g2_o21ai_1 _11488_ (.B1(_02493_),
    .Y(_04054_),
    .A1(_04052_),
    .A2(_04053_));
 sg13g2_and2_1 _11489_ (.A(_04051_),
    .B(_04054_),
    .X(_04055_));
 sg13g2_nand2_1 _11490_ (.Y(_04056_),
    .A(net522),
    .B(_04055_));
 sg13g2_o21ai_1 _11491_ (.B1(_04056_),
    .Y(_04057_),
    .A1(net522),
    .A2(_04048_));
 sg13g2_inv_1 _11492_ (.Y(_04058_),
    .A(_04057_));
 sg13g2_a21oi_1 _11493_ (.A1(net164),
    .A2(_04047_),
    .Y(_04059_),
    .B1(_04058_));
 sg13g2_buf_2 _11494_ (.A(_04059_),
    .X(_04060_));
 sg13g2_nand3_1 _11495_ (.B(net141),
    .C(_03151_),
    .A(net165),
    .Y(_04061_));
 sg13g2_nor2_1 _11496_ (.A(net181),
    .B(_03151_),
    .Y(_04062_));
 sg13g2_nand2_1 _11497_ (.Y(_04063_),
    .A(_03637_),
    .B(_04062_));
 sg13g2_mux2_1 _11498_ (.A0(_04061_),
    .A1(_04063_),
    .S(_03150_),
    .X(_04064_));
 sg13g2_nand2_1 _11499_ (.Y(_04065_),
    .A(net184),
    .B(_02062_));
 sg13g2_mux2_1 _11500_ (.A0(net310),
    .A1(net174),
    .S(_04065_),
    .X(_04066_));
 sg13g2_buf_1 _11501_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[22] ),
    .X(_04067_));
 sg13g2_o21ai_1 _11502_ (.B1(net362),
    .Y(_04068_),
    .A1(net173),
    .A2(_02070_));
 sg13g2_a22oi_1 _11503_ (.Y(_04069_),
    .B1(_02062_),
    .B2(_04068_),
    .A2(net176),
    .A1(_04067_));
 sg13g2_o21ai_1 _11504_ (.B1(_04069_),
    .Y(_04070_),
    .A1(_02090_),
    .A2(_04066_));
 sg13g2_and4_1 _11505_ (.A(net175),
    .B(net141),
    .C(_03151_),
    .D(_03128_),
    .X(_04071_));
 sg13g2_nor2b_1 _11506_ (.A(net141),
    .B_N(_04062_),
    .Y(_04072_));
 sg13g2_nor3_1 _11507_ (.A(_04070_),
    .B(_04071_),
    .C(_04072_),
    .Y(_04073_));
 sg13g2_nand3_1 _11508_ (.B(_04064_),
    .C(_04073_),
    .A(net525),
    .Y(_04074_));
 sg13g2_nand2_1 _11509_ (.Y(_04075_),
    .A(net524),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[22] ));
 sg13g2_nand2b_1 _11510_ (.Y(_04076_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[22] ),
    .A_N(net524));
 sg13g2_nand3_1 _11511_ (.B(_04075_),
    .C(_04076_),
    .A(net444),
    .Y(_04077_));
 sg13g2_mux2_1 _11512_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[20] ),
    .S(net595),
    .X(_04078_));
 sg13g2_buf_1 _11513_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[20] ),
    .X(_04079_));
 sg13g2_o21ai_1 _11514_ (.B1(net415),
    .Y(_04080_),
    .A1(net173),
    .A2(_02239_));
 sg13g2_nand3_1 _11515_ (.B(net207),
    .C(_02237_),
    .A(net177),
    .Y(_04081_));
 sg13g2_o21ai_1 _11516_ (.B1(net213),
    .Y(_04082_),
    .A1(net263),
    .A2(_02048_));
 sg13g2_a21oi_1 _11517_ (.A1(_04081_),
    .A2(_04082_),
    .Y(_04083_),
    .B1(_02054_));
 sg13g2_a221oi_1 _11518_ (.B2(_04080_),
    .C1(_04083_),
    .B1(_02237_),
    .A1(_04079_),
    .Y(_04084_),
    .A2(net176));
 sg13g2_nand2_1 _11519_ (.Y(_04085_),
    .A(net522),
    .B(_04084_));
 sg13g2_o21ai_1 _11520_ (.B1(_04085_),
    .Y(_04086_),
    .A1(net525),
    .A2(_04078_));
 sg13g2_nor2_1 _11521_ (.A(_03362_),
    .B(_03727_),
    .Y(_04087_));
 sg13g2_o21ai_1 _11522_ (.B1(_04087_),
    .Y(_04088_),
    .A1(_03353_),
    .A2(_03360_));
 sg13g2_nand2_1 _11523_ (.Y(_04089_),
    .A(_03362_),
    .B(net164));
 sg13g2_or3_1 _11524_ (.A(_03353_),
    .B(_03360_),
    .C(_04089_),
    .X(_04090_));
 sg13g2_nand3_1 _11525_ (.B(_04088_),
    .C(_04090_),
    .A(_04086_),
    .Y(_04091_));
 sg13g2_buf_1 _11526_ (.A(_04091_),
    .X(_04092_));
 sg13g2_a221oi_1 _11527_ (.B2(_04077_),
    .C1(_04092_),
    .B1(_04074_),
    .A1(_03581_),
    .Y(_04093_),
    .A2(net521));
 sg13g2_nor4_1 _11528_ (.A(_02049_),
    .B(_02064_),
    .C(_02489_),
    .D(net414),
    .Y(_04094_));
 sg13g2_a21o_1 _11529_ (.A2(_04093_),
    .A1(_04060_),
    .B1(_04094_),
    .X(_04095_));
 sg13g2_buf_1 _11530_ (.A(_04095_),
    .X(_04096_));
 sg13g2_and4_1 _11531_ (.A(_03673_),
    .B(_03788_),
    .C(_04046_),
    .D(_04096_),
    .X(_04097_));
 sg13g2_nand2_1 _11532_ (.Y(_04098_),
    .A(_03573_),
    .B(_04097_));
 sg13g2_inv_1 _11533_ (.Y(_04099_),
    .A(_03835_));
 sg13g2_buf_1 _11534_ (.A(\soc_I.spi_div_ready ),
    .X(_04100_));
 sg13g2_nor3_1 _11535_ (.A(\soc_I.spi0_I.ready_ctrl ),
    .B(\soc_I.spi0_I.ready_xfer ),
    .C(net618),
    .Y(_04101_));
 sg13g2_buf_1 _11536_ (.A(\soc_I.div_ready ),
    .X(_04102_));
 sg13g2_buf_1 _11537_ (.A(\soc_I.uart_tx_ready ),
    .X(_04103_));
 sg13g2_inv_1 _11538_ (.Y(_04104_),
    .A(_04103_));
 sg13g2_buf_1 _11539_ (.A(\soc_I.rx_uart_i.data_rd ),
    .X(_04105_));
 sg13g2_inv_1 _11540_ (.Y(_04106_),
    .A(_04105_));
 sg13g2_nand2_1 _11541_ (.Y(_04107_),
    .A(net594),
    .B(_04106_));
 sg13g2_nor3_1 _11542_ (.A(_04102_),
    .B(\soc_I.cycle_cnt_ready ),
    .C(_04107_),
    .Y(_04108_));
 sg13g2_nand3_1 _11543_ (.B(_04101_),
    .C(_04108_),
    .A(_00049_),
    .Y(_04109_));
 sg13g2_buf_1 _11544_ (.A(_04109_),
    .X(_04110_));
 sg13g2_inv_1 _11545_ (.Y(_04111_),
    .A(_04110_));
 sg13g2_and3_1 _11546_ (.X(_04112_),
    .A(_03573_),
    .B(_04099_),
    .C(_04111_));
 sg13g2_or2_1 _11547_ (.X(_04113_),
    .B(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[13] ),
    .A(net446));
 sg13g2_buf_1 _11548_ (.A(_04113_),
    .X(_04114_));
 sg13g2_nor3_1 _11549_ (.A(net447),
    .B(net414),
    .C(_04114_),
    .Y(_04115_));
 sg13g2_buf_2 _11550_ (.A(_04115_),
    .X(_04116_));
 sg13g2_nand2_1 _11551_ (.Y(_04117_),
    .A(_03551_),
    .B(_03560_));
 sg13g2_a21oi_1 _11552_ (.A1(_03531_),
    .A2(_03533_),
    .Y(_04118_),
    .B1(_04117_));
 sg13g2_nand2_1 _11553_ (.Y(_04119_),
    .A(_03735_),
    .B(_03736_));
 sg13g2_and3_1 _11554_ (.X(_04120_),
    .A(_03743_),
    .B(_04119_),
    .C(_03734_));
 sg13g2_nand2_1 _11555_ (.Y(_04121_),
    .A(_04033_),
    .B(_04036_));
 sg13g2_a21oi_2 _11556_ (.B1(_04121_),
    .Y(_04122_),
    .A2(_03458_),
    .A1(net159));
 sg13g2_nor4_2 _11557_ (.A(_04017_),
    .B(_04018_),
    .C(_04020_),
    .Y(_04123_),
    .D(_04028_));
 sg13g2_and2_1 _11558_ (.A(_04122_),
    .B(_04123_),
    .X(_04124_));
 sg13g2_a21o_1 _11559_ (.A2(_03378_),
    .A1(net159),
    .B1(_03912_),
    .X(_04125_));
 sg13g2_nand4_1 _11560_ (.B(_03899_),
    .C(_03801_),
    .A(_01791_),
    .Y(_04126_),
    .D(_03845_));
 sg13g2_nor3_1 _11561_ (.A(_03827_),
    .B(_04125_),
    .C(_04126_),
    .Y(_04127_));
 sg13g2_and4_1 _11562_ (.A(_04120_),
    .B(_04124_),
    .C(_03954_),
    .D(_04127_),
    .X(_04128_));
 sg13g2_o21ai_1 _11563_ (.B1(net159),
    .Y(_04129_),
    .A1(_03318_),
    .A2(_03321_));
 sg13g2_and2_1 _11564_ (.A(_03396_),
    .B(_03778_),
    .X(_04130_));
 sg13g2_nand4_1 _11565_ (.B(_03766_),
    .C(_03769_),
    .A(_03398_),
    .Y(_04131_),
    .D(_04130_));
 sg13g2_nand2_1 _11566_ (.Y(_04132_),
    .A(net172),
    .B(_03778_));
 sg13g2_a21oi_1 _11567_ (.A1(_04131_),
    .A2(_04132_),
    .Y(_04133_),
    .B1(_03645_));
 sg13g2_nand4_1 _11568_ (.B(_04128_),
    .C(_04129_),
    .A(_03721_),
    .Y(_04134_),
    .D(_04133_));
 sg13g2_nand3_1 _11569_ (.B(_03684_),
    .C(_03691_),
    .A(_03681_),
    .Y(_04135_));
 sg13g2_o21ai_1 _11570_ (.B1(_04084_),
    .Y(_04136_),
    .A1(net172),
    .A2(_03363_));
 sg13g2_xor2_1 _11571_ (.B(_03389_),
    .A(_03735_),
    .X(_04137_));
 sg13g2_inv_1 _11572_ (.Y(_04138_),
    .A(_04006_));
 sg13g2_a21oi_1 _11573_ (.A1(_03546_),
    .A2(_04137_),
    .Y(_04139_),
    .B1(_04138_));
 sg13g2_and2_1 _11574_ (.A(_03384_),
    .B(_03866_),
    .X(_04140_));
 sg13g2_a21o_1 _11575_ (.A2(_03858_),
    .A1(_03857_),
    .B1(_03860_),
    .X(_04141_));
 sg13g2_o21ai_1 _11576_ (.B1(net165),
    .Y(_04142_),
    .A1(_03384_),
    .A2(_04141_));
 sg13g2_a21oi_1 _11577_ (.A1(_03545_),
    .A2(_03882_),
    .Y(_04143_),
    .B1(_03876_));
 sg13g2_o21ai_1 _11578_ (.B1(_04143_),
    .Y(_04144_),
    .A1(_04140_),
    .A2(_04142_));
 sg13g2_nor4_2 _11579_ (.A(net172),
    .B(_03241_),
    .C(_03242_),
    .Y(_04145_),
    .D(_03245_));
 sg13g2_nor3_1 _11580_ (.A(_04144_),
    .B(_03928_),
    .C(_04145_),
    .Y(_04146_));
 sg13g2_nand4_1 _11581_ (.B(_03600_),
    .C(_04139_),
    .A(_03592_),
    .Y(_04147_),
    .D(_04146_));
 sg13g2_or3_1 _11582_ (.A(_03344_),
    .B(_03326_),
    .C(_03699_),
    .X(_04148_));
 sg13g2_nand3_1 _11583_ (.B(_04148_),
    .C(_03698_),
    .A(_03706_),
    .Y(_04149_));
 sg13g2_nand2_1 _11584_ (.Y(_04150_),
    .A(_03988_),
    .B(_03981_));
 sg13g2_or3_1 _11585_ (.A(_04149_),
    .B(_03976_),
    .C(_04150_),
    .X(_04151_));
 sg13g2_or4_1 _11586_ (.A(_04135_),
    .B(_04136_),
    .C(_04147_),
    .D(_04151_),
    .X(_04152_));
 sg13g2_nor4_1 _11587_ (.A(net172),
    .B(_03219_),
    .C(_03222_),
    .D(_03230_),
    .Y(_04153_));
 sg13g2_and2_1 _11588_ (.A(net175),
    .B(_03219_),
    .X(_04154_));
 sg13g2_mux2_1 _11589_ (.A0(_04153_),
    .A1(_04154_),
    .S(_03237_),
    .X(_04155_));
 sg13g2_a21oi_1 _11590_ (.A1(net213),
    .A2(net211),
    .Y(_04156_),
    .B1(_03616_));
 sg13g2_buf_1 _11591_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[27] ),
    .X(_04157_));
 sg13g2_nand2_1 _11592_ (.Y(_04158_),
    .A(_04157_),
    .B(net166));
 sg13g2_o21ai_1 _11593_ (.B1(_04158_),
    .Y(_04159_),
    .A1(_02542_),
    .A2(_04156_));
 sg13g2_nand3_1 _11594_ (.B(net207),
    .C(_02589_),
    .A(net167),
    .Y(_04160_));
 sg13g2_o21ai_1 _11595_ (.B1(net213),
    .Y(_04161_),
    .A1(net263),
    .A2(_02542_));
 sg13g2_a21oi_1 _11596_ (.A1(_04160_),
    .A2(_04161_),
    .Y(_04162_),
    .B1(_02591_));
 sg13g2_nor2_1 _11597_ (.A(net172),
    .B(_03494_),
    .Y(_04163_));
 sg13g2_nor4_2 _11598_ (.A(_04155_),
    .B(_04159_),
    .C(_04162_),
    .Y(_04164_),
    .D(_04163_));
 sg13g2_mux2_1 _11599_ (.A0(_03682_),
    .A1(_03683_),
    .S(_03121_),
    .X(_04165_));
 sg13g2_buf_1 _11600_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[26] ),
    .X(_04166_));
 sg13g2_o21ai_1 _11601_ (.B1(net362),
    .Y(_04167_),
    .A1(net174),
    .A2(_02555_));
 sg13g2_nand3_1 _11602_ (.B(net207),
    .C(net264),
    .A(net167),
    .Y(_04168_));
 sg13g2_o21ai_1 _11603_ (.B1(net213),
    .Y(_04169_),
    .A1(net263),
    .A2(_02606_));
 sg13g2_a21oi_1 _11604_ (.A1(_04168_),
    .A2(_04169_),
    .Y(_04170_),
    .B1(_02604_));
 sg13g2_a221oi_1 _11605_ (.B2(_04167_),
    .C1(_04170_),
    .B1(net264),
    .A1(_04166_),
    .Y(_04171_),
    .A2(net166));
 sg13g2_nand3_1 _11606_ (.B(_04165_),
    .C(_04171_),
    .A(_04164_),
    .Y(_04172_));
 sg13g2_a21o_1 _11607_ (.A2(_03524_),
    .A1(_03521_),
    .B1(_03944_),
    .X(_04173_));
 sg13g2_inv_1 _11608_ (.Y(_04174_),
    .A(_03663_));
 sg13g2_a21oi_1 _11609_ (.A1(_03546_),
    .A2(_03216_),
    .Y(_04175_),
    .B1(_04174_));
 sg13g2_nand3_1 _11610_ (.B(_04173_),
    .C(_04175_),
    .A(_03761_),
    .Y(_04176_));
 sg13g2_xnor2_1 _11611_ (.Y(_04177_),
    .A(net142),
    .B(_03036_));
 sg13g2_o21ai_1 _11612_ (.B1(_04055_),
    .Y(_04178_),
    .A1(_03944_),
    .A2(_04177_));
 sg13g2_nand2_1 _11613_ (.Y(_04179_),
    .A(_04064_),
    .B(_04073_));
 sg13g2_nand3_1 _11614_ (.B(_02986_),
    .C(_02988_),
    .A(net159),
    .Y(_04180_));
 sg13g2_or4_1 _11615_ (.A(net172),
    .B(_02827_),
    .C(_02986_),
    .D(_02988_),
    .X(_04181_));
 sg13g2_nand3_1 _11616_ (.B(_02827_),
    .C(_02988_),
    .A(net159),
    .Y(_04182_));
 sg13g2_nand4_1 _11617_ (.B(_04180_),
    .C(_04181_),
    .A(_03620_),
    .Y(_04183_),
    .D(_04182_));
 sg13g2_or2_1 _11618_ (.X(_04184_),
    .B(_04183_),
    .A(_04179_));
 sg13g2_or4_1 _11619_ (.A(_04172_),
    .B(_04176_),
    .C(_04178_),
    .D(_04184_),
    .X(_04185_));
 sg13g2_nor4_1 _11620_ (.A(_01594_),
    .B(_04134_),
    .C(_04152_),
    .D(_04185_),
    .Y(_04186_));
 sg13g2_nand3b_1 _11621_ (.B(_04118_),
    .C(_04186_),
    .Y(_04187_),
    .A_N(_03529_));
 sg13g2_buf_2 _11622_ (.A(_04187_),
    .X(_04188_));
 sg13g2_nor2b_1 _11623_ (.A(_03807_),
    .B_N(_03962_),
    .Y(_04189_));
 sg13g2_nor2_2 _11624_ (.A(\soc_I.spi0_I.ready_ctrl ),
    .B(\soc_I.spi0_I.ready_xfer ),
    .Y(_04190_));
 sg13g2_nand2_1 _11625_ (.Y(_04191_),
    .A(net447),
    .B(net414));
 sg13g2_nor2_1 _11626_ (.A(\soc_I.kianv_I.datapath_unit_I.DataLatched[26] ),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[27] ),
    .Y(_04192_));
 sg13g2_nor3_1 _11627_ (.A(net446),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[26] ),
    .C(\soc_I.kianv_I.datapath_unit_I.ALUOut[27] ),
    .Y(_04193_));
 sg13g2_a21oi_1 _11628_ (.A1(net446),
    .A2(_04192_),
    .Y(_04194_),
    .B1(_04193_));
 sg13g2_nor3_1 _11629_ (.A(net525),
    .B(_01559_),
    .C(_04194_),
    .Y(_04195_));
 sg13g2_nor3_1 _11630_ (.A(_02551_),
    .B(_02544_),
    .C(net445),
    .Y(_04196_));
 sg13g2_nor2_1 _11631_ (.A(_04195_),
    .B(_04196_),
    .Y(_04197_));
 sg13g2_o21ai_1 _11632_ (.B1(_04197_),
    .Y(_04198_),
    .A1(_04191_),
    .A2(_04172_));
 sg13g2_buf_2 _11633_ (.A(_04198_),
    .X(_04199_));
 sg13g2_nand2_1 _11634_ (.Y(_04200_),
    .A(_03990_),
    .B(_03994_));
 sg13g2_nand2_1 _11635_ (.Y(_04201_),
    .A(_03997_),
    .B(_04043_));
 sg13g2_and3_1 _11636_ (.X(_04202_),
    .A(_04200_),
    .B(_03921_),
    .C(_04201_));
 sg13g2_o21ai_1 _11637_ (.B1(_04057_),
    .Y(_04203_),
    .A1(_03727_),
    .A2(_04177_));
 sg13g2_or2_1 _11638_ (.X(_04204_),
    .B(_03670_),
    .A(_02489_));
 sg13g2_o21ai_1 _11639_ (.B1(_04204_),
    .Y(_04205_),
    .A1(_03669_),
    .A2(_04203_));
 sg13g2_nand2_1 _11640_ (.Y(_04206_),
    .A(_04074_),
    .B(_04077_));
 sg13g2_buf_1 _11641_ (.A(_04206_),
    .X(_04207_));
 sg13g2_nand2_1 _11642_ (.Y(_04208_),
    .A(net414),
    .B(_04092_));
 sg13g2_nand3_1 _11643_ (.B(_02064_),
    .C(net457),
    .A(_02049_),
    .Y(_04209_));
 sg13g2_o21ai_1 _11644_ (.B1(_04209_),
    .Y(_04210_),
    .A1(net112),
    .A2(_04208_));
 sg13g2_and4_1 _11645_ (.A(_04199_),
    .B(_04202_),
    .C(_04205_),
    .D(_04210_),
    .X(_04211_));
 sg13g2_nand4_1 _11646_ (.B(_04189_),
    .C(_04190_),
    .A(_03788_),
    .Y(_04212_),
    .D(_04211_));
 sg13g2_a21oi_2 _11647_ (.B1(_04212_),
    .Y(_04213_),
    .A2(_04188_),
    .A1(_04116_));
 sg13g2_nor2b_1 _11648_ (.A(_03753_),
    .B_N(_03763_),
    .Y(_04214_));
 sg13g2_buf_1 _11649_ (.A(_04214_),
    .X(_04215_));
 sg13g2_nor2_1 _11650_ (.A(_02514_),
    .B(net414),
    .Y(_04216_));
 sg13g2_a21oi_1 _11651_ (.A1(net414),
    .A2(net88),
    .Y(_04217_),
    .B1(_04216_));
 sg13g2_a21o_1 _11652_ (.A2(_03654_),
    .A1(_03652_),
    .B1(_04217_),
    .X(_04218_));
 sg13g2_nand2_1 _11653_ (.Y(_04219_),
    .A(_04199_),
    .B(_04218_));
 sg13g2_a221oi_1 _11654_ (.B2(_04213_),
    .C1(_04219_),
    .B1(_04112_),
    .A1(_03672_),
    .Y(_04220_),
    .A2(_04098_));
 sg13g2_buf_1 _11655_ (.A(_04220_),
    .X(_04221_));
 sg13g2_nand3_1 _11656_ (.B(_03671_),
    .C(_04096_),
    .A(_04199_),
    .Y(_04222_));
 sg13g2_buf_2 _11657_ (.A(_04222_),
    .X(_04223_));
 sg13g2_nor2_1 _11658_ (.A(_04110_),
    .B(_04223_),
    .Y(_04224_));
 sg13g2_buf_1 _11659_ (.A(_01557_),
    .X(_04225_));
 sg13g2_buf_2 _11660_ (.A(\soc_I.uart_lsr_rdy ),
    .X(_04226_));
 sg13g2_nor4_1 _11661_ (.A(net593),
    .B(_04226_),
    .C(_03835_),
    .D(_03854_),
    .Y(_04227_));
 sg13g2_and3_1 _11662_ (.X(_04228_),
    .A(_04202_),
    .B(_04189_),
    .C(_04227_));
 sg13g2_a21oi_1 _11663_ (.A1(_04224_),
    .A2(_04228_),
    .Y(_04229_),
    .B1(net76));
 sg13g2_a21oi_1 _11664_ (.A1(_03752_),
    .A2(_03751_),
    .Y(_04230_),
    .B1(_03786_));
 sg13g2_nand2_1 _11665_ (.Y(_04231_),
    .A(_03655_),
    .B(_04230_));
 sg13g2_a21oi_1 _11666_ (.A1(_04116_),
    .A2(_04188_),
    .Y(_04232_),
    .B1(_04231_));
 sg13g2_and3_1 _11667_ (.X(_04233_),
    .A(_04199_),
    .B(_03671_),
    .C(_04096_));
 sg13g2_buf_1 _11668_ (.A(_04233_),
    .X(_04234_));
 sg13g2_nand3_1 _11669_ (.B(_04111_),
    .C(_04234_),
    .A(_04046_),
    .Y(_04235_));
 sg13g2_nand2_1 _11670_ (.Y(_04236_),
    .A(net76),
    .B(_04235_));
 sg13g2_nand3b_1 _11671_ (.B(_04232_),
    .C(_04236_),
    .Y(_04237_),
    .A_N(_04229_));
 sg13g2_buf_1 _11672_ (.A(_04237_),
    .X(_04238_));
 sg13g2_nand4_1 _11673_ (.B(_03807_),
    .C(_03962_),
    .A(_03921_),
    .Y(_04239_),
    .D(_04044_));
 sg13g2_buf_1 _11674_ (.A(_04239_),
    .X(_04240_));
 sg13g2_nor2_1 _11675_ (.A(\soc_I.cpu_mem_addr[1] ),
    .B(_04240_),
    .Y(_04241_));
 sg13g2_nand3_1 _11676_ (.B(_04234_),
    .C(_04241_),
    .A(_03788_),
    .Y(_04242_));
 sg13g2_a21oi_1 _11677_ (.A1(_04116_),
    .A2(_04188_),
    .Y(_04243_),
    .B1(_04242_));
 sg13g2_nand2_1 _11678_ (.Y(_04244_),
    .A(_02282_),
    .B(net457));
 sg13g2_o21ai_1 _11679_ (.B1(_04244_),
    .Y(_04245_),
    .A1(_01560_),
    .A2(_03832_));
 sg13g2_nand3b_1 _11680_ (.B(_03854_),
    .C(_04245_),
    .Y(_04246_),
    .A_N(\soc_I.cycle_cnt_ready ));
 sg13g2_or3_1 _11681_ (.A(\soc_I.pwm_ready ),
    .B(_03854_),
    .C(_04245_),
    .X(_04247_));
 sg13g2_a21oi_1 _11682_ (.A1(_04246_),
    .A2(_04247_),
    .Y(_04248_),
    .B1(_04110_));
 sg13g2_and2_1 _11683_ (.A(_03573_),
    .B(_04248_),
    .X(_04249_));
 sg13g2_inv_1 _11684_ (.Y(_04250_),
    .A(_04100_));
 sg13g2_nand4_1 _11685_ (.B(_04199_),
    .C(_04205_),
    .A(_04250_),
    .Y(_04251_),
    .D(_04210_));
 sg13g2_o21ai_1 _11686_ (.B1(_04251_),
    .Y(_04252_),
    .A1(_04102_),
    .A2(_04223_));
 sg13g2_nor3_1 _11687_ (.A(_03855_),
    .B(_04110_),
    .C(_04240_),
    .Y(_04253_));
 sg13g2_and3_1 _11688_ (.X(_04254_),
    .A(_03574_),
    .B(_04252_),
    .C(_04253_));
 sg13g2_a22oi_1 _11689_ (.Y(_04255_),
    .B1(_04254_),
    .B2(_04232_),
    .A2(_04249_),
    .A1(_04243_));
 sg13g2_buf_1 _11690_ (.A(_04255_),
    .X(_04256_));
 sg13g2_nand3_1 _11691_ (.B(_04238_),
    .C(_04256_),
    .A(_04221_),
    .Y(_04257_));
 sg13g2_buf_1 _11692_ (.A(net444),
    .X(_04258_));
 sg13g2_a21oi_1 _11693_ (.A1(_00048_),
    .A2(_04257_),
    .Y(_04259_),
    .B1(_04258_));
 sg13g2_buf_2 _11694_ (.A(_04259_),
    .X(_04260_));
 sg13g2_nand2_1 _11695_ (.Y(_04261_),
    .A(_00053_),
    .B(_03536_));
 sg13g2_o21ai_1 _11696_ (.B1(_04261_),
    .Y(_04262_),
    .A1(_03580_),
    .A2(_04260_));
 sg13g2_buf_2 _11697_ (.A(_04262_),
    .X(_04263_));
 sg13g2_buf_8 _11698_ (.A(_04263_),
    .X(_04264_));
 sg13g2_nor4_1 _11699_ (.A(net455),
    .B(_01842_),
    .C(_03579_),
    .D(net27),
    .Y(_00012_));
 sg13g2_inv_1 _11700_ (.Y(_04265_),
    .A(_03576_));
 sg13g2_buf_1 _11701_ (.A(_04265_),
    .X(_04266_));
 sg13g2_buf_2 _11702_ (.A(net520),
    .X(_04267_));
 sg13g2_nor2_1 _11703_ (.A(net413),
    .B(_04267_),
    .Y(_04268_));
 sg13g2_inv_1 _11704_ (.Y(_04269_),
    .A(_00048_));
 sg13g2_and3_1 _11705_ (.X(_04270_),
    .A(_04221_),
    .B(_04238_),
    .C(_04256_));
 sg13g2_buf_2 _11706_ (.A(_04270_),
    .X(_04271_));
 sg13g2_nor2_2 _11707_ (.A(_04269_),
    .B(_04271_),
    .Y(_04272_));
 sg13g2_buf_1 _11708_ (.A(_00057_),
    .X(_04273_));
 sg13g2_nor2b_1 _11709_ (.A(net616),
    .B_N(_01576_),
    .Y(_04274_));
 sg13g2_and2_1 _11710_ (.A(\soc_I.kianv_I.Instr[0] ),
    .B(\soc_I.kianv_I.Instr[1] ),
    .X(_04275_));
 sg13g2_o21ai_1 _11711_ (.B1(_03575_),
    .Y(_04276_),
    .A1(net628),
    .A2(_02420_));
 sg13g2_and2_1 _11712_ (.A(net600),
    .B(net601),
    .X(_04277_));
 sg13g2_a22oi_1 _11713_ (.Y(_04278_),
    .B1(_04276_),
    .B2(_04277_),
    .A2(_01689_),
    .A1(_01642_));
 sg13g2_nand3_1 _11714_ (.B(_01655_),
    .C(_04278_),
    .A(_04275_),
    .Y(_04279_));
 sg13g2_a21o_1 _11715_ (.A2(_04279_),
    .A1(_04274_),
    .B1(_01562_),
    .X(_04280_));
 sg13g2_a21oi_1 _11716_ (.A1(_01648_),
    .A2(_04280_),
    .Y(_04281_),
    .B1(_01561_));
 sg13g2_a21oi_1 _11717_ (.A1(_00053_),
    .A2(net166),
    .Y(_04282_),
    .B1(_04281_));
 sg13g2_nor3_1 _11718_ (.A(net616),
    .B(_04114_),
    .C(_04282_),
    .Y(_04283_));
 sg13g2_o21ai_1 _11719_ (.B1(_04283_),
    .Y(_04284_),
    .A1(net521),
    .A2(_04272_));
 sg13g2_a21o_1 _11720_ (.A2(_04268_),
    .A1(_04264_),
    .B1(_04284_),
    .X(_00007_));
 sg13g2_inv_1 _11721_ (.Y(_04285_),
    .A(_04273_));
 sg13g2_nand2_1 _11722_ (.Y(_04286_),
    .A(net632),
    .B(net592));
 sg13g2_or3_1 _11723_ (.A(net628),
    .B(_01692_),
    .C(_04286_),
    .X(_04287_));
 sg13g2_buf_1 _11724_ (.A(_04287_),
    .X(_04288_));
 sg13g2_nor2_1 _11725_ (.A(_01811_),
    .B(_04288_),
    .Y(_04289_));
 sg13g2_and2_1 _11726_ (.A(_01565_),
    .B(net523),
    .X(_04290_));
 sg13g2_mux2_1 _11727_ (.A0(_04289_),
    .A1(_04290_),
    .S(net27),
    .X(_00011_));
 sg13g2_buf_1 _11728_ (.A(\soc_I.qqspi_I.xfer_cycles[0] ),
    .X(_04291_));
 sg13g2_nor2_1 _11729_ (.A(_04291_),
    .B(\soc_I.qqspi_I.xfer_cycles[1] ),
    .Y(_04292_));
 sg13g2_buf_1 _11730_ (.A(\soc_I.qqspi_I.xfer_cycles[3] ),
    .X(_04293_));
 sg13g2_buf_1 _11731_ (.A(\soc_I.qqspi_I.xfer_cycles[2] ),
    .X(_04294_));
 sg13g2_nor4_1 _11732_ (.A(_04293_),
    .B(_04294_),
    .C(\soc_I.qqspi_I.xfer_cycles[5] ),
    .D(\soc_I.qqspi_I.xfer_cycles[4] ),
    .Y(_04295_));
 sg13g2_and2_1 _11733_ (.A(_04292_),
    .B(_04295_),
    .X(_04296_));
 sg13g2_buf_1 _11734_ (.A(_04296_),
    .X(_04297_));
 sg13g2_buf_1 _11735_ (.A(net443),
    .X(_04298_));
 sg13g2_buf_1 _11736_ (.A(net412),
    .X(_04299_));
 sg13g2_buf_1 _11737_ (.A(net361),
    .X(_04300_));
 sg13g2_nand2_1 _11738_ (.Y(_04301_),
    .A(\soc_I.qqspi_I.state[3] ),
    .B(net592));
 sg13g2_buf_2 _11739_ (.A(\soc_I.qqspi_I.state[5] ),
    .X(_04302_));
 sg13g2_buf_1 _11740_ (.A(_04302_),
    .X(_04303_));
 sg13g2_buf_1 _11741_ (.A(net591),
    .X(_04304_));
 sg13g2_buf_1 _11742_ (.A(net596),
    .X(_04305_));
 sg13g2_nand3_1 _11743_ (.B(net518),
    .C(net336),
    .A(net519),
    .Y(_04306_));
 sg13g2_o21ai_1 _11744_ (.B1(_04306_),
    .Y(_00021_),
    .A1(net336),
    .A2(_04301_));
 sg13g2_buf_1 _11745_ (.A(\soc_I.qqspi_I.state[4] ),
    .X(_04307_));
 sg13g2_buf_1 _11746_ (.A(_04292_),
    .X(_04308_));
 sg13g2_buf_1 _11747_ (.A(_04295_),
    .X(_04309_));
 sg13g2_nand2_1 _11748_ (.Y(_04310_),
    .A(net517),
    .B(net516));
 sg13g2_buf_1 _11749_ (.A(_04310_),
    .X(_04311_));
 sg13g2_buf_1 _11750_ (.A(_04311_),
    .X(_04312_));
 sg13g2_buf_1 _11751_ (.A(net360),
    .X(_04313_));
 sg13g2_nand2_1 _11752_ (.Y(_04314_),
    .A(_04307_),
    .B(net335));
 sg13g2_buf_1 _11753_ (.A(\soc_I.qqspi_I.state[0] ),
    .X(_04315_));
 sg13g2_inv_1 _11754_ (.Y(_04316_),
    .A(_04315_));
 sg13g2_and2_1 _11755_ (.A(_04116_),
    .B(_04188_),
    .X(_04317_));
 sg13g2_buf_1 _11756_ (.A(_04317_),
    .X(_04318_));
 sg13g2_and2_1 _11757_ (.A(_04199_),
    .B(_04205_),
    .X(_04319_));
 sg13g2_inv_1 _11758_ (.Y(_04320_),
    .A(_02665_));
 sg13g2_buf_1 _11759_ (.A(_01560_),
    .X(_04321_));
 sg13g2_nand3_1 _11760_ (.B(_04320_),
    .C(net411),
    .A(_03783_),
    .Y(_04322_));
 sg13g2_buf_1 _11761_ (.A(net414),
    .X(_04323_));
 sg13g2_nand3_1 _11762_ (.B(_03650_),
    .C(_04215_),
    .A(net359),
    .Y(_04324_));
 sg13g2_buf_1 _11763_ (.A(\soc_I.qqspi_I.ready ),
    .X(_04325_));
 sg13g2_a21oi_1 _11764_ (.A1(_04322_),
    .A2(_04324_),
    .Y(_04326_),
    .B1(net615));
 sg13g2_nand2_2 _11765_ (.Y(_04327_),
    .A(_04319_),
    .B(_04326_));
 sg13g2_inv_1 _11766_ (.Y(_04328_),
    .A(_02527_));
 sg13g2_nand3_1 _11767_ (.B(_02658_),
    .C(net411),
    .A(_04328_),
    .Y(_04329_));
 sg13g2_buf_1 _11768_ (.A(_03607_),
    .X(_04330_));
 sg13g2_a21o_1 _11769_ (.A2(net164),
    .A1(_02989_),
    .B1(_03623_),
    .X(_04331_));
 sg13g2_buf_1 _11770_ (.A(_04331_),
    .X(_04332_));
 sg13g2_nand3_1 _11771_ (.B(net111),
    .C(_04332_),
    .A(net359),
    .Y(_04333_));
 sg13g2_nand2_1 _11772_ (.Y(_04334_),
    .A(_02074_),
    .B(net457));
 sg13g2_o21ai_1 _11773_ (.B1(_04334_),
    .Y(_04335_),
    .A1(net411),
    .A2(_03714_));
 sg13g2_a21o_1 _11774_ (.A2(_04333_),
    .A1(_04329_),
    .B1(_04335_),
    .X(_04336_));
 sg13g2_nor3_1 _11775_ (.A(_03581_),
    .B(_04330_),
    .C(_04332_),
    .Y(_04337_));
 sg13g2_nor3_1 _11776_ (.A(_01556_),
    .B(_04328_),
    .C(_02658_),
    .Y(_04338_));
 sg13g2_o21ai_1 _11777_ (.B1(net521),
    .Y(_04339_),
    .A1(_04337_),
    .A2(_04338_));
 sg13g2_a21o_1 _11778_ (.A2(_04339_),
    .A1(_04336_),
    .B1(_04269_),
    .X(_04340_));
 sg13g2_buf_1 _11779_ (.A(_04340_),
    .X(_04341_));
 sg13g2_nor4_1 _11780_ (.A(_04316_),
    .B(_04318_),
    .C(_04327_),
    .D(_04341_),
    .Y(_04342_));
 sg13g2_nand2_1 _11781_ (.Y(_04343_),
    .A(net336),
    .B(_04342_));
 sg13g2_a21oi_1 _11782_ (.A1(_04314_),
    .A2(_04343_),
    .Y(_00022_),
    .B1(net616));
 sg13g2_buf_2 _11783_ (.A(\soc_I.qqspi_I.state[6] ),
    .X(_04344_));
 sg13g2_and3_1 _11784_ (.X(_04345_),
    .A(net593),
    .B(_04344_),
    .C(net361));
 sg13g2_a21oi_1 _11785_ (.A1(_04304_),
    .A2(net335),
    .Y(_04346_),
    .B1(_04345_));
 sg13g2_buf_1 _11786_ (.A(\soc_I.qqspi_I.state[1] ),
    .X(_04347_));
 sg13g2_nand3_1 _11787_ (.B(net518),
    .C(net336),
    .A(_04347_),
    .Y(_04348_));
 sg13g2_o21ai_1 _11788_ (.B1(_04348_),
    .Y(_00023_),
    .A1(net616),
    .A2(_04346_));
 sg13g2_nand2_1 _11789_ (.Y(_04349_),
    .A(_04344_),
    .B(net592));
 sg13g2_buf_1 _11790_ (.A(\soc_I.qqspi_I.state[2] ),
    .X(_04350_));
 sg13g2_nand3_1 _11791_ (.B(_04305_),
    .C(net361),
    .A(_04350_),
    .Y(_04351_));
 sg13g2_o21ai_1 _11792_ (.B1(_04351_),
    .Y(_00024_),
    .A1(_04300_),
    .A2(_04349_));
 sg13g2_nand2_1 _11793_ (.Y(_04352_),
    .A(_04347_),
    .B(net335));
 sg13g2_nand3_1 _11794_ (.B(_04344_),
    .C(net361),
    .A(net521),
    .Y(_04353_));
 sg13g2_a21oi_1 _11795_ (.A1(_04352_),
    .A2(_04353_),
    .Y(_00019_),
    .B1(net616));
 sg13g2_nand2_1 _11796_ (.Y(_04354_),
    .A(_04350_),
    .B(net592));
 sg13g2_nand3_1 _11797_ (.B(_04307_),
    .C(net361),
    .A(net518),
    .Y(_04355_));
 sg13g2_o21ai_1 _11798_ (.B1(_04355_),
    .Y(_00020_),
    .A1(net336),
    .A2(_04354_));
 sg13g2_buf_1 _11799_ (.A(_04318_),
    .X(_04356_));
 sg13g2_buf_1 _11800_ (.A(_04311_),
    .X(_04357_));
 sg13g2_buf_1 _11801_ (.A(net358),
    .X(_04358_));
 sg13g2_nor4_1 _11802_ (.A(_04356_),
    .B(net334),
    .C(_04327_),
    .D(_04341_),
    .Y(_04359_));
 sg13g2_nand3_1 _11803_ (.B(\soc_I.qqspi_I.state[3] ),
    .C(net443),
    .A(_03576_),
    .Y(_04360_));
 sg13g2_buf_1 _11804_ (.A(_04360_),
    .X(_04361_));
 sg13g2_buf_1 _11805_ (.A(_04361_),
    .X(_04362_));
 sg13g2_and2_1 _11806_ (.A(net592),
    .B(_04362_),
    .X(_04363_));
 sg13g2_o21ai_1 _11807_ (.B1(_04363_),
    .Y(_00018_),
    .A1(_04316_),
    .A2(_04359_));
 sg13g2_nor3_1 _11808_ (.A(net455),
    .B(_01689_),
    .C(_04286_),
    .Y(_04364_));
 sg13g2_inv_1 _11809_ (.Y(_04365_),
    .A(_01563_));
 sg13g2_nor2_1 _11810_ (.A(_04365_),
    .B(_04267_),
    .Y(_04366_));
 sg13g2_mux2_1 _11811_ (.A0(_04364_),
    .A1(_04366_),
    .S(net27),
    .X(_00010_));
 sg13g2_nand4_1 _11812_ (.B(_01562_),
    .C(net592),
    .A(_01730_),
    .Y(_04367_),
    .D(_01965_));
 sg13g2_nand3_1 _11813_ (.B(net518),
    .C(_04272_),
    .A(_01556_),
    .Y(_04368_));
 sg13g2_o21ai_1 _11814_ (.B1(_04368_),
    .Y(_00009_),
    .A1(_04264_),
    .A2(_04367_));
 sg13g2_nand4_1 _11815_ (.B(net627),
    .C(_02536_),
    .A(_01730_),
    .Y(_04369_),
    .D(_04274_));
 sg13g2_nor2_1 _11816_ (.A(net27),
    .B(_04369_),
    .Y(_00008_));
 sg13g2_nand4_1 _11817_ (.B(_01562_),
    .C(net592),
    .A(_01650_),
    .Y(_04370_),
    .D(_01965_));
 sg13g2_buf_1 _11818_ (.A(net596),
    .X(_04371_));
 sg13g2_nand3_1 _11819_ (.B(net515),
    .C(_04272_),
    .A(net593),
    .Y(_04372_));
 sg13g2_o21ai_1 _11820_ (.B1(_04372_),
    .Y(_00017_),
    .A1(net27),
    .A2(_04370_));
 sg13g2_nand3_1 _11821_ (.B(net632),
    .C(_04275_),
    .A(_01642_),
    .Y(_04373_));
 sg13g2_o21ai_1 _11822_ (.B1(_04365_),
    .Y(_04374_),
    .A1(_01689_),
    .A2(_04373_));
 sg13g2_and2_1 _11823_ (.A(net592),
    .B(_04374_),
    .X(_04375_));
 sg13g2_and2_1 _11824_ (.A(_01577_),
    .B(net523),
    .X(_04376_));
 sg13g2_mux2_1 _11825_ (.A0(_04375_),
    .A1(_04376_),
    .S(net27),
    .X(_00016_));
 sg13g2_nor2_1 _11826_ (.A(net413),
    .B(net616),
    .Y(_04377_));
 sg13g2_o21ai_1 _11827_ (.B1(net523),
    .Y(_04378_),
    .A1(_01562_),
    .A2(net632));
 sg13g2_inv_1 _11828_ (.Y(_04379_),
    .A(_04378_));
 sg13g2_mux2_1 _11829_ (.A0(_04377_),
    .A1(_04379_),
    .S(_04263_),
    .X(_00015_));
 sg13g2_inv_1 _11830_ (.Y(_04380_),
    .A(_02420_));
 sg13g2_nor4_1 _11831_ (.A(net629),
    .B(_04380_),
    .C(_01651_),
    .D(_04288_),
    .Y(_04381_));
 sg13g2_and2_1 _11832_ (.A(_01564_),
    .B(net523),
    .X(_04382_));
 sg13g2_mux2_1 _11833_ (.A0(_04381_),
    .A1(_04382_),
    .S(_04263_),
    .X(_00014_));
 sg13g2_nor4_1 _11834_ (.A(net627),
    .B(_01669_),
    .C(net27),
    .D(_04288_),
    .Y(_00013_));
 sg13g2_nor3_1 _11835_ (.A(_03581_),
    .B(net616),
    .C(_04272_),
    .Y(_00004_));
 sg13g2_nor3_1 _11836_ (.A(_01577_),
    .B(_01863_),
    .C(_01632_),
    .Y(_04383_));
 sg13g2_nor3_1 _11837_ (.A(net616),
    .B(net27),
    .C(_04383_),
    .Y(_00006_));
 sg13g2_and4_1 _11838_ (.A(_01965_),
    .B(_04261_),
    .C(_04274_),
    .D(_04279_),
    .X(_00005_));
 sg13g2_buf_1 _11839_ (.A(_00052_),
    .X(_04384_));
 sg13g2_nand2b_1 _11840_ (.Y(_04385_),
    .B(_03536_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_ready ));
 sg13g2_buf_1 _11841_ (.A(_04385_),
    .X(_04386_));
 sg13g2_a21o_1 _11842_ (.A2(_04386_),
    .A1(_04384_),
    .B1(_04265_),
    .X(_04387_));
 sg13g2_buf_2 _11843_ (.A(_04387_),
    .X(_04388_));
 sg13g2_buf_1 _11844_ (.A(_04388_),
    .X(_04389_));
 sg13g2_buf_1 _11845_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_state ),
    .X(_04390_));
 sg13g2_inv_2 _11846_ (.Y(_04391_),
    .A(_04390_));
 sg13g2_nand2_1 _11847_ (.Y(_04392_),
    .A(net325),
    .B(_01734_));
 sg13g2_buf_1 _11848_ (.A(_04392_),
    .X(_04393_));
 sg13g2_buf_1 _11849_ (.A(_04393_),
    .X(_04394_));
 sg13g2_buf_1 _11850_ (.A(_04390_),
    .X(_04395_));
 sg13g2_and2_1 _11851_ (.A(_01777_),
    .B(net590),
    .X(_04396_));
 sg13g2_a22oi_1 _11852_ (.Y(_04397_),
    .B1(_04394_),
    .B2(_04396_),
    .A2(_01715_),
    .A1(_04391_));
 sg13g2_buf_1 _11853_ (.A(_04388_),
    .X(_04398_));
 sg13g2_nand2_1 _11854_ (.Y(_04399_),
    .A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[0] ),
    .B(_04398_));
 sg13g2_o21ai_1 _11855_ (.B1(_04399_),
    .Y(_00361_),
    .A1(net138),
    .A2(_04397_));
 sg13g2_buf_1 _11856_ (.A(_04395_),
    .X(_04400_));
 sg13g2_mux2_1 _11857_ (.A0(_03872_),
    .A1(_04000_),
    .S(_04394_),
    .X(_04401_));
 sg13g2_buf_1 _11858_ (.A(_04390_),
    .X(_04402_));
 sg13g2_buf_1 _11859_ (.A(net589),
    .X(_04403_));
 sg13g2_nor2_1 _11860_ (.A(net513),
    .B(_01998_),
    .Y(_04404_));
 sg13g2_a21oi_1 _11861_ (.A1(_04400_),
    .A2(_04401_),
    .Y(_04405_),
    .B1(_04404_));
 sg13g2_nand2_1 _11862_ (.Y(_04406_),
    .A(_04024_),
    .B(net137));
 sg13g2_o21ai_1 _11863_ (.B1(_04406_),
    .Y(_00362_),
    .A1(net138),
    .A2(_04405_));
 sg13g2_mux2_1 _11864_ (.A0(_04024_),
    .A1(_03906_),
    .S(net206),
    .X(_04407_));
 sg13g2_nor2_1 _11865_ (.A(net513),
    .B(_01984_),
    .Y(_04408_));
 sg13g2_a21oi_1 _11866_ (.A1(net514),
    .A2(_04407_),
    .Y(_04409_),
    .B1(_04408_));
 sg13g2_nand2_1 _11867_ (.Y(_04410_),
    .A(_04000_),
    .B(net137));
 sg13g2_o21ai_1 _11868_ (.B1(_04410_),
    .Y(_00363_),
    .A1(_04389_),
    .A2(_04409_));
 sg13g2_mux2_1 _11869_ (.A0(_04000_),
    .A1(_03963_),
    .S(net206),
    .X(_04411_));
 sg13g2_nor2_1 _11870_ (.A(net513),
    .B(_02837_),
    .Y(_04412_));
 sg13g2_a21oi_1 _11871_ (.A1(net514),
    .A2(_04411_),
    .Y(_04413_),
    .B1(_04412_));
 sg13g2_nand2_1 _11872_ (.Y(_04414_),
    .A(_03906_),
    .B(net137));
 sg13g2_o21ai_1 _11873_ (.B1(_04414_),
    .Y(_00364_),
    .A1(_04389_),
    .A2(_04413_));
 sg13g2_mux2_1 _11874_ (.A0(_03906_),
    .A1(_03982_),
    .S(net206),
    .X(_04415_));
 sg13g2_nor2_1 _11875_ (.A(net513),
    .B(_02173_),
    .Y(_04416_));
 sg13g2_a21oi_1 _11876_ (.A1(net514),
    .A2(_04415_),
    .Y(_04417_),
    .B1(_04416_));
 sg13g2_nand2_1 _11877_ (.Y(_04418_),
    .A(_03963_),
    .B(net137));
 sg13g2_o21ai_1 _11878_ (.B1(_04418_),
    .Y(_00365_),
    .A1(net138),
    .A2(_04417_));
 sg13g2_mux2_1 _11879_ (.A0(_03963_),
    .A1(_03922_),
    .S(net206),
    .X(_04419_));
 sg13g2_nor2_1 _11880_ (.A(net513),
    .B(_01892_),
    .Y(_04420_));
 sg13g2_a21oi_1 _11881_ (.A1(net514),
    .A2(_04419_),
    .Y(_04421_),
    .B1(_04420_));
 sg13g2_nand2_1 _11882_ (.Y(_04422_),
    .A(_03982_),
    .B(net137));
 sg13g2_o21ai_1 _11883_ (.B1(_04422_),
    .Y(_00366_),
    .A1(net138),
    .A2(_04421_));
 sg13g2_mux2_1 _11884_ (.A0(_03982_),
    .A1(_03687_),
    .S(net206),
    .X(_04423_));
 sg13g2_nor2_1 _11885_ (.A(net513),
    .B(_02185_),
    .Y(_04424_));
 sg13g2_a21oi_1 _11886_ (.A1(net514),
    .A2(_04423_),
    .Y(_04425_),
    .B1(_04424_));
 sg13g2_nand2_1 _11887_ (.Y(_04426_),
    .A(_03922_),
    .B(net137));
 sg13g2_o21ai_1 _11888_ (.B1(_04426_),
    .Y(_00367_),
    .A1(net138),
    .A2(_04425_));
 sg13g2_mux2_1 _11889_ (.A0(_03922_),
    .A1(_03715_),
    .S(net206),
    .X(_04427_));
 sg13g2_nor2_1 _11890_ (.A(net513),
    .B(_02217_),
    .Y(_04428_));
 sg13g2_a21oi_1 _11891_ (.A1(net514),
    .A2(_04427_),
    .Y(_04429_),
    .B1(_04428_));
 sg13g2_nand2_1 _11892_ (.Y(_04430_),
    .A(_03687_),
    .B(net137));
 sg13g2_o21ai_1 _11893_ (.B1(_04430_),
    .Y(_00368_),
    .A1(net138),
    .A2(_04429_));
 sg13g2_mux2_1 _11894_ (.A0(_03687_),
    .A1(_03674_),
    .S(net206),
    .X(_04431_));
 sg13g2_buf_1 _11895_ (.A(net589),
    .X(_04432_));
 sg13g2_nor2_1 _11896_ (.A(_04432_),
    .B(_02205_),
    .Y(_04433_));
 sg13g2_a21oi_1 _11897_ (.A1(net514),
    .A2(_04431_),
    .Y(_04434_),
    .B1(_04433_));
 sg13g2_nand2_1 _11898_ (.Y(_04435_),
    .A(_03715_),
    .B(net137));
 sg13g2_o21ai_1 _11899_ (.B1(_04435_),
    .Y(_00369_),
    .A1(net138),
    .A2(_04434_));
 sg13g2_mux2_1 _11900_ (.A0(_03715_),
    .A1(_03737_),
    .S(net206),
    .X(_04436_));
 sg13g2_nor2_1 _11901_ (.A(net512),
    .B(_02124_),
    .Y(_04437_));
 sg13g2_a21oi_1 _11902_ (.A1(net514),
    .A2(_04436_),
    .Y(_04438_),
    .B1(_04437_));
 sg13g2_buf_1 _11903_ (.A(_04388_),
    .X(_04439_));
 sg13g2_nand2_1 _11904_ (.Y(_04440_),
    .A(_03674_),
    .B(_04439_));
 sg13g2_o21ai_1 _11905_ (.B1(_04440_),
    .Y(_00370_),
    .A1(net138),
    .A2(_04438_));
 sg13g2_buf_1 _11906_ (.A(_04388_),
    .X(_04441_));
 sg13g2_buf_1 _11907_ (.A(net590),
    .X(_04442_));
 sg13g2_buf_1 _11908_ (.A(_04393_),
    .X(_04443_));
 sg13g2_mux2_1 _11909_ (.A0(_03674_),
    .A1(_04079_),
    .S(_04443_),
    .X(_04444_));
 sg13g2_nor2_1 _11910_ (.A(net512),
    .B(_02226_),
    .Y(_04445_));
 sg13g2_a21oi_1 _11911_ (.A1(_04442_),
    .A2(_04444_),
    .Y(_04446_),
    .B1(_04445_));
 sg13g2_nand2_1 _11912_ (.Y(_04447_),
    .A(_03737_),
    .B(net136));
 sg13g2_o21ai_1 _11913_ (.B1(_04447_),
    .Y(_00371_),
    .A1(_04441_),
    .A2(_04446_));
 sg13g2_mux2_1 _11914_ (.A0(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[0] ),
    .A1(_03838_),
    .S(_04443_),
    .X(_04448_));
 sg13g2_nor2_1 _11915_ (.A(_04432_),
    .B(_01775_),
    .Y(_04449_));
 sg13g2_a21oi_1 _11916_ (.A1(_04442_),
    .A2(_04448_),
    .Y(_04450_),
    .B1(_04449_));
 sg13g2_nand2_1 _11917_ (.Y(_04451_),
    .A(_01777_),
    .B(_04439_));
 sg13g2_o21ai_1 _11918_ (.B1(_04451_),
    .Y(_00372_),
    .A1(_04441_),
    .A2(_04450_));
 sg13g2_mux2_1 _11919_ (.A0(_03737_),
    .A1(_03771_),
    .S(net205),
    .X(_04452_));
 sg13g2_nor2_1 _11920_ (.A(net512),
    .B(_02054_),
    .Y(_04453_));
 sg13g2_a21oi_1 _11921_ (.A1(net511),
    .A2(_04452_),
    .Y(_04454_),
    .B1(_04453_));
 sg13g2_nand2_1 _11922_ (.Y(_04455_),
    .A(_04079_),
    .B(net136));
 sg13g2_o21ai_1 _11923_ (.B1(_04455_),
    .Y(_00373_),
    .A1(net135),
    .A2(_04454_));
 sg13g2_mux2_1 _11924_ (.A0(_04079_),
    .A1(_04067_),
    .S(net205),
    .X(_04456_));
 sg13g2_nor2_1 _11925_ (.A(net512),
    .B(_02255_),
    .Y(_04457_));
 sg13g2_a21oi_1 _11926_ (.A1(net511),
    .A2(_04456_),
    .Y(_04458_),
    .B1(_04457_));
 sg13g2_nand2_1 _11927_ (.Y(_04459_),
    .A(_03771_),
    .B(net136));
 sg13g2_o21ai_1 _11928_ (.B1(_04459_),
    .Y(_00374_),
    .A1(net135),
    .A2(_04458_));
 sg13g2_mux2_1 _11929_ (.A0(_03771_),
    .A1(_03700_),
    .S(net205),
    .X(_04460_));
 sg13g2_nor2_1 _11930_ (.A(net512),
    .B(_02090_),
    .Y(_04461_));
 sg13g2_a21oi_1 _11931_ (.A1(net511),
    .A2(_04460_),
    .Y(_04462_),
    .B1(_04461_));
 sg13g2_nand2_1 _11932_ (.Y(_04463_),
    .A(_04067_),
    .B(net136));
 sg13g2_o21ai_1 _11933_ (.B1(_04463_),
    .Y(_00375_),
    .A1(net135),
    .A2(_04462_));
 sg13g2_mux2_1 _11934_ (.A0(_04067_),
    .A1(_04049_),
    .S(net205),
    .X(_04464_));
 sg13g2_nor2_1 _11935_ (.A(net512),
    .B(_02092_),
    .Y(_04465_));
 sg13g2_a21oi_1 _11936_ (.A1(net511),
    .A2(_04464_),
    .Y(_04466_),
    .B1(_04465_));
 sg13g2_nand2_1 _11937_ (.Y(_04467_),
    .A(_03700_),
    .B(net136));
 sg13g2_o21ai_1 _11938_ (.B1(_04467_),
    .Y(_00376_),
    .A1(net135),
    .A2(_04466_));
 sg13g2_buf_1 _11939_ (.A(net589),
    .X(_04468_));
 sg13g2_buf_1 _11940_ (.A(net589),
    .X(_04469_));
 sg13g2_and2_1 _11941_ (.A(net325),
    .B(_01734_),
    .X(_04470_));
 sg13g2_buf_2 _11942_ (.A(_04470_),
    .X(_04471_));
 sg13g2_nand2_1 _11943_ (.Y(_04472_),
    .A(_03700_),
    .B(_04471_));
 sg13g2_buf_1 _11944_ (.A(_04393_),
    .X(_04473_));
 sg13g2_nand2_1 _11945_ (.Y(_04474_),
    .A(_03658_),
    .B(net204));
 sg13g2_nand3_1 _11946_ (.B(_04472_),
    .C(_04474_),
    .A(net509),
    .Y(_04475_));
 sg13g2_o21ai_1 _11947_ (.B1(_04475_),
    .Y(_04476_),
    .A1(net510),
    .A2(_02493_));
 sg13g2_nand2_1 _11948_ (.Y(_04477_),
    .A(_04049_),
    .B(net136));
 sg13g2_o21ai_1 _11949_ (.B1(_04477_),
    .Y(_00377_),
    .A1(net135),
    .A2(_04476_));
 sg13g2_mux2_1 _11950_ (.A0(_04049_),
    .A1(_04166_),
    .S(net205),
    .X(_04478_));
 sg13g2_nor2_1 _11951_ (.A(net512),
    .B(_02503_),
    .Y(_04479_));
 sg13g2_a21oi_1 _11952_ (.A1(net511),
    .A2(_04478_),
    .Y(_04480_),
    .B1(_04479_));
 sg13g2_nand2_1 _11953_ (.Y(_04481_),
    .A(_03658_),
    .B(net136));
 sg13g2_o21ai_1 _11954_ (.B1(_04481_),
    .Y(_00378_),
    .A1(net135),
    .A2(_04480_));
 sg13g2_mux2_1 _11955_ (.A0(_03658_),
    .A1(_04157_),
    .S(net205),
    .X(_04482_));
 sg13g2_nor2_1 _11956_ (.A(net512),
    .B(_02604_),
    .Y(_04483_));
 sg13g2_a21oi_1 _11957_ (.A1(net511),
    .A2(_04482_),
    .Y(_04484_),
    .B1(_04483_));
 sg13g2_nand2_1 _11958_ (.Y(_04485_),
    .A(_04166_),
    .B(net136));
 sg13g2_o21ai_1 _11959_ (.B1(_04485_),
    .Y(_00379_),
    .A1(net135),
    .A2(_04484_));
 sg13g2_mux2_1 _11960_ (.A0(_04166_),
    .A1(_03755_),
    .S(net205),
    .X(_04486_));
 sg13g2_nor2_1 _11961_ (.A(net509),
    .B(_02591_),
    .Y(_04487_));
 sg13g2_a21oi_1 _11962_ (.A1(net511),
    .A2(_04486_),
    .Y(_04488_),
    .B1(_04487_));
 sg13g2_buf_1 _11963_ (.A(_04388_),
    .X(_04489_));
 sg13g2_nand2_1 _11964_ (.Y(_04490_),
    .A(_04157_),
    .B(net134));
 sg13g2_o21ai_1 _11965_ (.B1(_04490_),
    .Y(_00380_),
    .A1(net135),
    .A2(_04488_));
 sg13g2_buf_1 _11966_ (.A(_04388_),
    .X(_04491_));
 sg13g2_mux2_1 _11967_ (.A0(_04157_),
    .A1(_03595_),
    .S(net205),
    .X(_04492_));
 sg13g2_nor2_1 _11968_ (.A(net509),
    .B(_02517_),
    .Y(_04493_));
 sg13g2_a21oi_1 _11969_ (.A1(net511),
    .A2(_04492_),
    .Y(_04494_),
    .B1(_04493_));
 sg13g2_nand2_1 _11970_ (.Y(_04495_),
    .A(_03755_),
    .B(net134));
 sg13g2_o21ai_1 _11971_ (.B1(_04495_),
    .Y(_00381_),
    .A1(net133),
    .A2(_04494_));
 sg13g2_nand2_1 _11972_ (.Y(_04496_),
    .A(_03755_),
    .B(_04471_));
 sg13g2_nand2_1 _11973_ (.Y(_04497_),
    .A(_03631_),
    .B(net204));
 sg13g2_nand3_1 _11974_ (.B(_04496_),
    .C(_04497_),
    .A(net509),
    .Y(_04498_));
 sg13g2_o21ai_1 _11975_ (.B1(_04498_),
    .Y(_04499_),
    .A1(net510),
    .A2(_02612_));
 sg13g2_nand2_1 _11976_ (.Y(_04500_),
    .A(_03595_),
    .B(net134));
 sg13g2_o21ai_1 _11977_ (.B1(_04500_),
    .Y(_00382_),
    .A1(net133),
    .A2(_04499_));
 sg13g2_mux2_1 _11978_ (.A0(_01777_),
    .A1(_03823_),
    .S(net204),
    .X(_04501_));
 sg13g2_nor2_1 _11979_ (.A(net509),
    .B(_02299_),
    .Y(_04502_));
 sg13g2_a21oi_1 _11980_ (.A1(net510),
    .A2(_04501_),
    .Y(_04503_),
    .B1(_04502_));
 sg13g2_nand2_1 _11981_ (.Y(_04504_),
    .A(_03838_),
    .B(net134));
 sg13g2_o21ai_1 _11982_ (.B1(_04504_),
    .Y(_00383_),
    .A1(net133),
    .A2(_04503_));
 sg13g2_mux2_1 _11983_ (.A0(_03595_),
    .A1(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[31] ),
    .S(net204),
    .X(_04505_));
 sg13g2_nor2_1 _11984_ (.A(net509),
    .B(net208),
    .Y(_04506_));
 sg13g2_a21oi_1 _11985_ (.A1(net510),
    .A2(_04505_),
    .Y(_04507_),
    .B1(_04506_));
 sg13g2_nand2_1 _11986_ (.Y(_04508_),
    .A(_03631_),
    .B(net134));
 sg13g2_o21ai_1 _11987_ (.B1(_04508_),
    .Y(_00384_),
    .A1(net133),
    .A2(_04507_));
 sg13g2_nand2_1 _11988_ (.Y(_04509_),
    .A(_04391_),
    .B(_04386_));
 sg13g2_nand4_1 _11989_ (.B(_01766_),
    .C(_03005_),
    .A(net589),
    .Y(_04510_),
    .D(net315));
 sg13g2_nand3_1 _11990_ (.B(_04509_),
    .C(_04510_),
    .A(net596),
    .Y(_04511_));
 sg13g2_and2_1 _11991_ (.A(_03631_),
    .B(net590),
    .X(_04512_));
 sg13g2_a22oi_1 _11992_ (.Y(_04513_),
    .B1(_04471_),
    .B2(_04512_),
    .A2(_02696_),
    .A1(_04391_));
 sg13g2_nand2_1 _11993_ (.Y(_04514_),
    .A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[31] ),
    .B(_04511_));
 sg13g2_o21ai_1 _11994_ (.B1(_04514_),
    .Y(_00385_),
    .A1(_04511_),
    .A2(_04513_));
 sg13g2_nand2_1 _11995_ (.Y(_04515_),
    .A(_03838_),
    .B(_04471_));
 sg13g2_nand2_1 _11996_ (.Y(_04516_),
    .A(_03792_),
    .B(net204));
 sg13g2_nand3_1 _11997_ (.B(_04515_),
    .C(_04516_),
    .A(net590),
    .Y(_04517_));
 sg13g2_o21ai_1 _11998_ (.B1(_04517_),
    .Y(_04518_),
    .A1(net510),
    .A2(net266));
 sg13g2_nand2_1 _11999_ (.Y(_04519_),
    .A(_03823_),
    .B(net134));
 sg13g2_o21ai_1 _12000_ (.B1(_04519_),
    .Y(_00386_),
    .A1(net133),
    .A2(_04518_));
 sg13g2_mux2_1 _12001_ (.A0(_03823_),
    .A1(_03949_),
    .S(net204),
    .X(_04520_));
 sg13g2_nor2_1 _12002_ (.A(net509),
    .B(_02401_),
    .Y(_04521_));
 sg13g2_a21oi_1 _12003_ (.A1(net510),
    .A2(_04520_),
    .Y(_04522_),
    .B1(_04521_));
 sg13g2_nand2_1 _12004_ (.Y(_04523_),
    .A(_03792_),
    .B(net134));
 sg13g2_o21ai_1 _12005_ (.B1(_04523_),
    .Y(_00387_),
    .A1(net133),
    .A2(_04522_));
 sg13g2_mux2_1 _12006_ (.A0(_03792_),
    .A1(_03890_),
    .S(net204),
    .X(_04524_));
 sg13g2_nor2_1 _12007_ (.A(net509),
    .B(_02432_),
    .Y(_04525_));
 sg13g2_a21oi_1 _12008_ (.A1(net510),
    .A2(_04524_),
    .Y(_04526_),
    .B1(_04525_));
 sg13g2_nand2_1 _12009_ (.Y(_04527_),
    .A(_03949_),
    .B(net134));
 sg13g2_o21ai_1 _12010_ (.B1(_04527_),
    .Y(_00388_),
    .A1(net133),
    .A2(_04526_));
 sg13g2_mux2_1 _12011_ (.A0(_03949_),
    .A1(_03934_),
    .S(net204),
    .X(_04528_));
 sg13g2_nor2_1 _12012_ (.A(_04469_),
    .B(_02867_),
    .Y(_04529_));
 sg13g2_a21oi_1 _12013_ (.A1(net510),
    .A2(_04528_),
    .Y(_04530_),
    .B1(_04529_));
 sg13g2_nand2_1 _12014_ (.Y(_04531_),
    .A(_03890_),
    .B(_04489_));
 sg13g2_o21ai_1 _12015_ (.B1(_04531_),
    .Y(_00389_),
    .A1(net133),
    .A2(_04530_));
 sg13g2_nand2_1 _12016_ (.Y(_04532_),
    .A(_03890_),
    .B(_04471_));
 sg13g2_nand2_1 _12017_ (.Y(_04533_),
    .A(_04034_),
    .B(_04473_));
 sg13g2_nand3_1 _12018_ (.B(_04532_),
    .C(_04533_),
    .A(net590),
    .Y(_04534_));
 sg13g2_o21ai_1 _12019_ (.B1(_04534_),
    .Y(_04535_),
    .A1(_04468_),
    .A2(_02334_));
 sg13g2_nand2_1 _12020_ (.Y(_04536_),
    .A(_03934_),
    .B(_04489_));
 sg13g2_o21ai_1 _12021_ (.B1(_04536_),
    .Y(_00390_),
    .A1(_04491_),
    .A2(_04535_));
 sg13g2_nand2_1 _12022_ (.Y(_04537_),
    .A(_03934_),
    .B(_04471_));
 sg13g2_nand2_1 _12023_ (.Y(_04538_),
    .A(_03872_),
    .B(_04393_));
 sg13g2_nand3_1 _12024_ (.B(_04537_),
    .C(_04538_),
    .A(net590),
    .Y(_04539_));
 sg13g2_o21ai_1 _12025_ (.B1(_04539_),
    .Y(_04540_),
    .A1(net513),
    .A2(_02925_));
 sg13g2_nand2_1 _12026_ (.Y(_04541_),
    .A(_04034_),
    .B(_04388_));
 sg13g2_o21ai_1 _12027_ (.B1(_04541_),
    .Y(_00391_),
    .A1(_04491_),
    .A2(_04540_));
 sg13g2_mux2_1 _12028_ (.A0(_04034_),
    .A1(_04024_),
    .S(_04473_),
    .X(_04542_));
 sg13g2_nor2_1 _12029_ (.A(_04469_),
    .B(_02935_),
    .Y(_04543_));
 sg13g2_a21oi_1 _12030_ (.A1(_04468_),
    .A2(_04542_),
    .Y(_04544_),
    .B1(_04543_));
 sg13g2_nand2_1 _12031_ (.Y(_04545_),
    .A(_03872_),
    .B(_04388_));
 sg13g2_o21ai_1 _12032_ (.B1(_04545_),
    .Y(_00392_),
    .A1(_04398_),
    .A2(_04544_));
 sg13g2_buf_1 _12033_ (.A(net447),
    .X(_04546_));
 sg13g2_nor2b_1 _12034_ (.A(_03529_),
    .B_N(_04118_),
    .Y(_04547_));
 sg13g2_a21o_1 _12035_ (.A2(_04547_),
    .A1(_04546_),
    .B1(_03569_),
    .X(_04548_));
 sg13g2_buf_2 _12036_ (.A(_04548_),
    .X(_04549_));
 sg13g2_buf_1 _12037_ (.A(_04549_),
    .X(_04550_));
 sg13g2_buf_1 _12038_ (.A(net446),
    .X(_04551_));
 sg13g2_nor2_1 _12039_ (.A(net409),
    .B(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[13] ),
    .Y(_04552_));
 sg13g2_nor3_2 _12040_ (.A(_02273_),
    .B(_02289_),
    .C(_04552_),
    .Y(_04553_));
 sg13g2_nor2_1 _12041_ (.A(net626),
    .B(net625),
    .Y(_04554_));
 sg13g2_nand3_1 _12042_ (.B(_04553_),
    .C(_04554_),
    .A(\soc_I.kianv_I.Instr[11] ),
    .Y(_04555_));
 sg13g2_buf_1 _12043_ (.A(_04555_),
    .X(_04556_));
 sg13g2_buf_1 _12044_ (.A(_04556_),
    .X(_04557_));
 sg13g2_buf_1 _12045_ (.A(net304),
    .X(_04558_));
 sg13g2_buf_1 _12046_ (.A(_04556_),
    .X(_04559_));
 sg13g2_nand2_1 _12047_ (.Y(_04560_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ),
    .B(net303));
 sg13g2_o21ai_1 _12048_ (.B1(_04560_),
    .Y(_00394_),
    .A1(_04550_),
    .A2(net261));
 sg13g2_buf_1 _12049_ (.A(net304),
    .X(_04561_));
 sg13g2_nor2_1 _12050_ (.A(_03657_),
    .B(_04123_),
    .Y(_04562_));
 sg13g2_a21oi_1 _12051_ (.A1(net413),
    .A2(_04039_),
    .Y(_04563_),
    .B1(_04562_));
 sg13g2_buf_1 _12052_ (.A(_04563_),
    .X(_04564_));
 sg13g2_buf_1 _12053_ (.A(net117),
    .X(_04565_));
 sg13g2_nand2_1 _12054_ (.Y(_04566_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ),
    .B(_04559_));
 sg13g2_o21ai_1 _12055_ (.B1(_04566_),
    .Y(_00395_),
    .A1(_04561_),
    .A2(net110));
 sg13g2_buf_1 _12056_ (.A(net129),
    .X(_04567_));
 sg13g2_buf_1 _12057_ (.A(_04556_),
    .X(_04568_));
 sg13g2_mux2_1 _12058_ (.A0(net127),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ),
    .S(net302),
    .X(_00396_));
 sg13g2_buf_1 _12059_ (.A(net131),
    .X(_04569_));
 sg13g2_nand2_1 _12060_ (.Y(_04570_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ),
    .B(net303));
 sg13g2_o21ai_1 _12061_ (.B1(_04570_),
    .Y(_00397_),
    .A1(net126),
    .A2(net261));
 sg13g2_nor2b_1 _12062_ (.A(net446),
    .B_N(\soc_I.kianv_I.datapath_unit_I.ALUOut[13] ),
    .Y(_04571_));
 sg13g2_a21oi_1 _12063_ (.A1(_04551_),
    .A2(\soc_I.kianv_I.datapath_unit_I.DataLatched[13] ),
    .Y(_04572_),
    .B1(_04571_));
 sg13g2_nand2_1 _12064_ (.Y(_04573_),
    .A(net447),
    .B(_03976_));
 sg13g2_o21ai_1 _12065_ (.B1(_04573_),
    .Y(_04574_),
    .A1(_03565_),
    .A2(_04572_));
 sg13g2_buf_1 _12066_ (.A(_04574_),
    .X(_04575_));
 sg13g2_buf_1 _12067_ (.A(net99),
    .X(_04576_));
 sg13g2_mux2_1 _12068_ (.A0(net87),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ),
    .S(net302),
    .X(_00398_));
 sg13g2_mux2_1 _12069_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[14] ),
    .S(net409),
    .X(_04577_));
 sg13g2_nand2_1 _12070_ (.Y(_04578_),
    .A(_03981_),
    .B(_03989_));
 sg13g2_o21ai_1 _12071_ (.B1(_04578_),
    .Y(_04579_),
    .A1(_04546_),
    .A2(_04577_));
 sg13g2_buf_1 _12072_ (.A(_04579_),
    .X(_04580_));
 sg13g2_buf_1 _12073_ (.A(net98),
    .X(_04581_));
 sg13g2_nand2_1 _12074_ (.Y(_04582_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ),
    .B(_04559_));
 sg13g2_o21ai_1 _12075_ (.B1(_04582_),
    .Y(_00399_),
    .A1(_04561_),
    .A2(net86));
 sg13g2_buf_1 _12076_ (.A(net130),
    .X(_04583_));
 sg13g2_nand2_1 _12077_ (.Y(_04584_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15] ),
    .B(net303));
 sg13g2_o21ai_1 _12078_ (.B1(_04584_),
    .Y(_00400_),
    .A1(net125),
    .A2(net261));
 sg13g2_mux2_1 _12079_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[16] ),
    .S(net409),
    .X(_04585_));
 sg13g2_and2_1 _12080_ (.A(_03684_),
    .B(_03691_),
    .X(_04586_));
 sg13g2_nor2_1 _12081_ (.A(net413),
    .B(_04586_),
    .Y(_04587_));
 sg13g2_a21oi_1 _12082_ (.A1(_04258_),
    .A2(_04585_),
    .Y(_04588_),
    .B1(_04587_));
 sg13g2_buf_1 _12083_ (.A(_04588_),
    .X(_04589_));
 sg13g2_buf_1 _12084_ (.A(net85),
    .X(_04590_));
 sg13g2_nand2_1 _12085_ (.Y(_04591_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ),
    .B(net303));
 sg13g2_o21ai_1 _12086_ (.B1(_04591_),
    .Y(_00401_),
    .A1(net302),
    .A2(net78));
 sg13g2_buf_1 _12087_ (.A(net121),
    .X(_04592_));
 sg13g2_nand2_1 _12088_ (.Y(_04593_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ),
    .B(net303));
 sg13g2_o21ai_1 _12089_ (.B1(_04593_),
    .Y(_00402_),
    .A1(net109),
    .A2(net261));
 sg13g2_mux2_1 _12090_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[18] ),
    .S(net409),
    .X(_04594_));
 sg13g2_nand2_1 _12091_ (.Y(_04595_),
    .A(net410),
    .B(_03681_));
 sg13g2_o21ai_1 _12092_ (.B1(_04595_),
    .Y(_04596_),
    .A1(net410),
    .A2(_04594_));
 sg13g2_buf_1 _12093_ (.A(_04596_),
    .X(_04597_));
 sg13g2_buf_1 _12094_ (.A(net97),
    .X(_04598_));
 sg13g2_nand2_1 _12095_ (.Y(_04599_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ),
    .B(net303));
 sg13g2_o21ai_1 _12096_ (.B1(_04599_),
    .Y(_00403_),
    .A1(net302),
    .A2(net84));
 sg13g2_buf_1 _12097_ (.A(net120),
    .X(_04600_));
 sg13g2_buf_1 _12098_ (.A(_04556_),
    .X(_04601_));
 sg13g2_nand2_1 _12099_ (.Y(_04602_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ),
    .B(_04601_));
 sg13g2_o21ai_1 _12100_ (.B1(_04602_),
    .Y(_00404_),
    .A1(net108),
    .A2(_04558_));
 sg13g2_buf_1 _12101_ (.A(_01800_),
    .X(_04603_));
 sg13g2_buf_1 _12102_ (.A(net124),
    .X(_04604_));
 sg13g2_nand2_1 _12103_ (.Y(_04605_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ),
    .B(_04601_));
 sg13g2_o21ai_1 _12104_ (.B1(_04605_),
    .Y(_00405_),
    .A1(net116),
    .A2(_04558_));
 sg13g2_buf_1 _12105_ (.A(_04092_),
    .X(_04606_));
 sg13g2_buf_1 _12106_ (.A(net96),
    .X(_04607_));
 sg13g2_mux2_1 _12107_ (.A0(net83),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ),
    .S(_04568_),
    .X(_00406_));
 sg13g2_a21oi_1 _12108_ (.A1(net164),
    .A2(_03770_),
    .Y(_04608_),
    .B1(_03781_));
 sg13g2_buf_2 _12109_ (.A(_04608_),
    .X(_04609_));
 sg13g2_buf_1 _12110_ (.A(_04609_),
    .X(_04610_));
 sg13g2_nand2_1 _12111_ (.Y(_04611_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ),
    .B(net301));
 sg13g2_o21ai_1 _12112_ (.B1(_04611_),
    .Y(_00407_),
    .A1(net95),
    .A2(net261));
 sg13g2_buf_1 _12113_ (.A(net112),
    .X(_04612_));
 sg13g2_nand2_1 _12114_ (.Y(_04613_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ),
    .B(net301));
 sg13g2_o21ai_1 _12115_ (.B1(_04613_),
    .Y(_00408_),
    .A1(net94),
    .A2(net261));
 sg13g2_buf_1 _12116_ (.A(net122),
    .X(_04614_));
 sg13g2_nand2_1 _12117_ (.Y(_04615_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ),
    .B(net301));
 sg13g2_o21ai_1 _12118_ (.B1(_04615_),
    .Y(_00409_),
    .A1(net107),
    .A2(net261));
 sg13g2_buf_1 _12119_ (.A(_04060_),
    .X(_04616_));
 sg13g2_nand2_1 _12120_ (.Y(_04617_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ),
    .B(net301));
 sg13g2_o21ai_1 _12121_ (.B1(_04617_),
    .Y(_00410_),
    .A1(net82),
    .A2(net261));
 sg13g2_nand2_1 _12122_ (.Y(_04618_),
    .A(_03656_),
    .B(_03667_));
 sg13g2_buf_2 _12123_ (.A(_04618_),
    .X(_04619_));
 sg13g2_buf_1 _12124_ (.A(_04619_),
    .X(_04620_));
 sg13g2_mux2_1 _12125_ (.A0(net81),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25] ),
    .S(net302),
    .X(_00411_));
 sg13g2_nand2_1 _12126_ (.Y(_04621_),
    .A(_04165_),
    .B(_04171_));
 sg13g2_nand2_1 _12127_ (.Y(_04622_),
    .A(net409),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[26] ));
 sg13g2_nand2b_1 _12128_ (.Y(_04623_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[26] ),
    .A_N(net409));
 sg13g2_a21oi_1 _12129_ (.A1(_04622_),
    .A2(_04623_),
    .Y(_04624_),
    .B1(net410));
 sg13g2_a21oi_1 _12130_ (.A1(net410),
    .A2(_04621_),
    .Y(_04625_),
    .B1(_04624_));
 sg13g2_buf_2 _12131_ (.A(_04625_),
    .X(_04626_));
 sg13g2_buf_1 _12132_ (.A(_04626_),
    .X(_04627_));
 sg13g2_nand2_1 _12133_ (.Y(_04628_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ),
    .B(net301));
 sg13g2_o21ai_1 _12134_ (.B1(_04628_),
    .Y(_00412_),
    .A1(net302),
    .A2(net80));
 sg13g2_mux2_1 _12135_ (.A0(\soc_I.kianv_I.datapath_unit_I.ALUOut[27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[27] ),
    .S(net409),
    .X(_04629_));
 sg13g2_nor2_1 _12136_ (.A(net413),
    .B(_04164_),
    .Y(_04630_));
 sg13g2_a21oi_1 _12137_ (.A1(net413),
    .A2(_04629_),
    .Y(_04631_),
    .B1(_04630_));
 sg13g2_buf_2 _12138_ (.A(_04631_),
    .X(_04632_));
 sg13g2_buf_1 _12139_ (.A(_04632_),
    .X(_04633_));
 sg13g2_nand2_1 _12140_ (.Y(_04634_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ),
    .B(net301));
 sg13g2_o21ai_1 _12141_ (.B1(_04634_),
    .Y(_00413_),
    .A1(net302),
    .A2(net79));
 sg13g2_buf_1 _12142_ (.A(net88),
    .X(_04635_));
 sg13g2_nand2_1 _12143_ (.Y(_04636_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ),
    .B(net301));
 sg13g2_o21ai_1 _12144_ (.B1(_04636_),
    .Y(_00414_),
    .A1(net77),
    .A2(net260));
 sg13g2_buf_1 _12145_ (.A(net111),
    .X(_04637_));
 sg13g2_nand2_1 _12146_ (.Y(_04638_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ),
    .B(net301));
 sg13g2_o21ai_1 _12147_ (.B1(_04638_),
    .Y(_00415_),
    .A1(net93),
    .A2(net260));
 sg13g2_inv_1 _12148_ (.Y(_04639_),
    .A(_03851_));
 sg13g2_buf_1 _12149_ (.A(_04639_),
    .X(_04640_));
 sg13g2_buf_1 _12150_ (.A(net106),
    .X(_04641_));
 sg13g2_nand2_1 _12151_ (.Y(_04642_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ),
    .B(net304));
 sg13g2_o21ai_1 _12152_ (.B1(_04642_),
    .Y(_00416_),
    .A1(net92),
    .A2(net260));
 sg13g2_buf_1 _12153_ (.A(net113),
    .X(_04643_));
 sg13g2_nand2_1 _12154_ (.Y(_04644_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ),
    .B(net304));
 sg13g2_o21ai_1 _12155_ (.B1(_04644_),
    .Y(_00417_),
    .A1(net91),
    .A2(net260));
 sg13g2_buf_1 _12156_ (.A(_03625_),
    .X(_04645_));
 sg13g2_nand2_1 _12157_ (.Y(_04646_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31] ),
    .B(net304));
 sg13g2_o21ai_1 _12158_ (.B1(_04646_),
    .Y(_00418_),
    .A1(net105),
    .A2(net260));
 sg13g2_buf_1 _12159_ (.A(net118),
    .X(_04647_));
 sg13g2_nand2_1 _12160_ (.Y(_04648_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ),
    .B(net304));
 sg13g2_o21ai_1 _12161_ (.B1(_04648_),
    .Y(_00419_),
    .A1(net104),
    .A2(net260));
 sg13g2_buf_1 _12162_ (.A(net119),
    .X(_04649_));
 sg13g2_nand2_1 _12163_ (.Y(_04650_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ),
    .B(_04557_));
 sg13g2_o21ai_1 _12164_ (.B1(_04650_),
    .Y(_00420_),
    .A1(net103),
    .A2(net260));
 sg13g2_a21o_1 _12165_ (.A2(_03386_),
    .A1(net159),
    .B1(_03953_),
    .X(_04651_));
 sg13g2_nand2_1 _12166_ (.Y(_04652_),
    .A(_04551_),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[5] ));
 sg13g2_nand2b_1 _12167_ (.Y(_04653_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[5] ),
    .A_N(_03567_));
 sg13g2_a21oi_1 _12168_ (.A1(_04652_),
    .A2(_04653_),
    .Y(_04654_),
    .B1(net447));
 sg13g2_a21oi_1 _12169_ (.A1(net410),
    .A2(_04651_),
    .Y(_04655_),
    .B1(_04654_));
 sg13g2_buf_1 _12170_ (.A(_04655_),
    .X(_04656_));
 sg13g2_buf_1 _12171_ (.A(net123),
    .X(_04657_));
 sg13g2_nand2_1 _12172_ (.Y(_04658_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ),
    .B(net304));
 sg13g2_o21ai_1 _12173_ (.B1(_04658_),
    .Y(_00421_),
    .A1(_04568_),
    .A2(net115));
 sg13g2_a21o_1 _12174_ (.A2(_03899_),
    .A1(net410),
    .B1(_03901_),
    .X(_04659_));
 sg13g2_buf_2 _12175_ (.A(_04659_),
    .X(_04660_));
 sg13g2_buf_1 _12176_ (.A(_04660_),
    .X(_04661_));
 sg13g2_nand2_1 _12177_ (.Y(_04662_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6] ),
    .B(_04557_));
 sg13g2_o21ai_1 _12178_ (.B1(_04662_),
    .Y(_00422_),
    .A1(net102),
    .A2(net260));
 sg13g2_o21ai_1 _12179_ (.B1(_03940_),
    .Y(_04663_),
    .A1(net172),
    .A2(_03493_));
 sg13g2_nand2_1 _12180_ (.Y(_04664_),
    .A(net409),
    .B(\soc_I.kianv_I.datapath_unit_I.DataLatched[7] ));
 sg13g2_nand2b_1 _12181_ (.Y(_04665_),
    .B(\soc_I.kianv_I.datapath_unit_I.ALUOut[7] ),
    .A_N(net446));
 sg13g2_a21oi_1 _12182_ (.A1(_04664_),
    .A2(_04665_),
    .Y(_04666_),
    .B1(_03565_));
 sg13g2_a21oi_1 _12183_ (.A1(net410),
    .A2(_04663_),
    .Y(_04667_),
    .B1(_04666_));
 sg13g2_buf_1 _12184_ (.A(_04667_),
    .X(_04668_));
 sg13g2_buf_1 _12185_ (.A(net101),
    .X(_04669_));
 sg13g2_nand2_1 _12186_ (.Y(_04670_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ),
    .B(net304));
 sg13g2_o21ai_1 _12187_ (.B1(_04670_),
    .Y(_00423_),
    .A1(net302),
    .A2(net90));
 sg13g2_nand2_1 _12188_ (.Y(_04671_),
    .A(net413),
    .B(_04040_));
 sg13g2_o21ai_1 _12189_ (.B1(_04671_),
    .Y(_04672_),
    .A1(net413),
    .A2(_04122_));
 sg13g2_buf_1 _12190_ (.A(_04672_),
    .X(_04673_));
 sg13g2_buf_1 _12191_ (.A(net100),
    .X(_04674_));
 sg13g2_mux2_1 _12192_ (.A0(net89),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ),
    .S(net303),
    .X(_00424_));
 sg13g2_buf_1 _12193_ (.A(net128),
    .X(_04675_));
 sg13g2_mux2_1 _12194_ (.A0(net114),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9] ),
    .S(net303),
    .X(_00425_));
 sg13g2_nand2_1 _12195_ (.Y(_04676_),
    .A(_02289_),
    .B(_04114_));
 sg13g2_nor2_1 _12196_ (.A(_02273_),
    .B(_04676_),
    .Y(_04677_));
 sg13g2_nor2b_1 _12197_ (.A(net625),
    .B_N(net626),
    .Y(_04678_));
 sg13g2_nand2_1 _12198_ (.Y(_04679_),
    .A(_04677_),
    .B(_04678_));
 sg13g2_buf_1 _12199_ (.A(_04679_),
    .X(_04680_));
 sg13g2_buf_1 _12200_ (.A(_04680_),
    .X(_04681_));
 sg13g2_buf_1 _12201_ (.A(net259),
    .X(_04682_));
 sg13g2_buf_1 _12202_ (.A(_04680_),
    .X(_04683_));
 sg13g2_nand2_1 _12203_ (.Y(_04684_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ),
    .B(net258));
 sg13g2_o21ai_1 _12204_ (.B1(_04684_),
    .Y(_00426_),
    .A1(net75),
    .A2(net203));
 sg13g2_nand2_1 _12205_ (.Y(_04685_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ),
    .B(net258));
 sg13g2_o21ai_1 _12206_ (.B1(_04685_),
    .Y(_00427_),
    .A1(net110),
    .A2(net203));
 sg13g2_buf_1 _12207_ (.A(_04680_),
    .X(_04686_));
 sg13g2_mux2_1 _12208_ (.A0(net127),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ),
    .S(net257),
    .X(_00428_));
 sg13g2_nand2_1 _12209_ (.Y(_04687_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ),
    .B(net258));
 sg13g2_o21ai_1 _12210_ (.B1(_04687_),
    .Y(_00429_),
    .A1(net126),
    .A2(net203));
 sg13g2_mux2_1 _12211_ (.A0(_04576_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ),
    .S(net257),
    .X(_00430_));
 sg13g2_nand2_1 _12212_ (.Y(_04688_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ),
    .B(net258));
 sg13g2_o21ai_1 _12213_ (.B1(_04688_),
    .Y(_00431_),
    .A1(net86),
    .A2(net203));
 sg13g2_nand2_1 _12214_ (.Y(_04689_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ),
    .B(net258));
 sg13g2_o21ai_1 _12215_ (.B1(_04689_),
    .Y(_00432_),
    .A1(_04583_),
    .A2(_04682_));
 sg13g2_nand2_1 _12216_ (.Y(_04690_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ),
    .B(net258));
 sg13g2_o21ai_1 _12217_ (.B1(_04690_),
    .Y(_00433_),
    .A1(net78),
    .A2(_04682_));
 sg13g2_nand2_1 _12218_ (.Y(_04691_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ),
    .B(net258));
 sg13g2_o21ai_1 _12219_ (.B1(_04691_),
    .Y(_00434_),
    .A1(net109),
    .A2(net203));
 sg13g2_nand2_1 _12220_ (.Y(_04692_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ),
    .B(net258));
 sg13g2_o21ai_1 _12221_ (.B1(_04692_),
    .Y(_00435_),
    .A1(net84),
    .A2(net203));
 sg13g2_buf_1 _12222_ (.A(_04680_),
    .X(_04693_));
 sg13g2_nand2_1 _12223_ (.Y(_04694_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ),
    .B(_04693_));
 sg13g2_o21ai_1 _12224_ (.B1(_04694_),
    .Y(_00436_),
    .A1(net108),
    .A2(net203));
 sg13g2_nand2_1 _12225_ (.Y(_04695_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ),
    .B(_04693_));
 sg13g2_o21ai_1 _12226_ (.B1(_04695_),
    .Y(_00437_),
    .A1(net116),
    .A2(net203));
 sg13g2_mux2_1 _12227_ (.A0(_04607_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ),
    .S(_04686_),
    .X(_00438_));
 sg13g2_buf_1 _12228_ (.A(net259),
    .X(_04696_));
 sg13g2_nand2_1 _12229_ (.Y(_04697_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ),
    .B(net256));
 sg13g2_o21ai_1 _12230_ (.B1(_04697_),
    .Y(_00439_),
    .A1(_04610_),
    .A2(_04696_));
 sg13g2_nand2_1 _12231_ (.Y(_04698_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ),
    .B(net256));
 sg13g2_o21ai_1 _12232_ (.B1(_04698_),
    .Y(_00440_),
    .A1(_04612_),
    .A2(net202));
 sg13g2_nand2_1 _12233_ (.Y(_04699_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ),
    .B(net256));
 sg13g2_o21ai_1 _12234_ (.B1(_04699_),
    .Y(_00441_),
    .A1(net107),
    .A2(net202));
 sg13g2_nand2_1 _12235_ (.Y(_04700_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ),
    .B(net256));
 sg13g2_o21ai_1 _12236_ (.B1(_04700_),
    .Y(_00442_),
    .A1(net82),
    .A2(net202));
 sg13g2_mux2_1 _12237_ (.A0(_04620_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ),
    .S(net257),
    .X(_00443_));
 sg13g2_nand2_1 _12238_ (.Y(_04701_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ),
    .B(net256));
 sg13g2_o21ai_1 _12239_ (.B1(_04701_),
    .Y(_00444_),
    .A1(_04627_),
    .A2(net202));
 sg13g2_nand2_1 _12240_ (.Y(_04702_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ),
    .B(net256));
 sg13g2_o21ai_1 _12241_ (.B1(_04702_),
    .Y(_00445_),
    .A1(_04633_),
    .A2(net202));
 sg13g2_nand2_1 _12242_ (.Y(_04703_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ),
    .B(net256));
 sg13g2_o21ai_1 _12243_ (.B1(_04703_),
    .Y(_00446_),
    .A1(net77),
    .A2(net202));
 sg13g2_nand2_1 _12244_ (.Y(_04704_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ),
    .B(net256));
 sg13g2_o21ai_1 _12245_ (.B1(_04704_),
    .Y(_00447_),
    .A1(_04637_),
    .A2(net202));
 sg13g2_nand2_1 _12246_ (.Y(_04705_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ),
    .B(net259));
 sg13g2_o21ai_1 _12247_ (.B1(_04705_),
    .Y(_00448_),
    .A1(net92),
    .A2(net202));
 sg13g2_nand2_1 _12248_ (.Y(_04706_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ),
    .B(net259));
 sg13g2_o21ai_1 _12249_ (.B1(_04706_),
    .Y(_00449_),
    .A1(net91),
    .A2(_04696_));
 sg13g2_nand2_1 _12250_ (.Y(_04707_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ),
    .B(net259));
 sg13g2_o21ai_1 _12251_ (.B1(_04707_),
    .Y(_00450_),
    .A1(_04645_),
    .A2(net257));
 sg13g2_nand2_1 _12252_ (.Y(_04708_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ),
    .B(net259));
 sg13g2_o21ai_1 _12253_ (.B1(_04708_),
    .Y(_00451_),
    .A1(net104),
    .A2(net257));
 sg13g2_nand2_1 _12254_ (.Y(_04709_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ),
    .B(net259));
 sg13g2_o21ai_1 _12255_ (.B1(_04709_),
    .Y(_00452_),
    .A1(_04649_),
    .A2(net257));
 sg13g2_nand2_1 _12256_ (.Y(_04710_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ),
    .B(net259));
 sg13g2_o21ai_1 _12257_ (.B1(_04710_),
    .Y(_00453_),
    .A1(net115),
    .A2(net257));
 sg13g2_nand2_1 _12258_ (.Y(_04711_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ),
    .B(_04681_));
 sg13g2_o21ai_1 _12259_ (.B1(_04711_),
    .Y(_00454_),
    .A1(_04661_),
    .A2(net257));
 sg13g2_nand2_1 _12260_ (.Y(_04712_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ),
    .B(_04681_));
 sg13g2_o21ai_1 _12261_ (.B1(_04712_),
    .Y(_00455_),
    .A1(_04669_),
    .A2(_04686_));
 sg13g2_mux2_1 _12262_ (.A0(_04674_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ),
    .S(_04683_),
    .X(_00456_));
 sg13g2_mux2_1 _12263_ (.A0(net114),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ),
    .S(_04683_),
    .X(_00457_));
 sg13g2_nand3_1 _12264_ (.B(net625),
    .C(_04677_),
    .A(net626),
    .Y(_04713_));
 sg13g2_buf_1 _12265_ (.A(_04713_),
    .X(_04714_));
 sg13g2_buf_1 _12266_ (.A(_04714_),
    .X(_04715_));
 sg13g2_buf_1 _12267_ (.A(net255),
    .X(_04716_));
 sg13g2_buf_1 _12268_ (.A(_04714_),
    .X(_04717_));
 sg13g2_nand2_1 _12269_ (.Y(_04718_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ),
    .B(net254));
 sg13g2_o21ai_1 _12270_ (.B1(_04718_),
    .Y(_00458_),
    .A1(net75),
    .A2(net201));
 sg13g2_nand2_1 _12271_ (.Y(_04719_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ),
    .B(net254));
 sg13g2_o21ai_1 _12272_ (.B1(_04719_),
    .Y(_00459_),
    .A1(net110),
    .A2(net201));
 sg13g2_buf_1 _12273_ (.A(_04714_),
    .X(_04720_));
 sg13g2_mux2_1 _12274_ (.A0(_04567_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ),
    .S(net253),
    .X(_00460_));
 sg13g2_nand2_1 _12275_ (.Y(_04721_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ),
    .B(net254));
 sg13g2_o21ai_1 _12276_ (.B1(_04721_),
    .Y(_00461_),
    .A1(net126),
    .A2(net201));
 sg13g2_mux2_1 _12277_ (.A0(net87),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ),
    .S(_04720_),
    .X(_00462_));
 sg13g2_nand2_1 _12278_ (.Y(_04722_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ),
    .B(net254));
 sg13g2_o21ai_1 _12279_ (.B1(_04722_),
    .Y(_00463_),
    .A1(net86),
    .A2(net201));
 sg13g2_nand2_1 _12280_ (.Y(_04723_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ),
    .B(net254));
 sg13g2_o21ai_1 _12281_ (.B1(_04723_),
    .Y(_00464_),
    .A1(net125),
    .A2(_04716_));
 sg13g2_nand2_1 _12282_ (.Y(_04724_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ),
    .B(net254));
 sg13g2_o21ai_1 _12283_ (.B1(_04724_),
    .Y(_00465_),
    .A1(net78),
    .A2(_04716_));
 sg13g2_nand2_1 _12284_ (.Y(_04725_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ),
    .B(net254));
 sg13g2_o21ai_1 _12285_ (.B1(_04725_),
    .Y(_00466_),
    .A1(net109),
    .A2(net201));
 sg13g2_nand2_1 _12286_ (.Y(_04726_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ),
    .B(net254));
 sg13g2_o21ai_1 _12287_ (.B1(_04726_),
    .Y(_00467_),
    .A1(net84),
    .A2(net201));
 sg13g2_buf_1 _12288_ (.A(_04714_),
    .X(_04727_));
 sg13g2_nand2_1 _12289_ (.Y(_04728_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ),
    .B(_04727_));
 sg13g2_o21ai_1 _12290_ (.B1(_04728_),
    .Y(_00468_),
    .A1(net108),
    .A2(net201));
 sg13g2_nand2_1 _12291_ (.Y(_04729_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ),
    .B(_04727_));
 sg13g2_o21ai_1 _12292_ (.B1(_04729_),
    .Y(_00469_),
    .A1(_04604_),
    .A2(net201));
 sg13g2_mux2_1 _12293_ (.A0(_04607_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ),
    .S(net253),
    .X(_00470_));
 sg13g2_buf_1 _12294_ (.A(net255),
    .X(_04730_));
 sg13g2_nand2_1 _12295_ (.Y(_04731_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ),
    .B(net252));
 sg13g2_o21ai_1 _12296_ (.B1(_04731_),
    .Y(_00471_),
    .A1(_04610_),
    .A2(net200));
 sg13g2_nand2_1 _12297_ (.Y(_04732_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ),
    .B(net252));
 sg13g2_o21ai_1 _12298_ (.B1(_04732_),
    .Y(_00472_),
    .A1(_04612_),
    .A2(net200));
 sg13g2_nand2_1 _12299_ (.Y(_04733_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ),
    .B(net252));
 sg13g2_o21ai_1 _12300_ (.B1(_04733_),
    .Y(_00473_),
    .A1(net107),
    .A2(net200));
 sg13g2_nand2_1 _12301_ (.Y(_04734_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ),
    .B(net252));
 sg13g2_o21ai_1 _12302_ (.B1(_04734_),
    .Y(_00474_),
    .A1(net82),
    .A2(net200));
 sg13g2_mux2_1 _12303_ (.A0(_04620_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ),
    .S(net253),
    .X(_00475_));
 sg13g2_nand2_1 _12304_ (.Y(_04735_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ),
    .B(net252));
 sg13g2_o21ai_1 _12305_ (.B1(_04735_),
    .Y(_00476_),
    .A1(_04627_),
    .A2(net200));
 sg13g2_nand2_1 _12306_ (.Y(_04736_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ),
    .B(net252));
 sg13g2_o21ai_1 _12307_ (.B1(_04736_),
    .Y(_00477_),
    .A1(_04633_),
    .A2(net200));
 sg13g2_nand2_1 _12308_ (.Y(_04737_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ),
    .B(net252));
 sg13g2_o21ai_1 _12309_ (.B1(_04737_),
    .Y(_00478_),
    .A1(_04635_),
    .A2(_04730_));
 sg13g2_nand2_1 _12310_ (.Y(_04738_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ),
    .B(net252));
 sg13g2_o21ai_1 _12311_ (.B1(_04738_),
    .Y(_00479_),
    .A1(net93),
    .A2(net200));
 sg13g2_nand2_1 _12312_ (.Y(_04739_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ),
    .B(net255));
 sg13g2_o21ai_1 _12313_ (.B1(_04739_),
    .Y(_00480_),
    .A1(_04641_),
    .A2(net200));
 sg13g2_nand2_1 _12314_ (.Y(_04740_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ),
    .B(net255));
 sg13g2_o21ai_1 _12315_ (.B1(_04740_),
    .Y(_00481_),
    .A1(net91),
    .A2(_04730_));
 sg13g2_nand2_1 _12316_ (.Y(_04741_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ),
    .B(net255));
 sg13g2_o21ai_1 _12317_ (.B1(_04741_),
    .Y(_00482_),
    .A1(_04645_),
    .A2(net253));
 sg13g2_nand2_1 _12318_ (.Y(_04742_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ),
    .B(net255));
 sg13g2_o21ai_1 _12319_ (.B1(_04742_),
    .Y(_00483_),
    .A1(net104),
    .A2(net253));
 sg13g2_nand2_1 _12320_ (.Y(_04743_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ),
    .B(net255));
 sg13g2_o21ai_1 _12321_ (.B1(_04743_),
    .Y(_00484_),
    .A1(_04649_),
    .A2(net253));
 sg13g2_nand2_1 _12322_ (.Y(_04744_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ),
    .B(net255));
 sg13g2_o21ai_1 _12323_ (.B1(_04744_),
    .Y(_00485_),
    .A1(_04657_),
    .A2(net253));
 sg13g2_nand2_1 _12324_ (.Y(_04745_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ),
    .B(_04715_));
 sg13g2_o21ai_1 _12325_ (.B1(_04745_),
    .Y(_00486_),
    .A1(_04661_),
    .A2(net253));
 sg13g2_nand2_1 _12326_ (.Y(_04746_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ),
    .B(_04715_));
 sg13g2_o21ai_1 _12327_ (.B1(_04746_),
    .Y(_00487_),
    .A1(_04669_),
    .A2(_04720_));
 sg13g2_mux2_1 _12328_ (.A0(_04674_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ),
    .S(_04717_),
    .X(_00488_));
 sg13g2_mux2_1 _12329_ (.A0(net114),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ),
    .S(_04717_),
    .X(_00489_));
 sg13g2_inv_1 _12330_ (.Y(_04747_),
    .A(_02273_));
 sg13g2_nor2_1 _12331_ (.A(_04747_),
    .B(_04676_),
    .Y(_04748_));
 sg13g2_nand2_1 _12332_ (.Y(_04749_),
    .A(_04554_),
    .B(_04748_));
 sg13g2_buf_1 _12333_ (.A(_04749_),
    .X(_04750_));
 sg13g2_buf_1 _12334_ (.A(_04750_),
    .X(_04751_));
 sg13g2_buf_1 _12335_ (.A(net251),
    .X(_04752_));
 sg13g2_buf_1 _12336_ (.A(_04750_),
    .X(_04753_));
 sg13g2_nand2_1 _12337_ (.Y(_04754_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ),
    .B(net250));
 sg13g2_o21ai_1 _12338_ (.B1(_04754_),
    .Y(_00490_),
    .A1(net75),
    .A2(net199));
 sg13g2_nand2_1 _12339_ (.Y(_04755_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ),
    .B(net250));
 sg13g2_o21ai_1 _12340_ (.B1(_04755_),
    .Y(_00491_),
    .A1(net110),
    .A2(net199));
 sg13g2_buf_1 _12341_ (.A(_04750_),
    .X(_04756_));
 sg13g2_mux2_1 _12342_ (.A0(net127),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ),
    .S(net249),
    .X(_00492_));
 sg13g2_nand2_1 _12343_ (.Y(_04757_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ),
    .B(net250));
 sg13g2_o21ai_1 _12344_ (.B1(_04757_),
    .Y(_00493_),
    .A1(net126),
    .A2(net199));
 sg13g2_mux2_1 _12345_ (.A0(net87),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ),
    .S(net249),
    .X(_00494_));
 sg13g2_nand2_1 _12346_ (.Y(_04758_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ),
    .B(net250));
 sg13g2_o21ai_1 _12347_ (.B1(_04758_),
    .Y(_00495_),
    .A1(net86),
    .A2(net199));
 sg13g2_nand2_1 _12348_ (.Y(_04759_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ),
    .B(net250));
 sg13g2_o21ai_1 _12349_ (.B1(_04759_),
    .Y(_00496_),
    .A1(net125),
    .A2(_04752_));
 sg13g2_nand2_1 _12350_ (.Y(_04760_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ),
    .B(net250));
 sg13g2_o21ai_1 _12351_ (.B1(_04760_),
    .Y(_00497_),
    .A1(net78),
    .A2(_04752_));
 sg13g2_nand2_1 _12352_ (.Y(_04761_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ),
    .B(net250));
 sg13g2_o21ai_1 _12353_ (.B1(_04761_),
    .Y(_00498_),
    .A1(net109),
    .A2(net199));
 sg13g2_nand2_1 _12354_ (.Y(_04762_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ),
    .B(net250));
 sg13g2_o21ai_1 _12355_ (.B1(_04762_),
    .Y(_00499_),
    .A1(net84),
    .A2(net199));
 sg13g2_buf_1 _12356_ (.A(_04750_),
    .X(_04763_));
 sg13g2_nand2_1 _12357_ (.Y(_04764_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19] ),
    .B(_04763_));
 sg13g2_o21ai_1 _12358_ (.B1(_04764_),
    .Y(_00500_),
    .A1(net108),
    .A2(net199));
 sg13g2_nand2_1 _12359_ (.Y(_04765_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ),
    .B(_04763_));
 sg13g2_o21ai_1 _12360_ (.B1(_04765_),
    .Y(_00501_),
    .A1(net116),
    .A2(net199));
 sg13g2_mux2_1 _12361_ (.A0(net83),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ),
    .S(_04756_),
    .X(_00502_));
 sg13g2_buf_1 _12362_ (.A(net251),
    .X(_04766_));
 sg13g2_nand2_1 _12363_ (.Y(_04767_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ),
    .B(net248));
 sg13g2_o21ai_1 _12364_ (.B1(_04767_),
    .Y(_00503_),
    .A1(net95),
    .A2(net198));
 sg13g2_nand2_1 _12365_ (.Y(_04768_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ),
    .B(net248));
 sg13g2_o21ai_1 _12366_ (.B1(_04768_),
    .Y(_00504_),
    .A1(net94),
    .A2(net198));
 sg13g2_nand2_1 _12367_ (.Y(_04769_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ),
    .B(net248));
 sg13g2_o21ai_1 _12368_ (.B1(_04769_),
    .Y(_00505_),
    .A1(net107),
    .A2(net198));
 sg13g2_nand2_1 _12369_ (.Y(_04770_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ),
    .B(net248));
 sg13g2_o21ai_1 _12370_ (.B1(_04770_),
    .Y(_00506_),
    .A1(net82),
    .A2(net198));
 sg13g2_mux2_1 _12371_ (.A0(net81),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ),
    .S(net249),
    .X(_00507_));
 sg13g2_nand2_1 _12372_ (.Y(_04771_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ),
    .B(net248));
 sg13g2_o21ai_1 _12373_ (.B1(_04771_),
    .Y(_00508_),
    .A1(net80),
    .A2(net198));
 sg13g2_nand2_1 _12374_ (.Y(_04772_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ),
    .B(net248));
 sg13g2_o21ai_1 _12375_ (.B1(_04772_),
    .Y(_00509_),
    .A1(net79),
    .A2(net198));
 sg13g2_nand2_1 _12376_ (.Y(_04773_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ),
    .B(net248));
 sg13g2_o21ai_1 _12377_ (.B1(_04773_),
    .Y(_00510_),
    .A1(net77),
    .A2(net198));
 sg13g2_nand2_1 _12378_ (.Y(_04774_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ),
    .B(net248));
 sg13g2_o21ai_1 _12379_ (.B1(_04774_),
    .Y(_00511_),
    .A1(net93),
    .A2(net198));
 sg13g2_nand2_1 _12380_ (.Y(_04775_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ),
    .B(net251));
 sg13g2_o21ai_1 _12381_ (.B1(_04775_),
    .Y(_00512_),
    .A1(net92),
    .A2(_04766_));
 sg13g2_nand2_1 _12382_ (.Y(_04776_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ),
    .B(net251));
 sg13g2_o21ai_1 _12383_ (.B1(_04776_),
    .Y(_00513_),
    .A1(net91),
    .A2(_04766_));
 sg13g2_nand2_1 _12384_ (.Y(_04777_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ),
    .B(net251));
 sg13g2_o21ai_1 _12385_ (.B1(_04777_),
    .Y(_00514_),
    .A1(net105),
    .A2(net249));
 sg13g2_nand2_1 _12386_ (.Y(_04778_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ),
    .B(net251));
 sg13g2_o21ai_1 _12387_ (.B1(_04778_),
    .Y(_00515_),
    .A1(net104),
    .A2(net249));
 sg13g2_nand2_1 _12388_ (.Y(_04779_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ),
    .B(net251));
 sg13g2_o21ai_1 _12389_ (.B1(_04779_),
    .Y(_00516_),
    .A1(net103),
    .A2(net249));
 sg13g2_nand2_1 _12390_ (.Y(_04780_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ),
    .B(net251));
 sg13g2_o21ai_1 _12391_ (.B1(_04780_),
    .Y(_00517_),
    .A1(net115),
    .A2(net249));
 sg13g2_nand2_1 _12392_ (.Y(_04781_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ),
    .B(_04751_));
 sg13g2_o21ai_1 _12393_ (.B1(_04781_),
    .Y(_00518_),
    .A1(net102),
    .A2(net249));
 sg13g2_nand2_1 _12394_ (.Y(_04782_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ),
    .B(_04751_));
 sg13g2_o21ai_1 _12395_ (.B1(_04782_),
    .Y(_00519_),
    .A1(net90),
    .A2(_04756_));
 sg13g2_mux2_1 _12396_ (.A0(net89),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ),
    .S(_04753_),
    .X(_00520_));
 sg13g2_mux2_1 _12397_ (.A0(net114),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ),
    .S(_04753_),
    .X(_00521_));
 sg13g2_nor2_1 _12398_ (.A(net626),
    .B(_01703_),
    .Y(_04783_));
 sg13g2_nand2_1 _12399_ (.Y(_04784_),
    .A(_04748_),
    .B(_04783_));
 sg13g2_buf_1 _12400_ (.A(_04784_),
    .X(_04785_));
 sg13g2_buf_1 _12401_ (.A(_04785_),
    .X(_04786_));
 sg13g2_buf_1 _12402_ (.A(net247),
    .X(_04787_));
 sg13g2_buf_1 _12403_ (.A(_04785_),
    .X(_04788_));
 sg13g2_nand2_1 _12404_ (.Y(_04789_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ),
    .B(net246));
 sg13g2_o21ai_1 _12405_ (.B1(_04789_),
    .Y(_00522_),
    .A1(net75),
    .A2(net197));
 sg13g2_nand2_1 _12406_ (.Y(_04790_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ),
    .B(net246));
 sg13g2_o21ai_1 _12407_ (.B1(_04790_),
    .Y(_00523_),
    .A1(net110),
    .A2(net197));
 sg13g2_buf_1 _12408_ (.A(_04785_),
    .X(_04791_));
 sg13g2_mux2_1 _12409_ (.A0(net127),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ),
    .S(net245),
    .X(_00524_));
 sg13g2_nand2_1 _12410_ (.Y(_04792_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ),
    .B(net246));
 sg13g2_o21ai_1 _12411_ (.B1(_04792_),
    .Y(_00525_),
    .A1(net126),
    .A2(net197));
 sg13g2_mux2_1 _12412_ (.A0(net87),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ),
    .S(net245),
    .X(_00526_));
 sg13g2_nand2_1 _12413_ (.Y(_04793_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ),
    .B(net246));
 sg13g2_o21ai_1 _12414_ (.B1(_04793_),
    .Y(_00527_),
    .A1(net86),
    .A2(net197));
 sg13g2_nand2_1 _12415_ (.Y(_04794_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ),
    .B(net246));
 sg13g2_o21ai_1 _12416_ (.B1(_04794_),
    .Y(_00528_),
    .A1(net125),
    .A2(_04787_));
 sg13g2_nand2_1 _12417_ (.Y(_04795_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ),
    .B(net246));
 sg13g2_o21ai_1 _12418_ (.B1(_04795_),
    .Y(_00529_),
    .A1(net78),
    .A2(_04787_));
 sg13g2_nand2_1 _12419_ (.Y(_04796_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ),
    .B(net246));
 sg13g2_o21ai_1 _12420_ (.B1(_04796_),
    .Y(_00530_),
    .A1(net109),
    .A2(net197));
 sg13g2_nand2_1 _12421_ (.Y(_04797_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ),
    .B(net246));
 sg13g2_o21ai_1 _12422_ (.B1(_04797_),
    .Y(_00531_),
    .A1(net84),
    .A2(net197));
 sg13g2_buf_1 _12423_ (.A(_04785_),
    .X(_04798_));
 sg13g2_nand2_1 _12424_ (.Y(_04799_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ),
    .B(_04798_));
 sg13g2_o21ai_1 _12425_ (.B1(_04799_),
    .Y(_00532_),
    .A1(net108),
    .A2(net197));
 sg13g2_nand2_1 _12426_ (.Y(_04800_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ),
    .B(_04798_));
 sg13g2_o21ai_1 _12427_ (.B1(_04800_),
    .Y(_00533_),
    .A1(net116),
    .A2(net197));
 sg13g2_mux2_1 _12428_ (.A0(net83),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ),
    .S(_04791_),
    .X(_00534_));
 sg13g2_buf_1 _12429_ (.A(net247),
    .X(_04801_));
 sg13g2_nand2_1 _12430_ (.Y(_04802_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ),
    .B(net244));
 sg13g2_o21ai_1 _12431_ (.B1(_04802_),
    .Y(_00535_),
    .A1(net95),
    .A2(net196));
 sg13g2_nand2_1 _12432_ (.Y(_04803_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ),
    .B(net244));
 sg13g2_o21ai_1 _12433_ (.B1(_04803_),
    .Y(_00536_),
    .A1(net94),
    .A2(net196));
 sg13g2_nand2_1 _12434_ (.Y(_04804_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ),
    .B(net244));
 sg13g2_o21ai_1 _12435_ (.B1(_04804_),
    .Y(_00537_),
    .A1(_04614_),
    .A2(net196));
 sg13g2_nand2_1 _12436_ (.Y(_04805_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ),
    .B(net244));
 sg13g2_o21ai_1 _12437_ (.B1(_04805_),
    .Y(_00538_),
    .A1(_04616_),
    .A2(net196));
 sg13g2_mux2_1 _12438_ (.A0(net81),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ),
    .S(net245),
    .X(_00539_));
 sg13g2_nand2_1 _12439_ (.Y(_04806_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ),
    .B(net244));
 sg13g2_o21ai_1 _12440_ (.B1(_04806_),
    .Y(_00540_),
    .A1(net80),
    .A2(net196));
 sg13g2_nand2_1 _12441_ (.Y(_04807_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ),
    .B(net244));
 sg13g2_o21ai_1 _12442_ (.B1(_04807_),
    .Y(_00541_),
    .A1(net79),
    .A2(net196));
 sg13g2_nand2_1 _12443_ (.Y(_04808_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ),
    .B(net244));
 sg13g2_o21ai_1 _12444_ (.B1(_04808_),
    .Y(_00542_),
    .A1(net77),
    .A2(net196));
 sg13g2_nand2_1 _12445_ (.Y(_04809_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ),
    .B(net244));
 sg13g2_o21ai_1 _12446_ (.B1(_04809_),
    .Y(_00543_),
    .A1(net93),
    .A2(net196));
 sg13g2_nand2_1 _12447_ (.Y(_04810_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ),
    .B(net247));
 sg13g2_o21ai_1 _12448_ (.B1(_04810_),
    .Y(_00544_),
    .A1(net92),
    .A2(_04801_));
 sg13g2_nand2_1 _12449_ (.Y(_04811_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ),
    .B(net247));
 sg13g2_o21ai_1 _12450_ (.B1(_04811_),
    .Y(_00545_),
    .A1(_04643_),
    .A2(_04801_));
 sg13g2_nand2_1 _12451_ (.Y(_04812_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ),
    .B(net247));
 sg13g2_o21ai_1 _12452_ (.B1(_04812_),
    .Y(_00546_),
    .A1(net105),
    .A2(net245));
 sg13g2_nand2_1 _12453_ (.Y(_04813_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ),
    .B(net247));
 sg13g2_o21ai_1 _12454_ (.B1(_04813_),
    .Y(_00547_),
    .A1(_04647_),
    .A2(net245));
 sg13g2_nand2_1 _12455_ (.Y(_04814_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ),
    .B(_04786_));
 sg13g2_o21ai_1 _12456_ (.B1(_04814_),
    .Y(_00548_),
    .A1(net103),
    .A2(net245));
 sg13g2_nand2_1 _12457_ (.Y(_04815_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ),
    .B(net247));
 sg13g2_o21ai_1 _12458_ (.B1(_04815_),
    .Y(_00549_),
    .A1(_04657_),
    .A2(net245));
 sg13g2_nand2_1 _12459_ (.Y(_04816_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ),
    .B(_04786_));
 sg13g2_o21ai_1 _12460_ (.B1(_04816_),
    .Y(_00550_),
    .A1(net102),
    .A2(net245));
 sg13g2_nand2_1 _12461_ (.Y(_04817_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ),
    .B(net247));
 sg13g2_o21ai_1 _12462_ (.B1(_04817_),
    .Y(_00551_),
    .A1(net90),
    .A2(_04791_));
 sg13g2_mux2_1 _12463_ (.A0(net89),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ),
    .S(_04788_),
    .X(_00552_));
 sg13g2_mux2_1 _12464_ (.A0(_04675_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ),
    .S(_04788_),
    .X(_00553_));
 sg13g2_nand2_1 _12465_ (.Y(_04818_),
    .A(_04678_),
    .B(_04748_));
 sg13g2_buf_1 _12466_ (.A(_04818_),
    .X(_04819_));
 sg13g2_buf_1 _12467_ (.A(_04819_),
    .X(_04820_));
 sg13g2_buf_1 _12468_ (.A(net243),
    .X(_04821_));
 sg13g2_buf_1 _12469_ (.A(_04819_),
    .X(_04822_));
 sg13g2_nand2_1 _12470_ (.Y(_04823_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ),
    .B(net242));
 sg13g2_o21ai_1 _12471_ (.B1(_04823_),
    .Y(_00554_),
    .A1(net75),
    .A2(net195));
 sg13g2_nand2_1 _12472_ (.Y(_04824_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ),
    .B(net242));
 sg13g2_o21ai_1 _12473_ (.B1(_04824_),
    .Y(_00555_),
    .A1(net110),
    .A2(net195));
 sg13g2_buf_1 _12474_ (.A(_04819_),
    .X(_04825_));
 sg13g2_mux2_1 _12475_ (.A0(net127),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ),
    .S(net241),
    .X(_00556_));
 sg13g2_nand2_1 _12476_ (.Y(_04826_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ),
    .B(net242));
 sg13g2_o21ai_1 _12477_ (.B1(_04826_),
    .Y(_00557_),
    .A1(net126),
    .A2(net195));
 sg13g2_mux2_1 _12478_ (.A0(net87),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ),
    .S(net241),
    .X(_00558_));
 sg13g2_nand2_1 _12479_ (.Y(_04827_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ),
    .B(net242));
 sg13g2_o21ai_1 _12480_ (.B1(_04827_),
    .Y(_00559_),
    .A1(net86),
    .A2(net195));
 sg13g2_nand2_1 _12481_ (.Y(_04828_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ),
    .B(net242));
 sg13g2_o21ai_1 _12482_ (.B1(_04828_),
    .Y(_00560_),
    .A1(net125),
    .A2(_04821_));
 sg13g2_nand2_1 _12483_ (.Y(_04829_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ),
    .B(net242));
 sg13g2_o21ai_1 _12484_ (.B1(_04829_),
    .Y(_00561_),
    .A1(net78),
    .A2(_04821_));
 sg13g2_nand2_1 _12485_ (.Y(_04830_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ),
    .B(net242));
 sg13g2_o21ai_1 _12486_ (.B1(_04830_),
    .Y(_00562_),
    .A1(net109),
    .A2(net195));
 sg13g2_nand2_1 _12487_ (.Y(_04831_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ),
    .B(net242));
 sg13g2_o21ai_1 _12488_ (.B1(_04831_),
    .Y(_00563_),
    .A1(net84),
    .A2(net195));
 sg13g2_buf_1 _12489_ (.A(_04819_),
    .X(_04832_));
 sg13g2_nand2_1 _12490_ (.Y(_04833_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ),
    .B(_04832_));
 sg13g2_o21ai_1 _12491_ (.B1(_04833_),
    .Y(_00564_),
    .A1(net108),
    .A2(net195));
 sg13g2_nand2_1 _12492_ (.Y(_04834_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ),
    .B(_04832_));
 sg13g2_o21ai_1 _12493_ (.B1(_04834_),
    .Y(_00565_),
    .A1(net116),
    .A2(net195));
 sg13g2_mux2_1 _12494_ (.A0(net83),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ),
    .S(_04825_),
    .X(_00566_));
 sg13g2_buf_1 _12495_ (.A(net243),
    .X(_04835_));
 sg13g2_nand2_1 _12496_ (.Y(_04836_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ),
    .B(net240));
 sg13g2_o21ai_1 _12497_ (.B1(_04836_),
    .Y(_00567_),
    .A1(net95),
    .A2(net194));
 sg13g2_nand2_1 _12498_ (.Y(_04837_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ),
    .B(net240));
 sg13g2_o21ai_1 _12499_ (.B1(_04837_),
    .Y(_00568_),
    .A1(net94),
    .A2(net194));
 sg13g2_nand2_1 _12500_ (.Y(_04838_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ),
    .B(net240));
 sg13g2_o21ai_1 _12501_ (.B1(_04838_),
    .Y(_00569_),
    .A1(_04614_),
    .A2(net194));
 sg13g2_nand2_1 _12502_ (.Y(_04839_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ),
    .B(net240));
 sg13g2_o21ai_1 _12503_ (.B1(_04839_),
    .Y(_00570_),
    .A1(_04616_),
    .A2(net194));
 sg13g2_mux2_1 _12504_ (.A0(net81),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ),
    .S(net241),
    .X(_00571_));
 sg13g2_nand2_1 _12505_ (.Y(_04840_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ),
    .B(net240));
 sg13g2_o21ai_1 _12506_ (.B1(_04840_),
    .Y(_00572_),
    .A1(net80),
    .A2(net194));
 sg13g2_nand2_1 _12507_ (.Y(_04841_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ),
    .B(net240));
 sg13g2_o21ai_1 _12508_ (.B1(_04841_),
    .Y(_00573_),
    .A1(net79),
    .A2(net194));
 sg13g2_nand2_1 _12509_ (.Y(_04842_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ),
    .B(net240));
 sg13g2_o21ai_1 _12510_ (.B1(_04842_),
    .Y(_00574_),
    .A1(net77),
    .A2(_04835_));
 sg13g2_nand2_1 _12511_ (.Y(_04843_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ),
    .B(net240));
 sg13g2_o21ai_1 _12512_ (.B1(_04843_),
    .Y(_00575_),
    .A1(_04637_),
    .A2(net194));
 sg13g2_nand2_1 _12513_ (.Y(_04844_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ),
    .B(net243));
 sg13g2_o21ai_1 _12514_ (.B1(_04844_),
    .Y(_00576_),
    .A1(_04641_),
    .A2(net194));
 sg13g2_nand2_1 _12515_ (.Y(_04845_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ),
    .B(net243));
 sg13g2_o21ai_1 _12516_ (.B1(_04845_),
    .Y(_00577_),
    .A1(_04643_),
    .A2(_04835_));
 sg13g2_nand2_1 _12517_ (.Y(_04846_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ),
    .B(net243));
 sg13g2_o21ai_1 _12518_ (.B1(_04846_),
    .Y(_00578_),
    .A1(net105),
    .A2(net241));
 sg13g2_nand2_1 _12519_ (.Y(_04847_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ),
    .B(net243));
 sg13g2_o21ai_1 _12520_ (.B1(_04847_),
    .Y(_00579_),
    .A1(_04647_),
    .A2(net241));
 sg13g2_nand2_1 _12521_ (.Y(_04848_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ),
    .B(net243));
 sg13g2_o21ai_1 _12522_ (.B1(_04848_),
    .Y(_00580_),
    .A1(net103),
    .A2(net241));
 sg13g2_nand2_1 _12523_ (.Y(_04849_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ),
    .B(net243));
 sg13g2_o21ai_1 _12524_ (.B1(_04849_),
    .Y(_00581_),
    .A1(net115),
    .A2(net241));
 sg13g2_nand2_1 _12525_ (.Y(_04850_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ),
    .B(_04820_));
 sg13g2_o21ai_1 _12526_ (.B1(_04850_),
    .Y(_00582_),
    .A1(net102),
    .A2(net241));
 sg13g2_nand2_1 _12527_ (.Y(_04851_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ),
    .B(_04820_));
 sg13g2_o21ai_1 _12528_ (.B1(_04851_),
    .Y(_00583_),
    .A1(net90),
    .A2(_04825_));
 sg13g2_mux2_1 _12529_ (.A0(net89),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ),
    .S(_04822_),
    .X(_00584_));
 sg13g2_mux2_1 _12530_ (.A0(_04675_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ),
    .S(_04822_),
    .X(_00585_));
 sg13g2_nand3_1 _12531_ (.B(net625),
    .C(_04748_),
    .A(net626),
    .Y(_04852_));
 sg13g2_buf_1 _12532_ (.A(_04852_),
    .X(_04853_));
 sg13g2_buf_1 _12533_ (.A(_04853_),
    .X(_04854_));
 sg13g2_buf_1 _12534_ (.A(net239),
    .X(_04855_));
 sg13g2_buf_1 _12535_ (.A(_04853_),
    .X(_04856_));
 sg13g2_nand2_1 _12536_ (.Y(_04857_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ),
    .B(net238));
 sg13g2_o21ai_1 _12537_ (.B1(_04857_),
    .Y(_00586_),
    .A1(net75),
    .A2(net193));
 sg13g2_nand2_1 _12538_ (.Y(_04858_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ),
    .B(net238));
 sg13g2_o21ai_1 _12539_ (.B1(_04858_),
    .Y(_00587_),
    .A1(net110),
    .A2(net193));
 sg13g2_buf_1 _12540_ (.A(_04853_),
    .X(_04859_));
 sg13g2_mux2_1 _12541_ (.A0(net127),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ),
    .S(net237),
    .X(_00588_));
 sg13g2_nand2_1 _12542_ (.Y(_04860_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ),
    .B(net238));
 sg13g2_o21ai_1 _12543_ (.B1(_04860_),
    .Y(_00589_),
    .A1(net126),
    .A2(net193));
 sg13g2_mux2_1 _12544_ (.A0(net87),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ),
    .S(net237),
    .X(_00590_));
 sg13g2_nand2_1 _12545_ (.Y(_04861_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ),
    .B(net238));
 sg13g2_o21ai_1 _12546_ (.B1(_04861_),
    .Y(_00591_),
    .A1(net86),
    .A2(net193));
 sg13g2_nand2_1 _12547_ (.Y(_04862_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ),
    .B(net238));
 sg13g2_o21ai_1 _12548_ (.B1(_04862_),
    .Y(_00592_),
    .A1(net125),
    .A2(_04855_));
 sg13g2_nand2_1 _12549_ (.Y(_04863_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ),
    .B(net238));
 sg13g2_o21ai_1 _12550_ (.B1(_04863_),
    .Y(_00593_),
    .A1(net78),
    .A2(_04855_));
 sg13g2_nand2_1 _12551_ (.Y(_04864_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ),
    .B(net238));
 sg13g2_o21ai_1 _12552_ (.B1(_04864_),
    .Y(_00594_),
    .A1(net109),
    .A2(net193));
 sg13g2_nand2_1 _12553_ (.Y(_04865_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ),
    .B(net238));
 sg13g2_o21ai_1 _12554_ (.B1(_04865_),
    .Y(_00595_),
    .A1(net84),
    .A2(net193));
 sg13g2_buf_1 _12555_ (.A(_04853_),
    .X(_04866_));
 sg13g2_nand2_1 _12556_ (.Y(_04867_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ),
    .B(_04866_));
 sg13g2_o21ai_1 _12557_ (.B1(_04867_),
    .Y(_00596_),
    .A1(net108),
    .A2(net193));
 sg13g2_nand2_1 _12558_ (.Y(_04868_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ),
    .B(_04866_));
 sg13g2_o21ai_1 _12559_ (.B1(_04868_),
    .Y(_00597_),
    .A1(net116),
    .A2(net193));
 sg13g2_mux2_1 _12560_ (.A0(net83),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ),
    .S(_04859_),
    .X(_00598_));
 sg13g2_buf_1 _12561_ (.A(net239),
    .X(_04869_));
 sg13g2_nand2_1 _12562_ (.Y(_04870_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ),
    .B(net236));
 sg13g2_o21ai_1 _12563_ (.B1(_04870_),
    .Y(_00599_),
    .A1(net95),
    .A2(net192));
 sg13g2_nand2_1 _12564_ (.Y(_04871_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ),
    .B(net236));
 sg13g2_o21ai_1 _12565_ (.B1(_04871_),
    .Y(_00600_),
    .A1(net94),
    .A2(net192));
 sg13g2_nand2_1 _12566_ (.Y(_04872_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ),
    .B(net236));
 sg13g2_o21ai_1 _12567_ (.B1(_04872_),
    .Y(_00601_),
    .A1(net107),
    .A2(net192));
 sg13g2_nand2_1 _12568_ (.Y(_04873_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ),
    .B(net236));
 sg13g2_o21ai_1 _12569_ (.B1(_04873_),
    .Y(_00602_),
    .A1(net82),
    .A2(net192));
 sg13g2_mux2_1 _12570_ (.A0(net81),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ),
    .S(net237),
    .X(_00603_));
 sg13g2_nand2_1 _12571_ (.Y(_04874_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ),
    .B(net236));
 sg13g2_o21ai_1 _12572_ (.B1(_04874_),
    .Y(_00604_),
    .A1(net80),
    .A2(net192));
 sg13g2_nand2_1 _12573_ (.Y(_04875_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ),
    .B(net236));
 sg13g2_o21ai_1 _12574_ (.B1(_04875_),
    .Y(_00605_),
    .A1(net79),
    .A2(net192));
 sg13g2_nand2_1 _12575_ (.Y(_04876_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ),
    .B(net236));
 sg13g2_o21ai_1 _12576_ (.B1(_04876_),
    .Y(_00606_),
    .A1(_04635_),
    .A2(_04869_));
 sg13g2_nand2_1 _12577_ (.Y(_04877_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ),
    .B(net236));
 sg13g2_o21ai_1 _12578_ (.B1(_04877_),
    .Y(_00607_),
    .A1(net93),
    .A2(net192));
 sg13g2_nand2_1 _12579_ (.Y(_04878_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ),
    .B(net239));
 sg13g2_o21ai_1 _12580_ (.B1(_04878_),
    .Y(_00608_),
    .A1(net92),
    .A2(net192));
 sg13g2_nand2_1 _12581_ (.Y(_04879_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ),
    .B(net239));
 sg13g2_o21ai_1 _12582_ (.B1(_04879_),
    .Y(_00609_),
    .A1(net91),
    .A2(_04869_));
 sg13g2_nand2_1 _12583_ (.Y(_04880_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ),
    .B(net239));
 sg13g2_o21ai_1 _12584_ (.B1(_04880_),
    .Y(_00610_),
    .A1(net105),
    .A2(net237));
 sg13g2_nand2_1 _12585_ (.Y(_04881_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ),
    .B(net239));
 sg13g2_o21ai_1 _12586_ (.B1(_04881_),
    .Y(_00611_),
    .A1(net104),
    .A2(net237));
 sg13g2_nand2_1 _12587_ (.Y(_04882_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ),
    .B(net239));
 sg13g2_o21ai_1 _12588_ (.B1(_04882_),
    .Y(_00612_),
    .A1(net103),
    .A2(net237));
 sg13g2_nand2_1 _12589_ (.Y(_04883_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ),
    .B(net239));
 sg13g2_o21ai_1 _12590_ (.B1(_04883_),
    .Y(_00613_),
    .A1(net115),
    .A2(net237));
 sg13g2_nand2_1 _12591_ (.Y(_04884_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ),
    .B(_04854_));
 sg13g2_o21ai_1 _12592_ (.B1(_04884_),
    .Y(_00614_),
    .A1(net102),
    .A2(net237));
 sg13g2_nand2_1 _12593_ (.Y(_04885_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ),
    .B(_04854_));
 sg13g2_o21ai_1 _12594_ (.B1(_04885_),
    .Y(_00615_),
    .A1(net90),
    .A2(_04859_));
 sg13g2_mux2_1 _12595_ (.A0(net89),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8] ),
    .S(_04856_),
    .X(_00616_));
 sg13g2_mux2_1 _12596_ (.A0(net114),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ),
    .S(_04856_),
    .X(_00617_));
 sg13g2_nand2_1 _12597_ (.Y(_04886_),
    .A(_04553_),
    .B(_04783_));
 sg13g2_buf_1 _12598_ (.A(_04886_),
    .X(_04887_));
 sg13g2_buf_1 _12599_ (.A(_04887_),
    .X(_04888_));
 sg13g2_buf_1 _12600_ (.A(net300),
    .X(_04889_));
 sg13g2_buf_1 _12601_ (.A(_04887_),
    .X(_04890_));
 sg13g2_nand2_1 _12602_ (.Y(_04891_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ),
    .B(net299));
 sg13g2_o21ai_1 _12603_ (.B1(_04891_),
    .Y(_00618_),
    .A1(_04550_),
    .A2(net235));
 sg13g2_nand2_1 _12604_ (.Y(_04892_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ),
    .B(net299));
 sg13g2_o21ai_1 _12605_ (.B1(_04892_),
    .Y(_00619_),
    .A1(_04565_),
    .A2(net235));
 sg13g2_buf_1 _12606_ (.A(_04887_),
    .X(_04893_));
 sg13g2_mux2_1 _12607_ (.A0(_04567_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ),
    .S(net298),
    .X(_00620_));
 sg13g2_nand2_1 _12608_ (.Y(_04894_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ),
    .B(net299));
 sg13g2_o21ai_1 _12609_ (.B1(_04894_),
    .Y(_00621_),
    .A1(_04569_),
    .A2(net235));
 sg13g2_mux2_1 _12610_ (.A0(_04576_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ),
    .S(net298),
    .X(_00622_));
 sg13g2_nand2_1 _12611_ (.Y(_04895_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ),
    .B(_04890_));
 sg13g2_o21ai_1 _12612_ (.B1(_04895_),
    .Y(_00623_),
    .A1(_04581_),
    .A2(net235));
 sg13g2_nand2_1 _12613_ (.Y(_04896_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ),
    .B(net299));
 sg13g2_o21ai_1 _12614_ (.B1(_04896_),
    .Y(_00624_),
    .A1(net125),
    .A2(_04889_));
 sg13g2_nand2_1 _12615_ (.Y(_04897_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ),
    .B(net299));
 sg13g2_o21ai_1 _12616_ (.B1(_04897_),
    .Y(_00625_),
    .A1(net78),
    .A2(_04889_));
 sg13g2_nand2_1 _12617_ (.Y(_04898_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ),
    .B(net299));
 sg13g2_o21ai_1 _12618_ (.B1(_04898_),
    .Y(_00626_),
    .A1(_04592_),
    .A2(net235));
 sg13g2_nand2_1 _12619_ (.Y(_04899_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ),
    .B(net299));
 sg13g2_o21ai_1 _12620_ (.B1(_04899_),
    .Y(_00627_),
    .A1(_04598_),
    .A2(net235));
 sg13g2_buf_1 _12621_ (.A(_04887_),
    .X(_04900_));
 sg13g2_nand2_1 _12622_ (.Y(_04901_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ),
    .B(_04900_));
 sg13g2_o21ai_1 _12623_ (.B1(_04901_),
    .Y(_00628_),
    .A1(_04600_),
    .A2(net235));
 sg13g2_nand2_1 _12624_ (.Y(_04902_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ),
    .B(_04900_));
 sg13g2_o21ai_1 _12625_ (.B1(_04902_),
    .Y(_00629_),
    .A1(net116),
    .A2(net235));
 sg13g2_mux2_1 _12626_ (.A0(net83),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ),
    .S(_04893_),
    .X(_00630_));
 sg13g2_buf_1 _12627_ (.A(net300),
    .X(_04903_));
 sg13g2_nand2_1 _12628_ (.Y(_04904_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ),
    .B(net297));
 sg13g2_o21ai_1 _12629_ (.B1(_04904_),
    .Y(_00631_),
    .A1(net95),
    .A2(_04903_));
 sg13g2_nand2_1 _12630_ (.Y(_04905_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ),
    .B(net297));
 sg13g2_o21ai_1 _12631_ (.B1(_04905_),
    .Y(_00632_),
    .A1(net94),
    .A2(net234));
 sg13g2_nand2_1 _12632_ (.Y(_04906_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ),
    .B(net297));
 sg13g2_o21ai_1 _12633_ (.B1(_04906_),
    .Y(_00633_),
    .A1(net107),
    .A2(net234));
 sg13g2_nand2_1 _12634_ (.Y(_04907_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ),
    .B(net297));
 sg13g2_o21ai_1 _12635_ (.B1(_04907_),
    .Y(_00634_),
    .A1(net82),
    .A2(net234));
 sg13g2_mux2_1 _12636_ (.A0(net81),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ),
    .S(net298),
    .X(_00635_));
 sg13g2_nand2_1 _12637_ (.Y(_04908_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ),
    .B(net297));
 sg13g2_o21ai_1 _12638_ (.B1(_04908_),
    .Y(_00636_),
    .A1(net80),
    .A2(net234));
 sg13g2_nand2_1 _12639_ (.Y(_04909_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ),
    .B(net297));
 sg13g2_o21ai_1 _12640_ (.B1(_04909_),
    .Y(_00637_),
    .A1(net79),
    .A2(net234));
 sg13g2_nand2_1 _12641_ (.Y(_04910_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ),
    .B(net297));
 sg13g2_o21ai_1 _12642_ (.B1(_04910_),
    .Y(_00638_),
    .A1(net77),
    .A2(net234));
 sg13g2_nand2_1 _12643_ (.Y(_04911_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ),
    .B(net297));
 sg13g2_o21ai_1 _12644_ (.B1(_04911_),
    .Y(_00639_),
    .A1(net93),
    .A2(net234));
 sg13g2_nand2_1 _12645_ (.Y(_04912_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ),
    .B(net300));
 sg13g2_o21ai_1 _12646_ (.B1(_04912_),
    .Y(_00640_),
    .A1(net92),
    .A2(_04903_));
 sg13g2_nand2_1 _12647_ (.Y(_04913_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ),
    .B(net300));
 sg13g2_o21ai_1 _12648_ (.B1(_04913_),
    .Y(_00641_),
    .A1(net91),
    .A2(net234));
 sg13g2_nand2_1 _12649_ (.Y(_04914_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ),
    .B(net300));
 sg13g2_o21ai_1 _12650_ (.B1(_04914_),
    .Y(_00642_),
    .A1(net105),
    .A2(net298));
 sg13g2_nand2_1 _12651_ (.Y(_04915_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ),
    .B(net300));
 sg13g2_o21ai_1 _12652_ (.B1(_04915_),
    .Y(_00643_),
    .A1(net104),
    .A2(net298));
 sg13g2_nand2_1 _12653_ (.Y(_04916_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ),
    .B(net300));
 sg13g2_o21ai_1 _12654_ (.B1(_04916_),
    .Y(_00644_),
    .A1(net103),
    .A2(net298));
 sg13g2_nand2_1 _12655_ (.Y(_04917_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ),
    .B(net300));
 sg13g2_o21ai_1 _12656_ (.B1(_04917_),
    .Y(_00645_),
    .A1(net115),
    .A2(net298));
 sg13g2_nand2_1 _12657_ (.Y(_04918_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ),
    .B(_04888_));
 sg13g2_o21ai_1 _12658_ (.B1(_04918_),
    .Y(_00646_),
    .A1(net102),
    .A2(net298));
 sg13g2_nand2_1 _12659_ (.Y(_04919_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ),
    .B(_04888_));
 sg13g2_o21ai_1 _12660_ (.B1(_04919_),
    .Y(_00647_),
    .A1(net90),
    .A2(_04893_));
 sg13g2_mux2_1 _12661_ (.A0(net89),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ),
    .S(_04890_),
    .X(_00648_));
 sg13g2_mux2_1 _12662_ (.A0(net114),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ),
    .S(net299),
    .X(_00649_));
 sg13g2_nand2_1 _12663_ (.Y(_04920_),
    .A(_04553_),
    .B(_04678_));
 sg13g2_buf_1 _12664_ (.A(_04920_),
    .X(_04921_));
 sg13g2_buf_1 _12665_ (.A(_04921_),
    .X(_04922_));
 sg13g2_buf_1 _12666_ (.A(net296),
    .X(_04923_));
 sg13g2_buf_1 _12667_ (.A(_04921_),
    .X(_04924_));
 sg13g2_nand2_1 _12668_ (.Y(_04925_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ),
    .B(net295));
 sg13g2_o21ai_1 _12669_ (.B1(_04925_),
    .Y(_00650_),
    .A1(net75),
    .A2(net233));
 sg13g2_nand2_1 _12670_ (.Y(_04926_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ),
    .B(net295));
 sg13g2_o21ai_1 _12671_ (.B1(_04926_),
    .Y(_00651_),
    .A1(_04565_),
    .A2(net233));
 sg13g2_buf_1 _12672_ (.A(_04921_),
    .X(_04927_));
 sg13g2_mux2_1 _12673_ (.A0(net127),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ),
    .S(_04927_),
    .X(_00652_));
 sg13g2_nand2_1 _12674_ (.Y(_04928_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ),
    .B(net295));
 sg13g2_o21ai_1 _12675_ (.B1(_04928_),
    .Y(_00653_),
    .A1(_04569_),
    .A2(net233));
 sg13g2_mux2_1 _12676_ (.A0(net87),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ),
    .S(net294),
    .X(_00654_));
 sg13g2_nand2_1 _12677_ (.Y(_04929_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ),
    .B(net295));
 sg13g2_o21ai_1 _12678_ (.B1(_04929_),
    .Y(_00655_),
    .A1(_04581_),
    .A2(net233));
 sg13g2_nand2_1 _12679_ (.Y(_04930_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ),
    .B(net295));
 sg13g2_o21ai_1 _12680_ (.B1(_04930_),
    .Y(_00656_),
    .A1(_04583_),
    .A2(_04923_));
 sg13g2_nand2_1 _12681_ (.Y(_04931_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ),
    .B(net295));
 sg13g2_o21ai_1 _12682_ (.B1(_04931_),
    .Y(_00657_),
    .A1(_04590_),
    .A2(_04923_));
 sg13g2_nand2_1 _12683_ (.Y(_04932_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ),
    .B(net295));
 sg13g2_o21ai_1 _12684_ (.B1(_04932_),
    .Y(_00658_),
    .A1(_04592_),
    .A2(net233));
 sg13g2_nand2_1 _12685_ (.Y(_04933_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ),
    .B(net295));
 sg13g2_o21ai_1 _12686_ (.B1(_04933_),
    .Y(_00659_),
    .A1(_04598_),
    .A2(net233));
 sg13g2_buf_1 _12687_ (.A(_04921_),
    .X(_04934_));
 sg13g2_nand2_1 _12688_ (.Y(_04935_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ),
    .B(_04934_));
 sg13g2_o21ai_1 _12689_ (.B1(_04935_),
    .Y(_00660_),
    .A1(_04600_),
    .A2(net233));
 sg13g2_nand2_1 _12690_ (.Y(_04936_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ),
    .B(_04934_));
 sg13g2_o21ai_1 _12691_ (.B1(_04936_),
    .Y(_00661_),
    .A1(_04604_),
    .A2(net233));
 sg13g2_mux2_1 _12692_ (.A0(net83),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ),
    .S(_04927_),
    .X(_00662_));
 sg13g2_buf_1 _12693_ (.A(net296),
    .X(_04937_));
 sg13g2_nand2_1 _12694_ (.Y(_04938_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ),
    .B(net293));
 sg13g2_o21ai_1 _12695_ (.B1(_04938_),
    .Y(_00663_),
    .A1(net95),
    .A2(_04937_));
 sg13g2_nand2_1 _12696_ (.Y(_04939_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ),
    .B(net293));
 sg13g2_o21ai_1 _12697_ (.B1(_04939_),
    .Y(_00664_),
    .A1(net94),
    .A2(net232));
 sg13g2_nand2_1 _12698_ (.Y(_04940_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ),
    .B(net293));
 sg13g2_o21ai_1 _12699_ (.B1(_04940_),
    .Y(_00665_),
    .A1(net107),
    .A2(net232));
 sg13g2_nand2_1 _12700_ (.Y(_04941_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ),
    .B(net293));
 sg13g2_o21ai_1 _12701_ (.B1(_04941_),
    .Y(_00666_),
    .A1(net82),
    .A2(net232));
 sg13g2_mux2_1 _12702_ (.A0(net81),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ),
    .S(net294),
    .X(_00667_));
 sg13g2_nand2_1 _12703_ (.Y(_04942_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ),
    .B(net293));
 sg13g2_o21ai_1 _12704_ (.B1(_04942_),
    .Y(_00668_),
    .A1(net80),
    .A2(net232));
 sg13g2_nand2_1 _12705_ (.Y(_04943_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ),
    .B(net293));
 sg13g2_o21ai_1 _12706_ (.B1(_04943_),
    .Y(_00669_),
    .A1(net79),
    .A2(net232));
 sg13g2_nand2_1 _12707_ (.Y(_04944_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ),
    .B(net293));
 sg13g2_o21ai_1 _12708_ (.B1(_04944_),
    .Y(_00670_),
    .A1(net77),
    .A2(net232));
 sg13g2_nand2_1 _12709_ (.Y(_04945_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ),
    .B(net293));
 sg13g2_o21ai_1 _12710_ (.B1(_04945_),
    .Y(_00671_),
    .A1(net93),
    .A2(net232));
 sg13g2_nand2_1 _12711_ (.Y(_04946_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ),
    .B(net296));
 sg13g2_o21ai_1 _12712_ (.B1(_04946_),
    .Y(_00672_),
    .A1(net92),
    .A2(_04937_));
 sg13g2_nand2_1 _12713_ (.Y(_04947_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ),
    .B(net296));
 sg13g2_o21ai_1 _12714_ (.B1(_04947_),
    .Y(_00673_),
    .A1(net91),
    .A2(net232));
 sg13g2_nand2_1 _12715_ (.Y(_04948_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ),
    .B(net296));
 sg13g2_o21ai_1 _12716_ (.B1(_04948_),
    .Y(_00674_),
    .A1(net105),
    .A2(net294));
 sg13g2_nand2_1 _12717_ (.Y(_04949_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ),
    .B(net296));
 sg13g2_o21ai_1 _12718_ (.B1(_04949_),
    .Y(_00675_),
    .A1(net104),
    .A2(net294));
 sg13g2_nand2_1 _12719_ (.Y(_04950_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ),
    .B(net296));
 sg13g2_o21ai_1 _12720_ (.B1(_04950_),
    .Y(_00676_),
    .A1(net103),
    .A2(net294));
 sg13g2_nand2_1 _12721_ (.Y(_04951_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ),
    .B(net296));
 sg13g2_o21ai_1 _12722_ (.B1(_04951_),
    .Y(_00677_),
    .A1(net115),
    .A2(net294));
 sg13g2_nand2_1 _12723_ (.Y(_04952_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ),
    .B(_04922_));
 sg13g2_o21ai_1 _12724_ (.B1(_04952_),
    .Y(_00678_),
    .A1(net102),
    .A2(net294));
 sg13g2_nand2_1 _12725_ (.Y(_04953_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ),
    .B(_04922_));
 sg13g2_o21ai_1 _12726_ (.B1(_04953_),
    .Y(_00679_),
    .A1(net90),
    .A2(net294));
 sg13g2_mux2_1 _12727_ (.A0(net89),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ),
    .S(_04924_),
    .X(_00680_));
 sg13g2_mux2_1 _12728_ (.A0(net114),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ),
    .S(_04924_),
    .X(_00681_));
 sg13g2_nand3_1 _12729_ (.B(net625),
    .C(_04553_),
    .A(net626),
    .Y(_04954_));
 sg13g2_buf_1 _12730_ (.A(_04954_),
    .X(_04955_));
 sg13g2_buf_1 _12731_ (.A(_04955_),
    .X(_04956_));
 sg13g2_buf_1 _12732_ (.A(net292),
    .X(_04957_));
 sg13g2_buf_1 _12733_ (.A(_04955_),
    .X(_04958_));
 sg13g2_nand2_1 _12734_ (.Y(_04959_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ),
    .B(net291));
 sg13g2_o21ai_1 _12735_ (.B1(_04959_),
    .Y(_00682_),
    .A1(net75),
    .A2(net231));
 sg13g2_nand2_1 _12736_ (.Y(_04960_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ),
    .B(net291));
 sg13g2_o21ai_1 _12737_ (.B1(_04960_),
    .Y(_00683_),
    .A1(net110),
    .A2(net231));
 sg13g2_buf_1 _12738_ (.A(_04955_),
    .X(_04961_));
 sg13g2_mux2_1 _12739_ (.A0(net127),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ),
    .S(_04961_),
    .X(_00684_));
 sg13g2_nand2_1 _12740_ (.Y(_04962_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ),
    .B(net291));
 sg13g2_o21ai_1 _12741_ (.B1(_04962_),
    .Y(_00685_),
    .A1(net126),
    .A2(net231));
 sg13g2_mux2_1 _12742_ (.A0(net87),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ),
    .S(_04961_),
    .X(_00686_));
 sg13g2_nand2_1 _12743_ (.Y(_04963_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ),
    .B(net291));
 sg13g2_o21ai_1 _12744_ (.B1(_04963_),
    .Y(_00687_),
    .A1(net86),
    .A2(net231));
 sg13g2_nand2_1 _12745_ (.Y(_04964_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ),
    .B(net291));
 sg13g2_o21ai_1 _12746_ (.B1(_04964_),
    .Y(_00688_),
    .A1(net125),
    .A2(_04957_));
 sg13g2_nand2_1 _12747_ (.Y(_04965_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ),
    .B(net291));
 sg13g2_o21ai_1 _12748_ (.B1(_04965_),
    .Y(_00689_),
    .A1(_04590_),
    .A2(_04957_));
 sg13g2_nand2_1 _12749_ (.Y(_04966_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ),
    .B(net291));
 sg13g2_o21ai_1 _12750_ (.B1(_04966_),
    .Y(_00690_),
    .A1(net109),
    .A2(net231));
 sg13g2_nand2_1 _12751_ (.Y(_04967_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ),
    .B(net291));
 sg13g2_o21ai_1 _12752_ (.B1(_04967_),
    .Y(_00691_),
    .A1(net84),
    .A2(net231));
 sg13g2_buf_1 _12753_ (.A(_04955_),
    .X(_04968_));
 sg13g2_nand2_1 _12754_ (.Y(_04969_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ),
    .B(_04968_));
 sg13g2_o21ai_1 _12755_ (.B1(_04969_),
    .Y(_00692_),
    .A1(net108),
    .A2(net231));
 sg13g2_nand2_1 _12756_ (.Y(_04970_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ),
    .B(_04968_));
 sg13g2_o21ai_1 _12757_ (.B1(_04970_),
    .Y(_00693_),
    .A1(net116),
    .A2(net231));
 sg13g2_mux2_1 _12758_ (.A0(net83),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ),
    .S(net290),
    .X(_00694_));
 sg13g2_buf_1 _12759_ (.A(net292),
    .X(_04971_));
 sg13g2_nand2_1 _12760_ (.Y(_04972_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ),
    .B(net289));
 sg13g2_o21ai_1 _12761_ (.B1(_04972_),
    .Y(_00695_),
    .A1(net95),
    .A2(_04971_));
 sg13g2_nand2_1 _12762_ (.Y(_04973_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ),
    .B(net289));
 sg13g2_o21ai_1 _12763_ (.B1(_04973_),
    .Y(_00696_),
    .A1(net94),
    .A2(net230));
 sg13g2_nand2_1 _12764_ (.Y(_04974_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ),
    .B(net289));
 sg13g2_o21ai_1 _12765_ (.B1(_04974_),
    .Y(_00697_),
    .A1(net107),
    .A2(net230));
 sg13g2_nand2_1 _12766_ (.Y(_04975_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ),
    .B(net289));
 sg13g2_o21ai_1 _12767_ (.B1(_04975_),
    .Y(_00698_),
    .A1(net82),
    .A2(net230));
 sg13g2_mux2_1 _12768_ (.A0(net81),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ),
    .S(net290),
    .X(_00699_));
 sg13g2_nand2_1 _12769_ (.Y(_04976_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ),
    .B(net289));
 sg13g2_o21ai_1 _12770_ (.B1(_04976_),
    .Y(_00700_),
    .A1(net80),
    .A2(net230));
 sg13g2_nand2_1 _12771_ (.Y(_04977_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ),
    .B(net289));
 sg13g2_o21ai_1 _12772_ (.B1(_04977_),
    .Y(_00701_),
    .A1(net79),
    .A2(net230));
 sg13g2_nand2_1 _12773_ (.Y(_04978_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ),
    .B(net289));
 sg13g2_o21ai_1 _12774_ (.B1(_04978_),
    .Y(_00702_),
    .A1(net77),
    .A2(net230));
 sg13g2_nand2_1 _12775_ (.Y(_04979_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ),
    .B(net289));
 sg13g2_o21ai_1 _12776_ (.B1(_04979_),
    .Y(_00703_),
    .A1(net93),
    .A2(net230));
 sg13g2_nand2_1 _12777_ (.Y(_04980_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ),
    .B(net292));
 sg13g2_o21ai_1 _12778_ (.B1(_04980_),
    .Y(_00704_),
    .A1(net92),
    .A2(_04971_));
 sg13g2_nand2_1 _12779_ (.Y(_04981_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ),
    .B(net292));
 sg13g2_o21ai_1 _12780_ (.B1(_04981_),
    .Y(_00705_),
    .A1(net91),
    .A2(net230));
 sg13g2_nand2_1 _12781_ (.Y(_04982_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ),
    .B(net292));
 sg13g2_o21ai_1 _12782_ (.B1(_04982_),
    .Y(_00706_),
    .A1(net105),
    .A2(net290));
 sg13g2_nand2_1 _12783_ (.Y(_04983_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ),
    .B(net292));
 sg13g2_o21ai_1 _12784_ (.B1(_04983_),
    .Y(_00707_),
    .A1(net104),
    .A2(net290));
 sg13g2_nand2_1 _12785_ (.Y(_04984_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ),
    .B(net292));
 sg13g2_o21ai_1 _12786_ (.B1(_04984_),
    .Y(_00708_),
    .A1(net103),
    .A2(net290));
 sg13g2_nand2_1 _12787_ (.Y(_04985_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ),
    .B(net292));
 sg13g2_o21ai_1 _12788_ (.B1(_04985_),
    .Y(_00709_),
    .A1(net115),
    .A2(net290));
 sg13g2_nand2_1 _12789_ (.Y(_04986_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ),
    .B(_04956_));
 sg13g2_o21ai_1 _12790_ (.B1(_04986_),
    .Y(_00710_),
    .A1(net102),
    .A2(net290));
 sg13g2_nand2_1 _12791_ (.Y(_04987_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ),
    .B(_04956_));
 sg13g2_o21ai_1 _12792_ (.B1(_04987_),
    .Y(_00711_),
    .A1(net90),
    .A2(net290));
 sg13g2_mux2_1 _12793_ (.A0(net89),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ),
    .S(_04958_),
    .X(_00712_));
 sg13g2_mux2_1 _12794_ (.A0(net114),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ),
    .S(_04958_),
    .X(_00713_));
 sg13g2_nor3_2 _12795_ (.A(_04747_),
    .B(_02289_),
    .C(_04552_),
    .Y(_04988_));
 sg13g2_nand2_1 _12796_ (.Y(_04989_),
    .A(_04554_),
    .B(_04988_));
 sg13g2_buf_1 _12797_ (.A(_04989_),
    .X(_04990_));
 sg13g2_buf_1 _12798_ (.A(_04990_),
    .X(_04991_));
 sg13g2_buf_1 _12799_ (.A(net288),
    .X(_04992_));
 sg13g2_buf_1 _12800_ (.A(_04990_),
    .X(_04993_));
 sg13g2_nand2_1 _12801_ (.Y(_04994_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ),
    .B(net287));
 sg13g2_o21ai_1 _12802_ (.B1(_04994_),
    .Y(_00714_),
    .A1(_04549_),
    .A2(net229));
 sg13g2_nand2_1 _12803_ (.Y(_04995_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ),
    .B(net287));
 sg13g2_o21ai_1 _12804_ (.B1(_04995_),
    .Y(_00715_),
    .A1(net117),
    .A2(net229));
 sg13g2_buf_1 _12805_ (.A(_04990_),
    .X(_04996_));
 sg13g2_mux2_1 _12806_ (.A0(net129),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ),
    .S(net286),
    .X(_00716_));
 sg13g2_nand2_1 _12807_ (.Y(_04997_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ),
    .B(net287));
 sg13g2_o21ai_1 _12808_ (.B1(_04997_),
    .Y(_00717_),
    .A1(net131),
    .A2(net229));
 sg13g2_mux2_1 _12809_ (.A0(net99),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ),
    .S(_04996_),
    .X(_00718_));
 sg13g2_nand2_1 _12810_ (.Y(_04998_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ),
    .B(_04993_));
 sg13g2_o21ai_1 _12811_ (.B1(_04998_),
    .Y(_00719_),
    .A1(net98),
    .A2(net229));
 sg13g2_nand2_1 _12812_ (.Y(_04999_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ),
    .B(net287));
 sg13g2_o21ai_1 _12813_ (.B1(_04999_),
    .Y(_00720_),
    .A1(net130),
    .A2(_04992_));
 sg13g2_nand2_1 _12814_ (.Y(_05000_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ),
    .B(net287));
 sg13g2_o21ai_1 _12815_ (.B1(_05000_),
    .Y(_00721_),
    .A1(net85),
    .A2(net229));
 sg13g2_nand2_1 _12816_ (.Y(_05001_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ),
    .B(net287));
 sg13g2_o21ai_1 _12817_ (.B1(_05001_),
    .Y(_00722_),
    .A1(net121),
    .A2(_04992_));
 sg13g2_nand2_1 _12818_ (.Y(_05002_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ),
    .B(net287));
 sg13g2_o21ai_1 _12819_ (.B1(_05002_),
    .Y(_00723_),
    .A1(net97),
    .A2(net229));
 sg13g2_buf_1 _12820_ (.A(_04990_),
    .X(_05003_));
 sg13g2_nand2_1 _12821_ (.Y(_05004_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ),
    .B(_05003_));
 sg13g2_o21ai_1 _12822_ (.B1(_05004_),
    .Y(_00724_),
    .A1(net120),
    .A2(net229));
 sg13g2_nand2_1 _12823_ (.Y(_05005_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ),
    .B(_05003_));
 sg13g2_o21ai_1 _12824_ (.B1(_05005_),
    .Y(_00725_),
    .A1(net124),
    .A2(net229));
 sg13g2_mux2_1 _12825_ (.A0(net96),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ),
    .S(_04996_),
    .X(_00726_));
 sg13g2_buf_1 _12826_ (.A(net288),
    .X(_05006_));
 sg13g2_nand2_1 _12827_ (.Y(_05007_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ),
    .B(net285));
 sg13g2_o21ai_1 _12828_ (.B1(_05007_),
    .Y(_00727_),
    .A1(_04609_),
    .A2(_05006_));
 sg13g2_nand2_1 _12829_ (.Y(_05008_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ),
    .B(net285));
 sg13g2_o21ai_1 _12830_ (.B1(_05008_),
    .Y(_00728_),
    .A1(net112),
    .A2(net228));
 sg13g2_nand2_1 _12831_ (.Y(_05009_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ),
    .B(net285));
 sg13g2_o21ai_1 _12832_ (.B1(_05009_),
    .Y(_00729_),
    .A1(net122),
    .A2(net228));
 sg13g2_nand2_1 _12833_ (.Y(_05010_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ),
    .B(net285));
 sg13g2_o21ai_1 _12834_ (.B1(_05010_),
    .Y(_00730_),
    .A1(_04060_),
    .A2(net228));
 sg13g2_mux2_1 _12835_ (.A0(_04619_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ),
    .S(net286),
    .X(_00731_));
 sg13g2_nand2_1 _12836_ (.Y(_05011_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ),
    .B(net285));
 sg13g2_o21ai_1 _12837_ (.B1(_05011_),
    .Y(_00732_),
    .A1(_04626_),
    .A2(net228));
 sg13g2_nand2_1 _12838_ (.Y(_05012_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ),
    .B(net285));
 sg13g2_o21ai_1 _12839_ (.B1(_05012_),
    .Y(_00733_),
    .A1(_04632_),
    .A2(net228));
 sg13g2_nand2_1 _12840_ (.Y(_05013_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ),
    .B(net285));
 sg13g2_o21ai_1 _12841_ (.B1(_05013_),
    .Y(_00734_),
    .A1(net88),
    .A2(net228));
 sg13g2_nand2_1 _12842_ (.Y(_05014_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ),
    .B(net285));
 sg13g2_o21ai_1 _12843_ (.B1(_05014_),
    .Y(_00735_),
    .A1(net111),
    .A2(net228));
 sg13g2_nand2_1 _12844_ (.Y(_05015_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ),
    .B(net288));
 sg13g2_o21ai_1 _12845_ (.B1(_05015_),
    .Y(_00736_),
    .A1(net106),
    .A2(net228));
 sg13g2_nand2_1 _12846_ (.Y(_05016_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ),
    .B(net288));
 sg13g2_o21ai_1 _12847_ (.B1(_05016_),
    .Y(_00737_),
    .A1(net113),
    .A2(_05006_));
 sg13g2_nand2_1 _12848_ (.Y(_05017_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ),
    .B(net288));
 sg13g2_o21ai_1 _12849_ (.B1(_05017_),
    .Y(_00738_),
    .A1(_03625_),
    .A2(net286));
 sg13g2_nand2_1 _12850_ (.Y(_05018_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ),
    .B(net288));
 sg13g2_o21ai_1 _12851_ (.B1(_05018_),
    .Y(_00739_),
    .A1(net118),
    .A2(net286));
 sg13g2_nand2_1 _12852_ (.Y(_05019_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ),
    .B(_04991_));
 sg13g2_o21ai_1 _12853_ (.B1(_05019_),
    .Y(_00740_),
    .A1(net119),
    .A2(net286));
 sg13g2_nand2_1 _12854_ (.Y(_05020_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ),
    .B(net288));
 sg13g2_o21ai_1 _12855_ (.B1(_05020_),
    .Y(_00741_),
    .A1(net123),
    .A2(net286));
 sg13g2_nand2_1 _12856_ (.Y(_05021_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ),
    .B(_04991_));
 sg13g2_o21ai_1 _12857_ (.B1(_05021_),
    .Y(_00742_),
    .A1(_04660_),
    .A2(net286));
 sg13g2_nand2_1 _12858_ (.Y(_05022_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ),
    .B(net288));
 sg13g2_o21ai_1 _12859_ (.B1(_05022_),
    .Y(_00743_),
    .A1(net101),
    .A2(net286));
 sg13g2_mux2_1 _12860_ (.A0(net100),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ),
    .S(net287),
    .X(_00744_));
 sg13g2_mux2_1 _12861_ (.A0(net128),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ),
    .S(_04993_),
    .X(_00745_));
 sg13g2_nand2_1 _12862_ (.Y(_05023_),
    .A(_04783_),
    .B(_04988_));
 sg13g2_buf_1 _12863_ (.A(_05023_),
    .X(_05024_));
 sg13g2_buf_1 _12864_ (.A(_05024_),
    .X(_05025_));
 sg13g2_buf_1 _12865_ (.A(net284),
    .X(_05026_));
 sg13g2_buf_1 _12866_ (.A(_05024_),
    .X(_05027_));
 sg13g2_nand2_1 _12867_ (.Y(_05028_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ),
    .B(net283));
 sg13g2_o21ai_1 _12868_ (.B1(_05028_),
    .Y(_00746_),
    .A1(_04549_),
    .A2(net227));
 sg13g2_nand2_1 _12869_ (.Y(_05029_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ),
    .B(net283));
 sg13g2_o21ai_1 _12870_ (.B1(_05029_),
    .Y(_00747_),
    .A1(_04564_),
    .A2(net227));
 sg13g2_buf_1 _12871_ (.A(_05024_),
    .X(_05030_));
 sg13g2_mux2_1 _12872_ (.A0(net129),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ),
    .S(net282),
    .X(_00748_));
 sg13g2_nand2_1 _12873_ (.Y(_05031_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ),
    .B(net283));
 sg13g2_o21ai_1 _12874_ (.B1(_05031_),
    .Y(_00749_),
    .A1(net131),
    .A2(net227));
 sg13g2_mux2_1 _12875_ (.A0(net99),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ),
    .S(_05030_),
    .X(_00750_));
 sg13g2_nand2_1 _12876_ (.Y(_05032_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ),
    .B(_05027_));
 sg13g2_o21ai_1 _12877_ (.B1(_05032_),
    .Y(_00751_),
    .A1(_04580_),
    .A2(net227));
 sg13g2_nand2_1 _12878_ (.Y(_05033_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ),
    .B(net283));
 sg13g2_o21ai_1 _12879_ (.B1(_05033_),
    .Y(_00752_),
    .A1(net130),
    .A2(_05026_));
 sg13g2_nand2_1 _12880_ (.Y(_05034_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ),
    .B(net283));
 sg13g2_o21ai_1 _12881_ (.B1(_05034_),
    .Y(_00753_),
    .A1(net85),
    .A2(_05026_));
 sg13g2_nand2_1 _12882_ (.Y(_05035_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ),
    .B(net283));
 sg13g2_o21ai_1 _12883_ (.B1(_05035_),
    .Y(_00754_),
    .A1(net121),
    .A2(net227));
 sg13g2_nand2_1 _12884_ (.Y(_05036_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ),
    .B(net283));
 sg13g2_o21ai_1 _12885_ (.B1(_05036_),
    .Y(_00755_),
    .A1(net97),
    .A2(net227));
 sg13g2_buf_1 _12886_ (.A(_05024_),
    .X(_05037_));
 sg13g2_nand2_1 _12887_ (.Y(_05038_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ),
    .B(_05037_));
 sg13g2_o21ai_1 _12888_ (.B1(_05038_),
    .Y(_00756_),
    .A1(net120),
    .A2(net227));
 sg13g2_nand2_1 _12889_ (.Y(_05039_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ),
    .B(_05037_));
 sg13g2_o21ai_1 _12890_ (.B1(_05039_),
    .Y(_00757_),
    .A1(net124),
    .A2(net227));
 sg13g2_mux2_1 _12891_ (.A0(net96),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ),
    .S(_05030_),
    .X(_00758_));
 sg13g2_buf_1 _12892_ (.A(net284),
    .X(_05040_));
 sg13g2_nand2_1 _12893_ (.Y(_05041_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ),
    .B(net281));
 sg13g2_o21ai_1 _12894_ (.B1(_05041_),
    .Y(_00759_),
    .A1(_04609_),
    .A2(net226));
 sg13g2_nand2_1 _12895_ (.Y(_05042_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ),
    .B(net281));
 sg13g2_o21ai_1 _12896_ (.B1(_05042_),
    .Y(_00760_),
    .A1(net112),
    .A2(net226));
 sg13g2_nand2_1 _12897_ (.Y(_05043_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ),
    .B(net281));
 sg13g2_o21ai_1 _12898_ (.B1(_05043_),
    .Y(_00761_),
    .A1(net122),
    .A2(net226));
 sg13g2_nand2_1 _12899_ (.Y(_05044_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ),
    .B(net281));
 sg13g2_o21ai_1 _12900_ (.B1(_05044_),
    .Y(_00762_),
    .A1(_04060_),
    .A2(net226));
 sg13g2_mux2_1 _12901_ (.A0(_04619_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ),
    .S(net282),
    .X(_00763_));
 sg13g2_nand2_1 _12902_ (.Y(_05045_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ),
    .B(net281));
 sg13g2_o21ai_1 _12903_ (.B1(_05045_),
    .Y(_00764_),
    .A1(_04626_),
    .A2(net226));
 sg13g2_nand2_1 _12904_ (.Y(_05046_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ),
    .B(net281));
 sg13g2_o21ai_1 _12905_ (.B1(_05046_),
    .Y(_00765_),
    .A1(_04632_),
    .A2(net226));
 sg13g2_nand2_1 _12906_ (.Y(_05047_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ),
    .B(net281));
 sg13g2_o21ai_1 _12907_ (.B1(_05047_),
    .Y(_00766_),
    .A1(net88),
    .A2(_05040_));
 sg13g2_nand2_1 _12908_ (.Y(_05048_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ),
    .B(net281));
 sg13g2_o21ai_1 _12909_ (.B1(_05048_),
    .Y(_00767_),
    .A1(net111),
    .A2(net226));
 sg13g2_nand2_1 _12910_ (.Y(_05049_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ),
    .B(net284));
 sg13g2_o21ai_1 _12911_ (.B1(_05049_),
    .Y(_00768_),
    .A1(net106),
    .A2(net226));
 sg13g2_nand2_1 _12912_ (.Y(_05050_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ),
    .B(net284));
 sg13g2_o21ai_1 _12913_ (.B1(_05050_),
    .Y(_00769_),
    .A1(net113),
    .A2(_05040_));
 sg13g2_nand2_1 _12914_ (.Y(_05051_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ),
    .B(net284));
 sg13g2_o21ai_1 _12915_ (.B1(_05051_),
    .Y(_00770_),
    .A1(_03625_),
    .A2(net282));
 sg13g2_nand2_1 _12916_ (.Y(_05052_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ),
    .B(net284));
 sg13g2_o21ai_1 _12917_ (.B1(_05052_),
    .Y(_00771_),
    .A1(net118),
    .A2(net282));
 sg13g2_nand2_1 _12918_ (.Y(_05053_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ),
    .B(net284));
 sg13g2_o21ai_1 _12919_ (.B1(_05053_),
    .Y(_00772_),
    .A1(net119),
    .A2(net282));
 sg13g2_nand2_1 _12920_ (.Y(_05054_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ),
    .B(net284));
 sg13g2_o21ai_1 _12921_ (.B1(_05054_),
    .Y(_00773_),
    .A1(net123),
    .A2(net282));
 sg13g2_nand2_1 _12922_ (.Y(_05055_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ),
    .B(_05025_));
 sg13g2_o21ai_1 _12923_ (.B1(_05055_),
    .Y(_00774_),
    .A1(_04660_),
    .A2(net282));
 sg13g2_nand2_1 _12924_ (.Y(_05056_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ),
    .B(_05025_));
 sg13g2_o21ai_1 _12925_ (.B1(_05056_),
    .Y(_00775_),
    .A1(net101),
    .A2(net282));
 sg13g2_mux2_1 _12926_ (.A0(net100),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ),
    .S(net283),
    .X(_00776_));
 sg13g2_mux2_1 _12927_ (.A0(net128),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ),
    .S(_05027_),
    .X(_00777_));
 sg13g2_nand2_1 _12928_ (.Y(_05057_),
    .A(_04678_),
    .B(_04988_));
 sg13g2_buf_1 _12929_ (.A(_05057_),
    .X(_05058_));
 sg13g2_buf_1 _12930_ (.A(_05058_),
    .X(_05059_));
 sg13g2_buf_1 _12931_ (.A(net280),
    .X(_05060_));
 sg13g2_buf_1 _12932_ (.A(_05058_),
    .X(_05061_));
 sg13g2_nand2_1 _12933_ (.Y(_05062_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ),
    .B(net279));
 sg13g2_o21ai_1 _12934_ (.B1(_05062_),
    .Y(_00778_),
    .A1(_04549_),
    .A2(net225));
 sg13g2_nand2_1 _12935_ (.Y(_05063_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ),
    .B(net279));
 sg13g2_o21ai_1 _12936_ (.B1(_05063_),
    .Y(_00779_),
    .A1(net117),
    .A2(net225));
 sg13g2_buf_1 _12937_ (.A(_05058_),
    .X(_05064_));
 sg13g2_mux2_1 _12938_ (.A0(net129),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ),
    .S(net278),
    .X(_00780_));
 sg13g2_nand2_1 _12939_ (.Y(_05065_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ),
    .B(net279));
 sg13g2_o21ai_1 _12940_ (.B1(_05065_),
    .Y(_00781_),
    .A1(net131),
    .A2(net225));
 sg13g2_mux2_1 _12941_ (.A0(net99),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ),
    .S(_05064_),
    .X(_00782_));
 sg13g2_nand2_1 _12942_ (.Y(_05066_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ),
    .B(net279));
 sg13g2_o21ai_1 _12943_ (.B1(_05066_),
    .Y(_00783_),
    .A1(net98),
    .A2(net225));
 sg13g2_nand2_1 _12944_ (.Y(_05067_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ),
    .B(net279));
 sg13g2_o21ai_1 _12945_ (.B1(_05067_),
    .Y(_00784_),
    .A1(net130),
    .A2(_05060_));
 sg13g2_nand2_1 _12946_ (.Y(_05068_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ),
    .B(net279));
 sg13g2_o21ai_1 _12947_ (.B1(_05068_),
    .Y(_00785_),
    .A1(net85),
    .A2(_05060_));
 sg13g2_nand2_1 _12948_ (.Y(_05069_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ),
    .B(net279));
 sg13g2_o21ai_1 _12949_ (.B1(_05069_),
    .Y(_00786_),
    .A1(net121),
    .A2(net225));
 sg13g2_nand2_1 _12950_ (.Y(_05070_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ),
    .B(net279));
 sg13g2_o21ai_1 _12951_ (.B1(_05070_),
    .Y(_00787_),
    .A1(net97),
    .A2(net225));
 sg13g2_buf_1 _12952_ (.A(_05058_),
    .X(_05071_));
 sg13g2_nand2_1 _12953_ (.Y(_05072_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ),
    .B(_05071_));
 sg13g2_o21ai_1 _12954_ (.B1(_05072_),
    .Y(_00788_),
    .A1(net120),
    .A2(net225));
 sg13g2_nand2_1 _12955_ (.Y(_05073_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ),
    .B(_05071_));
 sg13g2_o21ai_1 _12956_ (.B1(_05073_),
    .Y(_00789_),
    .A1(net124),
    .A2(net225));
 sg13g2_mux2_1 _12957_ (.A0(net96),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ),
    .S(_05064_),
    .X(_00790_));
 sg13g2_buf_1 _12958_ (.A(net280),
    .X(_05074_));
 sg13g2_nand2_1 _12959_ (.Y(_05075_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ),
    .B(net277));
 sg13g2_o21ai_1 _12960_ (.B1(_05075_),
    .Y(_00791_),
    .A1(_04609_),
    .A2(net224));
 sg13g2_nand2_1 _12961_ (.Y(_05076_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ),
    .B(net277));
 sg13g2_o21ai_1 _12962_ (.B1(_05076_),
    .Y(_00792_),
    .A1(net112),
    .A2(net224));
 sg13g2_nand2_1 _12963_ (.Y(_05077_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ),
    .B(net277));
 sg13g2_o21ai_1 _12964_ (.B1(_05077_),
    .Y(_00793_),
    .A1(net122),
    .A2(net224));
 sg13g2_nand2_1 _12965_ (.Y(_05078_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ),
    .B(net277));
 sg13g2_o21ai_1 _12966_ (.B1(_05078_),
    .Y(_00794_),
    .A1(_04060_),
    .A2(net224));
 sg13g2_mux2_1 _12967_ (.A0(_04619_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ),
    .S(net278),
    .X(_00795_));
 sg13g2_nand2_1 _12968_ (.Y(_05079_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ),
    .B(net277));
 sg13g2_o21ai_1 _12969_ (.B1(_05079_),
    .Y(_00796_),
    .A1(_04626_),
    .A2(net224));
 sg13g2_nand2_1 _12970_ (.Y(_05080_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ),
    .B(net277));
 sg13g2_o21ai_1 _12971_ (.B1(_05080_),
    .Y(_00797_),
    .A1(_04632_),
    .A2(net224));
 sg13g2_nand2_1 _12972_ (.Y(_05081_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ),
    .B(net277));
 sg13g2_o21ai_1 _12973_ (.B1(_05081_),
    .Y(_00798_),
    .A1(net88),
    .A2(_05074_));
 sg13g2_nand2_1 _12974_ (.Y(_05082_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ),
    .B(net277));
 sg13g2_o21ai_1 _12975_ (.B1(_05082_),
    .Y(_00799_),
    .A1(net111),
    .A2(net224));
 sg13g2_nand2_1 _12976_ (.Y(_05083_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ),
    .B(net280));
 sg13g2_o21ai_1 _12977_ (.B1(_05083_),
    .Y(_00800_),
    .A1(net106),
    .A2(net224));
 sg13g2_nand2_1 _12978_ (.Y(_05084_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ),
    .B(net280));
 sg13g2_o21ai_1 _12979_ (.B1(_05084_),
    .Y(_00801_),
    .A1(net113),
    .A2(_05074_));
 sg13g2_nand2_1 _12980_ (.Y(_05085_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ),
    .B(net280));
 sg13g2_o21ai_1 _12981_ (.B1(_05085_),
    .Y(_00802_),
    .A1(_03625_),
    .A2(net278));
 sg13g2_nand2_1 _12982_ (.Y(_05086_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ),
    .B(net280));
 sg13g2_o21ai_1 _12983_ (.B1(_05086_),
    .Y(_00803_),
    .A1(net118),
    .A2(net278));
 sg13g2_nand2_1 _12984_ (.Y(_05087_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ),
    .B(net280));
 sg13g2_o21ai_1 _12985_ (.B1(_05087_),
    .Y(_00804_),
    .A1(net119),
    .A2(net278));
 sg13g2_nand2_1 _12986_ (.Y(_05088_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ),
    .B(net280));
 sg13g2_o21ai_1 _12987_ (.B1(_05088_),
    .Y(_00805_),
    .A1(net123),
    .A2(net278));
 sg13g2_nand2_1 _12988_ (.Y(_05089_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ),
    .B(_05059_));
 sg13g2_o21ai_1 _12989_ (.B1(_05089_),
    .Y(_00806_),
    .A1(_04660_),
    .A2(net278));
 sg13g2_nand2_1 _12990_ (.Y(_05090_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ),
    .B(_05059_));
 sg13g2_o21ai_1 _12991_ (.B1(_05090_),
    .Y(_00807_),
    .A1(net101),
    .A2(net278));
 sg13g2_mux2_1 _12992_ (.A0(net100),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ),
    .S(_05061_),
    .X(_00808_));
 sg13g2_mux2_1 _12993_ (.A0(net128),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ),
    .S(_05061_),
    .X(_00809_));
 sg13g2_nand3_1 _12994_ (.B(net625),
    .C(_04988_),
    .A(net626),
    .Y(_05091_));
 sg13g2_buf_1 _12995_ (.A(_05091_),
    .X(_05092_));
 sg13g2_buf_1 _12996_ (.A(_05092_),
    .X(_05093_));
 sg13g2_buf_1 _12997_ (.A(net276),
    .X(_05094_));
 sg13g2_buf_1 _12998_ (.A(_05092_),
    .X(_05095_));
 sg13g2_nand2_1 _12999_ (.Y(_05096_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ),
    .B(net275));
 sg13g2_o21ai_1 _13000_ (.B1(_05096_),
    .Y(_00810_),
    .A1(_04549_),
    .A2(net223));
 sg13g2_nand2_1 _13001_ (.Y(_05097_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ),
    .B(net275));
 sg13g2_o21ai_1 _13002_ (.B1(_05097_),
    .Y(_00811_),
    .A1(net117),
    .A2(net223));
 sg13g2_buf_1 _13003_ (.A(_05092_),
    .X(_05098_));
 sg13g2_mux2_1 _13004_ (.A0(net129),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ),
    .S(_05098_),
    .X(_00812_));
 sg13g2_nand2_1 _13005_ (.Y(_05099_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ),
    .B(net275));
 sg13g2_o21ai_1 _13006_ (.B1(_05099_),
    .Y(_00813_),
    .A1(net131),
    .A2(net223));
 sg13g2_mux2_1 _13007_ (.A0(net99),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ),
    .S(net274),
    .X(_00814_));
 sg13g2_nand2_1 _13008_ (.Y(_05100_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ),
    .B(net275));
 sg13g2_o21ai_1 _13009_ (.B1(_05100_),
    .Y(_00815_),
    .A1(net98),
    .A2(net223));
 sg13g2_nand2_1 _13010_ (.Y(_05101_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ),
    .B(net275));
 sg13g2_o21ai_1 _13011_ (.B1(_05101_),
    .Y(_00816_),
    .A1(net130),
    .A2(_05094_));
 sg13g2_nand2_1 _13012_ (.Y(_05102_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ),
    .B(net275));
 sg13g2_o21ai_1 _13013_ (.B1(_05102_),
    .Y(_00817_),
    .A1(net85),
    .A2(_05094_));
 sg13g2_nand2_1 _13014_ (.Y(_05103_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ),
    .B(net275));
 sg13g2_o21ai_1 _13015_ (.B1(_05103_),
    .Y(_00818_),
    .A1(net121),
    .A2(net223));
 sg13g2_nand2_1 _13016_ (.Y(_05104_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ),
    .B(net275));
 sg13g2_o21ai_1 _13017_ (.B1(_05104_),
    .Y(_00819_),
    .A1(net97),
    .A2(net223));
 sg13g2_buf_1 _13018_ (.A(_05092_),
    .X(_05105_));
 sg13g2_nand2_1 _13019_ (.Y(_05106_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ),
    .B(_05105_));
 sg13g2_o21ai_1 _13020_ (.B1(_05106_),
    .Y(_00820_),
    .A1(net120),
    .A2(net223));
 sg13g2_nand2_1 _13021_ (.Y(_05107_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ),
    .B(_05105_));
 sg13g2_o21ai_1 _13022_ (.B1(_05107_),
    .Y(_00821_),
    .A1(net124),
    .A2(net223));
 sg13g2_mux2_1 _13023_ (.A0(net96),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ),
    .S(_05098_),
    .X(_00822_));
 sg13g2_buf_1 _13024_ (.A(net276),
    .X(_05108_));
 sg13g2_nand2_1 _13025_ (.Y(_05109_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ),
    .B(net273));
 sg13g2_o21ai_1 _13026_ (.B1(_05109_),
    .Y(_00823_),
    .A1(_04609_),
    .A2(net222));
 sg13g2_nand2_1 _13027_ (.Y(_05110_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ),
    .B(net273));
 sg13g2_o21ai_1 _13028_ (.B1(_05110_),
    .Y(_00824_),
    .A1(net112),
    .A2(net222));
 sg13g2_nand2_1 _13029_ (.Y(_05111_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ),
    .B(net273));
 sg13g2_o21ai_1 _13030_ (.B1(_05111_),
    .Y(_00825_),
    .A1(net122),
    .A2(net222));
 sg13g2_nand2_1 _13031_ (.Y(_05112_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ),
    .B(net273));
 sg13g2_o21ai_1 _13032_ (.B1(_05112_),
    .Y(_00826_),
    .A1(_04060_),
    .A2(net222));
 sg13g2_mux2_1 _13033_ (.A0(_04619_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ),
    .S(net274),
    .X(_00827_));
 sg13g2_nand2_1 _13034_ (.Y(_05113_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ),
    .B(net273));
 sg13g2_o21ai_1 _13035_ (.B1(_05113_),
    .Y(_00828_),
    .A1(_04626_),
    .A2(net222));
 sg13g2_nand2_1 _13036_ (.Y(_05114_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ),
    .B(net273));
 sg13g2_o21ai_1 _13037_ (.B1(_05114_),
    .Y(_00829_),
    .A1(_04632_),
    .A2(net222));
 sg13g2_nand2_1 _13038_ (.Y(_05115_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ),
    .B(net273));
 sg13g2_o21ai_1 _13039_ (.B1(_05115_),
    .Y(_00830_),
    .A1(net88),
    .A2(_05108_));
 sg13g2_nand2_1 _13040_ (.Y(_05116_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ),
    .B(net273));
 sg13g2_o21ai_1 _13041_ (.B1(_05116_),
    .Y(_00831_),
    .A1(net111),
    .A2(net222));
 sg13g2_nand2_1 _13042_ (.Y(_05117_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ),
    .B(net276));
 sg13g2_o21ai_1 _13043_ (.B1(_05117_),
    .Y(_00832_),
    .A1(net106),
    .A2(net222));
 sg13g2_nand2_1 _13044_ (.Y(_05118_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ),
    .B(net276));
 sg13g2_o21ai_1 _13045_ (.B1(_05118_),
    .Y(_00833_),
    .A1(net113),
    .A2(_05108_));
 sg13g2_nand2_1 _13046_ (.Y(_05119_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ),
    .B(net276));
 sg13g2_o21ai_1 _13047_ (.B1(_05119_),
    .Y(_00834_),
    .A1(_03625_),
    .A2(net274));
 sg13g2_nand2_1 _13048_ (.Y(_05120_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ),
    .B(net276));
 sg13g2_o21ai_1 _13049_ (.B1(_05120_),
    .Y(_00835_),
    .A1(net118),
    .A2(net274));
 sg13g2_nand2_1 _13050_ (.Y(_05121_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ),
    .B(net276));
 sg13g2_o21ai_1 _13051_ (.B1(_05121_),
    .Y(_00836_),
    .A1(net119),
    .A2(net274));
 sg13g2_nand2_1 _13052_ (.Y(_05122_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ),
    .B(net276));
 sg13g2_o21ai_1 _13053_ (.B1(_05122_),
    .Y(_00837_),
    .A1(net123),
    .A2(net274));
 sg13g2_nand2_1 _13054_ (.Y(_05123_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ),
    .B(_05093_));
 sg13g2_o21ai_1 _13055_ (.B1(_05123_),
    .Y(_00838_),
    .A1(_04660_),
    .A2(net274));
 sg13g2_nand2_1 _13056_ (.Y(_05124_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ),
    .B(_05093_));
 sg13g2_o21ai_1 _13057_ (.B1(_05124_),
    .Y(_00839_),
    .A1(net101),
    .A2(net274));
 sg13g2_mux2_1 _13058_ (.A0(net100),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ),
    .S(_05095_),
    .X(_00840_));
 sg13g2_mux2_1 _13059_ (.A0(net128),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ),
    .S(_05095_),
    .X(_00841_));
 sg13g2_nand2_1 _13060_ (.Y(_05125_),
    .A(_04554_),
    .B(_04677_));
 sg13g2_buf_1 _13061_ (.A(_05125_),
    .X(_05126_));
 sg13g2_buf_1 _13062_ (.A(_05126_),
    .X(_05127_));
 sg13g2_buf_1 _13063_ (.A(net221),
    .X(_05128_));
 sg13g2_buf_1 _13064_ (.A(_05126_),
    .X(_05129_));
 sg13g2_nand2_1 _13065_ (.Y(_05130_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ),
    .B(net220));
 sg13g2_o21ai_1 _13066_ (.B1(_05130_),
    .Y(_00842_),
    .A1(_04549_),
    .A2(net191));
 sg13g2_nand2_1 _13067_ (.Y(_05131_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ),
    .B(net220));
 sg13g2_o21ai_1 _13068_ (.B1(_05131_),
    .Y(_00843_),
    .A1(net117),
    .A2(net191));
 sg13g2_buf_1 _13069_ (.A(_05126_),
    .X(_05132_));
 sg13g2_mux2_1 _13070_ (.A0(net129),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ),
    .S(net219),
    .X(_00844_));
 sg13g2_nand2_1 _13071_ (.Y(_05133_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ),
    .B(net220));
 sg13g2_o21ai_1 _13072_ (.B1(_05133_),
    .Y(_00845_),
    .A1(net131),
    .A2(net191));
 sg13g2_mux2_1 _13073_ (.A0(net99),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ),
    .S(net219),
    .X(_00846_));
 sg13g2_nand2_1 _13074_ (.Y(_05134_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ),
    .B(net220));
 sg13g2_o21ai_1 _13075_ (.B1(_05134_),
    .Y(_00847_),
    .A1(net98),
    .A2(net191));
 sg13g2_nand2_1 _13076_ (.Y(_05135_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ),
    .B(net220));
 sg13g2_o21ai_1 _13077_ (.B1(_05135_),
    .Y(_00848_),
    .A1(net130),
    .A2(_05128_));
 sg13g2_nand2_1 _13078_ (.Y(_05136_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ),
    .B(net220));
 sg13g2_o21ai_1 _13079_ (.B1(_05136_),
    .Y(_00849_),
    .A1(net85),
    .A2(_05128_));
 sg13g2_nand2_1 _13080_ (.Y(_05137_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ),
    .B(net220));
 sg13g2_o21ai_1 _13081_ (.B1(_05137_),
    .Y(_00850_),
    .A1(net121),
    .A2(net191));
 sg13g2_nand2_1 _13082_ (.Y(_05138_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ),
    .B(net220));
 sg13g2_o21ai_1 _13083_ (.B1(_05138_),
    .Y(_00851_),
    .A1(net97),
    .A2(net191));
 sg13g2_buf_1 _13084_ (.A(_05126_),
    .X(_05139_));
 sg13g2_nand2_1 _13085_ (.Y(_05140_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ),
    .B(_05139_));
 sg13g2_o21ai_1 _13086_ (.B1(_05140_),
    .Y(_00852_),
    .A1(net120),
    .A2(net191));
 sg13g2_nand2_1 _13087_ (.Y(_05141_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ),
    .B(_05139_));
 sg13g2_o21ai_1 _13088_ (.B1(_05141_),
    .Y(_00853_),
    .A1(net124),
    .A2(net191));
 sg13g2_mux2_1 _13089_ (.A0(net96),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ),
    .S(_05132_),
    .X(_00854_));
 sg13g2_buf_1 _13090_ (.A(net221),
    .X(_05142_));
 sg13g2_nand2_1 _13091_ (.Y(_05143_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ),
    .B(net218));
 sg13g2_o21ai_1 _13092_ (.B1(_05143_),
    .Y(_00855_),
    .A1(_04609_),
    .A2(_05142_));
 sg13g2_nand2_1 _13093_ (.Y(_05144_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ),
    .B(net218));
 sg13g2_o21ai_1 _13094_ (.B1(_05144_),
    .Y(_00856_),
    .A1(net112),
    .A2(net190));
 sg13g2_nand2_1 _13095_ (.Y(_05145_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ),
    .B(net218));
 sg13g2_o21ai_1 _13096_ (.B1(_05145_),
    .Y(_00857_),
    .A1(net122),
    .A2(net190));
 sg13g2_nand2_1 _13097_ (.Y(_05146_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ),
    .B(net218));
 sg13g2_o21ai_1 _13098_ (.B1(_05146_),
    .Y(_00858_),
    .A1(_04060_),
    .A2(net190));
 sg13g2_mux2_1 _13099_ (.A0(_04619_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ),
    .S(net219),
    .X(_00859_));
 sg13g2_nand2_1 _13100_ (.Y(_05147_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ),
    .B(net218));
 sg13g2_o21ai_1 _13101_ (.B1(_05147_),
    .Y(_00860_),
    .A1(_04626_),
    .A2(net190));
 sg13g2_nand2_1 _13102_ (.Y(_05148_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ),
    .B(net218));
 sg13g2_o21ai_1 _13103_ (.B1(_05148_),
    .Y(_00861_),
    .A1(_04632_),
    .A2(net190));
 sg13g2_nand2_1 _13104_ (.Y(_05149_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ),
    .B(net218));
 sg13g2_o21ai_1 _13105_ (.B1(_05149_),
    .Y(_00862_),
    .A1(net88),
    .A2(net190));
 sg13g2_nand2_1 _13106_ (.Y(_05150_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ),
    .B(net218));
 sg13g2_o21ai_1 _13107_ (.B1(_05150_),
    .Y(_00863_),
    .A1(net111),
    .A2(net190));
 sg13g2_nand2_1 _13108_ (.Y(_05151_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ),
    .B(net221));
 sg13g2_o21ai_1 _13109_ (.B1(_05151_),
    .Y(_00864_),
    .A1(net106),
    .A2(net190));
 sg13g2_nand2_1 _13110_ (.Y(_05152_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ),
    .B(net221));
 sg13g2_o21ai_1 _13111_ (.B1(_05152_),
    .Y(_00865_),
    .A1(net113),
    .A2(_05142_));
 sg13g2_nand2_1 _13112_ (.Y(_05153_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ),
    .B(net221));
 sg13g2_o21ai_1 _13113_ (.B1(_05153_),
    .Y(_00866_),
    .A1(_03625_),
    .A2(net219));
 sg13g2_nand2_1 _13114_ (.Y(_05154_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ),
    .B(net221));
 sg13g2_o21ai_1 _13115_ (.B1(_05154_),
    .Y(_00867_),
    .A1(net118),
    .A2(net219));
 sg13g2_nand2_1 _13116_ (.Y(_05155_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ),
    .B(net221));
 sg13g2_o21ai_1 _13117_ (.B1(_05155_),
    .Y(_00868_),
    .A1(net119),
    .A2(net219));
 sg13g2_nand2_1 _13118_ (.Y(_05156_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ),
    .B(net221));
 sg13g2_o21ai_1 _13119_ (.B1(_05156_),
    .Y(_00869_),
    .A1(net123),
    .A2(net219));
 sg13g2_nand2_1 _13120_ (.Y(_05157_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ),
    .B(_05127_));
 sg13g2_o21ai_1 _13121_ (.B1(_05157_),
    .Y(_00870_),
    .A1(_04660_),
    .A2(net219));
 sg13g2_nand2_1 _13122_ (.Y(_05158_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ),
    .B(_05127_));
 sg13g2_o21ai_1 _13123_ (.B1(_05158_),
    .Y(_00871_),
    .A1(net101),
    .A2(_05132_));
 sg13g2_mux2_1 _13124_ (.A0(net100),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ),
    .S(_05129_),
    .X(_00872_));
 sg13g2_mux2_1 _13125_ (.A0(_03888_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ),
    .S(_05129_),
    .X(_00873_));
 sg13g2_nand2_1 _13126_ (.Y(_05159_),
    .A(_04677_),
    .B(_04783_));
 sg13g2_buf_1 _13127_ (.A(_05159_),
    .X(_05160_));
 sg13g2_buf_1 _13128_ (.A(_05160_),
    .X(_05161_));
 sg13g2_buf_1 _13129_ (.A(net217),
    .X(_05162_));
 sg13g2_buf_1 _13130_ (.A(_05160_),
    .X(_05163_));
 sg13g2_nand2_1 _13131_ (.Y(_05164_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ),
    .B(net216));
 sg13g2_o21ai_1 _13132_ (.B1(_05164_),
    .Y(_00874_),
    .A1(_04549_),
    .A2(net189));
 sg13g2_nand2_1 _13133_ (.Y(_05165_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ),
    .B(net216));
 sg13g2_o21ai_1 _13134_ (.B1(_05165_),
    .Y(_00875_),
    .A1(net117),
    .A2(net189));
 sg13g2_buf_1 _13135_ (.A(_05160_),
    .X(_05166_));
 sg13g2_mux2_1 _13136_ (.A0(net129),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ),
    .S(net215),
    .X(_00876_));
 sg13g2_nand2_1 _13137_ (.Y(_05167_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ),
    .B(net216));
 sg13g2_o21ai_1 _13138_ (.B1(_05167_),
    .Y(_00877_),
    .A1(_03917_),
    .A2(net189));
 sg13g2_mux2_1 _13139_ (.A0(net99),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ),
    .S(net215),
    .X(_00878_));
 sg13g2_nand2_1 _13140_ (.Y(_05168_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ),
    .B(net216));
 sg13g2_o21ai_1 _13141_ (.B1(_05168_),
    .Y(_00879_),
    .A1(net98),
    .A2(net189));
 sg13g2_nand2_1 _13142_ (.Y(_05169_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ),
    .B(net216));
 sg13g2_o21ai_1 _13143_ (.B1(_05169_),
    .Y(_00880_),
    .A1(net130),
    .A2(_05162_));
 sg13g2_nand2_1 _13144_ (.Y(_05170_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ),
    .B(net216));
 sg13g2_o21ai_1 _13145_ (.B1(_05170_),
    .Y(_00881_),
    .A1(net85),
    .A2(_05162_));
 sg13g2_nand2_1 _13146_ (.Y(_05171_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ),
    .B(net216));
 sg13g2_o21ai_1 _13147_ (.B1(_05171_),
    .Y(_00882_),
    .A1(net121),
    .A2(net189));
 sg13g2_nand2_1 _13148_ (.Y(_05172_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ),
    .B(net216));
 sg13g2_o21ai_1 _13149_ (.B1(_05172_),
    .Y(_00883_),
    .A1(net97),
    .A2(net189));
 sg13g2_buf_1 _13150_ (.A(_05160_),
    .X(_05173_));
 sg13g2_nand2_1 _13151_ (.Y(_05174_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ),
    .B(_05173_));
 sg13g2_o21ai_1 _13152_ (.B1(_05174_),
    .Y(_00884_),
    .A1(net120),
    .A2(net189));
 sg13g2_nand2_1 _13153_ (.Y(_05175_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ),
    .B(_05173_));
 sg13g2_o21ai_1 _13154_ (.B1(_05175_),
    .Y(_00885_),
    .A1(net124),
    .A2(net189));
 sg13g2_mux2_1 _13155_ (.A0(net96),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ),
    .S(_05166_),
    .X(_00886_));
 sg13g2_buf_1 _13156_ (.A(net217),
    .X(_05176_));
 sg13g2_nand2_1 _13157_ (.Y(_05177_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ),
    .B(net214));
 sg13g2_o21ai_1 _13158_ (.B1(_05177_),
    .Y(_00887_),
    .A1(_04609_),
    .A2(net188));
 sg13g2_nand2_1 _13159_ (.Y(_05178_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ),
    .B(net214));
 sg13g2_o21ai_1 _13160_ (.B1(_05178_),
    .Y(_00888_),
    .A1(net112),
    .A2(net188));
 sg13g2_nand2_1 _13161_ (.Y(_05179_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ),
    .B(net214));
 sg13g2_o21ai_1 _13162_ (.B1(_05179_),
    .Y(_00889_),
    .A1(net122),
    .A2(net188));
 sg13g2_nand2_1 _13163_ (.Y(_05180_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ),
    .B(net214));
 sg13g2_o21ai_1 _13164_ (.B1(_05180_),
    .Y(_00890_),
    .A1(_04060_),
    .A2(net188));
 sg13g2_mux2_1 _13165_ (.A0(_04619_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ),
    .S(net215),
    .X(_00891_));
 sg13g2_nand2_1 _13166_ (.Y(_05181_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ),
    .B(net214));
 sg13g2_o21ai_1 _13167_ (.B1(_05181_),
    .Y(_00892_),
    .A1(_04626_),
    .A2(net188));
 sg13g2_nand2_1 _13168_ (.Y(_05182_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ),
    .B(net214));
 sg13g2_o21ai_1 _13169_ (.B1(_05182_),
    .Y(_00893_),
    .A1(_04632_),
    .A2(net188));
 sg13g2_nand2_1 _13170_ (.Y(_05183_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ),
    .B(net214));
 sg13g2_o21ai_1 _13171_ (.B1(_05183_),
    .Y(_00894_),
    .A1(net88),
    .A2(_05176_));
 sg13g2_nand2_1 _13172_ (.Y(_05184_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ),
    .B(net214));
 sg13g2_o21ai_1 _13173_ (.B1(_05184_),
    .Y(_00895_),
    .A1(net111),
    .A2(net188));
 sg13g2_nand2_1 _13174_ (.Y(_05185_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ),
    .B(net217));
 sg13g2_o21ai_1 _13175_ (.B1(_05185_),
    .Y(_00896_),
    .A1(net106),
    .A2(net188));
 sg13g2_nand2_1 _13176_ (.Y(_05186_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ),
    .B(net217));
 sg13g2_o21ai_1 _13177_ (.B1(_05186_),
    .Y(_00897_),
    .A1(net113),
    .A2(_05176_));
 sg13g2_nand2_1 _13178_ (.Y(_05187_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ),
    .B(net217));
 sg13g2_o21ai_1 _13179_ (.B1(_05187_),
    .Y(_00898_),
    .A1(_03625_),
    .A2(net215));
 sg13g2_nand2_1 _13180_ (.Y(_05188_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ),
    .B(net217));
 sg13g2_o21ai_1 _13181_ (.B1(_05188_),
    .Y(_00899_),
    .A1(net118),
    .A2(net215));
 sg13g2_nand2_1 _13182_ (.Y(_05189_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ),
    .B(net217));
 sg13g2_o21ai_1 _13183_ (.B1(_05189_),
    .Y(_00900_),
    .A1(net119),
    .A2(net215));
 sg13g2_nand2_1 _13184_ (.Y(_05190_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ),
    .B(net217));
 sg13g2_o21ai_1 _13185_ (.B1(_05190_),
    .Y(_00901_),
    .A1(net123),
    .A2(net215));
 sg13g2_nand2_1 _13186_ (.Y(_05191_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ),
    .B(_05161_));
 sg13g2_o21ai_1 _13187_ (.B1(_05191_),
    .Y(_00902_),
    .A1(_04660_),
    .A2(net215));
 sg13g2_nand2_1 _13188_ (.Y(_05192_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ),
    .B(_05161_));
 sg13g2_o21ai_1 _13189_ (.B1(_05192_),
    .Y(_00903_),
    .A1(net101),
    .A2(_05166_));
 sg13g2_mux2_1 _13190_ (.A0(net100),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ),
    .S(_05163_),
    .X(_00904_));
 sg13g2_mux2_1 _13191_ (.A0(net128),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ),
    .S(_05163_),
    .X(_00905_));
 sg13g2_buf_1 _13192_ (.A(net333),
    .X(_05193_));
 sg13g2_buf_1 _13193_ (.A(\soc_I.qqspi_I.spi_buf[0] ),
    .X(_05194_));
 sg13g2_nor3_1 _13194_ (.A(_04318_),
    .B(_04327_),
    .C(_04336_),
    .Y(_05195_));
 sg13g2_buf_1 _13195_ (.A(_05195_),
    .X(_05196_));
 sg13g2_buf_1 _13196_ (.A(_05196_),
    .X(_05197_));
 sg13g2_buf_1 _13197_ (.A(net66),
    .X(_05198_));
 sg13g2_buf_1 _13198_ (.A(net66),
    .X(_05199_));
 sg13g2_buf_1 _13199_ (.A(\soc_I.qqspi_I.spi_buf[24] ),
    .X(_05200_));
 sg13g2_nor2b_1 _13200_ (.A(net63),
    .B_N(_05200_),
    .Y(_05201_));
 sg13g2_a21oi_1 _13201_ (.A1(_05194_),
    .A2(net64),
    .Y(_05202_),
    .B1(_05201_));
 sg13g2_buf_1 _13202_ (.A(_04361_),
    .X(_05203_));
 sg13g2_nand2_1 _13203_ (.Y(_05204_),
    .A(\soc_I.qqspi_I.rdata[0] ),
    .B(net332));
 sg13g2_o21ai_1 _13204_ (.B1(_05204_),
    .Y(_00927_),
    .A1(net322),
    .A2(_05202_));
 sg13g2_buf_1 _13205_ (.A(\soc_I.qqspi_I.spi_buf[10] ),
    .X(_05205_));
 sg13g2_buf_1 _13206_ (.A(\soc_I.qqspi_I.spi_buf[18] ),
    .X(_05206_));
 sg13g2_nor2b_1 _13207_ (.A(net63),
    .B_N(_05206_),
    .Y(_05207_));
 sg13g2_a21oi_1 _13208_ (.A1(_05205_),
    .A2(net64),
    .Y(_05208_),
    .B1(_05207_));
 sg13g2_nand2_1 _13209_ (.Y(_05209_),
    .A(\soc_I.qqspi_I.rdata[10] ),
    .B(net332));
 sg13g2_o21ai_1 _13210_ (.B1(_05209_),
    .Y(_00928_),
    .A1(net322),
    .A2(_05208_));
 sg13g2_buf_1 _13211_ (.A(\soc_I.qqspi_I.spi_buf[11] ),
    .X(_05210_));
 sg13g2_buf_1 _13212_ (.A(\soc_I.qqspi_I.spi_buf[19] ),
    .X(_05211_));
 sg13g2_nor2b_1 _13213_ (.A(net63),
    .B_N(_05211_),
    .Y(_05212_));
 sg13g2_a21oi_1 _13214_ (.A1(_05210_),
    .A2(net64),
    .Y(_05213_),
    .B1(_05212_));
 sg13g2_nand2_1 _13215_ (.Y(_05214_),
    .A(\soc_I.qqspi_I.rdata[11] ),
    .B(_05203_));
 sg13g2_o21ai_1 _13216_ (.B1(_05214_),
    .Y(_00929_),
    .A1(net322),
    .A2(_05213_));
 sg13g2_buf_1 _13217_ (.A(\soc_I.qqspi_I.spi_buf[12] ),
    .X(_05215_));
 sg13g2_buf_1 _13218_ (.A(\soc_I.qqspi_I.spi_buf[20] ),
    .X(_05216_));
 sg13g2_nor2b_1 _13219_ (.A(net63),
    .B_N(_05216_),
    .Y(_05217_));
 sg13g2_a21oi_1 _13220_ (.A1(_05215_),
    .A2(_05198_),
    .Y(_05218_),
    .B1(_05217_));
 sg13g2_nand2_1 _13221_ (.Y(_05219_),
    .A(\soc_I.qqspi_I.rdata[12] ),
    .B(_05203_));
 sg13g2_o21ai_1 _13222_ (.B1(_05219_),
    .Y(_00930_),
    .A1(_05193_),
    .A2(_05218_));
 sg13g2_buf_1 _13223_ (.A(\soc_I.qqspi_I.spi_buf[13] ),
    .X(_05220_));
 sg13g2_buf_1 _13224_ (.A(\soc_I.qqspi_I.spi_buf[21] ),
    .X(_05221_));
 sg13g2_nor2b_1 _13225_ (.A(net63),
    .B_N(_05221_),
    .Y(_05222_));
 sg13g2_a21oi_1 _13226_ (.A1(_05220_),
    .A2(net64),
    .Y(_05223_),
    .B1(_05222_));
 sg13g2_nand2_1 _13227_ (.Y(_05224_),
    .A(\soc_I.qqspi_I.rdata[13] ),
    .B(net332));
 sg13g2_o21ai_1 _13228_ (.B1(_05224_),
    .Y(_00931_),
    .A1(net322),
    .A2(_05223_));
 sg13g2_buf_1 _13229_ (.A(\soc_I.qqspi_I.spi_buf[14] ),
    .X(_05225_));
 sg13g2_buf_1 _13230_ (.A(\soc_I.qqspi_I.spi_buf[22] ),
    .X(_05226_));
 sg13g2_nor2b_1 _13231_ (.A(net63),
    .B_N(_05226_),
    .Y(_05227_));
 sg13g2_a21oi_1 _13232_ (.A1(_05225_),
    .A2(net64),
    .Y(_05228_),
    .B1(_05227_));
 sg13g2_nand2_1 _13233_ (.Y(_05229_),
    .A(\soc_I.qqspi_I.rdata[14] ),
    .B(net332));
 sg13g2_o21ai_1 _13234_ (.B1(_05229_),
    .Y(_00932_),
    .A1(net322),
    .A2(_05228_));
 sg13g2_buf_1 _13235_ (.A(\soc_I.qqspi_I.spi_buf[15] ),
    .X(_05230_));
 sg13g2_buf_1 _13236_ (.A(\soc_I.qqspi_I.spi_buf[23] ),
    .X(_05231_));
 sg13g2_nor2b_1 _13237_ (.A(_05199_),
    .B_N(_05231_),
    .Y(_05232_));
 sg13g2_a21oi_1 _13238_ (.A1(_05230_),
    .A2(_05198_),
    .Y(_05233_),
    .B1(_05232_));
 sg13g2_nand2_1 _13239_ (.Y(_05234_),
    .A(\soc_I.qqspi_I.rdata[15] ),
    .B(net332));
 sg13g2_o21ai_1 _13240_ (.B1(_05234_),
    .Y(_00933_),
    .A1(_05193_),
    .A2(_05233_));
 sg13g2_buf_1 _13241_ (.A(\soc_I.qqspi_I.spi_buf[16] ),
    .X(_05235_));
 sg13g2_buf_1 _13242_ (.A(net66),
    .X(_05236_));
 sg13g2_buf_1 _13243_ (.A(\soc_I.qqspi_I.spi_buf[8] ),
    .X(_05237_));
 sg13g2_nor2b_1 _13244_ (.A(_05236_),
    .B_N(_05237_),
    .Y(_05238_));
 sg13g2_a21oi_1 _13245_ (.A1(_05235_),
    .A2(net64),
    .Y(_05239_),
    .B1(_05238_));
 sg13g2_nand2_1 _13246_ (.Y(_05240_),
    .A(\soc_I.qqspi_I.rdata[16] ),
    .B(net332));
 sg13g2_o21ai_1 _13247_ (.B1(_05240_),
    .Y(_00934_),
    .A1(net322),
    .A2(_05239_));
 sg13g2_buf_1 _13248_ (.A(\soc_I.qqspi_I.spi_buf[17] ),
    .X(_05241_));
 sg13g2_buf_1 _13249_ (.A(\soc_I.qqspi_I.spi_buf[9] ),
    .X(_05242_));
 sg13g2_nor2b_1 _13250_ (.A(net62),
    .B_N(_05242_),
    .Y(_05243_));
 sg13g2_a21oi_1 _13251_ (.A1(_05241_),
    .A2(net64),
    .Y(_05244_),
    .B1(_05243_));
 sg13g2_buf_1 _13252_ (.A(net333),
    .X(_05245_));
 sg13g2_nand2_1 _13253_ (.Y(_05246_),
    .A(\soc_I.qqspi_I.rdata[17] ),
    .B(net321));
 sg13g2_o21ai_1 _13254_ (.B1(_05246_),
    .Y(_00935_),
    .A1(net322),
    .A2(_05244_));
 sg13g2_nor2b_1 _13255_ (.A(net62),
    .B_N(_05205_),
    .Y(_05247_));
 sg13g2_a21oi_1 _13256_ (.A1(_05206_),
    .A2(net64),
    .Y(_05248_),
    .B1(_05247_));
 sg13g2_nand2_1 _13257_ (.Y(_05249_),
    .A(\soc_I.qqspi_I.rdata[18] ),
    .B(net321));
 sg13g2_o21ai_1 _13258_ (.B1(_05249_),
    .Y(_00936_),
    .A1(net322),
    .A2(_05248_));
 sg13g2_buf_1 _13259_ (.A(net333),
    .X(_05250_));
 sg13g2_buf_1 _13260_ (.A(net66),
    .X(_05251_));
 sg13g2_nor2b_1 _13261_ (.A(net62),
    .B_N(_05210_),
    .Y(_05252_));
 sg13g2_a21oi_1 _13262_ (.A1(_05211_),
    .A2(net61),
    .Y(_05253_),
    .B1(_05252_));
 sg13g2_nand2_1 _13263_ (.Y(_05254_),
    .A(\soc_I.qqspi_I.rdata[19] ),
    .B(net321));
 sg13g2_o21ai_1 _13264_ (.B1(_05254_),
    .Y(_00937_),
    .A1(_05250_),
    .A2(_05253_));
 sg13g2_buf_1 _13265_ (.A(\soc_I.qqspi_I.spi_buf[1] ),
    .X(_05255_));
 sg13g2_buf_1 _13266_ (.A(\soc_I.qqspi_I.spi_buf[25] ),
    .X(_05256_));
 sg13g2_nor2b_1 _13267_ (.A(net62),
    .B_N(_05256_),
    .Y(_05257_));
 sg13g2_a21oi_1 _13268_ (.A1(_05255_),
    .A2(net61),
    .Y(_05258_),
    .B1(_05257_));
 sg13g2_nand2_1 _13269_ (.Y(_05259_),
    .A(\soc_I.qqspi_I.rdata[1] ),
    .B(net321));
 sg13g2_o21ai_1 _13270_ (.B1(_05259_),
    .Y(_00938_),
    .A1(net320),
    .A2(_05258_));
 sg13g2_nor2b_1 _13271_ (.A(net62),
    .B_N(_05215_),
    .Y(_05260_));
 sg13g2_a21oi_1 _13272_ (.A1(_05216_),
    .A2(net61),
    .Y(_05261_),
    .B1(_05260_));
 sg13g2_nand2_1 _13273_ (.Y(_05262_),
    .A(\soc_I.qqspi_I.rdata[20] ),
    .B(net321));
 sg13g2_o21ai_1 _13274_ (.B1(_05262_),
    .Y(_00939_),
    .A1(net320),
    .A2(_05261_));
 sg13g2_nor2b_1 _13275_ (.A(net62),
    .B_N(_05220_),
    .Y(_05263_));
 sg13g2_a21oi_1 _13276_ (.A1(_05221_),
    .A2(net61),
    .Y(_05264_),
    .B1(_05263_));
 sg13g2_nand2_1 _13277_ (.Y(_05265_),
    .A(\soc_I.qqspi_I.rdata[21] ),
    .B(_05245_));
 sg13g2_o21ai_1 _13278_ (.B1(_05265_),
    .Y(_00940_),
    .A1(_05250_),
    .A2(_05264_));
 sg13g2_nor2b_1 _13279_ (.A(net62),
    .B_N(_05225_),
    .Y(_05266_));
 sg13g2_a21oi_1 _13280_ (.A1(_05226_),
    .A2(_05251_),
    .Y(_05267_),
    .B1(_05266_));
 sg13g2_nand2_1 _13281_ (.Y(_05268_),
    .A(\soc_I.qqspi_I.rdata[22] ),
    .B(net321));
 sg13g2_o21ai_1 _13282_ (.B1(_05268_),
    .Y(_00941_),
    .A1(net320),
    .A2(_05267_));
 sg13g2_nor2b_1 _13283_ (.A(_05236_),
    .B_N(_05230_),
    .Y(_05269_));
 sg13g2_a21oi_1 _13284_ (.A1(_05231_),
    .A2(net61),
    .Y(_05270_),
    .B1(_05269_));
 sg13g2_nand2_1 _13285_ (.Y(_05271_),
    .A(\soc_I.qqspi_I.rdata[23] ),
    .B(_05245_));
 sg13g2_o21ai_1 _13286_ (.B1(_05271_),
    .Y(_00942_),
    .A1(net320),
    .A2(_05270_));
 sg13g2_nor2b_1 _13287_ (.A(net62),
    .B_N(_05194_),
    .Y(_05272_));
 sg13g2_a21oi_1 _13288_ (.A1(_05200_),
    .A2(_05251_),
    .Y(_05273_),
    .B1(_05272_));
 sg13g2_nand2_1 _13289_ (.Y(_05274_),
    .A(\soc_I.qqspi_I.rdata[24] ),
    .B(net321));
 sg13g2_o21ai_1 _13290_ (.B1(_05274_),
    .Y(_00943_),
    .A1(net320),
    .A2(_05273_));
 sg13g2_buf_1 _13291_ (.A(_05196_),
    .X(_05275_));
 sg13g2_nor2b_1 _13292_ (.A(net65),
    .B_N(_05255_),
    .Y(_05276_));
 sg13g2_a21oi_1 _13293_ (.A1(_05256_),
    .A2(net61),
    .Y(_05277_),
    .B1(_05276_));
 sg13g2_nand2_1 _13294_ (.Y(_05278_),
    .A(\soc_I.qqspi_I.rdata[25] ),
    .B(net321));
 sg13g2_o21ai_1 _13295_ (.B1(_05278_),
    .Y(_00944_),
    .A1(net320),
    .A2(_05277_));
 sg13g2_buf_1 _13296_ (.A(\soc_I.qqspi_I.spi_buf[26] ),
    .X(_05279_));
 sg13g2_buf_1 _13297_ (.A(\soc_I.qqspi_I.spi_buf[2] ),
    .X(_05280_));
 sg13g2_nor2b_1 _13298_ (.A(net65),
    .B_N(_05280_),
    .Y(_05281_));
 sg13g2_a21oi_1 _13299_ (.A1(_05279_),
    .A2(net61),
    .Y(_05282_),
    .B1(_05281_));
 sg13g2_buf_1 _13300_ (.A(net333),
    .X(_05283_));
 sg13g2_nand2_1 _13301_ (.Y(_05284_),
    .A(\soc_I.qqspi_I.rdata[26] ),
    .B(net319));
 sg13g2_o21ai_1 _13302_ (.B1(_05284_),
    .Y(_00945_),
    .A1(net320),
    .A2(_05282_));
 sg13g2_buf_1 _13303_ (.A(\soc_I.qqspi_I.spi_buf[27] ),
    .X(_05285_));
 sg13g2_buf_1 _13304_ (.A(\soc_I.qqspi_I.spi_buf[3] ),
    .X(_05286_));
 sg13g2_nor2b_1 _13305_ (.A(net65),
    .B_N(_05286_),
    .Y(_05287_));
 sg13g2_a21oi_1 _13306_ (.A1(_05285_),
    .A2(net61),
    .Y(_05288_),
    .B1(_05287_));
 sg13g2_nand2_1 _13307_ (.Y(_05289_),
    .A(\soc_I.qqspi_I.rdata[27] ),
    .B(_05283_));
 sg13g2_o21ai_1 _13308_ (.B1(_05289_),
    .Y(_00946_),
    .A1(net320),
    .A2(_05288_));
 sg13g2_buf_1 _13309_ (.A(net333),
    .X(_05290_));
 sg13g2_buf_1 _13310_ (.A(\soc_I.qqspi_I.spi_buf[28] ),
    .X(_05291_));
 sg13g2_buf_1 _13311_ (.A(net66),
    .X(_05292_));
 sg13g2_buf_1 _13312_ (.A(\soc_I.qqspi_I.spi_buf[4] ),
    .X(_05293_));
 sg13g2_nor2b_1 _13313_ (.A(_05275_),
    .B_N(_05293_),
    .Y(_05294_));
 sg13g2_a21oi_1 _13314_ (.A1(_05291_),
    .A2(net60),
    .Y(_05295_),
    .B1(_05294_));
 sg13g2_nand2_1 _13315_ (.Y(_05296_),
    .A(\soc_I.qqspi_I.rdata[28] ),
    .B(net319));
 sg13g2_o21ai_1 _13316_ (.B1(_05296_),
    .Y(_00947_),
    .A1(net318),
    .A2(_05295_));
 sg13g2_buf_1 _13317_ (.A(\soc_I.qqspi_I.spi_buf[29] ),
    .X(_05297_));
 sg13g2_buf_1 _13318_ (.A(\soc_I.qqspi_I.spi_buf[5] ),
    .X(_05298_));
 sg13g2_nor2b_1 _13319_ (.A(net65),
    .B_N(_05298_),
    .Y(_05299_));
 sg13g2_a21oi_1 _13320_ (.A1(_05297_),
    .A2(net60),
    .Y(_05300_),
    .B1(_05299_));
 sg13g2_nand2_1 _13321_ (.Y(_05301_),
    .A(\soc_I.qqspi_I.rdata[29] ),
    .B(net319));
 sg13g2_o21ai_1 _13322_ (.B1(_05301_),
    .Y(_00948_),
    .A1(net318),
    .A2(_05300_));
 sg13g2_nor2b_1 _13323_ (.A(net65),
    .B_N(_05279_),
    .Y(_05302_));
 sg13g2_a21oi_1 _13324_ (.A1(_05280_),
    .A2(net60),
    .Y(_05303_),
    .B1(_05302_));
 sg13g2_nand2_1 _13325_ (.Y(_05304_),
    .A(\soc_I.qqspi_I.rdata[2] ),
    .B(net319));
 sg13g2_o21ai_1 _13326_ (.B1(_05304_),
    .Y(_00949_),
    .A1(net318),
    .A2(_05303_));
 sg13g2_buf_1 _13327_ (.A(\soc_I.qqspi_I.spi_buf[30] ),
    .X(_05305_));
 sg13g2_buf_1 _13328_ (.A(\soc_I.qqspi_I.spi_buf[6] ),
    .X(_05306_));
 sg13g2_nor2b_1 _13329_ (.A(net65),
    .B_N(_05306_),
    .Y(_05307_));
 sg13g2_a21oi_1 _13330_ (.A1(_05305_),
    .A2(net60),
    .Y(_05308_),
    .B1(_05307_));
 sg13g2_nand2_1 _13331_ (.Y(_05309_),
    .A(\soc_I.qqspi_I.rdata[30] ),
    .B(net319));
 sg13g2_o21ai_1 _13332_ (.B1(_05309_),
    .Y(_00950_),
    .A1(net318),
    .A2(_05308_));
 sg13g2_buf_1 _13333_ (.A(\soc_I.qqspi_I.spi_buf[31] ),
    .X(_05310_));
 sg13g2_buf_1 _13334_ (.A(\soc_I.qqspi_I.spi_buf[7] ),
    .X(_05311_));
 sg13g2_nor2b_1 _13335_ (.A(net65),
    .B_N(_05311_),
    .Y(_05312_));
 sg13g2_a21oi_1 _13336_ (.A1(_05310_),
    .A2(net60),
    .Y(_05313_),
    .B1(_05312_));
 sg13g2_nand2_1 _13337_ (.Y(_05314_),
    .A(\soc_I.qqspi_I.rdata[31] ),
    .B(net319));
 sg13g2_o21ai_1 _13338_ (.B1(_05314_),
    .Y(_00951_),
    .A1(net318),
    .A2(_05313_));
 sg13g2_nor2b_1 _13339_ (.A(net65),
    .B_N(_05285_),
    .Y(_05315_));
 sg13g2_a21oi_1 _13340_ (.A1(_05286_),
    .A2(net60),
    .Y(_05316_),
    .B1(_05315_));
 sg13g2_nand2_1 _13341_ (.Y(_05317_),
    .A(\soc_I.qqspi_I.rdata[3] ),
    .B(_05283_));
 sg13g2_o21ai_1 _13342_ (.B1(_05317_),
    .Y(_00952_),
    .A1(net318),
    .A2(_05316_));
 sg13g2_nor2b_1 _13343_ (.A(_05275_),
    .B_N(_05291_),
    .Y(_05318_));
 sg13g2_a21oi_1 _13344_ (.A1(_05293_),
    .A2(_05292_),
    .Y(_05319_),
    .B1(_05318_));
 sg13g2_nand2_1 _13345_ (.Y(_05320_),
    .A(\soc_I.qqspi_I.rdata[4] ),
    .B(net319));
 sg13g2_o21ai_1 _13346_ (.B1(_05320_),
    .Y(_00953_),
    .A1(_05290_),
    .A2(_05319_));
 sg13g2_nor2b_1 _13347_ (.A(net66),
    .B_N(_05297_),
    .Y(_05321_));
 sg13g2_a21oi_1 _13348_ (.A1(_05298_),
    .A2(_05292_),
    .Y(_05322_),
    .B1(_05321_));
 sg13g2_nand2_1 _13349_ (.Y(_05323_),
    .A(\soc_I.qqspi_I.rdata[5] ),
    .B(net319));
 sg13g2_o21ai_1 _13350_ (.B1(_05323_),
    .Y(_00954_),
    .A1(_05290_),
    .A2(_05322_));
 sg13g2_nor2b_1 _13351_ (.A(net66),
    .B_N(_05305_),
    .Y(_05324_));
 sg13g2_a21oi_1 _13352_ (.A1(_05306_),
    .A2(net60),
    .Y(_05325_),
    .B1(_05324_));
 sg13g2_nand2_1 _13353_ (.Y(_05326_),
    .A(\soc_I.qqspi_I.rdata[6] ),
    .B(net333));
 sg13g2_o21ai_1 _13354_ (.B1(_05326_),
    .Y(_00955_),
    .A1(net318),
    .A2(_05325_));
 sg13g2_nor2b_1 _13355_ (.A(net66),
    .B_N(_05310_),
    .Y(_05327_));
 sg13g2_a21oi_1 _13356_ (.A1(_05311_),
    .A2(net60),
    .Y(_05328_),
    .B1(_05327_));
 sg13g2_nand2_1 _13357_ (.Y(_05329_),
    .A(\soc_I.qqspi_I.rdata[7] ),
    .B(net333));
 sg13g2_o21ai_1 _13358_ (.B1(_05329_),
    .Y(_00956_),
    .A1(net318),
    .A2(_05328_));
 sg13g2_nor2b_1 _13359_ (.A(_05197_),
    .B_N(_05235_),
    .Y(_05330_));
 sg13g2_a21oi_1 _13360_ (.A1(_05237_),
    .A2(net63),
    .Y(_05331_),
    .B1(_05330_));
 sg13g2_nand2_1 _13361_ (.Y(_05332_),
    .A(\soc_I.qqspi_I.rdata[8] ),
    .B(_04362_));
 sg13g2_o21ai_1 _13362_ (.B1(_05332_),
    .Y(_00957_),
    .A1(net332),
    .A2(_05331_));
 sg13g2_nor2b_1 _13363_ (.A(_05197_),
    .B_N(_05241_),
    .Y(_05333_));
 sg13g2_a21oi_1 _13364_ (.A1(_05242_),
    .A2(net63),
    .Y(_05334_),
    .B1(_05333_));
 sg13g2_nand2_1 _13365_ (.Y(_05335_),
    .A(\soc_I.qqspi_I.rdata[9] ),
    .B(net333));
 sg13g2_o21ai_1 _13366_ (.B1(_05335_),
    .Y(_00958_),
    .A1(net332),
    .A2(_05334_));
 sg13g2_buf_2 _13367_ (.A(\soc_I.rx_uart_i.fifo_i.din[0] ),
    .X(_05336_));
 sg13g2_buf_1 _13368_ (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ),
    .X(_05337_));
 sg13g2_buf_1 _13369_ (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[2] ),
    .X(_05338_));
 sg13g2_buf_1 _13370_ (.A(\soc_I.rx_uart_i.fifo_i.cnt[4] ),
    .X(_05339_));
 sg13g2_buf_1 _13371_ (.A(\soc_I.rx_uart_i.fifo_i.cnt[1] ),
    .X(_05340_));
 sg13g2_buf_1 _13372_ (.A(\soc_I.rx_uart_i.fifo_i.cnt[0] ),
    .X(_05341_));
 sg13g2_buf_1 _13373_ (.A(\soc_I.rx_uart_i.fifo_i.cnt[2] ),
    .X(_05342_));
 sg13g2_nor4_2 _13374_ (.A(_05340_),
    .B(_05341_),
    .C(\soc_I.rx_uart_i.fifo_i.cnt[3] ),
    .Y(_05343_),
    .D(_05342_));
 sg13g2_buf_1 _13375_ (.A(\soc_I.rx_uart_i.ready ),
    .X(_05344_));
 sg13g2_inv_1 _13376_ (.Y(_05345_),
    .A(_05344_));
 sg13g2_a21o_1 _13377_ (.A2(_05343_),
    .A1(_05339_),
    .B1(_05345_),
    .X(_05346_));
 sg13g2_buf_1 _13378_ (.A(_05346_),
    .X(_05347_));
 sg13g2_nor3_1 _13379_ (.A(net614),
    .B(net613),
    .C(_05347_),
    .Y(_05348_));
 sg13g2_buf_1 _13380_ (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[1] ),
    .X(_05349_));
 sg13g2_buf_1 _13381_ (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[0] ),
    .X(_05350_));
 sg13g2_nor2_1 _13382_ (.A(_05349_),
    .B(_05350_),
    .Y(_05351_));
 sg13g2_and2_1 _13383_ (.A(_05348_),
    .B(_05351_),
    .X(_05352_));
 sg13g2_buf_4 _13384_ (.X(_05353_),
    .A(_05352_));
 sg13g2_mux2_1 _13385_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[0][0] ),
    .A1(_05336_),
    .S(_05353_),
    .X(_01017_));
 sg13g2_buf_2 _13386_ (.A(\soc_I.rx_uart_i.fifo_i.din[1] ),
    .X(_05354_));
 sg13g2_mux2_1 _13387_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[0][1] ),
    .A1(_05354_),
    .S(_05353_),
    .X(_01018_));
 sg13g2_buf_2 _13388_ (.A(\soc_I.rx_uart_i.fifo_i.din[2] ),
    .X(_05355_));
 sg13g2_mux2_1 _13389_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[0][2] ),
    .A1(_05355_),
    .S(_05353_),
    .X(_01019_));
 sg13g2_buf_2 _13390_ (.A(\soc_I.rx_uart_i.fifo_i.din[3] ),
    .X(_05356_));
 sg13g2_mux2_1 _13391_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[0][3] ),
    .A1(_05356_),
    .S(_05353_),
    .X(_01020_));
 sg13g2_buf_2 _13392_ (.A(\soc_I.rx_uart_i.fifo_i.din[4] ),
    .X(_05357_));
 sg13g2_mux2_1 _13393_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[0][4] ),
    .A1(_05357_),
    .S(_05353_),
    .X(_01021_));
 sg13g2_buf_2 _13394_ (.A(\soc_I.rx_uart_i.fifo_i.din[5] ),
    .X(_05358_));
 sg13g2_mux2_1 _13395_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[0][5] ),
    .A1(_05358_),
    .S(_05353_),
    .X(_01022_));
 sg13g2_buf_2 _13396_ (.A(\soc_I.rx_uart_i.fifo_i.din[6] ),
    .X(_05359_));
 sg13g2_mux2_1 _13397_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[0][6] ),
    .A1(_05359_),
    .S(_05353_),
    .X(_01023_));
 sg13g2_buf_2 _13398_ (.A(\soc_I.rx_uart_i.fifo_i.din[7] ),
    .X(_05360_));
 sg13g2_mux2_1 _13399_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[0][7] ),
    .A1(_05360_),
    .S(_05353_),
    .X(_01024_));
 sg13g2_buf_1 _13400_ (.A(_05336_),
    .X(_05361_));
 sg13g2_inv_1 _13401_ (.Y(_05362_),
    .A(_05337_));
 sg13g2_nor3_1 _13402_ (.A(_05362_),
    .B(net613),
    .C(_05347_),
    .Y(_05363_));
 sg13g2_nor2b_1 _13403_ (.A(_05350_),
    .B_N(_05349_),
    .Y(_05364_));
 sg13g2_nand2_1 _13404_ (.Y(_05365_),
    .A(_05363_),
    .B(_05364_));
 sg13g2_buf_4 _13405_ (.X(_05366_),
    .A(_05365_));
 sg13g2_mux2_1 _13406_ (.A0(net588),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[10][0] ),
    .S(_05366_),
    .X(_01025_));
 sg13g2_buf_1 _13407_ (.A(_05354_),
    .X(_05367_));
 sg13g2_mux2_1 _13408_ (.A0(net587),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[10][1] ),
    .S(_05366_),
    .X(_01026_));
 sg13g2_buf_1 _13409_ (.A(_05355_),
    .X(_05368_));
 sg13g2_mux2_1 _13410_ (.A0(net586),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[10][2] ),
    .S(_05366_),
    .X(_01027_));
 sg13g2_buf_1 _13411_ (.A(_05356_),
    .X(_05369_));
 sg13g2_mux2_1 _13412_ (.A0(net585),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[10][3] ),
    .S(_05366_),
    .X(_01028_));
 sg13g2_buf_1 _13413_ (.A(_05357_),
    .X(_05370_));
 sg13g2_mux2_1 _13414_ (.A0(net584),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[10][4] ),
    .S(_05366_),
    .X(_01029_));
 sg13g2_buf_1 _13415_ (.A(_05358_),
    .X(_05371_));
 sg13g2_mux2_1 _13416_ (.A0(net583),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[10][5] ),
    .S(_05366_),
    .X(_01030_));
 sg13g2_buf_1 _13417_ (.A(_05359_),
    .X(_05372_));
 sg13g2_mux2_1 _13418_ (.A0(net582),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[10][6] ),
    .S(_05366_),
    .X(_01031_));
 sg13g2_buf_1 _13419_ (.A(_05360_),
    .X(_05373_));
 sg13g2_mux2_1 _13420_ (.A0(_05373_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[10][7] ),
    .S(_05366_),
    .X(_01032_));
 sg13g2_nand2_1 _13421_ (.Y(_05374_),
    .A(_05349_),
    .B(_05350_));
 sg13g2_buf_1 _13422_ (.A(_05374_),
    .X(_05375_));
 sg13g2_nor4_1 _13423_ (.A(_05362_),
    .B(net613),
    .C(_05347_),
    .D(_05375_),
    .Y(_05376_));
 sg13g2_buf_4 _13424_ (.X(_05377_),
    .A(_05376_));
 sg13g2_mux2_1 _13425_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[11][0] ),
    .A1(_05336_),
    .S(_05377_),
    .X(_01033_));
 sg13g2_mux2_1 _13426_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[11][1] ),
    .A1(_05354_),
    .S(_05377_),
    .X(_01034_));
 sg13g2_mux2_1 _13427_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[11][2] ),
    .A1(_05355_),
    .S(_05377_),
    .X(_01035_));
 sg13g2_mux2_1 _13428_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[11][3] ),
    .A1(_05356_),
    .S(_05377_),
    .X(_01036_));
 sg13g2_mux2_1 _13429_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[11][4] ),
    .A1(_05357_),
    .S(_05377_),
    .X(_01037_));
 sg13g2_mux2_1 _13430_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[11][5] ),
    .A1(_05358_),
    .S(_05377_),
    .X(_01038_));
 sg13g2_mux2_1 _13431_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[11][6] ),
    .A1(_05359_),
    .S(_05377_),
    .X(_01039_));
 sg13g2_mux2_1 _13432_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[11][7] ),
    .A1(_05360_),
    .S(_05377_),
    .X(_01040_));
 sg13g2_a21oi_1 _13433_ (.A1(_05339_),
    .A2(_05343_),
    .Y(_05378_),
    .B1(_05345_));
 sg13g2_buf_1 _13434_ (.A(_05378_),
    .X(_05379_));
 sg13g2_nand4_1 _13435_ (.B(net613),
    .C(net442),
    .A(net614),
    .Y(_05380_),
    .D(_05351_));
 sg13g2_buf_4 _13436_ (.X(_05381_),
    .A(_05380_));
 sg13g2_mux2_1 _13437_ (.A0(net588),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[12][0] ),
    .S(_05381_),
    .X(_01041_));
 sg13g2_mux2_1 _13438_ (.A0(net587),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[12][1] ),
    .S(_05381_),
    .X(_01042_));
 sg13g2_mux2_1 _13439_ (.A0(net586),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[12][2] ),
    .S(_05381_),
    .X(_01043_));
 sg13g2_mux2_1 _13440_ (.A0(net585),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[12][3] ),
    .S(_05381_),
    .X(_01044_));
 sg13g2_mux2_1 _13441_ (.A0(net584),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[12][4] ),
    .S(_05381_),
    .X(_01045_));
 sg13g2_mux2_1 _13442_ (.A0(net583),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[12][5] ),
    .S(_05381_),
    .X(_01046_));
 sg13g2_mux2_1 _13443_ (.A0(net582),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[12][6] ),
    .S(_05381_),
    .X(_01047_));
 sg13g2_mux2_1 _13444_ (.A0(net581),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[12][7] ),
    .S(_05381_),
    .X(_01048_));
 sg13g2_nand3_1 _13445_ (.B(net613),
    .C(net442),
    .A(net614),
    .Y(_05382_));
 sg13g2_nor2b_1 _13446_ (.A(_05349_),
    .B_N(_05350_),
    .Y(_05383_));
 sg13g2_nand2b_1 _13447_ (.Y(_05384_),
    .B(_05383_),
    .A_N(_05382_));
 sg13g2_buf_4 _13448_ (.X(_05385_),
    .A(_05384_));
 sg13g2_mux2_1 _13449_ (.A0(net588),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][0] ),
    .S(_05385_),
    .X(_01049_));
 sg13g2_mux2_1 _13450_ (.A0(net587),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][1] ),
    .S(_05385_),
    .X(_01050_));
 sg13g2_mux2_1 _13451_ (.A0(net586),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][2] ),
    .S(_05385_),
    .X(_01051_));
 sg13g2_mux2_1 _13452_ (.A0(net585),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][3] ),
    .S(_05385_),
    .X(_01052_));
 sg13g2_mux2_1 _13453_ (.A0(net584),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][4] ),
    .S(_05385_),
    .X(_01053_));
 sg13g2_mux2_1 _13454_ (.A0(net583),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][5] ),
    .S(_05385_),
    .X(_01054_));
 sg13g2_mux2_1 _13455_ (.A0(net582),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][6] ),
    .S(_05385_),
    .X(_01055_));
 sg13g2_mux2_1 _13456_ (.A0(net581),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][7] ),
    .S(_05385_),
    .X(_01056_));
 sg13g2_nand4_1 _13457_ (.B(net613),
    .C(net442),
    .A(net614),
    .Y(_05386_),
    .D(_05364_));
 sg13g2_buf_4 _13458_ (.X(_05387_),
    .A(_05386_));
 sg13g2_mux2_1 _13459_ (.A0(net588),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[14][0] ),
    .S(_05387_),
    .X(_01057_));
 sg13g2_mux2_1 _13460_ (.A0(net587),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[14][1] ),
    .S(_05387_),
    .X(_01058_));
 sg13g2_mux2_1 _13461_ (.A0(net586),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[14][2] ),
    .S(_05387_),
    .X(_01059_));
 sg13g2_mux2_1 _13462_ (.A0(net585),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[14][3] ),
    .S(_05387_),
    .X(_01060_));
 sg13g2_mux2_1 _13463_ (.A0(net584),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[14][4] ),
    .S(_05387_),
    .X(_01061_));
 sg13g2_mux2_1 _13464_ (.A0(net583),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[14][5] ),
    .S(_05387_),
    .X(_01062_));
 sg13g2_mux2_1 _13465_ (.A0(net582),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[14][6] ),
    .S(_05387_),
    .X(_01063_));
 sg13g2_mux2_1 _13466_ (.A0(net581),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[14][7] ),
    .S(_05387_),
    .X(_01064_));
 sg13g2_or2_1 _13467_ (.X(_05388_),
    .B(_05382_),
    .A(_05375_));
 sg13g2_buf_4 _13468_ (.X(_05389_),
    .A(_05388_));
 sg13g2_mux2_1 _13469_ (.A0(net588),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][0] ),
    .S(_05389_),
    .X(_01065_));
 sg13g2_mux2_1 _13470_ (.A0(net587),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][1] ),
    .S(_05389_),
    .X(_01066_));
 sg13g2_mux2_1 _13471_ (.A0(net586),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][2] ),
    .S(_05389_),
    .X(_01067_));
 sg13g2_mux2_1 _13472_ (.A0(net585),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][3] ),
    .S(_05389_),
    .X(_01068_));
 sg13g2_mux2_1 _13473_ (.A0(net584),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][4] ),
    .S(_05389_),
    .X(_01069_));
 sg13g2_mux2_1 _13474_ (.A0(net583),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][5] ),
    .S(_05389_),
    .X(_01070_));
 sg13g2_mux2_1 _13475_ (.A0(net582),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][6] ),
    .S(_05389_),
    .X(_01071_));
 sg13g2_mux2_1 _13476_ (.A0(net581),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][7] ),
    .S(_05389_),
    .X(_01072_));
 sg13g2_and2_1 _13477_ (.A(_05348_),
    .B(_05383_),
    .X(_05390_));
 sg13g2_buf_4 _13478_ (.X(_05391_),
    .A(_05390_));
 sg13g2_mux2_1 _13479_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[1][0] ),
    .A1(_05336_),
    .S(_05391_),
    .X(_01073_));
 sg13g2_mux2_1 _13480_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[1][1] ),
    .A1(_05354_),
    .S(_05391_),
    .X(_01074_));
 sg13g2_mux2_1 _13481_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[1][2] ),
    .A1(_05355_),
    .S(_05391_),
    .X(_01075_));
 sg13g2_mux2_1 _13482_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[1][3] ),
    .A1(_05356_),
    .S(_05391_),
    .X(_01076_));
 sg13g2_mux2_1 _13483_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[1][4] ),
    .A1(_05357_),
    .S(_05391_),
    .X(_01077_));
 sg13g2_mux2_1 _13484_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[1][5] ),
    .A1(_05358_),
    .S(_05391_),
    .X(_01078_));
 sg13g2_mux2_1 _13485_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[1][6] ),
    .A1(_05359_),
    .S(_05391_),
    .X(_01079_));
 sg13g2_mux2_1 _13486_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[1][7] ),
    .A1(_05360_),
    .S(_05391_),
    .X(_01080_));
 sg13g2_and2_1 _13487_ (.A(_05348_),
    .B(_05364_),
    .X(_05392_));
 sg13g2_buf_4 _13488_ (.X(_05393_),
    .A(_05392_));
 sg13g2_mux2_1 _13489_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[2][0] ),
    .A1(_05336_),
    .S(_05393_),
    .X(_01081_));
 sg13g2_mux2_1 _13490_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[2][1] ),
    .A1(_05354_),
    .S(_05393_),
    .X(_01082_));
 sg13g2_mux2_1 _13491_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[2][2] ),
    .A1(_05355_),
    .S(_05393_),
    .X(_01083_));
 sg13g2_mux2_1 _13492_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[2][3] ),
    .A1(_05356_),
    .S(_05393_),
    .X(_01084_));
 sg13g2_mux2_1 _13493_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[2][4] ),
    .A1(_05357_),
    .S(_05393_),
    .X(_01085_));
 sg13g2_mux2_1 _13494_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[2][5] ),
    .A1(_05358_),
    .S(_05393_),
    .X(_01086_));
 sg13g2_mux2_1 _13495_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[2][6] ),
    .A1(_05359_),
    .S(_05393_),
    .X(_01087_));
 sg13g2_mux2_1 _13496_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[2][7] ),
    .A1(_05360_),
    .S(_05393_),
    .X(_01088_));
 sg13g2_nor4_1 _13497_ (.A(net614),
    .B(_05338_),
    .C(_05347_),
    .D(_05375_),
    .Y(_05394_));
 sg13g2_buf_4 _13498_ (.X(_05395_),
    .A(_05394_));
 sg13g2_mux2_1 _13499_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[3][0] ),
    .A1(_05336_),
    .S(_05395_),
    .X(_01089_));
 sg13g2_mux2_1 _13500_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[3][1] ),
    .A1(_05354_),
    .S(_05395_),
    .X(_01090_));
 sg13g2_mux2_1 _13501_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[3][2] ),
    .A1(_05355_),
    .S(_05395_),
    .X(_01091_));
 sg13g2_mux2_1 _13502_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[3][3] ),
    .A1(_05356_),
    .S(_05395_),
    .X(_01092_));
 sg13g2_mux2_1 _13503_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[3][4] ),
    .A1(_05357_),
    .S(_05395_),
    .X(_01093_));
 sg13g2_mux2_1 _13504_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[3][5] ),
    .A1(_05358_),
    .S(_05395_),
    .X(_01094_));
 sg13g2_mux2_1 _13505_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[3][6] ),
    .A1(_05359_),
    .S(_05395_),
    .X(_01095_));
 sg13g2_mux2_1 _13506_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[3][7] ),
    .A1(_05360_),
    .S(_05395_),
    .X(_01096_));
 sg13g2_nand2_1 _13507_ (.Y(_05396_),
    .A(net613),
    .B(net442));
 sg13g2_nor2_1 _13508_ (.A(net614),
    .B(_05396_),
    .Y(_05397_));
 sg13g2_nand2_1 _13509_ (.Y(_05398_),
    .A(_05351_),
    .B(_05397_));
 sg13g2_buf_4 _13510_ (.X(_05399_),
    .A(_05398_));
 sg13g2_mux2_1 _13511_ (.A0(net588),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[4][0] ),
    .S(_05399_),
    .X(_01097_));
 sg13g2_mux2_1 _13512_ (.A0(net587),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[4][1] ),
    .S(_05399_),
    .X(_01098_));
 sg13g2_mux2_1 _13513_ (.A0(net586),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[4][2] ),
    .S(_05399_),
    .X(_01099_));
 sg13g2_mux2_1 _13514_ (.A0(net585),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[4][3] ),
    .S(_05399_),
    .X(_01100_));
 sg13g2_mux2_1 _13515_ (.A0(net584),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[4][4] ),
    .S(_05399_),
    .X(_01101_));
 sg13g2_mux2_1 _13516_ (.A0(net583),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[4][5] ),
    .S(_05399_),
    .X(_01102_));
 sg13g2_mux2_1 _13517_ (.A0(net582),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[4][6] ),
    .S(_05399_),
    .X(_01103_));
 sg13g2_mux2_1 _13518_ (.A0(net581),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[4][7] ),
    .S(_05399_),
    .X(_01104_));
 sg13g2_nand2_1 _13519_ (.Y(_05400_),
    .A(_05383_),
    .B(_05397_));
 sg13g2_buf_4 _13520_ (.X(_05401_),
    .A(_05400_));
 sg13g2_mux2_1 _13521_ (.A0(net588),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][0] ),
    .S(_05401_),
    .X(_01105_));
 sg13g2_mux2_1 _13522_ (.A0(net587),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][1] ),
    .S(_05401_),
    .X(_01106_));
 sg13g2_mux2_1 _13523_ (.A0(net586),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][2] ),
    .S(_05401_),
    .X(_01107_));
 sg13g2_mux2_1 _13524_ (.A0(net585),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][3] ),
    .S(_05401_),
    .X(_01108_));
 sg13g2_mux2_1 _13525_ (.A0(_05370_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][4] ),
    .S(_05401_),
    .X(_01109_));
 sg13g2_mux2_1 _13526_ (.A0(net583),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][5] ),
    .S(_05401_),
    .X(_01110_));
 sg13g2_mux2_1 _13527_ (.A0(net582),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][6] ),
    .S(_05401_),
    .X(_01111_));
 sg13g2_mux2_1 _13528_ (.A0(net581),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][7] ),
    .S(_05401_),
    .X(_01112_));
 sg13g2_nand2_1 _13529_ (.Y(_05402_),
    .A(_05364_),
    .B(_05397_));
 sg13g2_buf_4 _13530_ (.X(_05403_),
    .A(_05402_));
 sg13g2_mux2_1 _13531_ (.A0(_05361_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[6][0] ),
    .S(_05403_),
    .X(_01113_));
 sg13g2_mux2_1 _13532_ (.A0(net587),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[6][1] ),
    .S(_05403_),
    .X(_01114_));
 sg13g2_mux2_1 _13533_ (.A0(net586),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[6][2] ),
    .S(_05403_),
    .X(_01115_));
 sg13g2_mux2_1 _13534_ (.A0(_05369_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[6][3] ),
    .S(_05403_),
    .X(_01116_));
 sg13g2_mux2_1 _13535_ (.A0(_05370_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[6][4] ),
    .S(_05403_),
    .X(_01117_));
 sg13g2_mux2_1 _13536_ (.A0(_05371_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[6][5] ),
    .S(_05403_),
    .X(_01118_));
 sg13g2_mux2_1 _13537_ (.A0(_05372_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[6][6] ),
    .S(_05403_),
    .X(_01119_));
 sg13g2_mux2_1 _13538_ (.A0(net581),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[6][7] ),
    .S(_05403_),
    .X(_01120_));
 sg13g2_nor3_1 _13539_ (.A(net614),
    .B(_05375_),
    .C(_05396_),
    .Y(_05404_));
 sg13g2_buf_1 _13540_ (.A(_05404_),
    .X(_05405_));
 sg13g2_mux2_1 _13541_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[7][0] ),
    .A1(_05336_),
    .S(net331),
    .X(_01121_));
 sg13g2_mux2_1 _13542_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[7][1] ),
    .A1(_05354_),
    .S(net331),
    .X(_01122_));
 sg13g2_mux2_1 _13543_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[7][2] ),
    .A1(_05355_),
    .S(net331),
    .X(_01123_));
 sg13g2_mux2_1 _13544_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[7][3] ),
    .A1(_05356_),
    .S(net331),
    .X(_01124_));
 sg13g2_mux2_1 _13545_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[7][4] ),
    .A1(_05357_),
    .S(_05405_),
    .X(_01125_));
 sg13g2_mux2_1 _13546_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[7][5] ),
    .A1(_05358_),
    .S(net331),
    .X(_01126_));
 sg13g2_mux2_1 _13547_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[7][6] ),
    .A1(_05359_),
    .S(net331),
    .X(_01127_));
 sg13g2_mux2_1 _13548_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[7][7] ),
    .A1(_05360_),
    .S(net331),
    .X(_01128_));
 sg13g2_nand2_1 _13549_ (.Y(_05406_),
    .A(_05351_),
    .B(_05363_));
 sg13g2_buf_4 _13550_ (.X(_05407_),
    .A(_05406_));
 sg13g2_mux2_1 _13551_ (.A0(_05361_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[8][0] ),
    .S(_05407_),
    .X(_01129_));
 sg13g2_mux2_1 _13552_ (.A0(_05367_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[8][1] ),
    .S(_05407_),
    .X(_01130_));
 sg13g2_mux2_1 _13553_ (.A0(_05368_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[8][2] ),
    .S(_05407_),
    .X(_01131_));
 sg13g2_mux2_1 _13554_ (.A0(_05369_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[8][3] ),
    .S(_05407_),
    .X(_01132_));
 sg13g2_mux2_1 _13555_ (.A0(net584),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[8][4] ),
    .S(_05407_),
    .X(_01133_));
 sg13g2_mux2_1 _13556_ (.A0(_05371_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[8][5] ),
    .S(_05407_),
    .X(_01134_));
 sg13g2_mux2_1 _13557_ (.A0(net582),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[8][6] ),
    .S(_05407_),
    .X(_01135_));
 sg13g2_mux2_1 _13558_ (.A0(_05373_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[8][7] ),
    .S(_05407_),
    .X(_01136_));
 sg13g2_nand2_1 _13559_ (.Y(_05408_),
    .A(_05363_),
    .B(_05383_));
 sg13g2_buf_4 _13560_ (.X(_05409_),
    .A(_05408_));
 sg13g2_mux2_1 _13561_ (.A0(net588),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][0] ),
    .S(_05409_),
    .X(_01137_));
 sg13g2_mux2_1 _13562_ (.A0(_05367_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][1] ),
    .S(_05409_),
    .X(_01138_));
 sg13g2_mux2_1 _13563_ (.A0(_05368_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][2] ),
    .S(_05409_),
    .X(_01139_));
 sg13g2_mux2_1 _13564_ (.A0(net585),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][3] ),
    .S(_05409_),
    .X(_01140_));
 sg13g2_mux2_1 _13565_ (.A0(net584),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][4] ),
    .S(_05409_),
    .X(_01141_));
 sg13g2_mux2_1 _13566_ (.A0(net583),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][5] ),
    .S(_05409_),
    .X(_01142_));
 sg13g2_mux2_1 _13567_ (.A0(_05372_),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][6] ),
    .S(_05409_),
    .X(_01143_));
 sg13g2_mux2_1 _13568_ (.A0(net581),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][7] ),
    .S(_05409_),
    .X(_01144_));
 sg13g2_buf_1 _13569_ (.A(\soc_I.rx_uart_i.bit_idx[2] ),
    .X(_05410_));
 sg13g2_buf_1 _13570_ (.A(\soc_I.rx_uart_i.state[0] ),
    .X(_05411_));
 sg13g2_buf_1 _13571_ (.A(_05411_),
    .X(_05412_));
 sg13g2_buf_2 _13572_ (.A(\soc_I.rx_uart_i.state[1] ),
    .X(_05413_));
 sg13g2_buf_1 _13573_ (.A(_00047_),
    .X(_05414_));
 sg13g2_nand2_2 _13574_ (.Y(_05415_),
    .A(_05413_),
    .B(net612));
 sg13g2_nor2_1 _13575_ (.A(net580),
    .B(_05415_),
    .Y(_05416_));
 sg13g2_nand2_2 _13576_ (.Y(_05417_),
    .A(_05410_),
    .B(_05416_));
 sg13g2_buf_1 _13577_ (.A(\soc_I.rx_uart_i.bit_idx[1] ),
    .X(_05418_));
 sg13g2_buf_2 _13578_ (.A(\soc_I.rx_uart_i.bit_idx[0] ),
    .X(_05419_));
 sg13g2_nand2_1 _13579_ (.Y(_05420_),
    .A(_05418_),
    .B(_05419_));
 sg13g2_nor2_1 _13580_ (.A(_05413_),
    .B(_05411_),
    .Y(_05421_));
 sg13g2_nor2b_1 _13581_ (.A(_05421_),
    .B_N(net612),
    .Y(_05422_));
 sg13g2_buf_1 _13582_ (.A(_05422_),
    .X(_05423_));
 sg13g2_buf_1 _13583_ (.A(net441),
    .X(_05424_));
 sg13g2_o21ai_1 _13584_ (.B1(net408),
    .Y(_05425_),
    .A1(_05417_),
    .A2(_05420_));
 sg13g2_inv_1 _13585_ (.Y(_05426_),
    .A(_05412_));
 sg13g2_buf_1 _13586_ (.A(\soc_I.rx_uart_i.rx_in_sync[2] ),
    .X(_05427_));
 sg13g2_o21ai_1 _13587_ (.B1(_05413_),
    .Y(_05428_),
    .A1(_05426_),
    .A2(net611));
 sg13g2_nor2b_1 _13588_ (.A(\soc_I.rx_uart_i.rx_in_sync[1] ),
    .B_N(net611),
    .Y(_05429_));
 sg13g2_nor3_1 _13589_ (.A(_05413_),
    .B(_05426_),
    .C(net611),
    .Y(_05430_));
 sg13g2_a21oi_1 _13590_ (.A1(_05426_),
    .A2(_05429_),
    .Y(_05431_),
    .B1(_05430_));
 sg13g2_nand2_1 _13591_ (.Y(_05432_),
    .A(net612),
    .B(_03577_));
 sg13g2_a21oi_2 _13592_ (.B1(_05432_),
    .Y(_05433_),
    .A2(_05431_),
    .A1(_05428_));
 sg13g2_mux2_1 _13593_ (.A0(\soc_I.rx_uart_i.return_state[0] ),
    .A1(_05425_),
    .S(_05433_),
    .X(_01151_));
 sg13g2_inv_1 _13594_ (.Y(_05434_),
    .A(\soc_I.rx_uart_i.return_state[1] ));
 sg13g2_xor2_1 _13595_ (.B(net580),
    .A(_05413_),
    .X(_05435_));
 sg13g2_nand3_1 _13596_ (.B(_05433_),
    .C(_05435_),
    .A(net612),
    .Y(_05436_));
 sg13g2_o21ai_1 _13597_ (.B1(_05436_),
    .Y(_01152_),
    .A1(_05434_),
    .A2(_05433_));
 sg13g2_buf_1 _13598_ (.A(\soc_I.tx_uart_i.state[1] ),
    .X(_05437_));
 sg13g2_buf_1 _13599_ (.A(\soc_I.tx_uart_i.state[0] ),
    .X(_05438_));
 sg13g2_nand2_1 _13600_ (.Y(_05439_),
    .A(_05437_),
    .B(_05438_));
 sg13g2_buf_1 _13601_ (.A(_05439_),
    .X(_05440_));
 sg13g2_buf_1 _13602_ (.A(net508),
    .X(_05441_));
 sg13g2_buf_1 _13603_ (.A(net440),
    .X(_05442_));
 sg13g2_nand3_1 _13604_ (.B(_04232_),
    .C(_04234_),
    .A(_04046_),
    .Y(_05443_));
 sg13g2_buf_1 _13605_ (.A(_05443_),
    .X(_05444_));
 sg13g2_nand2_1 _13606_ (.Y(_05445_),
    .A(_04225_),
    .B(net594));
 sg13g2_or3_1 _13607_ (.A(\soc_I.tx_uart_i.ready ),
    .B(\soc_I.cpu_mem_addr[0] ),
    .C(_05445_),
    .X(_05446_));
 sg13g2_nor2_1 _13608_ (.A(_05437_),
    .B(net610),
    .Y(_05447_));
 sg13g2_buf_1 _13609_ (.A(_05447_),
    .X(_05448_));
 sg13g2_o21ai_1 _13610_ (.B1(_05448_),
    .Y(_05449_),
    .A1(_05444_),
    .A2(_05446_));
 sg13g2_and2_1 _13611_ (.A(_04285_),
    .B(_05449_),
    .X(_05450_));
 sg13g2_buf_2 _13612_ (.A(_05450_),
    .X(_05451_));
 sg13g2_nand2_1 _13613_ (.Y(_05452_),
    .A(net407),
    .B(_05451_));
 sg13g2_buf_1 _13614_ (.A(_05437_),
    .X(_05453_));
 sg13g2_nor2_2 _13615_ (.A(_05444_),
    .B(_05446_),
    .Y(_05454_));
 sg13g2_nor2b_1 _13616_ (.A(_05454_),
    .B_N(_05448_),
    .Y(_05455_));
 sg13g2_buf_2 _13617_ (.A(\soc_I.tx_uart_i.bit_idx[0] ),
    .X(_05456_));
 sg13g2_buf_1 _13618_ (.A(\soc_I.tx_uart_i.bit_idx[1] ),
    .X(_05457_));
 sg13g2_inv_1 _13619_ (.Y(_05458_),
    .A(net610));
 sg13g2_nor2_1 _13620_ (.A(net579),
    .B(_05458_),
    .Y(_05459_));
 sg13g2_nand3_1 _13621_ (.B(_05457_),
    .C(_05459_),
    .A(_05456_),
    .Y(_05460_));
 sg13g2_nor2_1 _13622_ (.A(_00083_),
    .B(_05460_),
    .Y(_05461_));
 sg13g2_nor4_1 _13623_ (.A(net579),
    .B(_04273_),
    .C(_05455_),
    .D(_05461_),
    .Y(_05462_));
 sg13g2_a21o_1 _13624_ (.A2(_05452_),
    .A1(\soc_I.tx_uart_i.return_state[0] ),
    .B1(_05462_),
    .X(_01266_));
 sg13g2_mux2_1 _13625_ (.A0(_05461_),
    .A1(\soc_I.tx_uart_i.return_state[1] ),
    .S(_05452_),
    .X(_01267_));
 sg13g2_buf_1 _13626_ (.A(\soc_I.tx_uart_i.wait_states[0] ),
    .X(_05463_));
 sg13g2_inv_1 _13627_ (.Y(_05464_),
    .A(_05463_));
 sg13g2_buf_1 _13628_ (.A(_05451_),
    .X(_05465_));
 sg13g2_buf_1 _13629_ (.A(_05451_),
    .X(_05466_));
 sg13g2_inv_1 _13630_ (.Y(_05467_),
    .A(_05437_));
 sg13g2_buf_2 _13631_ (.A(\soc_I.div_reg[0] ),
    .X(_05468_));
 sg13g2_nor2_1 _13632_ (.A(_05467_),
    .B(_05458_),
    .Y(_05469_));
 sg13g2_buf_1 _13633_ (.A(_05469_),
    .X(_05470_));
 sg13g2_a22oi_1 _13634_ (.Y(_05471_),
    .B1(_05463_),
    .B2(net439),
    .A2(_05468_),
    .A1(_05467_));
 sg13g2_nand2_1 _13635_ (.Y(_05472_),
    .A(net58),
    .B(_05471_));
 sg13g2_o21ai_1 _13636_ (.B1(_05472_),
    .Y(_01280_),
    .A1(_05464_),
    .A2(net59));
 sg13g2_nand2_1 _13637_ (.Y(_05473_),
    .A(_05437_),
    .B(_05458_));
 sg13g2_buf_1 _13638_ (.A(_05473_),
    .X(_05474_));
 sg13g2_buf_1 _13639_ (.A(_05474_),
    .X(_05475_));
 sg13g2_buf_1 _13640_ (.A(\soc_I.tx_uart_i.wait_states[9] ),
    .X(_05476_));
 sg13g2_buf_1 _13641_ (.A(\soc_I.tx_uart_i.wait_states[8] ),
    .X(_05477_));
 sg13g2_nor3_1 _13642_ (.A(_05476_),
    .B(_05477_),
    .C(_05440_),
    .Y(_05478_));
 sg13g2_buf_1 _13643_ (.A(\soc_I.div_reg[8] ),
    .X(_05479_));
 sg13g2_buf_2 _13644_ (.A(\soc_I.div_reg[9] ),
    .X(_05480_));
 sg13g2_nor3_1 _13645_ (.A(net609),
    .B(_05480_),
    .C(_05470_),
    .Y(_05481_));
 sg13g2_buf_1 _13646_ (.A(\soc_I.tx_uart_i.wait_states[7] ),
    .X(_05482_));
 sg13g2_buf_1 _13647_ (.A(\soc_I.tx_uart_i.wait_states[6] ),
    .X(_05483_));
 sg13g2_nor3_1 _13648_ (.A(_05482_),
    .B(_05483_),
    .C(net508),
    .Y(_05484_));
 sg13g2_buf_2 _13649_ (.A(\soc_I.div_reg[6] ),
    .X(_05485_));
 sg13g2_buf_2 _13650_ (.A(\soc_I.div_reg[7] ),
    .X(_05486_));
 sg13g2_nor3_1 _13651_ (.A(_05485_),
    .B(_05486_),
    .C(net439),
    .Y(_05487_));
 sg13g2_buf_1 _13652_ (.A(\soc_I.tx_uart_i.wait_states[5] ),
    .X(_05488_));
 sg13g2_buf_1 _13653_ (.A(\soc_I.tx_uart_i.wait_states[4] ),
    .X(_05489_));
 sg13g2_nor3_1 _13654_ (.A(_05488_),
    .B(_05489_),
    .C(net508),
    .Y(_05490_));
 sg13g2_buf_2 _13655_ (.A(\soc_I.div_reg[4] ),
    .X(_05491_));
 sg13g2_buf_2 _13656_ (.A(\soc_I.div_reg[5] ),
    .X(_05492_));
 sg13g2_nor3_1 _13657_ (.A(_05491_),
    .B(_05492_),
    .C(net439),
    .Y(_05493_));
 sg13g2_buf_1 _13658_ (.A(\soc_I.tx_uart_i.wait_states[3] ),
    .X(_05494_));
 sg13g2_buf_1 _13659_ (.A(\soc_I.tx_uart_i.wait_states[2] ),
    .X(_05495_));
 sg13g2_nor3_1 _13660_ (.A(_05494_),
    .B(_05495_),
    .C(net508),
    .Y(_05496_));
 sg13g2_buf_2 _13661_ (.A(\soc_I.div_reg[2] ),
    .X(_05497_));
 sg13g2_buf_2 _13662_ (.A(\soc_I.div_reg[3] ),
    .X(_05498_));
 sg13g2_nor3_1 _13663_ (.A(_05497_),
    .B(_05498_),
    .C(net439),
    .Y(_05499_));
 sg13g2_buf_2 _13664_ (.A(\soc_I.div_reg[1] ),
    .X(_05500_));
 sg13g2_nor2_1 _13665_ (.A(_05468_),
    .B(_05500_),
    .Y(_05501_));
 sg13g2_buf_1 _13666_ (.A(\soc_I.tx_uart_i.wait_states[1] ),
    .X(_05502_));
 sg13g2_nor3_1 _13667_ (.A(_05463_),
    .B(_05502_),
    .C(net508),
    .Y(_05503_));
 sg13g2_a21oi_2 _13668_ (.B1(_05503_),
    .Y(_05504_),
    .A2(_05501_),
    .A1(net508));
 sg13g2_inv_1 _13669_ (.Y(_05505_),
    .A(_05504_));
 sg13g2_o21ai_1 _13670_ (.B1(_05505_),
    .Y(_05506_),
    .A1(_05496_),
    .A2(_05499_));
 sg13g2_buf_1 _13671_ (.A(_05506_),
    .X(_05507_));
 sg13g2_inv_1 _13672_ (.Y(_05508_),
    .A(_05507_));
 sg13g2_o21ai_1 _13673_ (.B1(_05508_),
    .Y(_05509_),
    .A1(_05490_),
    .A2(_05493_));
 sg13g2_buf_1 _13674_ (.A(_05509_),
    .X(_05510_));
 sg13g2_inv_1 _13675_ (.Y(_05511_),
    .A(_05510_));
 sg13g2_o21ai_1 _13676_ (.B1(_05511_),
    .Y(_05512_),
    .A1(_05484_),
    .A2(_05487_));
 sg13g2_buf_1 _13677_ (.A(_05512_),
    .X(_05513_));
 sg13g2_inv_1 _13678_ (.Y(_05514_),
    .A(_05513_));
 sg13g2_o21ai_1 _13679_ (.B1(_05514_),
    .Y(_05515_),
    .A1(_05478_),
    .A2(_05481_));
 sg13g2_buf_2 _13680_ (.A(\soc_I.div_reg[10] ),
    .X(_05516_));
 sg13g2_mux2_1 _13681_ (.A0(\soc_I.tx_uart_i.wait_states[10] ),
    .A1(_05516_),
    .S(net508),
    .X(_05517_));
 sg13g2_xnor2_1 _13682_ (.Y(_05518_),
    .A(_05515_),
    .B(_05517_));
 sg13g2_nor3_2 _13683_ (.A(_05468_),
    .B(_05500_),
    .C(_05497_),
    .Y(_05519_));
 sg13g2_nor2b_1 _13684_ (.A(_05498_),
    .B_N(_05519_),
    .Y(_05520_));
 sg13g2_nor2b_1 _13685_ (.A(_05491_),
    .B_N(_05520_),
    .Y(_05521_));
 sg13g2_nor2b_1 _13686_ (.A(_05492_),
    .B_N(_05521_),
    .Y(_05522_));
 sg13g2_nor2b_1 _13687_ (.A(_05485_),
    .B_N(_05522_),
    .Y(_05523_));
 sg13g2_nand2b_1 _13688_ (.Y(_05524_),
    .B(_05523_),
    .A_N(_05486_));
 sg13g2_buf_1 _13689_ (.A(_05524_),
    .X(_05525_));
 sg13g2_nor2_1 _13690_ (.A(net609),
    .B(_05525_),
    .Y(_05526_));
 sg13g2_xnor2_1 _13691_ (.Y(_05527_),
    .A(_05480_),
    .B(_05526_));
 sg13g2_buf_1 _13692_ (.A(_05474_),
    .X(_05528_));
 sg13g2_nor2_1 _13693_ (.A(_05527_),
    .B(_05528_),
    .Y(_05529_));
 sg13g2_a21oi_1 _13694_ (.A1(_05475_),
    .A2(_05518_),
    .Y(_05530_),
    .B1(_05529_));
 sg13g2_nor2_1 _13695_ (.A(\soc_I.tx_uart_i.wait_states[10] ),
    .B(net58),
    .Y(_05531_));
 sg13g2_a21oi_1 _13696_ (.A1(net59),
    .A2(_05530_),
    .Y(_01281_),
    .B1(_05531_));
 sg13g2_or2_1 _13697_ (.X(_05532_),
    .B(_05517_),
    .A(_05515_));
 sg13g2_buf_1 _13698_ (.A(_05532_),
    .X(_05533_));
 sg13g2_buf_1 _13699_ (.A(\soc_I.tx_uart_i.wait_states[11] ),
    .X(_05534_));
 sg13g2_buf_1 _13700_ (.A(\soc_I.div_reg[11] ),
    .X(_05535_));
 sg13g2_mux2_1 _13701_ (.A0(_05534_),
    .A1(net608),
    .S(_05441_),
    .X(_05536_));
 sg13g2_xnor2_1 _13702_ (.Y(_05537_),
    .A(_05533_),
    .B(_05536_));
 sg13g2_nor3_1 _13703_ (.A(net609),
    .B(_05480_),
    .C(_05525_),
    .Y(_05538_));
 sg13g2_xnor2_1 _13704_ (.Y(_05539_),
    .A(_05516_),
    .B(_05538_));
 sg13g2_nor2_1 _13705_ (.A(_05528_),
    .B(_05539_),
    .Y(_05540_));
 sg13g2_a21oi_1 _13706_ (.A1(_05475_),
    .A2(_05537_),
    .Y(_05541_),
    .B1(_05540_));
 sg13g2_nor2_1 _13707_ (.A(_05534_),
    .B(net58),
    .Y(_05542_));
 sg13g2_a21oi_1 _13708_ (.A1(net59),
    .A2(_05541_),
    .Y(_01282_),
    .B1(_05542_));
 sg13g2_buf_1 _13709_ (.A(\soc_I.tx_uart_i.wait_states[12] ),
    .X(_05543_));
 sg13g2_buf_2 _13710_ (.A(\soc_I.div_reg[12] ),
    .X(_05544_));
 sg13g2_nor2_1 _13711_ (.A(net608),
    .B(_05533_),
    .Y(_05545_));
 sg13g2_xor2_1 _13712_ (.B(_05545_),
    .A(_05544_),
    .X(_05546_));
 sg13g2_nor2_1 _13713_ (.A(_05534_),
    .B(_05533_),
    .Y(_05547_));
 sg13g2_xnor2_1 _13714_ (.Y(_05548_),
    .A(_05543_),
    .B(_05547_));
 sg13g2_nor2_1 _13715_ (.A(net407),
    .B(_05548_),
    .Y(_05549_));
 sg13g2_a21oi_1 _13716_ (.A1(net407),
    .A2(_05546_),
    .Y(_05550_),
    .B1(_05549_));
 sg13g2_nor2b_1 _13717_ (.A(_05516_),
    .B_N(_05538_),
    .Y(_05551_));
 sg13g2_nor2b_1 _13718_ (.A(_05551_),
    .B_N(net608),
    .Y(_05552_));
 sg13g2_nor2b_1 _13719_ (.A(net608),
    .B_N(_05551_),
    .Y(_05553_));
 sg13g2_nor3_1 _13720_ (.A(_05474_),
    .B(_05552_),
    .C(_05553_),
    .Y(_05554_));
 sg13g2_a21oi_1 _13721_ (.A1(net406),
    .A2(_05550_),
    .Y(_05555_),
    .B1(_05554_));
 sg13g2_mux2_1 _13722_ (.A0(_05543_),
    .A1(_05555_),
    .S(net59),
    .X(_01283_));
 sg13g2_nor3_1 _13723_ (.A(_05534_),
    .B(_05543_),
    .C(net508),
    .Y(_05556_));
 sg13g2_nor3_1 _13724_ (.A(net608),
    .B(_05544_),
    .C(net439),
    .Y(_05557_));
 sg13g2_inv_1 _13725_ (.Y(_05558_),
    .A(_05533_));
 sg13g2_o21ai_1 _13726_ (.B1(_05558_),
    .Y(_05559_),
    .A1(_05556_),
    .A2(_05557_));
 sg13g2_buf_2 _13727_ (.A(\soc_I.div_reg[13] ),
    .X(_05560_));
 sg13g2_mux2_1 _13728_ (.A0(\soc_I.tx_uart_i.wait_states[13] ),
    .A1(_05560_),
    .S(net440),
    .X(_05561_));
 sg13g2_xnor2_1 _13729_ (.Y(_05562_),
    .A(_05559_),
    .B(_05561_));
 sg13g2_nand2b_1 _13730_ (.Y(_05563_),
    .B(_05544_),
    .A_N(_05553_));
 sg13g2_nand2b_1 _13731_ (.Y(_05564_),
    .B(_05553_),
    .A_N(_05544_));
 sg13g2_a21oi_1 _13732_ (.A1(_05563_),
    .A2(_05564_),
    .Y(_05565_),
    .B1(net405));
 sg13g2_a21oi_1 _13733_ (.A1(net406),
    .A2(_05562_),
    .Y(_05566_),
    .B1(_05565_));
 sg13g2_nor2_1 _13734_ (.A(\soc_I.tx_uart_i.wait_states[13] ),
    .B(net58),
    .Y(_05567_));
 sg13g2_a21oi_1 _13735_ (.A1(net59),
    .A2(_05566_),
    .Y(_01284_),
    .B1(_05567_));
 sg13g2_buf_2 _13736_ (.A(\soc_I.div_reg[14] ),
    .X(_05568_));
 sg13g2_or2_1 _13737_ (.X(_05569_),
    .B(_05561_),
    .A(_05559_));
 sg13g2_buf_1 _13738_ (.A(_05569_),
    .X(_05570_));
 sg13g2_xnor2_1 _13739_ (.Y(_05571_),
    .A(_05568_),
    .B(_05570_));
 sg13g2_xnor2_1 _13740_ (.Y(_05572_),
    .A(_05560_),
    .B(_05564_));
 sg13g2_buf_1 _13741_ (.A(\soc_I.tx_uart_i.wait_states[14] ),
    .X(_05573_));
 sg13g2_nor2_1 _13742_ (.A(_05573_),
    .B(_05570_),
    .Y(_05574_));
 sg13g2_nand2_1 _13743_ (.Y(_05575_),
    .A(_05573_),
    .B(_05570_));
 sg13g2_nand3b_1 _13744_ (.B(net610),
    .C(_05575_),
    .Y(_05576_),
    .A_N(_05574_));
 sg13g2_o21ai_1 _13745_ (.B1(_05576_),
    .Y(_05577_),
    .A1(net610),
    .A2(_05572_));
 sg13g2_nand2_1 _13746_ (.Y(_05578_),
    .A(net579),
    .B(_05577_));
 sg13g2_o21ai_1 _13747_ (.B1(_05578_),
    .Y(_05579_),
    .A1(net579),
    .A2(_05571_));
 sg13g2_nor2_1 _13748_ (.A(_05573_),
    .B(_05451_),
    .Y(_05580_));
 sg13g2_a21oi_1 _13749_ (.A1(net59),
    .A2(_05579_),
    .Y(_01285_),
    .B1(_05580_));
 sg13g2_buf_2 _13750_ (.A(\soc_I.div_reg[15] ),
    .X(_05581_));
 sg13g2_nor2_1 _13751_ (.A(_05568_),
    .B(_05570_),
    .Y(_05582_));
 sg13g2_xor2_1 _13752_ (.B(_05582_),
    .A(_05581_),
    .X(_05583_));
 sg13g2_xnor2_1 _13753_ (.Y(_05584_),
    .A(\soc_I.tx_uart_i.wait_states[15] ),
    .B(_05574_));
 sg13g2_nor2_1 _13754_ (.A(net440),
    .B(_05584_),
    .Y(_05585_));
 sg13g2_a21oi_1 _13755_ (.A1(net407),
    .A2(_05583_),
    .Y(_05586_),
    .B1(_05585_));
 sg13g2_nor2_1 _13756_ (.A(_05560_),
    .B(_05564_),
    .Y(_05587_));
 sg13g2_xor2_1 _13757_ (.B(_05587_),
    .A(_05568_),
    .X(_05588_));
 sg13g2_nor2_1 _13758_ (.A(net405),
    .B(_05588_),
    .Y(_05589_));
 sg13g2_a21oi_1 _13759_ (.A1(net406),
    .A2(_05586_),
    .Y(_05590_),
    .B1(_05589_));
 sg13g2_mux2_1 _13760_ (.A0(\soc_I.tx_uart_i.wait_states[15] ),
    .A1(_05590_),
    .S(net59),
    .X(_01286_));
 sg13g2_xnor2_1 _13761_ (.Y(_05591_),
    .A(_05463_),
    .B(_05502_));
 sg13g2_mux2_1 _13762_ (.A0(_00060_),
    .A1(_05591_),
    .S(net610),
    .X(_05592_));
 sg13g2_xor2_1 _13763_ (.B(_05500_),
    .A(_05468_),
    .X(_05593_));
 sg13g2_nor2_1 _13764_ (.A(net579),
    .B(_05593_),
    .Y(_05594_));
 sg13g2_a21oi_1 _13765_ (.A1(net579),
    .A2(_05592_),
    .Y(_05595_),
    .B1(_05594_));
 sg13g2_nor2_1 _13766_ (.A(_05502_),
    .B(_05451_),
    .Y(_05596_));
 sg13g2_a21oi_1 _13767_ (.A1(net59),
    .A2(_05595_),
    .Y(_01287_),
    .B1(_05596_));
 sg13g2_mux2_1 _13768_ (.A0(_05495_),
    .A1(_05497_),
    .S(net440),
    .X(_05597_));
 sg13g2_xor2_1 _13769_ (.B(_05597_),
    .A(_05504_),
    .X(_05598_));
 sg13g2_nor2b_1 _13770_ (.A(net405),
    .B_N(_05593_),
    .Y(_05599_));
 sg13g2_a21oi_1 _13771_ (.A1(net406),
    .A2(_05598_),
    .Y(_05600_),
    .B1(_05599_));
 sg13g2_mux2_1 _13772_ (.A0(_05495_),
    .A1(_05600_),
    .S(net58),
    .X(_01288_));
 sg13g2_nor2_1 _13773_ (.A(_05497_),
    .B(_05504_),
    .Y(_05601_));
 sg13g2_xor2_1 _13774_ (.B(_05601_),
    .A(_05498_),
    .X(_05602_));
 sg13g2_nor2_1 _13775_ (.A(_05495_),
    .B(_05504_),
    .Y(_05603_));
 sg13g2_xnor2_1 _13776_ (.Y(_05604_),
    .A(_05494_),
    .B(_05603_));
 sg13g2_nand2_1 _13777_ (.Y(_05605_),
    .A(net439),
    .B(_05604_));
 sg13g2_o21ai_1 _13778_ (.B1(_05605_),
    .Y(_05606_),
    .A1(net439),
    .A2(_05602_));
 sg13g2_nor2b_1 _13779_ (.A(_05501_),
    .B_N(_05497_),
    .Y(_05607_));
 sg13g2_nor3_1 _13780_ (.A(_05519_),
    .B(net405),
    .C(_05607_),
    .Y(_05608_));
 sg13g2_a21oi_1 _13781_ (.A1(net406),
    .A2(_05606_),
    .Y(_05609_),
    .B1(_05608_));
 sg13g2_mux2_1 _13782_ (.A0(_05494_),
    .A1(_05609_),
    .S(_05466_),
    .X(_01289_));
 sg13g2_mux2_1 _13783_ (.A0(_05489_),
    .A1(_05491_),
    .S(net440),
    .X(_05610_));
 sg13g2_xnor2_1 _13784_ (.Y(_05611_),
    .A(_05507_),
    .B(_05610_));
 sg13g2_xnor2_1 _13785_ (.Y(_05612_),
    .A(_05498_),
    .B(_05519_));
 sg13g2_nor2_1 _13786_ (.A(net405),
    .B(_05612_),
    .Y(_05613_));
 sg13g2_a21oi_1 _13787_ (.A1(net406),
    .A2(_05611_),
    .Y(_05614_),
    .B1(_05613_));
 sg13g2_nor2_1 _13788_ (.A(_05489_),
    .B(_05451_),
    .Y(_05615_));
 sg13g2_a21oi_1 _13789_ (.A1(_05465_),
    .A2(_05614_),
    .Y(_01290_),
    .B1(_05615_));
 sg13g2_nor2_1 _13790_ (.A(_05491_),
    .B(_05507_),
    .Y(_05616_));
 sg13g2_xor2_1 _13791_ (.B(_05616_),
    .A(_05492_),
    .X(_05617_));
 sg13g2_nor2_1 _13792_ (.A(_05489_),
    .B(_05507_),
    .Y(_05618_));
 sg13g2_xnor2_1 _13793_ (.Y(_05619_),
    .A(_05488_),
    .B(_05618_));
 sg13g2_nor2_1 _13794_ (.A(net440),
    .B(_05619_),
    .Y(_05620_));
 sg13g2_a21oi_1 _13795_ (.A1(net407),
    .A2(_05617_),
    .Y(_05621_),
    .B1(_05620_));
 sg13g2_nor2b_1 _13796_ (.A(_05520_),
    .B_N(_05491_),
    .Y(_05622_));
 sg13g2_nor3_1 _13797_ (.A(_05521_),
    .B(_05474_),
    .C(_05622_),
    .Y(_05623_));
 sg13g2_a21oi_1 _13798_ (.A1(net406),
    .A2(_05621_),
    .Y(_05624_),
    .B1(_05623_));
 sg13g2_mux2_1 _13799_ (.A0(_05488_),
    .A1(_05624_),
    .S(net58),
    .X(_01291_));
 sg13g2_mux2_1 _13800_ (.A0(_05483_),
    .A1(_05485_),
    .S(net440),
    .X(_05625_));
 sg13g2_xnor2_1 _13801_ (.Y(_05626_),
    .A(_05510_),
    .B(_05625_));
 sg13g2_xnor2_1 _13802_ (.Y(_05627_),
    .A(_05492_),
    .B(_05521_));
 sg13g2_nor2_1 _13803_ (.A(net405),
    .B(_05627_),
    .Y(_05628_));
 sg13g2_a21oi_1 _13804_ (.A1(net406),
    .A2(_05626_),
    .Y(_05629_),
    .B1(_05628_));
 sg13g2_nor2_1 _13805_ (.A(_05483_),
    .B(_05451_),
    .Y(_05630_));
 sg13g2_a21oi_1 _13806_ (.A1(_05465_),
    .A2(_05629_),
    .Y(_01292_),
    .B1(_05630_));
 sg13g2_nor2_1 _13807_ (.A(_05485_),
    .B(_05510_),
    .Y(_05631_));
 sg13g2_xor2_1 _13808_ (.B(_05631_),
    .A(_05486_),
    .X(_05632_));
 sg13g2_nor2_1 _13809_ (.A(_05483_),
    .B(_05510_),
    .Y(_05633_));
 sg13g2_xnor2_1 _13810_ (.Y(_05634_),
    .A(_05482_),
    .B(_05633_));
 sg13g2_nor2_1 _13811_ (.A(net440),
    .B(_05634_),
    .Y(_05635_));
 sg13g2_a21oi_1 _13812_ (.A1(net407),
    .A2(_05632_),
    .Y(_05636_),
    .B1(_05635_));
 sg13g2_nor2b_1 _13813_ (.A(_05522_),
    .B_N(_05485_),
    .Y(_05637_));
 sg13g2_nor3_1 _13814_ (.A(_05523_),
    .B(_05474_),
    .C(_05637_),
    .Y(_05638_));
 sg13g2_a21oi_1 _13815_ (.A1(net405),
    .A2(_05636_),
    .Y(_05639_),
    .B1(_05638_));
 sg13g2_mux2_1 _13816_ (.A0(_05482_),
    .A1(_05639_),
    .S(net58),
    .X(_01293_));
 sg13g2_xnor2_1 _13817_ (.Y(_05640_),
    .A(_05477_),
    .B(_05513_));
 sg13g2_nand2b_1 _13818_ (.Y(_05641_),
    .B(_05486_),
    .A_N(_05523_));
 sg13g2_a21oi_1 _13819_ (.A1(_05525_),
    .A2(_05641_),
    .Y(_05642_),
    .B1(net610));
 sg13g2_a21oi_1 _13820_ (.A1(net610),
    .A2(_05640_),
    .Y(_05643_),
    .B1(_05642_));
 sg13g2_and2_1 _13821_ (.A(net609),
    .B(_05513_),
    .X(_05644_));
 sg13g2_nor2_1 _13822_ (.A(net609),
    .B(_05513_),
    .Y(_05645_));
 sg13g2_nor3_1 _13823_ (.A(_05453_),
    .B(_05644_),
    .C(_05645_),
    .Y(_05646_));
 sg13g2_a21oi_1 _13824_ (.A1(_05453_),
    .A2(_05643_),
    .Y(_05647_),
    .B1(_05646_));
 sg13g2_mux2_1 _13825_ (.A0(_05477_),
    .A1(_05647_),
    .S(_05466_),
    .X(_01294_));
 sg13g2_xor2_1 _13826_ (.B(_05645_),
    .A(_05480_),
    .X(_05648_));
 sg13g2_nor2_1 _13827_ (.A(_05477_),
    .B(_05513_),
    .Y(_05649_));
 sg13g2_xnor2_1 _13828_ (.Y(_05650_),
    .A(_05476_),
    .B(_05649_));
 sg13g2_nor2_1 _13829_ (.A(_05441_),
    .B(_05650_),
    .Y(_05651_));
 sg13g2_a21oi_1 _13830_ (.A1(_05442_),
    .A2(_05648_),
    .Y(_05652_),
    .B1(_05651_));
 sg13g2_and2_1 _13831_ (.A(net609),
    .B(_05525_),
    .X(_05653_));
 sg13g2_nor3_1 _13832_ (.A(_05526_),
    .B(_05474_),
    .C(_05653_),
    .Y(_05654_));
 sg13g2_a21oi_1 _13833_ (.A1(net405),
    .A2(_05652_),
    .Y(_05655_),
    .B1(_05654_));
 sg13g2_mux2_1 _13834_ (.A0(_05476_),
    .A1(_05655_),
    .S(net58),
    .X(_01295_));
 sg13g2_inv_1 _13835_ (.Y(_05656_),
    .A(_00091_));
 sg13g2_buf_1 _13836_ (.A(\soc_I.spi0_I.div[9] ),
    .X(_05657_));
 sg13g2_buf_1 _13837_ (.A(\soc_I.spi0_I.tick_cnt[9] ),
    .X(_05658_));
 sg13g2_buf_1 _13838_ (.A(\soc_I.spi0_I.div[8] ),
    .X(_05659_));
 sg13g2_buf_1 _13839_ (.A(\soc_I.spi0_I.div[6] ),
    .X(_05660_));
 sg13g2_buf_1 _13840_ (.A(\soc_I.spi0_I.div[4] ),
    .X(_05661_));
 sg13g2_buf_1 _13841_ (.A(\soc_I.spi0_I.div[0] ),
    .X(_05662_));
 sg13g2_buf_1 _13842_ (.A(\soc_I.spi0_I.div[1] ),
    .X(_05663_));
 sg13g2_buf_1 _13843_ (.A(\soc_I.spi0_I.div[2] ),
    .X(_05664_));
 sg13g2_nor4_2 _13844_ (.A(_05662_),
    .B(_05663_),
    .C(_05664_),
    .Y(_05665_),
    .D(\soc_I.spi0_I.div[3] ));
 sg13g2_nor2b_1 _13845_ (.A(_05661_),
    .B_N(_05665_),
    .Y(_05666_));
 sg13g2_nor2b_1 _13846_ (.A(\soc_I.spi0_I.div[5] ),
    .B_N(_05666_),
    .Y(_05667_));
 sg13g2_nor2b_1 _13847_ (.A(_05660_),
    .B_N(_05667_),
    .Y(_05668_));
 sg13g2_nor2b_1 _13848_ (.A(\soc_I.spi0_I.div[7] ),
    .B_N(_05668_),
    .Y(_05669_));
 sg13g2_nor2b_1 _13849_ (.A(_05659_),
    .B_N(_05669_),
    .Y(_05670_));
 sg13g2_xor2_1 _13850_ (.B(_05670_),
    .A(_05658_),
    .X(_05671_));
 sg13g2_nor3_1 _13851_ (.A(_05657_),
    .B(_05658_),
    .C(_05670_),
    .Y(_05672_));
 sg13g2_a21oi_1 _13852_ (.A1(_05657_),
    .A2(_05671_),
    .Y(_05673_),
    .B1(_05672_));
 sg13g2_buf_1 _13853_ (.A(\soc_I.spi0_I.div[10] ),
    .X(_05674_));
 sg13g2_xnor2_1 _13854_ (.Y(_05675_),
    .A(_05674_),
    .B(\soc_I.spi0_I.tick_cnt[10] ));
 sg13g2_nor2b_1 _13855_ (.A(_05657_),
    .B_N(_05670_),
    .Y(_05676_));
 sg13g2_a21oi_1 _13856_ (.A1(_05658_),
    .A2(_05676_),
    .Y(_05677_),
    .B1(_05675_));
 sg13g2_a21oi_1 _13857_ (.A1(_05673_),
    .A2(_05675_),
    .Y(_05678_),
    .B1(_05677_));
 sg13g2_nor2_1 _13858_ (.A(_05662_),
    .B(_05663_),
    .Y(_05679_));
 sg13g2_buf_1 _13859_ (.A(\soc_I.spi0_I.tick_cnt[2] ),
    .X(_05680_));
 sg13g2_nor2b_1 _13860_ (.A(_05680_),
    .B_N(_05664_),
    .Y(_05681_));
 sg13g2_nor2b_1 _13861_ (.A(_05664_),
    .B_N(_05680_),
    .Y(_05682_));
 sg13g2_xor2_1 _13862_ (.B(\soc_I.spi0_I.tick_cnt[3] ),
    .A(\soc_I.spi0_I.div[3] ),
    .X(_05683_));
 sg13g2_mux2_1 _13863_ (.A0(_05681_),
    .A1(_05682_),
    .S(_05683_),
    .X(_05684_));
 sg13g2_nor4_1 _13864_ (.A(_05679_),
    .B(_05681_),
    .C(_05683_),
    .D(_05682_),
    .Y(_05685_));
 sg13g2_a21oi_1 _13865_ (.A1(_05679_),
    .A2(_05684_),
    .Y(_05686_),
    .B1(_05685_));
 sg13g2_buf_1 _13866_ (.A(\soc_I.spi0_I.tick_cnt[0] ),
    .X(_05687_));
 sg13g2_buf_1 _13867_ (.A(\soc_I.spi0_I.tick_cnt[1] ),
    .X(_05688_));
 sg13g2_xnor2_1 _13868_ (.Y(_05689_),
    .A(_05663_),
    .B(_05688_));
 sg13g2_nor2_1 _13869_ (.A(_05662_),
    .B(_05689_),
    .Y(_05690_));
 sg13g2_nor2b_1 _13870_ (.A(_05687_),
    .B_N(_05662_),
    .Y(_05691_));
 sg13g2_a22oi_1 _13871_ (.Y(_05692_),
    .B1(_05691_),
    .B2(_05689_),
    .A2(_05690_),
    .A1(_05687_));
 sg13g2_nor4_1 _13872_ (.A(\soc_I.spi0_I.tick_cnt[16] ),
    .B(\soc_I.spi0_I.tick_cnt[17] ),
    .C(_05686_),
    .D(_05692_),
    .Y(_05693_));
 sg13g2_buf_1 _13873_ (.A(\soc_I.spi0_I.tick_cnt[8] ),
    .X(_05694_));
 sg13g2_xor2_1 _13874_ (.B(_05694_),
    .A(_05659_),
    .X(_05695_));
 sg13g2_xnor2_1 _13875_ (.Y(_05696_),
    .A(_05669_),
    .B(_05695_));
 sg13g2_buf_2 _13876_ (.A(\soc_I.spi0_I.tick_cnt[4] ),
    .X(_05697_));
 sg13g2_xor2_1 _13877_ (.B(_05665_),
    .A(_05697_),
    .X(_05698_));
 sg13g2_nor3_1 _13878_ (.A(_05661_),
    .B(_05697_),
    .C(_05665_),
    .Y(_05699_));
 sg13g2_a21oi_1 _13879_ (.A1(_05661_),
    .A2(_05698_),
    .Y(_05700_),
    .B1(_05699_));
 sg13g2_buf_1 _13880_ (.A(\soc_I.spi0_I.tick_cnt[5] ),
    .X(_05701_));
 sg13g2_xnor2_1 _13881_ (.Y(_05702_),
    .A(\soc_I.spi0_I.div[5] ),
    .B(_05701_));
 sg13g2_a21oi_1 _13882_ (.A1(_05697_),
    .A2(_05666_),
    .Y(_05703_),
    .B1(_05702_));
 sg13g2_a21oi_1 _13883_ (.A1(_05700_),
    .A2(_05702_),
    .Y(_05704_),
    .B1(_05703_));
 sg13g2_buf_2 _13884_ (.A(\soc_I.spi0_I.tick_cnt[6] ),
    .X(_05705_));
 sg13g2_xor2_1 _13885_ (.B(_05667_),
    .A(_05705_),
    .X(_05706_));
 sg13g2_nor3_1 _13886_ (.A(_05660_),
    .B(_05705_),
    .C(_05667_),
    .Y(_05707_));
 sg13g2_a21oi_1 _13887_ (.A1(_05660_),
    .A2(_05706_),
    .Y(_05708_),
    .B1(_05707_));
 sg13g2_xor2_1 _13888_ (.B(\soc_I.spi0_I.tick_cnt[7] ),
    .A(\soc_I.spi0_I.div[7] ),
    .X(_05709_));
 sg13g2_nand3_1 _13889_ (.B(_05668_),
    .C(_05709_),
    .A(_05705_),
    .Y(_05710_));
 sg13g2_o21ai_1 _13890_ (.B1(_05710_),
    .Y(_05711_),
    .A1(_05708_),
    .A2(_05709_));
 sg13g2_nand4_1 _13891_ (.B(_05696_),
    .C(_05704_),
    .A(_05693_),
    .Y(_05712_),
    .D(_05711_));
 sg13g2_buf_1 _13892_ (.A(\soc_I.spi0_I.div[11] ),
    .X(_05713_));
 sg13g2_buf_1 _13893_ (.A(\soc_I.spi0_I.div[12] ),
    .X(_05714_));
 sg13g2_nand2b_1 _13894_ (.Y(_05715_),
    .B(_05676_),
    .A_N(_05674_));
 sg13g2_buf_1 _13895_ (.A(_05715_),
    .X(_05716_));
 sg13g2_nor3_1 _13896_ (.A(_05713_),
    .B(_05714_),
    .C(_05716_),
    .Y(_05717_));
 sg13g2_buf_1 _13897_ (.A(\soc_I.spi0_I.div[13] ),
    .X(_05718_));
 sg13g2_xnor2_1 _13898_ (.Y(_05719_),
    .A(_05718_),
    .B(\soc_I.spi0_I.tick_cnt[13] ));
 sg13g2_xnor2_1 _13899_ (.Y(_05720_),
    .A(_05717_),
    .B(_05719_));
 sg13g2_nor2_1 _13900_ (.A(_05712_),
    .B(_05720_),
    .Y(_05721_));
 sg13g2_buf_1 _13901_ (.A(\soc_I.spi0_I.tick_cnt[11] ),
    .X(_05722_));
 sg13g2_inv_1 _13902_ (.Y(_05723_),
    .A(_05722_));
 sg13g2_nand2_1 _13903_ (.Y(_05724_),
    .A(_05723_),
    .B(_05716_));
 sg13g2_xnor2_1 _13904_ (.Y(_05725_),
    .A(_05722_),
    .B(_05716_));
 sg13g2_nand2_1 _13905_ (.Y(_05726_),
    .A(_05713_),
    .B(_05725_));
 sg13g2_o21ai_1 _13906_ (.B1(_05726_),
    .Y(_05727_),
    .A1(_05713_),
    .A2(_05724_));
 sg13g2_xnor2_1 _13907_ (.Y(_05728_),
    .A(_05714_),
    .B(\soc_I.spi0_I.tick_cnt[12] ));
 sg13g2_nor4_1 _13908_ (.A(_05713_),
    .B(_05723_),
    .C(_05716_),
    .D(_05728_),
    .Y(_05729_));
 sg13g2_a21o_1 _13909_ (.A2(_05728_),
    .A1(_05727_),
    .B1(_05729_),
    .X(_05730_));
 sg13g2_buf_1 _13910_ (.A(\soc_I.spi0_I.div[15] ),
    .X(_05731_));
 sg13g2_buf_1 _13911_ (.A(\soc_I.spi0_I.tick_cnt[15] ),
    .X(_05732_));
 sg13g2_xor2_1 _13912_ (.B(_05732_),
    .A(_05731_),
    .X(_05733_));
 sg13g2_buf_1 _13913_ (.A(\soc_I.spi0_I.div[14] ),
    .X(_05734_));
 sg13g2_buf_1 _13914_ (.A(\soc_I.spi0_I.tick_cnt[14] ),
    .X(_05735_));
 sg13g2_nor2b_1 _13915_ (.A(_05718_),
    .B_N(_05717_),
    .Y(_05736_));
 sg13g2_xor2_1 _13916_ (.B(_05736_),
    .A(_05735_),
    .X(_05737_));
 sg13g2_nor3_1 _13917_ (.A(_05734_),
    .B(_05735_),
    .C(_05736_),
    .Y(_05738_));
 sg13g2_a21oi_1 _13918_ (.A1(_05734_),
    .A2(_05737_),
    .Y(_05739_),
    .B1(_05738_));
 sg13g2_inv_1 _13919_ (.Y(_05740_),
    .A(_05732_));
 sg13g2_nor2b_1 _13920_ (.A(_05734_),
    .B_N(_05736_),
    .Y(_05741_));
 sg13g2_nand4_1 _13921_ (.B(_05731_),
    .C(_05740_),
    .A(_05735_),
    .Y(_05742_),
    .D(_05741_));
 sg13g2_o21ai_1 _13922_ (.B1(_05742_),
    .Y(_05743_),
    .A1(_05733_),
    .A2(_05739_));
 sg13g2_nand4_1 _13923_ (.B(_05721_),
    .C(_05730_),
    .A(_05678_),
    .Y(_05744_),
    .D(_05743_));
 sg13g2_buf_1 _13924_ (.A(\soc_I.spi0_I.xfer_cycles[3] ),
    .X(_05745_));
 sg13g2_buf_1 _13925_ (.A(\soc_I.spi0_I.xfer_cycles[4] ),
    .X(_05746_));
 sg13g2_or2_1 _13926_ (.X(_05747_),
    .B(\soc_I.spi0_I.xfer_cycles[1] ),
    .A(\soc_I.spi0_I.xfer_cycles[0] ));
 sg13g2_or2_1 _13927_ (.X(_05748_),
    .B(_05747_),
    .A(\soc_I.spi0_I.xfer_cycles[2] ));
 sg13g2_buf_1 _13928_ (.A(_05748_),
    .X(_05749_));
 sg13g2_or4_1 _13929_ (.A(_05745_),
    .B(\soc_I.spi0_I.xfer_cycles[5] ),
    .C(_05746_),
    .D(_05749_),
    .X(_05750_));
 sg13g2_buf_2 _13930_ (.A(_05750_),
    .X(_05751_));
 sg13g2_nand3_1 _13931_ (.B(_05744_),
    .C(_05751_),
    .A(_04285_),
    .Y(_05752_));
 sg13g2_buf_1 _13932_ (.A(_05752_),
    .X(_05753_));
 sg13g2_buf_1 _13933_ (.A(net149),
    .X(_05754_));
 sg13g2_nor2_1 _13934_ (.A(_05656_),
    .B(net143),
    .Y(_01206_));
 sg13g2_inv_1 _13935_ (.Y(_05755_),
    .A(\soc_I.spi0_I.tick_cnt[10] ));
 sg13g2_inv_1 _13936_ (.Y(_05756_),
    .A(\soc_I.spi0_I.tick_cnt[7] ));
 sg13g2_inv_1 _13937_ (.Y(_05757_),
    .A(\soc_I.spi0_I.tick_cnt[3] ));
 sg13g2_nand3_1 _13938_ (.B(_05688_),
    .C(_05680_),
    .A(_05687_),
    .Y(_05758_));
 sg13g2_nor2_2 _13939_ (.A(_05757_),
    .B(_05758_),
    .Y(_05759_));
 sg13g2_nand4_1 _13940_ (.B(_05701_),
    .C(_05705_),
    .A(_05697_),
    .Y(_05760_),
    .D(_05759_));
 sg13g2_nor2_1 _13941_ (.A(_05756_),
    .B(_05760_),
    .Y(_05761_));
 sg13g2_nand3_1 _13942_ (.B(_05658_),
    .C(_05761_),
    .A(_05694_),
    .Y(_05762_));
 sg13g2_xnor2_1 _13943_ (.Y(_05763_),
    .A(_05755_),
    .B(_05762_));
 sg13g2_nor2_1 _13944_ (.A(net143),
    .B(_05763_),
    .Y(_01207_));
 sg13g2_nor2_1 _13945_ (.A(_05755_),
    .B(_05762_),
    .Y(_05764_));
 sg13g2_xnor2_1 _13946_ (.Y(_05765_),
    .A(_05722_),
    .B(_05764_));
 sg13g2_nor2_1 _13947_ (.A(net143),
    .B(_05765_),
    .Y(_01208_));
 sg13g2_nand2_1 _13948_ (.Y(_05766_),
    .A(_05722_),
    .B(_05764_));
 sg13g2_xor2_1 _13949_ (.B(_05766_),
    .A(\soc_I.spi0_I.tick_cnt[12] ),
    .X(_05767_));
 sg13g2_nor2_1 _13950_ (.A(net143),
    .B(_05767_),
    .Y(_01209_));
 sg13g2_inv_1 _13951_ (.Y(_05768_),
    .A(\soc_I.spi0_I.tick_cnt[13] ));
 sg13g2_nand3_1 _13952_ (.B(\soc_I.spi0_I.tick_cnt[12] ),
    .C(_05764_),
    .A(_05722_),
    .Y(_05769_));
 sg13g2_xnor2_1 _13953_ (.Y(_05770_),
    .A(_05768_),
    .B(_05769_));
 sg13g2_nor2_1 _13954_ (.A(net143),
    .B(_05770_),
    .Y(_01210_));
 sg13g2_nor2_1 _13955_ (.A(_05768_),
    .B(_05769_),
    .Y(_05771_));
 sg13g2_xnor2_1 _13956_ (.Y(_05772_),
    .A(_05735_),
    .B(_05771_));
 sg13g2_nor2_1 _13957_ (.A(net143),
    .B(_05772_),
    .Y(_01211_));
 sg13g2_and3_1 _13958_ (.X(_05773_),
    .A(_05735_),
    .B(_05751_),
    .C(_05771_));
 sg13g2_buf_1 _13959_ (.A(_05773_),
    .X(_05774_));
 sg13g2_xnor2_1 _13960_ (.Y(_05775_),
    .A(_05732_),
    .B(_05774_));
 sg13g2_nor2_1 _13961_ (.A(net143),
    .B(_05775_),
    .Y(_01212_));
 sg13g2_nand2_1 _13962_ (.Y(_05776_),
    .A(_05732_),
    .B(_05774_));
 sg13g2_xor2_1 _13963_ (.B(_05776_),
    .A(\soc_I.spi0_I.tick_cnt[16] ),
    .X(_05777_));
 sg13g2_nor2_1 _13964_ (.A(net143),
    .B(_05777_),
    .Y(_01213_));
 sg13g2_nand3_1 _13965_ (.B(\soc_I.spi0_I.tick_cnt[16] ),
    .C(_05774_),
    .A(_05732_),
    .Y(_05778_));
 sg13g2_xor2_1 _13966_ (.B(_05778_),
    .A(\soc_I.spi0_I.tick_cnt[17] ),
    .X(_05779_));
 sg13g2_nor2_1 _13967_ (.A(_05754_),
    .B(_05779_),
    .Y(_01214_));
 sg13g2_xnor2_1 _13968_ (.Y(_05780_),
    .A(_05687_),
    .B(_05688_));
 sg13g2_nor2_1 _13969_ (.A(_05754_),
    .B(_05780_),
    .Y(_01215_));
 sg13g2_nand2_1 _13970_ (.Y(_05781_),
    .A(_05687_),
    .B(_05688_));
 sg13g2_xor2_1 _13971_ (.B(_05781_),
    .A(_05680_),
    .X(_05782_));
 sg13g2_nor2_1 _13972_ (.A(net149),
    .B(_05782_),
    .Y(_01216_));
 sg13g2_xnor2_1 _13973_ (.Y(_05783_),
    .A(_05757_),
    .B(_05758_));
 sg13g2_nor2_1 _13974_ (.A(net149),
    .B(_05783_),
    .Y(_01217_));
 sg13g2_xnor2_1 _13975_ (.Y(_05784_),
    .A(_05697_),
    .B(_05759_));
 sg13g2_nor2_1 _13976_ (.A(net149),
    .B(_05784_),
    .Y(_01218_));
 sg13g2_nand2_1 _13977_ (.Y(_05785_),
    .A(_05697_),
    .B(_05759_));
 sg13g2_xor2_1 _13978_ (.B(_05785_),
    .A(_05701_),
    .X(_05786_));
 sg13g2_nor2_1 _13979_ (.A(_05753_),
    .B(_05786_),
    .Y(_01219_));
 sg13g2_nand3_1 _13980_ (.B(_05701_),
    .C(_05759_),
    .A(_05697_),
    .Y(_05787_));
 sg13g2_xor2_1 _13981_ (.B(_05787_),
    .A(_05705_),
    .X(_05788_));
 sg13g2_nor2_1 _13982_ (.A(net149),
    .B(_05788_),
    .Y(_01220_));
 sg13g2_xnor2_1 _13983_ (.Y(_05789_),
    .A(_05756_),
    .B(_05760_));
 sg13g2_nor2_1 _13984_ (.A(net149),
    .B(_05789_),
    .Y(_01221_));
 sg13g2_xnor2_1 _13985_ (.Y(_05790_),
    .A(_05694_),
    .B(_05761_));
 sg13g2_nor2_1 _13986_ (.A(net149),
    .B(_05790_),
    .Y(_01222_));
 sg13g2_nand2_1 _13987_ (.Y(_05791_),
    .A(_05694_),
    .B(_05761_));
 sg13g2_xor2_1 _13988_ (.B(_05791_),
    .A(_05658_),
    .X(_05792_));
 sg13g2_nor2_1 _13989_ (.A(net149),
    .B(_05792_),
    .Y(_01223_));
 sg13g2_buf_1 _13990_ (.A(_00050_),
    .X(_05793_));
 sg13g2_nor2b_1 _13991_ (.A(_05339_),
    .B_N(_05343_),
    .Y(_05794_));
 sg13g2_buf_1 _13992_ (.A(_05794_),
    .X(_05795_));
 sg13g2_buf_1 _13993_ (.A(\soc_I.rx_uart_i.fifo_i.rd_ptr[0] ),
    .X(_05796_));
 sg13g2_o21ai_1 _13994_ (.B1(_05796_),
    .Y(_05797_),
    .A1(_05793_),
    .A2(_05795_));
 sg13g2_nor2_1 _13995_ (.A(_05793_),
    .B(_05795_),
    .Y(_05798_));
 sg13g2_buf_2 _13996_ (.A(_05798_),
    .X(_05799_));
 sg13g2_nand2b_1 _13997_ (.Y(_05800_),
    .B(_05799_),
    .A_N(_05796_));
 sg13g2_buf_1 _13998_ (.A(_04267_),
    .X(_05801_));
 sg13g2_a21oi_1 _13999_ (.A1(_05797_),
    .A2(_05800_),
    .Y(_00093_),
    .B1(net404));
 sg13g2_buf_1 _14000_ (.A(net520),
    .X(_05802_));
 sg13g2_buf_1 _14001_ (.A(net438),
    .X(_05803_));
 sg13g2_nand2_1 _14002_ (.Y(_05804_),
    .A(_05796_),
    .B(_05799_));
 sg13g2_xor2_1 _14003_ (.B(_05804_),
    .A(\soc_I.rx_uart_i.fifo_i.rd_ptr[1] ),
    .X(_05805_));
 sg13g2_nor2_1 _14004_ (.A(net403),
    .B(_05805_),
    .Y(_00094_));
 sg13g2_nand3_1 _14005_ (.B(\soc_I.rx_uart_i.fifo_i.rd_ptr[1] ),
    .C(_05799_),
    .A(_05796_),
    .Y(_05806_));
 sg13g2_xor2_1 _14006_ (.B(_05806_),
    .A(\soc_I.rx_uart_i.fifo_i.rd_ptr[2] ),
    .X(_05807_));
 sg13g2_nor2_1 _14007_ (.A(net403),
    .B(_05807_),
    .Y(_00095_));
 sg13g2_nand4_1 _14008_ (.B(\soc_I.rx_uart_i.fifo_i.rd_ptr[1] ),
    .C(\soc_I.rx_uart_i.fifo_i.rd_ptr[2] ),
    .A(_05796_),
    .Y(_05808_),
    .D(_05799_));
 sg13g2_xor2_1 _14009_ (.B(_05808_),
    .A(\soc_I.rx_uart_i.fifo_i.rd_ptr[3] ),
    .X(_05809_));
 sg13g2_nor2_1 _14010_ (.A(net403),
    .B(_05809_),
    .Y(_00096_));
 sg13g2_buf_1 _14011_ (.A(_03578_),
    .X(_05810_));
 sg13g2_and2_1 _14012_ (.A(net437),
    .B(_00087_),
    .X(_00097_));
 sg13g2_buf_1 _14013_ (.A(\soc_I.cycle_cnt[9] ),
    .X(_05811_));
 sg13g2_inv_1 _14014_ (.Y(_05812_),
    .A(\soc_I.cycle_cnt[8] ));
 sg13g2_buf_1 _14015_ (.A(\soc_I.cycle_cnt[6] ),
    .X(_05813_));
 sg13g2_buf_1 _14016_ (.A(\soc_I.cycle_cnt[0] ),
    .X(_05814_));
 sg13g2_buf_1 _14017_ (.A(\soc_I.cycle_cnt[1] ),
    .X(_05815_));
 sg13g2_buf_1 _14018_ (.A(\soc_I.cycle_cnt[2] ),
    .X(_05816_));
 sg13g2_and4_1 _14019_ (.A(_05814_),
    .B(_05815_),
    .C(_05816_),
    .D(\soc_I.cycle_cnt[3] ),
    .X(_05817_));
 sg13g2_and2_1 _14020_ (.A(\soc_I.cycle_cnt[4] ),
    .B(_05817_),
    .X(_05818_));
 sg13g2_and2_1 _14021_ (.A(\soc_I.cycle_cnt[5] ),
    .B(_05818_),
    .X(_05819_));
 sg13g2_buf_1 _14022_ (.A(_05819_),
    .X(_05820_));
 sg13g2_nand3_1 _14023_ (.B(\soc_I.cycle_cnt[7] ),
    .C(_05820_),
    .A(_05813_),
    .Y(_05821_));
 sg13g2_nor2_1 _14024_ (.A(_05812_),
    .B(_05821_),
    .Y(_05822_));
 sg13g2_nand2_1 _14025_ (.Y(_05823_),
    .A(_05811_),
    .B(_05822_));
 sg13g2_xor2_1 _14026_ (.B(_05823_),
    .A(\soc_I.cycle_cnt[10] ),
    .X(_05824_));
 sg13g2_nor2_1 _14027_ (.A(net403),
    .B(_05824_),
    .Y(_00098_));
 sg13g2_buf_1 _14028_ (.A(\soc_I.cycle_cnt[11] ),
    .X(_05825_));
 sg13g2_and3_1 _14029_ (.X(_05826_),
    .A(_05811_),
    .B(\soc_I.cycle_cnt[10] ),
    .C(_05822_));
 sg13g2_buf_1 _14030_ (.A(_05826_),
    .X(_05827_));
 sg13g2_xnor2_1 _14031_ (.Y(_05828_),
    .A(_05825_),
    .B(_05827_));
 sg13g2_nor2_1 _14032_ (.A(net403),
    .B(_05828_),
    .Y(_00099_));
 sg13g2_nand2_1 _14033_ (.Y(_05829_),
    .A(_05825_),
    .B(_05827_));
 sg13g2_xor2_1 _14034_ (.B(_05829_),
    .A(\soc_I.cycle_cnt[12] ),
    .X(_05830_));
 sg13g2_nor2_1 _14035_ (.A(net403),
    .B(_05830_),
    .Y(_00100_));
 sg13g2_inv_1 _14036_ (.Y(_05831_),
    .A(\soc_I.cycle_cnt[13] ));
 sg13g2_nand3_1 _14037_ (.B(\soc_I.cycle_cnt[12] ),
    .C(_05827_),
    .A(_05825_),
    .Y(_05832_));
 sg13g2_xnor2_1 _14038_ (.Y(_05833_),
    .A(_05831_),
    .B(_05832_));
 sg13g2_nor2_1 _14039_ (.A(net403),
    .B(_05833_),
    .Y(_00101_));
 sg13g2_buf_1 _14040_ (.A(\soc_I.cycle_cnt[14] ),
    .X(_05834_));
 sg13g2_nor2_2 _14041_ (.A(_05831_),
    .B(_05832_),
    .Y(_05835_));
 sg13g2_xnor2_1 _14042_ (.Y(_05836_),
    .A(_05834_),
    .B(_05835_));
 sg13g2_nor2_1 _14043_ (.A(net403),
    .B(_05836_),
    .Y(_00102_));
 sg13g2_buf_1 _14044_ (.A(\soc_I.cycle_cnt[15] ),
    .X(_05837_));
 sg13g2_nand2_1 _14045_ (.Y(_05838_),
    .A(_05834_),
    .B(_05835_));
 sg13g2_xor2_1 _14046_ (.B(_05838_),
    .A(_05837_),
    .X(_05839_));
 sg13g2_nor2_1 _14047_ (.A(_05803_),
    .B(_05839_),
    .Y(_00103_));
 sg13g2_nand3_1 _14048_ (.B(_05837_),
    .C(_05835_),
    .A(_05834_),
    .Y(_05840_));
 sg13g2_xor2_1 _14049_ (.B(_05840_),
    .A(\soc_I.cycle_cnt[16] ),
    .X(_05841_));
 sg13g2_nor2_1 _14050_ (.A(_05803_),
    .B(_05841_),
    .Y(_00104_));
 sg13g2_buf_1 _14051_ (.A(net438),
    .X(_05842_));
 sg13g2_inv_1 _14052_ (.Y(_05843_),
    .A(\soc_I.cycle_cnt[17] ));
 sg13g2_nand4_1 _14053_ (.B(_05837_),
    .C(\soc_I.cycle_cnt[16] ),
    .A(_05834_),
    .Y(_05844_),
    .D(_05835_));
 sg13g2_xnor2_1 _14054_ (.Y(_05845_),
    .A(_05843_),
    .B(_05844_));
 sg13g2_nor2_1 _14055_ (.A(_05842_),
    .B(_05845_),
    .Y(_00105_));
 sg13g2_buf_1 _14056_ (.A(\soc_I.cycle_cnt[18] ),
    .X(_05846_));
 sg13g2_nor2_1 _14057_ (.A(_05843_),
    .B(_05844_),
    .Y(_05847_));
 sg13g2_xnor2_1 _14058_ (.Y(_05848_),
    .A(_05846_),
    .B(_05847_));
 sg13g2_nor2_1 _14059_ (.A(net402),
    .B(_05848_),
    .Y(_00106_));
 sg13g2_nand2_1 _14060_ (.Y(_05849_),
    .A(_05846_),
    .B(_05847_));
 sg13g2_xor2_1 _14061_ (.B(_05849_),
    .A(\soc_I.cycle_cnt[19] ),
    .X(_05850_));
 sg13g2_nor2_1 _14062_ (.A(net402),
    .B(_05850_),
    .Y(_00107_));
 sg13g2_xnor2_1 _14063_ (.Y(_05851_),
    .A(_05814_),
    .B(_05815_));
 sg13g2_nor2_1 _14064_ (.A(_05842_),
    .B(_05851_),
    .Y(_00108_));
 sg13g2_inv_1 _14065_ (.Y(_05852_),
    .A(\soc_I.cycle_cnt[20] ));
 sg13g2_nand3_1 _14066_ (.B(\soc_I.cycle_cnt[19] ),
    .C(_05847_),
    .A(_05846_),
    .Y(_05853_));
 sg13g2_xnor2_1 _14067_ (.Y(_05854_),
    .A(_05852_),
    .B(_05853_));
 sg13g2_nor2_1 _14068_ (.A(net402),
    .B(_05854_),
    .Y(_00109_));
 sg13g2_buf_1 _14069_ (.A(\soc_I.cycle_cnt[21] ),
    .X(_05855_));
 sg13g2_nor2_1 _14070_ (.A(_05852_),
    .B(_05853_),
    .Y(_05856_));
 sg13g2_xnor2_1 _14071_ (.Y(_05857_),
    .A(_05855_),
    .B(_05856_));
 sg13g2_nor2_1 _14072_ (.A(net402),
    .B(_05857_),
    .Y(_00110_));
 sg13g2_nand2_1 _14073_ (.Y(_05858_),
    .A(_05855_),
    .B(_05856_));
 sg13g2_xor2_1 _14074_ (.B(_05858_),
    .A(\soc_I.cycle_cnt[22] ),
    .X(_05859_));
 sg13g2_nor2_1 _14075_ (.A(net402),
    .B(_05859_),
    .Y(_00111_));
 sg13g2_inv_1 _14076_ (.Y(_05860_),
    .A(\soc_I.cycle_cnt[23] ));
 sg13g2_nand3_1 _14077_ (.B(\soc_I.cycle_cnt[22] ),
    .C(_05856_),
    .A(_05855_),
    .Y(_05861_));
 sg13g2_xnor2_1 _14078_ (.Y(_05862_),
    .A(_05860_),
    .B(_05861_));
 sg13g2_nor2_1 _14079_ (.A(net402),
    .B(_05862_),
    .Y(_00112_));
 sg13g2_buf_1 _14080_ (.A(\soc_I.cycle_cnt[24] ),
    .X(_05863_));
 sg13g2_nor2_1 _14081_ (.A(_05860_),
    .B(_05861_),
    .Y(_05864_));
 sg13g2_xnor2_1 _14082_ (.Y(_05865_),
    .A(_05863_),
    .B(_05864_));
 sg13g2_nor2_1 _14083_ (.A(net402),
    .B(_05865_),
    .Y(_00113_));
 sg13g2_nand2_1 _14084_ (.Y(_05866_),
    .A(_05863_),
    .B(_05864_));
 sg13g2_xor2_1 _14085_ (.B(_05866_),
    .A(\soc_I.cycle_cnt[25] ),
    .X(_05867_));
 sg13g2_nor2_1 _14086_ (.A(net402),
    .B(_05867_),
    .Y(_00114_));
 sg13g2_buf_1 _14087_ (.A(net438),
    .X(_05868_));
 sg13g2_inv_1 _14088_ (.Y(_05869_),
    .A(\soc_I.cycle_cnt[26] ));
 sg13g2_nand3_1 _14089_ (.B(\soc_I.cycle_cnt[25] ),
    .C(_05864_),
    .A(_05863_),
    .Y(_05870_));
 sg13g2_xnor2_1 _14090_ (.Y(_05871_),
    .A(_05869_),
    .B(_05870_));
 sg13g2_nor2_1 _14091_ (.A(net401),
    .B(_05871_),
    .Y(_00115_));
 sg13g2_buf_1 _14092_ (.A(\soc_I.cycle_cnt[27] ),
    .X(_05872_));
 sg13g2_nor2_2 _14093_ (.A(_05869_),
    .B(_05870_),
    .Y(_05873_));
 sg13g2_xnor2_1 _14094_ (.Y(_05874_),
    .A(_05872_),
    .B(_05873_));
 sg13g2_nor2_1 _14095_ (.A(net401),
    .B(_05874_),
    .Y(_00116_));
 sg13g2_buf_1 _14096_ (.A(\soc_I.cycle_cnt[28] ),
    .X(_05875_));
 sg13g2_nand2_1 _14097_ (.Y(_05876_),
    .A(_05872_),
    .B(_05873_));
 sg13g2_xor2_1 _14098_ (.B(_05876_),
    .A(_05875_),
    .X(_05877_));
 sg13g2_nor2_1 _14099_ (.A(net401),
    .B(_05877_),
    .Y(_00117_));
 sg13g2_nand3_1 _14100_ (.B(_05875_),
    .C(_05873_),
    .A(_05872_),
    .Y(_05878_));
 sg13g2_xor2_1 _14101_ (.B(_05878_),
    .A(\soc_I.cycle_cnt[29] ),
    .X(_05879_));
 sg13g2_nor2_1 _14102_ (.A(net401),
    .B(_05879_),
    .Y(_00118_));
 sg13g2_nand2_1 _14103_ (.Y(_05880_),
    .A(_05814_),
    .B(_05815_));
 sg13g2_xor2_1 _14104_ (.B(_05880_),
    .A(_05816_),
    .X(_05881_));
 sg13g2_nor2_1 _14105_ (.A(net401),
    .B(_05881_),
    .Y(_00119_));
 sg13g2_inv_1 _14106_ (.Y(_05882_),
    .A(\soc_I.cycle_cnt[30] ));
 sg13g2_nand4_1 _14107_ (.B(_05875_),
    .C(\soc_I.cycle_cnt[29] ),
    .A(_05872_),
    .Y(_05883_),
    .D(_05873_));
 sg13g2_xnor2_1 _14108_ (.Y(_05884_),
    .A(_05882_),
    .B(_05883_));
 sg13g2_nor2_1 _14109_ (.A(net401),
    .B(_05884_),
    .Y(_00120_));
 sg13g2_nor2_1 _14110_ (.A(_05882_),
    .B(_05883_),
    .Y(_05885_));
 sg13g2_xnor2_1 _14111_ (.Y(_05886_),
    .A(\soc_I.cycle_cnt[31] ),
    .B(_05885_));
 sg13g2_nor2_1 _14112_ (.A(net401),
    .B(_05886_),
    .Y(_00121_));
 sg13g2_nand3_1 _14113_ (.B(_05815_),
    .C(_05816_),
    .A(_05814_),
    .Y(_05887_));
 sg13g2_xor2_1 _14114_ (.B(_05887_),
    .A(\soc_I.cycle_cnt[3] ),
    .X(_05888_));
 sg13g2_nor2_1 _14115_ (.A(net401),
    .B(_05888_),
    .Y(_00122_));
 sg13g2_xnor2_1 _14116_ (.Y(_05889_),
    .A(\soc_I.cycle_cnt[4] ),
    .B(_05817_));
 sg13g2_nor2_1 _14117_ (.A(_05868_),
    .B(_05889_),
    .Y(_00123_));
 sg13g2_xnor2_1 _14118_ (.Y(_05890_),
    .A(\soc_I.cycle_cnt[5] ),
    .B(_05818_));
 sg13g2_nor2_1 _14119_ (.A(_05868_),
    .B(_05890_),
    .Y(_00124_));
 sg13g2_buf_1 _14120_ (.A(net438),
    .X(_05891_));
 sg13g2_xnor2_1 _14121_ (.Y(_05892_),
    .A(_05813_),
    .B(_05820_));
 sg13g2_nor2_1 _14122_ (.A(net400),
    .B(_05892_),
    .Y(_00125_));
 sg13g2_nand2_1 _14123_ (.Y(_05893_),
    .A(_05813_),
    .B(_05820_));
 sg13g2_xor2_1 _14124_ (.B(_05893_),
    .A(\soc_I.cycle_cnt[7] ),
    .X(_05894_));
 sg13g2_nor2_1 _14125_ (.A(net400),
    .B(_05894_),
    .Y(_00126_));
 sg13g2_xnor2_1 _14126_ (.Y(_05895_),
    .A(_05812_),
    .B(_05821_));
 sg13g2_nor2_1 _14127_ (.A(_05891_),
    .B(_05895_),
    .Y(_00127_));
 sg13g2_xnor2_1 _14128_ (.Y(_05896_),
    .A(_05811_),
    .B(_05822_));
 sg13g2_nor2_1 _14129_ (.A(_05891_),
    .B(_05896_),
    .Y(_00128_));
 sg13g2_nand2_1 _14130_ (.Y(_05897_),
    .A(_04116_),
    .B(_04188_));
 sg13g2_buf_1 _14131_ (.A(_05897_),
    .X(_05898_));
 sg13g2_nand2_1 _14132_ (.Y(_05899_),
    .A(_03788_),
    .B(_05898_));
 sg13g2_or3_1 _14133_ (.A(\soc_I.cpu_mem_addr[1] ),
    .B(_04223_),
    .C(_04240_),
    .X(_05900_));
 sg13g2_nand2_1 _14134_ (.Y(_05901_),
    .A(net596),
    .B(net76));
 sg13g2_nor4_1 _14135_ (.A(_05899_),
    .B(_04246_),
    .C(_05900_),
    .D(_05901_),
    .Y(_00129_));
 sg13g2_buf_1 _14136_ (.A(_04102_),
    .X(_05902_));
 sg13g2_buf_1 _14137_ (.A(net578),
    .X(_05903_));
 sg13g2_buf_1 _14138_ (.A(net507),
    .X(_05904_));
 sg13g2_buf_1 _14139_ (.A(_05904_),
    .X(_05905_));
 sg13g2_or3_1 _14140_ (.A(_05899_),
    .B(_04223_),
    .C(_04240_),
    .X(_05906_));
 sg13g2_buf_1 _14141_ (.A(_05906_),
    .X(_05907_));
 sg13g2_or2_1 _14142_ (.X(_05908_),
    .B(_05901_),
    .A(_03855_));
 sg13g2_nor3_1 _14143_ (.A(net399),
    .B(_05907_),
    .C(_05908_),
    .Y(_00130_));
 sg13g2_buf_1 _14144_ (.A(net515),
    .X(_05909_));
 sg13g2_buf_1 _14145_ (.A(\soc_I.cpu_mem_wdata[0] ),
    .X(_05910_));
 sg13g2_buf_1 _14146_ (.A(net578),
    .X(_05911_));
 sg13g2_nor2_2 _14147_ (.A(\soc_I.cpu_mem_addr[0] ),
    .B(_03835_),
    .Y(_05912_));
 sg13g2_nand2_1 _14148_ (.Y(_05913_),
    .A(_04225_),
    .B(_05912_));
 sg13g2_or4_1 _14149_ (.A(net506),
    .B(_03851_),
    .C(_05907_),
    .D(_05913_),
    .X(_05914_));
 sg13g2_buf_1 _14150_ (.A(_05914_),
    .X(_05915_));
 sg13g2_buf_8 _14151_ (.A(_05915_),
    .X(_05916_));
 sg13g2_mux2_1 _14152_ (.A0(net607),
    .A1(_05468_),
    .S(net50),
    .X(_05917_));
 sg13g2_and2_1 _14153_ (.A(net435),
    .B(_05917_),
    .X(_00131_));
 sg13g2_buf_1 _14154_ (.A(_04266_),
    .X(_05918_));
 sg13g2_buf_1 _14155_ (.A(_05918_),
    .X(_05919_));
 sg13g2_buf_1 _14156_ (.A(_05915_),
    .X(_05920_));
 sg13g2_nor2b_1 _14157_ (.A(_05516_),
    .B_N(net49),
    .Y(_05921_));
 sg13g2_buf_1 _14158_ (.A(net50),
    .X(_05922_));
 sg13g2_nor2_1 _14159_ (.A(_01609_),
    .B(net630),
    .Y(_05923_));
 sg13g2_buf_2 _14160_ (.A(_05923_),
    .X(_05924_));
 sg13g2_mux2_1 _14161_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[10] ),
    .A1(net619),
    .S(_05924_),
    .X(_05925_));
 sg13g2_buf_1 _14162_ (.A(_05925_),
    .X(_05926_));
 sg13g2_nor2_1 _14163_ (.A(net43),
    .B(_05926_),
    .Y(_05927_));
 sg13g2_nor3_1 _14164_ (.A(net398),
    .B(_05921_),
    .C(_05927_),
    .Y(_00132_));
 sg13g2_nor2b_1 _14165_ (.A(net608),
    .B_N(net49),
    .Y(_05928_));
 sg13g2_buf_2 _14166_ (.A(\soc_I.cpu_mem_wdata[3] ),
    .X(_05929_));
 sg13g2_mux2_1 _14167_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[11] ),
    .A1(_05929_),
    .S(_05924_),
    .X(_05930_));
 sg13g2_buf_1 _14168_ (.A(_05930_),
    .X(_05931_));
 sg13g2_nor2_1 _14169_ (.A(_05922_),
    .B(_05931_),
    .Y(_05932_));
 sg13g2_nor3_1 _14170_ (.A(net398),
    .B(_05928_),
    .C(_05932_),
    .Y(_00133_));
 sg13g2_nor2b_1 _14171_ (.A(_05544_),
    .B_N(net49),
    .Y(_05933_));
 sg13g2_buf_8 _14172_ (.A(net50),
    .X(_05934_));
 sg13g2_buf_1 _14173_ (.A(\soc_I.cpu_mem_wdata[4] ),
    .X(_05935_));
 sg13g2_buf_1 _14174_ (.A(_05924_),
    .X(_05936_));
 sg13g2_mux2_1 _14175_ (.A0(_01856_),
    .A1(net606),
    .S(net397),
    .X(_05937_));
 sg13g2_nor2_1 _14176_ (.A(net42),
    .B(_05937_),
    .Y(_05938_));
 sg13g2_nor3_1 _14177_ (.A(net398),
    .B(_05933_),
    .C(_05938_),
    .Y(_00134_));
 sg13g2_buf_1 _14178_ (.A(_05918_),
    .X(_05939_));
 sg13g2_nor2b_1 _14179_ (.A(_05560_),
    .B_N(net49),
    .Y(_05940_));
 sg13g2_buf_2 _14180_ (.A(\soc_I.cpu_mem_wdata[5] ),
    .X(_05941_));
 sg13g2_mux2_1 _14181_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[13] ),
    .A1(_05941_),
    .S(_05924_),
    .X(_05942_));
 sg13g2_buf_1 _14182_ (.A(_05942_),
    .X(_05943_));
 sg13g2_nor2_1 _14183_ (.A(net42),
    .B(_05943_),
    .Y(_05944_));
 sg13g2_nor3_1 _14184_ (.A(net396),
    .B(_05940_),
    .C(_05944_),
    .Y(_00135_));
 sg13g2_nor2b_1 _14185_ (.A(_05568_),
    .B_N(net49),
    .Y(_05945_));
 sg13g2_buf_2 _14186_ (.A(\soc_I.cpu_mem_wdata[6] ),
    .X(_05946_));
 sg13g2_nor2_1 _14187_ (.A(_01893_),
    .B(_05924_),
    .Y(_05947_));
 sg13g2_a21o_1 _14188_ (.A2(net397),
    .A1(_05946_),
    .B1(_05947_),
    .X(_05948_));
 sg13g2_nor2_1 _14189_ (.A(_05934_),
    .B(_05948_),
    .Y(_05949_));
 sg13g2_nor3_1 _14190_ (.A(net396),
    .B(_05945_),
    .C(_05949_),
    .Y(_00136_));
 sg13g2_nor2b_1 _14191_ (.A(_05581_),
    .B_N(net49),
    .Y(_05950_));
 sg13g2_buf_1 _14192_ (.A(\soc_I.cpu_mem_wdata[7] ),
    .X(_05951_));
 sg13g2_mux2_1 _14193_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[15] ),
    .A1(net605),
    .S(_05924_),
    .X(_05952_));
 sg13g2_buf_1 _14194_ (.A(_05952_),
    .X(_05953_));
 sg13g2_nor2_1 _14195_ (.A(_05934_),
    .B(_05953_),
    .Y(_05954_));
 sg13g2_nor3_1 _14196_ (.A(net396),
    .B(_05950_),
    .C(_05954_),
    .Y(_00137_));
 sg13g2_nor2b_1 _14197_ (.A(\soc_I.div_reg[16] ),
    .B_N(_05920_),
    .Y(_05955_));
 sg13g2_buf_1 _14198_ (.A(_01609_),
    .X(_05956_));
 sg13g2_buf_1 _14199_ (.A(net505),
    .X(_05957_));
 sg13g2_mux2_1 _14200_ (.A0(net607),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[16] ),
    .S(net434),
    .X(_05958_));
 sg13g2_nor2_1 _14201_ (.A(net42),
    .B(_05958_),
    .Y(_05959_));
 sg13g2_nor3_1 _14202_ (.A(_05939_),
    .B(_05955_),
    .C(_05959_),
    .Y(_00138_));
 sg13g2_nor2b_1 _14203_ (.A(\soc_I.div_reg[17] ),
    .B_N(_05920_),
    .Y(_05960_));
 sg13g2_buf_1 _14204_ (.A(\soc_I.cpu_mem_wdata[1] ),
    .X(_05961_));
 sg13g2_mux2_1 _14205_ (.A0(net604),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[17] ),
    .S(net505),
    .X(_05962_));
 sg13g2_nor2_1 _14206_ (.A(net42),
    .B(_05962_),
    .Y(_05963_));
 sg13g2_nor3_1 _14207_ (.A(_05939_),
    .B(_05960_),
    .C(_05963_),
    .Y(_00139_));
 sg13g2_buf_1 _14208_ (.A(_05915_),
    .X(_05964_));
 sg13g2_nor2b_1 _14209_ (.A(\soc_I.div_reg[18] ),
    .B_N(_05964_),
    .Y(_05965_));
 sg13g2_mux2_1 _14210_ (.A0(net619),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[18] ),
    .S(net505),
    .X(_05966_));
 sg13g2_nor2_1 _14211_ (.A(net42),
    .B(_05966_),
    .Y(_05967_));
 sg13g2_nor3_1 _14212_ (.A(net396),
    .B(_05965_),
    .C(_05967_),
    .Y(_00140_));
 sg13g2_nor2b_1 _14213_ (.A(\soc_I.div_reg[19] ),
    .B_N(net48),
    .Y(_05968_));
 sg13g2_mux2_1 _14214_ (.A0(_05929_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[19] ),
    .S(net505),
    .X(_05969_));
 sg13g2_buf_1 _14215_ (.A(_05969_),
    .X(_05970_));
 sg13g2_nor2_1 _14216_ (.A(net42),
    .B(_05970_),
    .Y(_05971_));
 sg13g2_nor3_1 _14217_ (.A(net396),
    .B(_05968_),
    .C(_05971_),
    .Y(_00141_));
 sg13g2_mux2_1 _14218_ (.A0(net604),
    .A1(_05500_),
    .S(net50),
    .X(_05972_));
 sg13g2_and2_1 _14219_ (.A(net435),
    .B(_05972_),
    .X(_00142_));
 sg13g2_nor2b_1 _14220_ (.A(\soc_I.div_reg[20] ),
    .B_N(net48),
    .Y(_05973_));
 sg13g2_mux2_1 _14221_ (.A0(net606),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[20] ),
    .S(net434),
    .X(_05974_));
 sg13g2_nor2_1 _14222_ (.A(net42),
    .B(_05974_),
    .Y(_05975_));
 sg13g2_nor3_1 _14223_ (.A(net396),
    .B(_05973_),
    .C(_05975_),
    .Y(_00143_));
 sg13g2_nor2b_1 _14224_ (.A(\soc_I.div_reg[21] ),
    .B_N(net48),
    .Y(_05976_));
 sg13g2_mux2_1 _14225_ (.A0(_05941_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[21] ),
    .S(net505),
    .X(_05977_));
 sg13g2_buf_1 _14226_ (.A(_05977_),
    .X(_05978_));
 sg13g2_nor2_1 _14227_ (.A(net42),
    .B(_05978_),
    .Y(_05979_));
 sg13g2_nor3_1 _14228_ (.A(net396),
    .B(_05976_),
    .C(_05979_),
    .Y(_00144_));
 sg13g2_nor2b_1 _14229_ (.A(\soc_I.div_reg[22] ),
    .B_N(net48),
    .Y(_05980_));
 sg13g2_buf_8 _14230_ (.A(net50),
    .X(_05981_));
 sg13g2_inv_2 _14231_ (.Y(_05982_),
    .A(_05946_));
 sg13g2_nand2_1 _14232_ (.Y(_05983_),
    .A(_05956_),
    .B(\soc_I.kianv_I.datapath_unit_I.A2[22] ));
 sg13g2_o21ai_1 _14233_ (.B1(_05983_),
    .Y(_05984_),
    .A1(_05956_),
    .A2(_05982_));
 sg13g2_nor2_1 _14234_ (.A(_05981_),
    .B(_05984_),
    .Y(_05985_));
 sg13g2_nor3_1 _14235_ (.A(net396),
    .B(_05980_),
    .C(_05985_),
    .Y(_00145_));
 sg13g2_buf_1 _14236_ (.A(_05918_),
    .X(_05986_));
 sg13g2_nor2b_1 _14237_ (.A(\soc_I.div_reg[23] ),
    .B_N(net48),
    .Y(_05987_));
 sg13g2_mux2_1 _14238_ (.A0(net605),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[23] ),
    .S(net434),
    .X(_05988_));
 sg13g2_nor2_1 _14239_ (.A(net41),
    .B(_05988_),
    .Y(_05989_));
 sg13g2_nor3_1 _14240_ (.A(net395),
    .B(_05987_),
    .C(_05989_),
    .Y(_00146_));
 sg13g2_buf_1 _14241_ (.A(net630),
    .X(_05990_));
 sg13g2_nand2_1 _14242_ (.Y(_05991_),
    .A(net577),
    .B(_01936_));
 sg13g2_o21ai_1 _14243_ (.B1(_05991_),
    .Y(_05992_),
    .A1(net577),
    .A2(_01691_));
 sg13g2_mux2_1 _14244_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[24] ),
    .A1(_05992_),
    .S(net529),
    .X(_05993_));
 sg13g2_nand2b_1 _14245_ (.Y(_05994_),
    .B(_05993_),
    .A_N(net41));
 sg13g2_nand2_1 _14246_ (.Y(_05995_),
    .A(\soc_I.div_reg[24] ),
    .B(net43));
 sg13g2_a21oi_1 _14247_ (.A1(_05994_),
    .A2(_05995_),
    .Y(_00147_),
    .B1(net404));
 sg13g2_buf_1 _14248_ (.A(net577),
    .X(_05996_));
 sg13g2_nand2_1 _14249_ (.Y(_05997_),
    .A(net504),
    .B(_01952_));
 sg13g2_o21ai_1 _14250_ (.B1(_05997_),
    .Y(_05998_),
    .A1(net504),
    .A2(_00033_));
 sg13g2_mux2_1 _14251_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[25] ),
    .A1(_05998_),
    .S(net529),
    .X(_05999_));
 sg13g2_nand2b_1 _14252_ (.Y(_06000_),
    .B(_05999_),
    .A_N(net41));
 sg13g2_nand2_1 _14253_ (.Y(_06001_),
    .A(\soc_I.div_reg[25] ),
    .B(net43));
 sg13g2_buf_2 _14254_ (.A(net520),
    .X(_06002_));
 sg13g2_buf_1 _14255_ (.A(_06002_),
    .X(_06003_));
 sg13g2_a21oi_1 _14256_ (.A1(_06000_),
    .A2(_06001_),
    .Y(_00148_),
    .B1(net394));
 sg13g2_nor2b_1 _14257_ (.A(\soc_I.div_reg[26] ),
    .B_N(net48),
    .Y(_06004_));
 sg13g2_nor2_1 _14258_ (.A(_01840_),
    .B(\soc_I.kianv_I.datapath_unit_I.A2[10] ),
    .Y(_06005_));
 sg13g2_nor2b_1 _14259_ (.A(net577),
    .B_N(_00080_),
    .Y(_06006_));
 sg13g2_nor3_1 _14260_ (.A(net434),
    .B(_06005_),
    .C(_06006_),
    .Y(_06007_));
 sg13g2_a21o_1 _14261_ (.A2(\soc_I.kianv_I.datapath_unit_I.A2[26] ),
    .A1(net434),
    .B1(_06007_),
    .X(_06008_));
 sg13g2_buf_1 _14262_ (.A(_06008_),
    .X(_06009_));
 sg13g2_nor2_1 _14263_ (.A(_05981_),
    .B(_06009_),
    .Y(_06010_));
 sg13g2_nor3_1 _14264_ (.A(net395),
    .B(_06004_),
    .C(_06010_),
    .Y(_00149_));
 sg13g2_nand2_1 _14265_ (.Y(_06011_),
    .A(net577),
    .B(\soc_I.kianv_I.datapath_unit_I.A2[11] ));
 sg13g2_o21ai_1 _14266_ (.B1(_06011_),
    .Y(_06012_),
    .A1(_05990_),
    .A2(_00036_));
 sg13g2_nor2_1 _14267_ (.A(net434),
    .B(_06012_),
    .Y(_06013_));
 sg13g2_a21oi_1 _14268_ (.A1(net434),
    .A2(_02539_),
    .Y(_06014_),
    .B1(_06013_));
 sg13g2_nand2b_1 _14269_ (.Y(_06015_),
    .B(_06014_),
    .A_N(net41));
 sg13g2_nand2_1 _14270_ (.Y(_06016_),
    .A(\soc_I.div_reg[27] ),
    .B(net43));
 sg13g2_a21oi_1 _14271_ (.A1(_06015_),
    .A2(_06016_),
    .Y(_00150_),
    .B1(net394));
 sg13g2_nand2_1 _14272_ (.Y(_06017_),
    .A(net504),
    .B(_01856_));
 sg13g2_o21ai_1 _14273_ (.B1(_06017_),
    .Y(_06018_),
    .A1(net504),
    .A2(_00038_));
 sg13g2_mux2_1 _14274_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[28] ),
    .A1(_06018_),
    .S(net529),
    .X(_06019_));
 sg13g2_nand2b_1 _14275_ (.Y(_06020_),
    .B(_06019_),
    .A_N(net41));
 sg13g2_nand2_1 _14276_ (.Y(_06021_),
    .A(\soc_I.div_reg[28] ),
    .B(net43));
 sg13g2_a21oi_1 _14277_ (.A1(_06020_),
    .A2(_06021_),
    .Y(_00151_),
    .B1(net394));
 sg13g2_nand2_1 _14278_ (.Y(_06022_),
    .A(net577),
    .B(\soc_I.kianv_I.datapath_unit_I.A2[13] ));
 sg13g2_o21ai_1 _14279_ (.B1(_06022_),
    .Y(_06023_),
    .A1(net504),
    .A2(_00040_));
 sg13g2_mux2_1 _14280_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[29] ),
    .A1(_06023_),
    .S(net529),
    .X(_06024_));
 sg13g2_nand2b_1 _14281_ (.Y(_06025_),
    .B(_06024_),
    .A_N(net41));
 sg13g2_nand2_1 _14282_ (.Y(_06026_),
    .A(\soc_I.div_reg[29] ),
    .B(net43));
 sg13g2_a21oi_1 _14283_ (.A1(_06025_),
    .A2(_06026_),
    .Y(_00152_),
    .B1(net394));
 sg13g2_mux2_1 _14284_ (.A0(net619),
    .A1(_05497_),
    .S(net50),
    .X(_06027_));
 sg13g2_and2_1 _14285_ (.A(net435),
    .B(_06027_),
    .X(_00153_));
 sg13g2_nand2_1 _14286_ (.Y(_06028_),
    .A(net504),
    .B(\soc_I.kianv_I.datapath_unit_I.A2[14] ));
 sg13g2_o21ai_1 _14287_ (.B1(_06028_),
    .Y(_06029_),
    .A1(net504),
    .A2(_00042_));
 sg13g2_mux2_1 _14288_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[30] ),
    .A1(_06029_),
    .S(net529),
    .X(_06030_));
 sg13g2_nand2b_1 _14289_ (.Y(_06031_),
    .B(_06030_),
    .A_N(net49));
 sg13g2_nand2_1 _14290_ (.Y(_06032_),
    .A(\soc_I.div_reg[30] ),
    .B(net43));
 sg13g2_a21oi_1 _14291_ (.A1(_06031_),
    .A2(_06032_),
    .Y(_00154_),
    .B1(net394));
 sg13g2_nand2_1 _14292_ (.Y(_06033_),
    .A(net577),
    .B(\soc_I.kianv_I.datapath_unit_I.A2[15] ));
 sg13g2_o21ai_1 _14293_ (.B1(_06033_),
    .Y(_06034_),
    .A1(net577),
    .A2(_00044_));
 sg13g2_mux2_1 _14294_ (.A0(\soc_I.kianv_I.datapath_unit_I.A2[31] ),
    .A1(_06034_),
    .S(net529),
    .X(_06035_));
 sg13g2_nand2b_1 _14295_ (.Y(_06036_),
    .B(_06035_),
    .A_N(net49));
 sg13g2_nand2_1 _14296_ (.Y(_06037_),
    .A(\soc_I.div_reg[31] ),
    .B(net43));
 sg13g2_a21oi_1 _14297_ (.A1(_06036_),
    .A2(_06037_),
    .Y(_00155_),
    .B1(_06003_));
 sg13g2_mux2_1 _14298_ (.A0(_05929_),
    .A1(_05498_),
    .S(net50),
    .X(_06038_));
 sg13g2_and2_1 _14299_ (.A(net435),
    .B(_06038_),
    .X(_00156_));
 sg13g2_mux2_1 _14300_ (.A0(net606),
    .A1(_05491_),
    .S(net50),
    .X(_06039_));
 sg13g2_and2_1 _14301_ (.A(net435),
    .B(_06039_),
    .X(_00157_));
 sg13g2_mux2_1 _14302_ (.A0(_05941_),
    .A1(_05492_),
    .S(_05916_),
    .X(_06040_));
 sg13g2_and2_1 _14303_ (.A(_05909_),
    .B(_06040_),
    .X(_00158_));
 sg13g2_or2_1 _14304_ (.X(_06041_),
    .B(net48),
    .A(_05982_));
 sg13g2_nand2_1 _14305_ (.Y(_06042_),
    .A(_05485_),
    .B(_05922_));
 sg13g2_a21oi_1 _14306_ (.A1(_06041_),
    .A2(_06042_),
    .Y(_00159_),
    .B1(_06003_));
 sg13g2_mux2_1 _14307_ (.A0(net605),
    .A1(_05486_),
    .S(_05916_),
    .X(_06043_));
 sg13g2_and2_1 _14308_ (.A(_05909_),
    .B(_06043_),
    .X(_00160_));
 sg13g2_nor2b_1 _14309_ (.A(net609),
    .B_N(_05964_),
    .Y(_06044_));
 sg13g2_mux2_1 _14310_ (.A0(_01936_),
    .A1(net607),
    .S(_05936_),
    .X(_06045_));
 sg13g2_buf_1 _14311_ (.A(_06045_),
    .X(_06046_));
 sg13g2_nor2_1 _14312_ (.A(net41),
    .B(_06046_),
    .Y(_06047_));
 sg13g2_nor3_1 _14313_ (.A(_05986_),
    .B(_06044_),
    .C(_06047_),
    .Y(_00161_));
 sg13g2_nor2b_1 _14314_ (.A(_05480_),
    .B_N(net48),
    .Y(_06048_));
 sg13g2_mux2_1 _14315_ (.A0(_01952_),
    .A1(net604),
    .S(_05936_),
    .X(_06049_));
 sg13g2_nor2_1 _14316_ (.A(net41),
    .B(_06049_),
    .Y(_06050_));
 sg13g2_nor3_1 _14317_ (.A(_05986_),
    .B(_06048_),
    .C(_06050_),
    .Y(_00162_));
 sg13g2_buf_2 _14318_ (.A(\soc_I.kianv_I.Instr[15] ),
    .X(_06051_));
 sg13g2_buf_2 _14319_ (.A(_06051_),
    .X(_06052_));
 sg13g2_buf_2 _14320_ (.A(_06052_),
    .X(_06053_));
 sg13g2_nor4_1 _14321_ (.A(_02147_),
    .B(net620),
    .C(net621),
    .D(\soc_I.kianv_I.Instr[19] ),
    .Y(_06054_));
 sg13g2_nor2b_1 _14322_ (.A(net503),
    .B_N(_06054_),
    .Y(_06055_));
 sg13g2_buf_1 _14323_ (.A(_06055_),
    .X(_06056_));
 sg13g2_buf_1 _14324_ (.A(_06056_),
    .X(_06057_));
 sg13g2_buf_2 _14325_ (.A(_06052_),
    .X(_06058_));
 sg13g2_buf_1 _14326_ (.A(_02147_),
    .X(_06059_));
 sg13g2_buf_1 _14327_ (.A(_06059_),
    .X(_06060_));
 sg13g2_mux4_1 _14328_ (.S0(net502),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ),
    .S1(net501),
    .X(_06061_));
 sg13g2_buf_1 _14329_ (.A(_02147_),
    .X(_06062_));
 sg13g2_buf_1 _14330_ (.A(net576),
    .X(_06063_));
 sg13g2_mux4_1 _14331_ (.S0(net503),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ),
    .S1(net500),
    .X(_06064_));
 sg13g2_buf_2 _14332_ (.A(_06051_),
    .X(_06065_));
 sg13g2_buf_1 _14333_ (.A(_02147_),
    .X(_06066_));
 sg13g2_mux4_1 _14334_ (.S0(net575),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ),
    .S1(net574),
    .X(_06067_));
 sg13g2_buf_2 _14335_ (.A(_06052_),
    .X(_06068_));
 sg13g2_buf_1 _14336_ (.A(_06059_),
    .X(_06069_));
 sg13g2_mux4_1 _14337_ (.S0(net499),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ),
    .S1(net498),
    .X(_06070_));
 sg13g2_buf_2 _14338_ (.A(net620),
    .X(_06071_));
 sg13g2_buf_1 _14339_ (.A(net621),
    .X(_06072_));
 sg13g2_mux4_1 _14340_ (.S0(net573),
    .A0(_06061_),
    .A1(_06064_),
    .A2(_06067_),
    .A3(_06070_),
    .S1(net572),
    .X(_06073_));
 sg13g2_nor2b_1 _14341_ (.A(net357),
    .B_N(_06073_),
    .Y(_00163_));
 sg13g2_mux4_1 _14342_ (.S0(net502),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ),
    .S1(net501),
    .X(_06074_));
 sg13g2_mux4_1 _14343_ (.S0(net503),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ),
    .S1(net500),
    .X(_06075_));
 sg13g2_mux4_1 _14344_ (.S0(net575),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ),
    .S1(net574),
    .X(_06076_));
 sg13g2_mux4_1 _14345_ (.S0(net499),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ),
    .S1(net498),
    .X(_06077_));
 sg13g2_mux4_1 _14346_ (.S0(net573),
    .A0(_06074_),
    .A1(_06075_),
    .A2(_06076_),
    .A3(_06077_),
    .S1(net572),
    .X(_06078_));
 sg13g2_nor2b_1 _14347_ (.A(net357),
    .B_N(_06078_),
    .Y(_00164_));
 sg13g2_mux4_1 _14348_ (.S0(net502),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ),
    .S1(net501),
    .X(_06079_));
 sg13g2_mux4_1 _14349_ (.S0(net503),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ),
    .S1(net500),
    .X(_06080_));
 sg13g2_buf_2 _14350_ (.A(_06051_),
    .X(_06081_));
 sg13g2_mux4_1 _14351_ (.S0(net571),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ),
    .S1(net574),
    .X(_06082_));
 sg13g2_mux4_1 _14352_ (.S0(net499),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ),
    .S1(net498),
    .X(_06083_));
 sg13g2_mux4_1 _14353_ (.S0(net573),
    .A0(_06079_),
    .A1(_06080_),
    .A2(_06082_),
    .A3(_06083_),
    .S1(net572),
    .X(_06084_));
 sg13g2_nor2b_1 _14354_ (.A(net357),
    .B_N(_06084_),
    .Y(_00165_));
 sg13g2_mux4_1 _14355_ (.S0(net502),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ),
    .S1(net501),
    .X(_06085_));
 sg13g2_mux4_1 _14356_ (.S0(net503),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ),
    .S1(net500),
    .X(_06086_));
 sg13g2_buf_1 _14357_ (.A(_02147_),
    .X(_06087_));
 sg13g2_mux4_1 _14358_ (.S0(net571),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ),
    .S1(net570),
    .X(_06088_));
 sg13g2_mux4_1 _14359_ (.S0(net499),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ),
    .S1(net498),
    .X(_06089_));
 sg13g2_mux4_1 _14360_ (.S0(net573),
    .A0(_06085_),
    .A1(_06086_),
    .A2(_06088_),
    .A3(_06089_),
    .S1(net572),
    .X(_06090_));
 sg13g2_nor2b_1 _14361_ (.A(net357),
    .B_N(_06090_),
    .Y(_00166_));
 sg13g2_mux4_1 _14362_ (.S0(net502),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ),
    .S1(net501),
    .X(_06091_));
 sg13g2_mux4_1 _14363_ (.S0(net503),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ),
    .S1(net500),
    .X(_06092_));
 sg13g2_mux4_1 _14364_ (.S0(net571),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ),
    .S1(net570),
    .X(_06093_));
 sg13g2_buf_2 _14365_ (.A(_06051_),
    .X(_06094_));
 sg13g2_mux4_1 _14366_ (.S0(net569),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ),
    .S1(net498),
    .X(_06095_));
 sg13g2_mux4_1 _14367_ (.S0(net573),
    .A0(_06091_),
    .A1(_06092_),
    .A2(_06093_),
    .A3(_06095_),
    .S1(net572),
    .X(_06096_));
 sg13g2_nor2b_1 _14368_ (.A(net357),
    .B_N(_06096_),
    .Y(_00167_));
 sg13g2_mux4_1 _14369_ (.S0(net502),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ),
    .S1(net501),
    .X(_06097_));
 sg13g2_mux4_1 _14370_ (.S0(net503),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ),
    .S1(_06063_),
    .X(_06098_));
 sg13g2_mux4_1 _14371_ (.S0(net571),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ),
    .S1(net570),
    .X(_06099_));
 sg13g2_buf_1 _14372_ (.A(_06059_),
    .X(_06100_));
 sg13g2_mux4_1 _14373_ (.S0(net569),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ),
    .S1(net497),
    .X(_06101_));
 sg13g2_mux4_1 _14374_ (.S0(net573),
    .A0(_06097_),
    .A1(_06098_),
    .A2(_06099_),
    .A3(_06101_),
    .S1(_06072_),
    .X(_06102_));
 sg13g2_nor2b_1 _14375_ (.A(_06057_),
    .B_N(_06102_),
    .Y(_00168_));
 sg13g2_buf_2 _14376_ (.A(_06052_),
    .X(_06103_));
 sg13g2_mux4_1 _14377_ (.S0(net496),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ),
    .S1(net501),
    .X(_06104_));
 sg13g2_mux4_1 _14378_ (.S0(net503),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ),
    .S1(_06063_),
    .X(_06105_));
 sg13g2_mux4_1 _14379_ (.S0(net571),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ),
    .S1(net570),
    .X(_06106_));
 sg13g2_mux4_1 _14380_ (.S0(net569),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ),
    .S1(net497),
    .X(_06107_));
 sg13g2_mux4_1 _14381_ (.S0(_06071_),
    .A0(_06104_),
    .A1(_06105_),
    .A2(_06106_),
    .A3(_06107_),
    .S1(_06072_),
    .X(_06108_));
 sg13g2_nor2b_1 _14382_ (.A(_06057_),
    .B_N(_06108_),
    .Y(_00169_));
 sg13g2_buf_1 _14383_ (.A(_06059_),
    .X(_06109_));
 sg13g2_mux4_1 _14384_ (.S0(net496),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ),
    .S1(net495),
    .X(_06110_));
 sg13g2_mux4_1 _14385_ (.S0(_06053_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ),
    .S1(net500),
    .X(_06111_));
 sg13g2_mux4_1 _14386_ (.S0(_06081_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ),
    .S1(_06087_),
    .X(_06112_));
 sg13g2_mux4_1 _14387_ (.S0(net569),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ),
    .S1(net497),
    .X(_06113_));
 sg13g2_mux4_1 _14388_ (.S0(net573),
    .A0(_06110_),
    .A1(_06111_),
    .A2(_06112_),
    .A3(_06113_),
    .S1(net572),
    .X(_06114_));
 sg13g2_nor2b_1 _14389_ (.A(net357),
    .B_N(_06114_),
    .Y(_00170_));
 sg13g2_mux4_1 _14390_ (.S0(_06103_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ),
    .S1(_06109_),
    .X(_06115_));
 sg13g2_buf_2 _14391_ (.A(_06052_),
    .X(_06116_));
 sg13g2_mux4_1 _14392_ (.S0(_06116_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ),
    .S1(net500),
    .X(_06117_));
 sg13g2_mux4_1 _14393_ (.S0(_06081_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ),
    .S1(_06087_),
    .X(_06118_));
 sg13g2_mux4_1 _14394_ (.S0(_06094_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ),
    .S1(_06100_),
    .X(_06119_));
 sg13g2_mux4_1 _14395_ (.S0(net573),
    .A0(_06115_),
    .A1(_06117_),
    .A2(_06118_),
    .A3(_06119_),
    .S1(net572),
    .X(_06120_));
 sg13g2_nor2b_1 _14396_ (.A(net357),
    .B_N(_06120_),
    .Y(_00171_));
 sg13g2_mux4_1 _14397_ (.S0(net496),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ),
    .S1(net495),
    .X(_06121_));
 sg13g2_buf_1 _14398_ (.A(_06059_),
    .X(_06122_));
 sg13g2_mux4_1 _14399_ (.S0(net494),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ),
    .S1(net493),
    .X(_06123_));
 sg13g2_mux4_1 _14400_ (.S0(net571),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ),
    .S1(net570),
    .X(_06124_));
 sg13g2_mux4_1 _14401_ (.S0(net569),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ),
    .S1(net497),
    .X(_06125_));
 sg13g2_buf_2 _14402_ (.A(net620),
    .X(_06126_));
 sg13g2_buf_1 _14403_ (.A(net621),
    .X(_06127_));
 sg13g2_mux4_1 _14404_ (.S0(net568),
    .A0(_06121_),
    .A1(_06123_),
    .A2(_06124_),
    .A3(_06125_),
    .S1(net567),
    .X(_06128_));
 sg13g2_nor2b_1 _14405_ (.A(net357),
    .B_N(_06128_),
    .Y(_00172_));
 sg13g2_buf_1 _14406_ (.A(_06056_),
    .X(_06129_));
 sg13g2_mux4_1 _14407_ (.S0(net496),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ),
    .S1(net495),
    .X(_06130_));
 sg13g2_mux4_1 _14408_ (.S0(net494),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ),
    .S1(net493),
    .X(_06131_));
 sg13g2_mux4_1 _14409_ (.S0(net571),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ),
    .S1(net570),
    .X(_06132_));
 sg13g2_mux4_1 _14410_ (.S0(net569),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ),
    .S1(net497),
    .X(_06133_));
 sg13g2_mux4_1 _14411_ (.S0(net568),
    .A0(_06130_),
    .A1(_06131_),
    .A2(_06132_),
    .A3(_06133_),
    .S1(net567),
    .X(_06134_));
 sg13g2_nor2b_1 _14412_ (.A(_06129_),
    .B_N(_06134_),
    .Y(_00173_));
 sg13g2_mux4_1 _14413_ (.S0(net496),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ),
    .S1(net495),
    .X(_06135_));
 sg13g2_mux4_1 _14414_ (.S0(net494),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ),
    .S1(_06122_),
    .X(_06136_));
 sg13g2_mux4_1 _14415_ (.S0(net571),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ),
    .S1(net570),
    .X(_06137_));
 sg13g2_mux4_1 _14416_ (.S0(net569),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ),
    .S1(net497),
    .X(_06138_));
 sg13g2_mux4_1 _14417_ (.S0(_06126_),
    .A0(_06135_),
    .A1(_06136_),
    .A2(_06137_),
    .A3(_06138_),
    .S1(_06127_),
    .X(_06139_));
 sg13g2_nor2b_1 _14418_ (.A(_06129_),
    .B_N(_06139_),
    .Y(_00174_));
 sg13g2_mux4_1 _14419_ (.S0(_06103_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ),
    .S1(_06109_),
    .X(_06140_));
 sg13g2_mux4_1 _14420_ (.S0(_06116_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ),
    .S1(_06122_),
    .X(_06141_));
 sg13g2_buf_2 _14421_ (.A(_06051_),
    .X(_06142_));
 sg13g2_mux4_1 _14422_ (.S0(_06142_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ),
    .S1(net570),
    .X(_06143_));
 sg13g2_mux4_1 _14423_ (.S0(net569),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ),
    .S1(_06100_),
    .X(_06144_));
 sg13g2_mux4_1 _14424_ (.S0(_06126_),
    .A0(_06140_),
    .A1(_06141_),
    .A2(_06143_),
    .A3(_06144_),
    .S1(_06127_),
    .X(_06145_));
 sg13g2_nor2b_1 _14425_ (.A(net356),
    .B_N(_06145_),
    .Y(_00175_));
 sg13g2_mux4_1 _14426_ (.S0(net496),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ),
    .S1(net495),
    .X(_06146_));
 sg13g2_mux4_1 _14427_ (.S0(net494),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ),
    .S1(net493),
    .X(_06147_));
 sg13g2_buf_1 _14428_ (.A(_02147_),
    .X(_06148_));
 sg13g2_mux4_1 _14429_ (.S0(net566),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ),
    .S1(net565),
    .X(_06149_));
 sg13g2_mux4_1 _14430_ (.S0(_06094_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ),
    .S1(net497),
    .X(_06150_));
 sg13g2_mux4_1 _14431_ (.S0(net568),
    .A0(_06146_),
    .A1(_06147_),
    .A2(_06149_),
    .A3(_06150_),
    .S1(net567),
    .X(_06151_));
 sg13g2_nor2b_1 _14432_ (.A(net356),
    .B_N(_06151_),
    .Y(_00176_));
 sg13g2_mux4_1 _14433_ (.S0(net496),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ),
    .S1(net495),
    .X(_06152_));
 sg13g2_mux4_1 _14434_ (.S0(net494),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ),
    .S1(net493),
    .X(_06153_));
 sg13g2_mux4_1 _14435_ (.S0(net566),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ),
    .S1(net565),
    .X(_06154_));
 sg13g2_buf_2 _14436_ (.A(_06051_),
    .X(_06155_));
 sg13g2_mux4_1 _14437_ (.S0(net564),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ),
    .S1(net497),
    .X(_06156_));
 sg13g2_mux4_1 _14438_ (.S0(net568),
    .A0(_06152_),
    .A1(_06153_),
    .A2(_06154_),
    .A3(_06156_),
    .S1(net567),
    .X(_06157_));
 sg13g2_nor2b_1 _14439_ (.A(net356),
    .B_N(_06157_),
    .Y(_00177_));
 sg13g2_mux4_1 _14440_ (.S0(net496),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ),
    .S1(net495),
    .X(_06158_));
 sg13g2_mux4_1 _14441_ (.S0(net494),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ),
    .S1(net493),
    .X(_06159_));
 sg13g2_mux4_1 _14442_ (.S0(net566),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ),
    .S1(net565),
    .X(_06160_));
 sg13g2_buf_1 _14443_ (.A(_02147_),
    .X(_06161_));
 sg13g2_mux4_1 _14444_ (.S0(net564),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ),
    .S1(net563),
    .X(_06162_));
 sg13g2_mux4_1 _14445_ (.S0(net568),
    .A0(_06158_),
    .A1(_06159_),
    .A2(_06160_),
    .A3(_06162_),
    .S1(net567),
    .X(_06163_));
 sg13g2_nor2b_1 _14446_ (.A(net356),
    .B_N(_06163_),
    .Y(_00178_));
 sg13g2_buf_2 _14447_ (.A(_06052_),
    .X(_06164_));
 sg13g2_mux4_1 _14448_ (.S0(net492),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ),
    .S1(net495),
    .X(_06165_));
 sg13g2_mux4_1 _14449_ (.S0(net494),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ),
    .S1(net493),
    .X(_06166_));
 sg13g2_mux4_1 _14450_ (.S0(net566),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ),
    .S1(net565),
    .X(_06167_));
 sg13g2_mux4_1 _14451_ (.S0(net564),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ),
    .S1(net563),
    .X(_06168_));
 sg13g2_mux4_1 _14452_ (.S0(net568),
    .A0(_06165_),
    .A1(_06166_),
    .A2(_06167_),
    .A3(_06168_),
    .S1(net567),
    .X(_06169_));
 sg13g2_nor2b_1 _14453_ (.A(net356),
    .B_N(_06169_),
    .Y(_00179_));
 sg13g2_buf_1 _14454_ (.A(_06059_),
    .X(_06170_));
 sg13g2_mux4_1 _14455_ (.S0(net492),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ),
    .S1(net491),
    .X(_06171_));
 sg13g2_mux4_1 _14456_ (.S0(net494),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ),
    .S1(net493),
    .X(_06172_));
 sg13g2_mux4_1 _14457_ (.S0(_06142_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ),
    .S1(_06148_),
    .X(_06173_));
 sg13g2_mux4_1 _14458_ (.S0(_06155_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ),
    .S1(_06161_),
    .X(_06174_));
 sg13g2_mux4_1 _14459_ (.S0(net568),
    .A0(_06171_),
    .A1(_06172_),
    .A2(_06173_),
    .A3(_06174_),
    .S1(net567),
    .X(_06175_));
 sg13g2_nor2b_1 _14460_ (.A(net356),
    .B_N(_06175_),
    .Y(_00180_));
 sg13g2_mux4_1 _14461_ (.S0(net492),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ),
    .S1(net491),
    .X(_06176_));
 sg13g2_buf_2 _14462_ (.A(_06052_),
    .X(_06177_));
 sg13g2_mux4_1 _14463_ (.S0(net490),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ),
    .S1(net493),
    .X(_06178_));
 sg13g2_mux4_1 _14464_ (.S0(net566),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ),
    .S1(net565),
    .X(_06179_));
 sg13g2_mux4_1 _14465_ (.S0(net564),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ),
    .S1(net563),
    .X(_06180_));
 sg13g2_mux4_1 _14466_ (.S0(net568),
    .A0(_06176_),
    .A1(_06178_),
    .A2(_06179_),
    .A3(_06180_),
    .S1(net567),
    .X(_06181_));
 sg13g2_nor2b_1 _14467_ (.A(net356),
    .B_N(_06181_),
    .Y(_00181_));
 sg13g2_mux4_1 _14468_ (.S0(net492),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ),
    .S1(net491),
    .X(_06182_));
 sg13g2_buf_1 _14469_ (.A(_06059_),
    .X(_06183_));
 sg13g2_mux4_1 _14470_ (.S0(net490),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ),
    .S1(net489),
    .X(_06184_));
 sg13g2_mux4_1 _14471_ (.S0(net566),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ),
    .S1(net565),
    .X(_06185_));
 sg13g2_mux4_1 _14472_ (.S0(net564),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ),
    .S1(net563),
    .X(_06186_));
 sg13g2_buf_2 _14473_ (.A(net620),
    .X(_06187_));
 sg13g2_buf_1 _14474_ (.A(net621),
    .X(_06188_));
 sg13g2_mux4_1 _14475_ (.S0(net562),
    .A0(_06182_),
    .A1(_06184_),
    .A2(_06185_),
    .A3(_06186_),
    .S1(net561),
    .X(_06189_));
 sg13g2_nor2b_1 _14476_ (.A(net356),
    .B_N(_06189_),
    .Y(_00182_));
 sg13g2_buf_1 _14477_ (.A(_06056_),
    .X(_06190_));
 sg13g2_mux4_1 _14478_ (.S0(net492),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ),
    .S1(net491),
    .X(_06191_));
 sg13g2_mux4_1 _14479_ (.S0(net490),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ),
    .S1(net489),
    .X(_06192_));
 sg13g2_mux4_1 _14480_ (.S0(net566),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ),
    .S1(net565),
    .X(_06193_));
 sg13g2_mux4_1 _14481_ (.S0(net564),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ),
    .S1(net563),
    .X(_06194_));
 sg13g2_mux4_1 _14482_ (.S0(net562),
    .A0(_06191_),
    .A1(_06192_),
    .A2(_06193_),
    .A3(_06194_),
    .S1(net561),
    .X(_06195_));
 sg13g2_nor2b_1 _14483_ (.A(net355),
    .B_N(_06195_),
    .Y(_00183_));
 sg13g2_mux4_1 _14484_ (.S0(net492),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ),
    .S1(net491),
    .X(_06196_));
 sg13g2_mux4_1 _14485_ (.S0(net490),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ),
    .S1(net489),
    .X(_06197_));
 sg13g2_mux4_1 _14486_ (.S0(net566),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ),
    .S1(net565),
    .X(_06198_));
 sg13g2_mux4_1 _14487_ (.S0(net564),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ),
    .S1(net563),
    .X(_06199_));
 sg13g2_mux4_1 _14488_ (.S0(net562),
    .A0(_06196_),
    .A1(_06197_),
    .A2(_06198_),
    .A3(_06199_),
    .S1(net561),
    .X(_06200_));
 sg13g2_nor2b_1 _14489_ (.A(net355),
    .B_N(_06200_),
    .Y(_00184_));
 sg13g2_mux4_1 _14490_ (.S0(_06164_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ),
    .S1(net491),
    .X(_06201_));
 sg13g2_mux4_1 _14491_ (.S0(net490),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ),
    .S1(net489),
    .X(_06202_));
 sg13g2_buf_2 _14492_ (.A(_06051_),
    .X(_06203_));
 sg13g2_mux4_1 _14493_ (.S0(net560),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ),
    .S1(_06148_),
    .X(_06204_));
 sg13g2_mux4_1 _14494_ (.S0(net564),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ),
    .S1(net563),
    .X(_06205_));
 sg13g2_mux4_1 _14495_ (.S0(net562),
    .A0(_06201_),
    .A1(_06202_),
    .A2(_06204_),
    .A3(_06205_),
    .S1(net561),
    .X(_06206_));
 sg13g2_nor2b_1 _14496_ (.A(net355),
    .B_N(_06206_),
    .Y(_00185_));
 sg13g2_mux4_1 _14497_ (.S0(net492),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ),
    .S1(net491),
    .X(_06207_));
 sg13g2_mux4_1 _14498_ (.S0(net490),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ),
    .S1(net489),
    .X(_06208_));
 sg13g2_mux4_1 _14499_ (.S0(net560),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ),
    .S1(net576),
    .X(_06209_));
 sg13g2_mux4_1 _14500_ (.S0(_06155_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ),
    .S1(net563),
    .X(_06210_));
 sg13g2_mux4_1 _14501_ (.S0(net562),
    .A0(_06207_),
    .A1(_06208_),
    .A2(_06209_),
    .A3(_06210_),
    .S1(net561),
    .X(_06211_));
 sg13g2_nor2b_1 _14502_ (.A(net355),
    .B_N(_06211_),
    .Y(_00186_));
 sg13g2_mux4_1 _14503_ (.S0(_06164_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ),
    .S1(net491),
    .X(_06212_));
 sg13g2_mux4_1 _14504_ (.S0(net490),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ),
    .S1(net489),
    .X(_06213_));
 sg13g2_mux4_1 _14505_ (.S0(net560),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ),
    .S1(net576),
    .X(_06214_));
 sg13g2_mux4_1 _14506_ (.S0(net575),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ),
    .S1(_06161_),
    .X(_06215_));
 sg13g2_mux4_1 _14507_ (.S0(net562),
    .A0(_06212_),
    .A1(_06213_),
    .A2(_06214_),
    .A3(_06215_),
    .S1(net561),
    .X(_06216_));
 sg13g2_nor2b_1 _14508_ (.A(_06190_),
    .B_N(_06216_),
    .Y(_00187_));
 sg13g2_mux4_1 _14509_ (.S0(net492),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ),
    .S1(_06170_),
    .X(_06217_));
 sg13g2_mux4_1 _14510_ (.S0(net490),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ),
    .S1(net489),
    .X(_06218_));
 sg13g2_mux4_1 _14511_ (.S0(net560),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ),
    .S1(net576),
    .X(_06219_));
 sg13g2_mux4_1 _14512_ (.S0(net575),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ),
    .S1(net574),
    .X(_06220_));
 sg13g2_mux4_1 _14513_ (.S0(net562),
    .A0(_06217_),
    .A1(_06218_),
    .A2(_06219_),
    .A3(_06220_),
    .S1(net561),
    .X(_06221_));
 sg13g2_nor2b_1 _14514_ (.A(_06190_),
    .B_N(_06221_),
    .Y(_00188_));
 sg13g2_mux4_1 _14515_ (.S0(net499),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ),
    .S1(_06170_),
    .X(_06222_));
 sg13g2_mux4_1 _14516_ (.S0(_06177_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ),
    .S1(net489),
    .X(_06223_));
 sg13g2_mux4_1 _14517_ (.S0(net560),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ),
    .S1(net576),
    .X(_06224_));
 sg13g2_mux4_1 _14518_ (.S0(net575),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ),
    .S1(net574),
    .X(_06225_));
 sg13g2_mux4_1 _14519_ (.S0(net562),
    .A0(_06222_),
    .A1(_06223_),
    .A2(_06224_),
    .A3(_06225_),
    .S1(net561),
    .X(_06226_));
 sg13g2_nor2b_1 _14520_ (.A(net355),
    .B_N(_06226_),
    .Y(_00189_));
 sg13g2_mux4_1 _14521_ (.S0(net499),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ),
    .S1(net498),
    .X(_06227_));
 sg13g2_mux4_1 _14522_ (.S0(_06177_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ),
    .S1(_06183_),
    .X(_06228_));
 sg13g2_mux4_1 _14523_ (.S0(net560),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ),
    .S1(net576),
    .X(_06229_));
 sg13g2_mux4_1 _14524_ (.S0(net575),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ),
    .S1(net574),
    .X(_06230_));
 sg13g2_mux4_1 _14525_ (.S0(_06187_),
    .A0(_06227_),
    .A1(_06228_),
    .A2(_06229_),
    .A3(_06230_),
    .S1(_06188_),
    .X(_06231_));
 sg13g2_nor2b_1 _14526_ (.A(net355),
    .B_N(_06231_),
    .Y(_00190_));
 sg13g2_mux4_1 _14527_ (.S0(net499),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ),
    .S1(net498),
    .X(_06232_));
 sg13g2_mux4_1 _14528_ (.S0(net502),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ),
    .S1(_06183_),
    .X(_06233_));
 sg13g2_mux4_1 _14529_ (.S0(net560),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ),
    .S1(net576),
    .X(_06234_));
 sg13g2_mux4_1 _14530_ (.S0(net575),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ),
    .S1(net574),
    .X(_06235_));
 sg13g2_mux4_1 _14531_ (.S0(_06187_),
    .A0(_06232_),
    .A1(_06233_),
    .A2(_06234_),
    .A3(_06235_),
    .S1(_06188_),
    .X(_06236_));
 sg13g2_nor2b_1 _14532_ (.A(net355),
    .B_N(_06236_),
    .Y(_00191_));
 sg13g2_mux4_1 _14533_ (.S0(net499),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ),
    .S1(net498),
    .X(_06237_));
 sg13g2_mux4_1 _14534_ (.S0(net502),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ),
    .S1(net501),
    .X(_06238_));
 sg13g2_mux4_1 _14535_ (.S0(net560),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ),
    .S1(net576),
    .X(_06239_));
 sg13g2_mux4_1 _14536_ (.S0(net575),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ),
    .S1(net574),
    .X(_06240_));
 sg13g2_mux4_1 _14537_ (.S0(net620),
    .A0(_06237_),
    .A1(_06238_),
    .A2(_06239_),
    .A3(_06240_),
    .S1(net621),
    .X(_06241_));
 sg13g2_nor2b_1 _14538_ (.A(net355),
    .B_N(_06241_),
    .Y(_00192_));
 sg13g2_mux4_1 _14539_ (.S0(_06068_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ),
    .S1(_06069_),
    .X(_06242_));
 sg13g2_mux4_1 _14540_ (.S0(_06058_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ),
    .S1(_06060_),
    .X(_06243_));
 sg13g2_mux4_1 _14541_ (.S0(_06203_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ),
    .S1(_06062_),
    .X(_06244_));
 sg13g2_mux4_1 _14542_ (.S0(_06065_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8] ),
    .S1(_06066_),
    .X(_06245_));
 sg13g2_mux4_1 _14543_ (.S0(net620),
    .A0(_06242_),
    .A1(_06243_),
    .A2(_06244_),
    .A3(_06245_),
    .S1(net621),
    .X(_06246_));
 sg13g2_nor2b_1 _14544_ (.A(_06056_),
    .B_N(_06246_),
    .Y(_00193_));
 sg13g2_mux4_1 _14545_ (.S0(_06068_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ),
    .S1(_06069_),
    .X(_06247_));
 sg13g2_mux4_1 _14546_ (.S0(_06058_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ),
    .S1(_06060_),
    .X(_06248_));
 sg13g2_mux4_1 _14547_ (.S0(_06203_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ),
    .S1(_06062_),
    .X(_06249_));
 sg13g2_mux4_1 _14548_ (.S0(_06065_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ),
    .S1(_06066_),
    .X(_06250_));
 sg13g2_mux4_1 _14549_ (.S0(_02131_),
    .A0(_06247_),
    .A1(_06248_),
    .A2(_06249_),
    .A3(_06250_),
    .S1(_02114_),
    .X(_06251_));
 sg13g2_nor2b_1 _14550_ (.A(_06056_),
    .B_N(_06251_),
    .Y(_00194_));
 sg13g2_buf_2 _14551_ (.A(\soc_I.kianv_I.Instr[20] ),
    .X(_06252_));
 sg13g2_buf_2 _14552_ (.A(_06252_),
    .X(_06253_));
 sg13g2_nor4_1 _14553_ (.A(net559),
    .B(_02031_),
    .C(_02081_),
    .D(\soc_I.kianv_I.Instr[24] ),
    .Y(_06254_));
 sg13g2_nor2b_1 _14554_ (.A(net622),
    .B_N(_06254_),
    .Y(_06255_));
 sg13g2_buf_1 _14555_ (.A(_06255_),
    .X(_06256_));
 sg13g2_buf_1 _14556_ (.A(_06256_),
    .X(_06257_));
 sg13g2_buf_2 _14557_ (.A(_06252_),
    .X(_06258_));
 sg13g2_buf_2 _14558_ (.A(_06258_),
    .X(_06259_));
 sg13g2_buf_1 _14559_ (.A(_02031_),
    .X(_06260_));
 sg13g2_buf_1 _14560_ (.A(_06260_),
    .X(_06261_));
 sg13g2_mux4_1 _14561_ (.S0(net488),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ),
    .S1(net487),
    .X(_06262_));
 sg13g2_buf_2 _14562_ (.A(_06258_),
    .X(_06263_));
 sg13g2_buf_2 _14563_ (.A(_02031_),
    .X(_06264_));
 sg13g2_buf_1 _14564_ (.A(net558),
    .X(_06265_));
 sg13g2_mux4_1 _14565_ (.S0(net486),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ),
    .S1(net485),
    .X(_06266_));
 sg13g2_buf_2 _14566_ (.A(_06252_),
    .X(_06267_));
 sg13g2_buf_1 _14567_ (.A(_02031_),
    .X(_06268_));
 sg13g2_mux4_1 _14568_ (.S0(net557),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ),
    .S1(net556),
    .X(_06269_));
 sg13g2_buf_2 _14569_ (.A(_06258_),
    .X(_06270_));
 sg13g2_buf_1 _14570_ (.A(_06260_),
    .X(_06271_));
 sg13g2_mux4_1 _14571_ (.S0(net484),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ),
    .S1(net483),
    .X(_06272_));
 sg13g2_buf_2 _14572_ (.A(net622),
    .X(_06273_));
 sg13g2_buf_1 _14573_ (.A(_02081_),
    .X(_06274_));
 sg13g2_mux4_1 _14574_ (.S0(net555),
    .A0(_06262_),
    .A1(_06266_),
    .A2(_06269_),
    .A3(_06272_),
    .S1(net554),
    .X(_06275_));
 sg13g2_nor2b_1 _14575_ (.A(net354),
    .B_N(_06275_),
    .Y(_00195_));
 sg13g2_mux4_1 _14576_ (.S0(net488),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ),
    .S1(net487),
    .X(_06276_));
 sg13g2_mux4_1 _14577_ (.S0(net486),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ),
    .S1(net485),
    .X(_06277_));
 sg13g2_mux4_1 _14578_ (.S0(net557),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ),
    .S1(net556),
    .X(_06278_));
 sg13g2_mux4_1 _14579_ (.S0(net484),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ),
    .S1(net483),
    .X(_06279_));
 sg13g2_mux4_1 _14580_ (.S0(net555),
    .A0(_06276_),
    .A1(_06277_),
    .A2(_06278_),
    .A3(_06279_),
    .S1(net554),
    .X(_06280_));
 sg13g2_nor2b_1 _14581_ (.A(net354),
    .B_N(_06280_),
    .Y(_00196_));
 sg13g2_mux4_1 _14582_ (.S0(net488),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ),
    .S1(net487),
    .X(_06281_));
 sg13g2_mux4_1 _14583_ (.S0(net486),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ),
    .S1(net485),
    .X(_06282_));
 sg13g2_mux4_1 _14584_ (.S0(net557),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ),
    .S1(net556),
    .X(_06283_));
 sg13g2_mux4_1 _14585_ (.S0(net484),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ),
    .S1(net483),
    .X(_06284_));
 sg13g2_mux4_1 _14586_ (.S0(net555),
    .A0(_06281_),
    .A1(_06282_),
    .A2(_06283_),
    .A3(_06284_),
    .S1(net554),
    .X(_06285_));
 sg13g2_nor2b_1 _14587_ (.A(net354),
    .B_N(_06285_),
    .Y(_00197_));
 sg13g2_mux4_1 _14588_ (.S0(net488),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ),
    .S1(net487),
    .X(_06286_));
 sg13g2_mux4_1 _14589_ (.S0(net486),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ),
    .S1(net485),
    .X(_06287_));
 sg13g2_buf_2 _14590_ (.A(_06252_),
    .X(_06288_));
 sg13g2_buf_1 _14591_ (.A(_02031_),
    .X(_06289_));
 sg13g2_mux4_1 _14592_ (.S0(net553),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ),
    .S1(net552),
    .X(_06290_));
 sg13g2_mux4_1 _14593_ (.S0(net484),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ),
    .S1(net483),
    .X(_06291_));
 sg13g2_mux4_1 _14594_ (.S0(net555),
    .A0(_06286_),
    .A1(_06287_),
    .A2(_06290_),
    .A3(_06291_),
    .S1(net554),
    .X(_06292_));
 sg13g2_nor2b_1 _14595_ (.A(net354),
    .B_N(_06292_),
    .Y(_00198_));
 sg13g2_mux4_1 _14596_ (.S0(net488),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ),
    .S1(net487),
    .X(_06293_));
 sg13g2_mux4_1 _14597_ (.S0(net486),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ),
    .S1(net485),
    .X(_06294_));
 sg13g2_mux4_1 _14598_ (.S0(net553),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ),
    .S1(net552),
    .X(_06295_));
 sg13g2_mux4_1 _14599_ (.S0(net484),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ),
    .S1(net483),
    .X(_06296_));
 sg13g2_mux4_1 _14600_ (.S0(net555),
    .A0(_06293_),
    .A1(_06294_),
    .A2(_06295_),
    .A3(_06296_),
    .S1(net554),
    .X(_06297_));
 sg13g2_nor2b_1 _14601_ (.A(net354),
    .B_N(_06297_),
    .Y(_00199_));
 sg13g2_mux4_1 _14602_ (.S0(net488),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ),
    .S1(net487),
    .X(_06298_));
 sg13g2_mux4_1 _14603_ (.S0(_06263_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ),
    .S1(_06265_),
    .X(_06299_));
 sg13g2_mux4_1 _14604_ (.S0(net553),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ),
    .S1(net552),
    .X(_06300_));
 sg13g2_buf_2 _14605_ (.A(_06252_),
    .X(_06301_));
 sg13g2_buf_1 _14606_ (.A(_06260_),
    .X(_06302_));
 sg13g2_mux4_1 _14607_ (.S0(net551),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ),
    .S1(net482),
    .X(_06303_));
 sg13g2_mux4_1 _14608_ (.S0(_06273_),
    .A0(_06298_),
    .A1(_06299_),
    .A2(_06300_),
    .A3(_06303_),
    .S1(_06274_),
    .X(_06304_));
 sg13g2_nor2b_1 _14609_ (.A(_06257_),
    .B_N(_06304_),
    .Y(_00200_));
 sg13g2_mux4_1 _14610_ (.S0(net488),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ),
    .S1(net487),
    .X(_06305_));
 sg13g2_mux4_1 _14611_ (.S0(_06263_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ),
    .S1(_06265_),
    .X(_06306_));
 sg13g2_mux4_1 _14612_ (.S0(net553),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ),
    .S1(net552),
    .X(_06307_));
 sg13g2_mux4_1 _14613_ (.S0(net551),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ),
    .S1(net482),
    .X(_06308_));
 sg13g2_mux4_1 _14614_ (.S0(_06273_),
    .A0(_06305_),
    .A1(_06306_),
    .A2(_06307_),
    .A3(_06308_),
    .S1(_06274_),
    .X(_06309_));
 sg13g2_nor2b_1 _14615_ (.A(net354),
    .B_N(_06309_),
    .Y(_00201_));
 sg13g2_buf_2 _14616_ (.A(_06258_),
    .X(_06310_));
 sg13g2_buf_1 _14617_ (.A(_06260_),
    .X(_06311_));
 sg13g2_mux4_1 _14618_ (.S0(net481),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ),
    .S1(net480),
    .X(_06312_));
 sg13g2_mux4_1 _14619_ (.S0(net486),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ),
    .S1(net485),
    .X(_06313_));
 sg13g2_mux4_1 _14620_ (.S0(_06288_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ),
    .S1(_06289_),
    .X(_06314_));
 sg13g2_mux4_1 _14621_ (.S0(net551),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ),
    .S1(net482),
    .X(_06315_));
 sg13g2_mux4_1 _14622_ (.S0(net555),
    .A0(_06312_),
    .A1(_06313_),
    .A2(_06314_),
    .A3(_06315_),
    .S1(net554),
    .X(_06316_));
 sg13g2_nor2b_1 _14623_ (.A(_06257_),
    .B_N(_06316_),
    .Y(_00202_));
 sg13g2_mux4_1 _14624_ (.S0(_06310_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ),
    .S1(_06311_),
    .X(_06317_));
 sg13g2_mux4_1 _14625_ (.S0(net486),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ),
    .S1(net485),
    .X(_06318_));
 sg13g2_mux4_1 _14626_ (.S0(_06288_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ),
    .S1(_06289_),
    .X(_06319_));
 sg13g2_mux4_1 _14627_ (.S0(_06301_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ),
    .S1(_06302_),
    .X(_06320_));
 sg13g2_mux4_1 _14628_ (.S0(net555),
    .A0(_06317_),
    .A1(_06318_),
    .A2(_06319_),
    .A3(_06320_),
    .S1(net554),
    .X(_06321_));
 sg13g2_nor2b_1 _14629_ (.A(net354),
    .B_N(_06321_),
    .Y(_00203_));
 sg13g2_mux4_1 _14630_ (.S0(net481),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ),
    .S1(net480),
    .X(_06322_));
 sg13g2_buf_2 _14631_ (.A(_06258_),
    .X(_06323_));
 sg13g2_buf_1 _14632_ (.A(_06260_),
    .X(_06324_));
 sg13g2_mux4_1 _14633_ (.S0(net479),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ),
    .S1(net478),
    .X(_06325_));
 sg13g2_mux4_1 _14634_ (.S0(net553),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ),
    .S1(net552),
    .X(_06326_));
 sg13g2_mux4_1 _14635_ (.S0(net551),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ),
    .S1(net482),
    .X(_06327_));
 sg13g2_buf_2 _14636_ (.A(net622),
    .X(_06328_));
 sg13g2_buf_1 _14637_ (.A(_02081_),
    .X(_06329_));
 sg13g2_mux4_1 _14638_ (.S0(net550),
    .A0(_06322_),
    .A1(_06325_),
    .A2(_06326_),
    .A3(_06327_),
    .S1(net549),
    .X(_06330_));
 sg13g2_nor2b_1 _14639_ (.A(net354),
    .B_N(_06330_),
    .Y(_00204_));
 sg13g2_buf_1 _14640_ (.A(_06256_),
    .X(_06331_));
 sg13g2_mux4_1 _14641_ (.S0(net481),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ),
    .S1(net480),
    .X(_06332_));
 sg13g2_mux4_1 _14642_ (.S0(net479),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ),
    .S1(net478),
    .X(_06333_));
 sg13g2_mux4_1 _14643_ (.S0(net553),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ),
    .S1(net552),
    .X(_06334_));
 sg13g2_mux4_1 _14644_ (.S0(net551),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ),
    .S1(net482),
    .X(_06335_));
 sg13g2_mux4_1 _14645_ (.S0(net550),
    .A0(_06332_),
    .A1(_06333_),
    .A2(_06334_),
    .A3(_06335_),
    .S1(net549),
    .X(_06336_));
 sg13g2_nor2b_1 _14646_ (.A(net353),
    .B_N(_06336_),
    .Y(_00205_));
 sg13g2_mux4_1 _14647_ (.S0(net481),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ),
    .S1(net480),
    .X(_06337_));
 sg13g2_mux4_1 _14648_ (.S0(_06323_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ),
    .S1(_06324_),
    .X(_06338_));
 sg13g2_mux4_1 _14649_ (.S0(net553),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ),
    .S1(net552),
    .X(_06339_));
 sg13g2_mux4_1 _14650_ (.S0(net551),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ),
    .S1(net482),
    .X(_06340_));
 sg13g2_mux4_1 _14651_ (.S0(_06328_),
    .A0(_06337_),
    .A1(_06338_),
    .A2(_06339_),
    .A3(_06340_),
    .S1(_06329_),
    .X(_06341_));
 sg13g2_nor2b_1 _14652_ (.A(_06331_),
    .B_N(_06341_),
    .Y(_00206_));
 sg13g2_mux4_1 _14653_ (.S0(_06310_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ),
    .S1(_06311_),
    .X(_06342_));
 sg13g2_mux4_1 _14654_ (.S0(_06323_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ),
    .S1(_06324_),
    .X(_06343_));
 sg13g2_mux4_1 _14655_ (.S0(net553),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ),
    .S1(net552),
    .X(_06344_));
 sg13g2_mux4_1 _14656_ (.S0(_06301_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ),
    .S1(_06302_),
    .X(_06345_));
 sg13g2_mux4_1 _14657_ (.S0(_06328_),
    .A0(_06342_),
    .A1(_06343_),
    .A2(_06344_),
    .A3(_06345_),
    .S1(_06329_),
    .X(_06346_));
 sg13g2_nor2b_1 _14658_ (.A(_06331_),
    .B_N(_06346_),
    .Y(_00207_));
 sg13g2_mux4_1 _14659_ (.S0(net481),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ),
    .S1(net480),
    .X(_06347_));
 sg13g2_mux4_1 _14660_ (.S0(net479),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ),
    .S1(net478),
    .X(_06348_));
 sg13g2_buf_2 _14661_ (.A(_06252_),
    .X(_06349_));
 sg13g2_buf_1 _14662_ (.A(_02031_),
    .X(_06350_));
 sg13g2_mux4_1 _14663_ (.S0(net548),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ),
    .S1(net547),
    .X(_06351_));
 sg13g2_mux4_1 _14664_ (.S0(net551),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ),
    .S1(net482),
    .X(_06352_));
 sg13g2_mux4_1 _14665_ (.S0(net550),
    .A0(_06347_),
    .A1(_06348_),
    .A2(_06351_),
    .A3(_06352_),
    .S1(net549),
    .X(_06353_));
 sg13g2_nor2b_1 _14666_ (.A(net353),
    .B_N(_06353_),
    .Y(_00208_));
 sg13g2_mux4_1 _14667_ (.S0(net481),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ),
    .S1(net480),
    .X(_06354_));
 sg13g2_mux4_1 _14668_ (.S0(net479),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ),
    .S1(net478),
    .X(_06355_));
 sg13g2_mux4_1 _14669_ (.S0(net548),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ),
    .S1(net547),
    .X(_06356_));
 sg13g2_mux4_1 _14670_ (.S0(net551),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ),
    .S1(net482),
    .X(_06357_));
 sg13g2_mux4_1 _14671_ (.S0(net550),
    .A0(_06354_),
    .A1(_06355_),
    .A2(_06356_),
    .A3(_06357_),
    .S1(net549),
    .X(_06358_));
 sg13g2_nor2b_1 _14672_ (.A(net353),
    .B_N(_06358_),
    .Y(_00209_));
 sg13g2_mux4_1 _14673_ (.S0(net481),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ),
    .S1(net480),
    .X(_06359_));
 sg13g2_mux4_1 _14674_ (.S0(net479),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ),
    .S1(net478),
    .X(_06360_));
 sg13g2_mux4_1 _14675_ (.S0(net548),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ),
    .S1(net547),
    .X(_06361_));
 sg13g2_buf_2 _14676_ (.A(_06252_),
    .X(_06362_));
 sg13g2_buf_1 _14677_ (.A(_02031_),
    .X(_06363_));
 sg13g2_mux4_1 _14678_ (.S0(net546),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ),
    .S1(net545),
    .X(_06364_));
 sg13g2_mux4_1 _14679_ (.S0(net550),
    .A0(_06359_),
    .A1(_06360_),
    .A2(_06361_),
    .A3(_06364_),
    .S1(net549),
    .X(_06365_));
 sg13g2_nor2b_1 _14680_ (.A(net353),
    .B_N(_06365_),
    .Y(_00210_));
 sg13g2_mux4_1 _14681_ (.S0(net481),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ),
    .S1(net480),
    .X(_06366_));
 sg13g2_mux4_1 _14682_ (.S0(net479),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ),
    .S1(net478),
    .X(_06367_));
 sg13g2_mux4_1 _14683_ (.S0(net548),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ),
    .S1(net547),
    .X(_06368_));
 sg13g2_mux4_1 _14684_ (.S0(net546),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ),
    .S1(net545),
    .X(_06369_));
 sg13g2_mux4_1 _14685_ (.S0(net550),
    .A0(_06366_),
    .A1(_06367_),
    .A2(_06368_),
    .A3(_06369_),
    .S1(net549),
    .X(_06370_));
 sg13g2_nor2b_1 _14686_ (.A(net353),
    .B_N(_06370_),
    .Y(_00211_));
 sg13g2_buf_2 _14687_ (.A(_06258_),
    .X(_06371_));
 sg13g2_buf_1 _14688_ (.A(_06260_),
    .X(_06372_));
 sg13g2_mux4_1 _14689_ (.S0(net477),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ),
    .S1(net476),
    .X(_06373_));
 sg13g2_mux4_1 _14690_ (.S0(net479),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ),
    .S1(net478),
    .X(_06374_));
 sg13g2_mux4_1 _14691_ (.S0(_06349_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ),
    .S1(_06350_),
    .X(_06375_));
 sg13g2_mux4_1 _14692_ (.S0(net546),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ),
    .S1(net545),
    .X(_06376_));
 sg13g2_mux4_1 _14693_ (.S0(net550),
    .A0(_06373_),
    .A1(_06374_),
    .A2(_06375_),
    .A3(_06376_),
    .S1(net549),
    .X(_06377_));
 sg13g2_nor2b_1 _14694_ (.A(net353),
    .B_N(_06377_),
    .Y(_00212_));
 sg13g2_mux4_1 _14695_ (.S0(net477),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ),
    .S1(net476),
    .X(_06378_));
 sg13g2_mux4_1 _14696_ (.S0(net479),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ),
    .S1(net478),
    .X(_06379_));
 sg13g2_mux4_1 _14697_ (.S0(net548),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ),
    .S1(net547),
    .X(_06380_));
 sg13g2_mux4_1 _14698_ (.S0(net546),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ),
    .S1(net545),
    .X(_06381_));
 sg13g2_mux4_1 _14699_ (.S0(net550),
    .A0(_06378_),
    .A1(_06379_),
    .A2(_06380_),
    .A3(_06381_),
    .S1(net549),
    .X(_06382_));
 sg13g2_nor2b_1 _14700_ (.A(net353),
    .B_N(_06382_),
    .Y(_00213_));
 sg13g2_mux4_1 _14701_ (.S0(net477),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ),
    .S1(net476),
    .X(_06383_));
 sg13g2_buf_2 _14702_ (.A(_06258_),
    .X(_06384_));
 sg13g2_buf_1 _14703_ (.A(_06260_),
    .X(_06385_));
 sg13g2_mux4_1 _14704_ (.S0(net475),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ),
    .S1(net474),
    .X(_06386_));
 sg13g2_mux4_1 _14705_ (.S0(net548),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ),
    .S1(net547),
    .X(_06387_));
 sg13g2_mux4_1 _14706_ (.S0(net546),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ),
    .S1(net545),
    .X(_06388_));
 sg13g2_buf_2 _14707_ (.A(net622),
    .X(_06389_));
 sg13g2_buf_1 _14708_ (.A(_02081_),
    .X(_06390_));
 sg13g2_mux4_1 _14709_ (.S0(net544),
    .A0(_06383_),
    .A1(_06386_),
    .A2(_06387_),
    .A3(_06388_),
    .S1(net543),
    .X(_06391_));
 sg13g2_nor2b_1 _14710_ (.A(net353),
    .B_N(_06391_),
    .Y(_00214_));
 sg13g2_buf_1 _14711_ (.A(_06256_),
    .X(_06392_));
 sg13g2_mux4_1 _14712_ (.S0(net477),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ),
    .S1(net476),
    .X(_06393_));
 sg13g2_mux4_1 _14713_ (.S0(net475),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ),
    .S1(net474),
    .X(_06394_));
 sg13g2_mux4_1 _14714_ (.S0(net548),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ),
    .S1(net547),
    .X(_06395_));
 sg13g2_mux4_1 _14715_ (.S0(net546),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ),
    .S1(net545),
    .X(_06396_));
 sg13g2_mux4_1 _14716_ (.S0(net544),
    .A0(_06393_),
    .A1(_06394_),
    .A2(_06395_),
    .A3(_06396_),
    .S1(net543),
    .X(_06397_));
 sg13g2_nor2b_1 _14717_ (.A(net352),
    .B_N(_06397_),
    .Y(_00215_));
 sg13g2_mux4_1 _14718_ (.S0(net477),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ),
    .S1(net476),
    .X(_06398_));
 sg13g2_mux4_1 _14719_ (.S0(net475),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ),
    .S1(net474),
    .X(_06399_));
 sg13g2_mux4_1 _14720_ (.S0(net548),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ),
    .S1(net547),
    .X(_06400_));
 sg13g2_mux4_1 _14721_ (.S0(net546),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ),
    .S1(net545),
    .X(_06401_));
 sg13g2_mux4_1 _14722_ (.S0(net544),
    .A0(_06398_),
    .A1(_06399_),
    .A2(_06400_),
    .A3(_06401_),
    .S1(net543),
    .X(_06402_));
 sg13g2_nor2b_1 _14723_ (.A(net352),
    .B_N(_06402_),
    .Y(_00216_));
 sg13g2_mux4_1 _14724_ (.S0(net477),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ),
    .S1(net476),
    .X(_06403_));
 sg13g2_mux4_1 _14725_ (.S0(net475),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ),
    .S1(net474),
    .X(_06404_));
 sg13g2_mux4_1 _14726_ (.S0(_06349_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ),
    .S1(_06350_),
    .X(_06405_));
 sg13g2_mux4_1 _14727_ (.S0(net546),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ),
    .S1(net545),
    .X(_06406_));
 sg13g2_mux4_1 _14728_ (.S0(net544),
    .A0(_06403_),
    .A1(_06404_),
    .A2(_06405_),
    .A3(_06406_),
    .S1(net543),
    .X(_06407_));
 sg13g2_nor2b_1 _14729_ (.A(net352),
    .B_N(_06407_),
    .Y(_00217_));
 sg13g2_mux4_1 _14730_ (.S0(_06371_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ),
    .S1(_06372_),
    .X(_06408_));
 sg13g2_mux4_1 _14731_ (.S0(net475),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ),
    .S1(net474),
    .X(_06409_));
 sg13g2_mux4_1 _14732_ (.S0(net559),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ),
    .S1(net558),
    .X(_06410_));
 sg13g2_mux4_1 _14733_ (.S0(_06362_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ),
    .S1(_06363_),
    .X(_06411_));
 sg13g2_mux4_1 _14734_ (.S0(net544),
    .A0(_06408_),
    .A1(_06409_),
    .A2(_06410_),
    .A3(_06411_),
    .S1(net543),
    .X(_06412_));
 sg13g2_nor2b_1 _14735_ (.A(net352),
    .B_N(_06412_),
    .Y(_00218_));
 sg13g2_mux4_1 _14736_ (.S0(net477),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ),
    .S1(net476),
    .X(_06413_));
 sg13g2_mux4_1 _14737_ (.S0(net475),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ),
    .S1(net474),
    .X(_06414_));
 sg13g2_mux4_1 _14738_ (.S0(net559),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ),
    .S1(net558),
    .X(_06415_));
 sg13g2_mux4_1 _14739_ (.S0(_06362_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ),
    .S1(_06363_),
    .X(_06416_));
 sg13g2_mux4_1 _14740_ (.S0(net544),
    .A0(_06413_),
    .A1(_06414_),
    .A2(_06415_),
    .A3(_06416_),
    .S1(net543),
    .X(_06417_));
 sg13g2_nor2b_1 _14741_ (.A(net352),
    .B_N(_06417_),
    .Y(_00219_));
 sg13g2_mux4_1 _14742_ (.S0(_06371_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ),
    .S1(_06372_),
    .X(_06418_));
 sg13g2_mux4_1 _14743_ (.S0(net475),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ),
    .S1(net474),
    .X(_06419_));
 sg13g2_mux4_1 _14744_ (.S0(net559),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ),
    .S1(net558),
    .X(_06420_));
 sg13g2_mux4_1 _14745_ (.S0(net557),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ),
    .S1(net556),
    .X(_06421_));
 sg13g2_mux4_1 _14746_ (.S0(net544),
    .A0(_06418_),
    .A1(_06419_),
    .A2(_06420_),
    .A3(_06421_),
    .S1(net543),
    .X(_06422_));
 sg13g2_nor2b_1 _14747_ (.A(net352),
    .B_N(_06422_),
    .Y(_00220_));
 sg13g2_mux4_1 _14748_ (.S0(net477),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ),
    .S1(net476),
    .X(_06423_));
 sg13g2_mux4_1 _14749_ (.S0(net475),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ),
    .S1(net474),
    .X(_06424_));
 sg13g2_mux4_1 _14750_ (.S0(net559),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ),
    .S1(net558),
    .X(_06425_));
 sg13g2_mux4_1 _14751_ (.S0(net557),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ),
    .S1(net556),
    .X(_06426_));
 sg13g2_mux4_1 _14752_ (.S0(net544),
    .A0(_06423_),
    .A1(_06424_),
    .A2(_06425_),
    .A3(_06426_),
    .S1(net543),
    .X(_06427_));
 sg13g2_nor2b_1 _14753_ (.A(net352),
    .B_N(_06427_),
    .Y(_00221_));
 sg13g2_mux4_1 _14754_ (.S0(net484),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ),
    .S1(net483),
    .X(_06428_));
 sg13g2_mux4_1 _14755_ (.S0(_06384_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ),
    .S1(_06385_),
    .X(_06429_));
 sg13g2_mux4_1 _14756_ (.S0(net559),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ),
    .S1(net558),
    .X(_06430_));
 sg13g2_mux4_1 _14757_ (.S0(net557),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ),
    .S1(net556),
    .X(_06431_));
 sg13g2_mux4_1 _14758_ (.S0(_06389_),
    .A0(_06428_),
    .A1(_06429_),
    .A2(_06430_),
    .A3(_06431_),
    .S1(_06390_),
    .X(_06432_));
 sg13g2_nor2b_1 _14759_ (.A(net352),
    .B_N(_06432_),
    .Y(_00222_));
 sg13g2_mux4_1 _14760_ (.S0(net484),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ),
    .S1(net483),
    .X(_06433_));
 sg13g2_mux4_1 _14761_ (.S0(_06384_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ),
    .S1(_06385_),
    .X(_06434_));
 sg13g2_mux4_1 _14762_ (.S0(net559),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ),
    .S1(net558),
    .X(_06435_));
 sg13g2_mux4_1 _14763_ (.S0(net557),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ),
    .S1(net556),
    .X(_06436_));
 sg13g2_mux4_1 _14764_ (.S0(_06389_),
    .A0(_06433_),
    .A1(_06434_),
    .A2(_06435_),
    .A3(_06436_),
    .S1(_06390_),
    .X(_06437_));
 sg13g2_nor2b_1 _14765_ (.A(_06392_),
    .B_N(_06437_),
    .Y(_00223_));
 sg13g2_mux4_1 _14766_ (.S0(net484),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ),
    .S1(net483),
    .X(_06438_));
 sg13g2_mux4_1 _14767_ (.S0(net488),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ),
    .S1(net487),
    .X(_06439_));
 sg13g2_mux4_1 _14768_ (.S0(net559),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ),
    .S1(net558),
    .X(_06440_));
 sg13g2_mux4_1 _14769_ (.S0(net557),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ),
    .S1(net556),
    .X(_06441_));
 sg13g2_mux4_1 _14770_ (.S0(net622),
    .A0(_06438_),
    .A1(_06439_),
    .A2(_06440_),
    .A3(_06441_),
    .S1(_02081_),
    .X(_06442_));
 sg13g2_nor2b_1 _14771_ (.A(_06392_),
    .B_N(_06442_),
    .Y(_00224_));
 sg13g2_mux4_1 _14772_ (.S0(_06270_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ),
    .S1(_06271_),
    .X(_06443_));
 sg13g2_mux4_1 _14773_ (.S0(_06259_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ),
    .S1(_06261_),
    .X(_06444_));
 sg13g2_mux4_1 _14774_ (.S0(_06253_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ),
    .S1(_06264_),
    .X(_06445_));
 sg13g2_mux4_1 _14775_ (.S0(_06267_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8] ),
    .S1(_06268_),
    .X(_06446_));
 sg13g2_mux4_1 _14776_ (.S0(net622),
    .A0(_06443_),
    .A1(_06444_),
    .A2(_06445_),
    .A3(_06446_),
    .S1(_02081_),
    .X(_06447_));
 sg13g2_nor2b_1 _14777_ (.A(_06256_),
    .B_N(_06447_),
    .Y(_00225_));
 sg13g2_mux4_1 _14778_ (.S0(_06270_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ),
    .S1(_06271_),
    .X(_06448_));
 sg13g2_mux4_1 _14779_ (.S0(_06259_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ),
    .S1(_06261_),
    .X(_06449_));
 sg13g2_mux4_1 _14780_ (.S0(_06253_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ),
    .S1(_06264_),
    .X(_06450_));
 sg13g2_mux4_1 _14781_ (.S0(_06267_),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ),
    .S1(_06268_),
    .X(_06451_));
 sg13g2_mux4_1 _14782_ (.S0(_02058_),
    .A0(_06448_),
    .A1(_06449_),
    .A2(_06450_),
    .A3(_06451_),
    .S1(_02081_),
    .X(_06452_));
 sg13g2_nor2b_1 _14783_ (.A(_06256_),
    .B_N(_06452_),
    .Y(_00226_));
 sg13g2_buf_1 _14784_ (.A(net74),
    .X(_06453_));
 sg13g2_nor2_1 _14785_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[0] ),
    .B(net71),
    .Y(_06454_));
 sg13g2_buf_1 _14786_ (.A(net74),
    .X(_06455_));
 sg13g2_and2_1 _14787_ (.A(_04547_),
    .B(net70),
    .X(_06456_));
 sg13g2_nor3_1 _14788_ (.A(net395),
    .B(_06454_),
    .C(_06456_),
    .Y(_00227_));
 sg13g2_nor2_1 _14789_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[10] ),
    .B(net71),
    .Y(_06457_));
 sg13g2_buf_1 _14790_ (.A(_05898_),
    .X(_06458_));
 sg13g2_nor2_1 _14791_ (.A(_04029_),
    .B(_06458_),
    .Y(_06459_));
 sg13g2_nor3_1 _14792_ (.A(net395),
    .B(_06457_),
    .C(_06459_),
    .Y(_00228_));
 sg13g2_nand2_1 _14793_ (.Y(_06460_),
    .A(_04139_),
    .B(net70));
 sg13g2_o21ai_1 _14794_ (.B1(_06460_),
    .Y(_06461_),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[11] ),
    .A2(net71));
 sg13g2_nor2_1 _14795_ (.A(net400),
    .B(_06461_),
    .Y(_00229_));
 sg13g2_buf_1 _14796_ (.A(net74),
    .X(_06462_));
 sg13g2_nor2_1 _14797_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[12] ),
    .B(net69),
    .Y(_06463_));
 sg13g2_nor2_1 _14798_ (.A(_04125_),
    .B(net73),
    .Y(_06464_));
 sg13g2_nor3_1 _14799_ (.A(net395),
    .B(_06463_),
    .C(_06464_),
    .Y(_00230_));
 sg13g2_nor2_1 _14800_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[13] ),
    .B(net69),
    .Y(_06465_));
 sg13g2_nor2_1 _14801_ (.A(_03976_),
    .B(_06458_),
    .Y(_06466_));
 sg13g2_nor3_1 _14802_ (.A(net395),
    .B(_06465_),
    .C(_06466_),
    .Y(_00231_));
 sg13g2_buf_1 _14803_ (.A(_05898_),
    .X(_06467_));
 sg13g2_a21o_1 _14804_ (.A2(_03981_),
    .A1(_03988_),
    .B1(_06467_),
    .X(_06468_));
 sg13g2_nand2_1 _14805_ (.Y(_06469_),
    .A(\soc_I.kianv_I.datapath_unit_I.ALUOut[14] ),
    .B(net72));
 sg13g2_a21oi_1 _14806_ (.A1(_06468_),
    .A2(_06469_),
    .Y(_00232_),
    .B1(net394));
 sg13g2_o21ai_1 _14807_ (.B1(net71),
    .Y(_06470_),
    .A1(_03928_),
    .A2(_04145_));
 sg13g2_nand2_1 _14808_ (.Y(_06471_),
    .A(\soc_I.kianv_I.datapath_unit_I.ALUOut[15] ),
    .B(net72));
 sg13g2_a21oi_1 _14809_ (.A1(_06470_),
    .A2(_06471_),
    .Y(_00233_),
    .B1(net394));
 sg13g2_nor2_1 _14810_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[16] ),
    .B(net69),
    .Y(_06472_));
 sg13g2_and2_1 _14811_ (.A(_04586_),
    .B(_06455_),
    .X(_06473_));
 sg13g2_nor3_1 _14812_ (.A(net395),
    .B(_06472_),
    .C(_06473_),
    .Y(_00234_));
 sg13g2_nor2_1 _14813_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[17] ),
    .B(net69),
    .Y(_06474_));
 sg13g2_nand2_1 _14814_ (.Y(_06475_),
    .A(_03721_),
    .B(_04129_));
 sg13g2_nor2_1 _14815_ (.A(_06475_),
    .B(net73),
    .Y(_06476_));
 sg13g2_nor3_1 _14816_ (.A(net395),
    .B(_06474_),
    .C(_06476_),
    .Y(_00235_));
 sg13g2_buf_1 _14817_ (.A(_05918_),
    .X(_06477_));
 sg13g2_nor2_1 _14818_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[18] ),
    .B(_06462_),
    .Y(_06478_));
 sg13g2_and2_1 _14819_ (.A(_03681_),
    .B(net70),
    .X(_06479_));
 sg13g2_nor3_1 _14820_ (.A(_06477_),
    .B(_06478_),
    .C(_06479_),
    .Y(_00236_));
 sg13g2_nor2_1 _14821_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[19] ),
    .B(net69),
    .Y(_06480_));
 sg13g2_and2_1 _14822_ (.A(_04120_),
    .B(net70),
    .X(_06481_));
 sg13g2_nor3_1 _14823_ (.A(net393),
    .B(_06480_),
    .C(_06481_),
    .Y(_00237_));
 sg13g2_nor2_1 _14824_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[1] ),
    .B(net69),
    .Y(_06482_));
 sg13g2_and2_1 _14825_ (.A(_01791_),
    .B(_06455_),
    .X(_06483_));
 sg13g2_nor3_1 _14826_ (.A(_06477_),
    .B(_06482_),
    .C(_06483_),
    .Y(_00238_));
 sg13g2_nand2_1 _14827_ (.Y(_06484_),
    .A(_04136_),
    .B(net71));
 sg13g2_nand2_1 _14828_ (.Y(_06485_),
    .A(\soc_I.kianv_I.datapath_unit_I.ALUOut[20] ),
    .B(net72));
 sg13g2_a21oi_1 _14829_ (.A1(_06484_),
    .A2(_06485_),
    .Y(_00239_),
    .B1(net394));
 sg13g2_nor2_1 _14830_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[21] ),
    .B(net69),
    .Y(_06486_));
 sg13g2_a21oi_1 _14831_ (.A1(_04131_),
    .A2(_04132_),
    .Y(_06487_),
    .B1(net72));
 sg13g2_nor3_1 _14832_ (.A(net393),
    .B(_06486_),
    .C(_06487_),
    .Y(_00240_));
 sg13g2_nor2_1 _14833_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[22] ),
    .B(_06462_),
    .Y(_06488_));
 sg13g2_nor2_1 _14834_ (.A(_04179_),
    .B(net73),
    .Y(_06489_));
 sg13g2_nor3_1 _14835_ (.A(net393),
    .B(_06488_),
    .C(_06489_),
    .Y(_00241_));
 sg13g2_nor2_1 _14836_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[23] ),
    .B(net69),
    .Y(_06490_));
 sg13g2_nor2_1 _14837_ (.A(_04149_),
    .B(net73),
    .Y(_06491_));
 sg13g2_nor3_1 _14838_ (.A(net393),
    .B(_06490_),
    .C(_06491_),
    .Y(_00242_));
 sg13g2_buf_1 _14839_ (.A(net74),
    .X(_06492_));
 sg13g2_nor2_1 _14840_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[24] ),
    .B(net68),
    .Y(_06493_));
 sg13g2_nor2_1 _14841_ (.A(_04178_),
    .B(net73),
    .Y(_06494_));
 sg13g2_nor3_1 _14842_ (.A(net393),
    .B(_06493_),
    .C(_06494_),
    .Y(_00243_));
 sg13g2_nand2_1 _14843_ (.Y(_06495_),
    .A(_04175_),
    .B(net70));
 sg13g2_o21ai_1 _14844_ (.B1(_06495_),
    .Y(_06496_),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[25] ),
    .A2(net71));
 sg13g2_nor2_1 _14845_ (.A(net400),
    .B(_06496_),
    .Y(_00244_));
 sg13g2_nor2_1 _14846_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[26] ),
    .B(net68),
    .Y(_06497_));
 sg13g2_nor2_1 _14847_ (.A(_04621_),
    .B(net73),
    .Y(_06498_));
 sg13g2_nor3_1 _14848_ (.A(net393),
    .B(_06497_),
    .C(_06498_),
    .Y(_00245_));
 sg13g2_nand2_1 _14849_ (.Y(_06499_),
    .A(_04164_),
    .B(net70));
 sg13g2_o21ai_1 _14850_ (.B1(_06499_),
    .Y(_06500_),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[27] ),
    .A2(net71));
 sg13g2_nor2_1 _14851_ (.A(net400),
    .B(_06500_),
    .Y(_00246_));
 sg13g2_buf_1 _14852_ (.A(net523),
    .X(_06501_));
 sg13g2_nand2b_1 _14853_ (.Y(_06502_),
    .B(_06467_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.ALUOut[28] ));
 sg13g2_nand3_1 _14854_ (.B(_04173_),
    .C(net68),
    .A(_03761_),
    .Y(_06503_));
 sg13g2_and3_1 _14855_ (.X(_00247_),
    .A(net433),
    .B(_06502_),
    .C(_06503_));
 sg13g2_nor2_1 _14856_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[29] ),
    .B(_06492_),
    .Y(_06504_));
 sg13g2_and3_1 _14857_ (.X(_06505_),
    .A(_03592_),
    .B(_03600_),
    .C(net70));
 sg13g2_nor3_1 _14858_ (.A(net393),
    .B(_06504_),
    .C(_06505_),
    .Y(_00248_));
 sg13g2_mux2_1 _14859_ (.A0(_03846_),
    .A1(_03845_),
    .S(net70),
    .X(_06506_));
 sg13g2_nor2_1 _14860_ (.A(net400),
    .B(_06506_),
    .Y(_00249_));
 sg13g2_nor2_1 _14861_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[30] ),
    .B(net68),
    .Y(_06507_));
 sg13g2_nor2_1 _14862_ (.A(_03645_),
    .B(net73),
    .Y(_06508_));
 sg13g2_nor3_1 _14863_ (.A(net393),
    .B(_06507_),
    .C(_06508_),
    .Y(_00250_));
 sg13g2_buf_1 _14864_ (.A(_05918_),
    .X(_06509_));
 sg13g2_nor2_1 _14865_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[31] ),
    .B(net68),
    .Y(_06510_));
 sg13g2_nor2_1 _14866_ (.A(_04183_),
    .B(net73),
    .Y(_06511_));
 sg13g2_nor3_1 _14867_ (.A(net392),
    .B(_06510_),
    .C(_06511_),
    .Y(_00251_));
 sg13g2_nor2_1 _14868_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[3] ),
    .B(net68),
    .Y(_06512_));
 sg13g2_nor2_1 _14869_ (.A(_03827_),
    .B(net72),
    .Y(_06513_));
 sg13g2_nor3_1 _14870_ (.A(net392),
    .B(_06512_),
    .C(_06513_),
    .Y(_00252_));
 sg13g2_nand2_1 _14871_ (.Y(_06514_),
    .A(_03801_),
    .B(net74));
 sg13g2_o21ai_1 _14872_ (.B1(_06514_),
    .Y(_06515_),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[4] ),
    .A2(net71));
 sg13g2_nor2_1 _14873_ (.A(net400),
    .B(_06515_),
    .Y(_00253_));
 sg13g2_nor2_1 _14874_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[5] ),
    .B(_06492_),
    .Y(_06516_));
 sg13g2_nor2_1 _14875_ (.A(_04651_),
    .B(net72),
    .Y(_06517_));
 sg13g2_nor3_1 _14876_ (.A(net392),
    .B(_06516_),
    .C(_06517_),
    .Y(_00254_));
 sg13g2_nand2_1 _14877_ (.Y(_06518_),
    .A(_03899_),
    .B(net74));
 sg13g2_o21ai_1 _14878_ (.B1(_06518_),
    .Y(_06519_),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[6] ),
    .A2(_06453_));
 sg13g2_nor2_1 _14879_ (.A(net400),
    .B(_06519_),
    .Y(_00255_));
 sg13g2_nor2_1 _14880_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[7] ),
    .B(net68),
    .Y(_06520_));
 sg13g2_nor2_1 _14881_ (.A(_04663_),
    .B(net72),
    .Y(_06521_));
 sg13g2_nor3_1 _14882_ (.A(net392),
    .B(_06520_),
    .C(_06521_),
    .Y(_00256_));
 sg13g2_buf_1 _14883_ (.A(net438),
    .X(_06522_));
 sg13g2_nand2_1 _14884_ (.Y(_06523_),
    .A(_04122_),
    .B(net74));
 sg13g2_o21ai_1 _14885_ (.B1(_06523_),
    .Y(_06524_),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[8] ),
    .A2(_06453_));
 sg13g2_nor2_1 _14886_ (.A(_06522_),
    .B(_06524_),
    .Y(_00257_));
 sg13g2_nor2_1 _14887_ (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[9] ),
    .B(net68),
    .Y(_06525_));
 sg13g2_nor2_1 _14888_ (.A(_04144_),
    .B(net72),
    .Y(_06526_));
 sg13g2_nor3_1 _14889_ (.A(net392),
    .B(_06525_),
    .C(_06526_),
    .Y(_00258_));
 sg13g2_buf_1 _14890_ (.A(_04260_),
    .X(_06527_));
 sg13g2_nor2_1 _14891_ (.A(\soc_I.kianv_I.Instr[0] ),
    .B(net47),
    .Y(_06528_));
 sg13g2_buf_1 _14892_ (.A(net615),
    .X(_06529_));
 sg13g2_buf_1 _14893_ (.A(net542),
    .X(_06530_));
 sg13g2_buf_1 _14894_ (.A(net473),
    .X(_06531_));
 sg13g2_nor2_1 _14895_ (.A(_04106_),
    .B(_05795_),
    .Y(_06532_));
 sg13g2_buf_1 _14896_ (.A(_06532_),
    .X(_06533_));
 sg13g2_buf_1 _14897_ (.A(net351),
    .X(_06534_));
 sg13g2_buf_4 _14898_ (.X(_06535_),
    .A(_00000_));
 sg13g2_buf_2 _14899_ (.A(_06535_),
    .X(_06536_));
 sg13g2_buf_2 _14900_ (.A(_00001_),
    .X(_06537_));
 sg13g2_buf_1 _14901_ (.A(_06537_),
    .X(_06538_));
 sg13g2_mux4_1 _14902_ (.S0(net541),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][0] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][0] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][0] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][0] ),
    .S1(net540),
    .X(_06539_));
 sg13g2_mux4_1 _14903_ (.S0(net541),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][0] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][0] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][0] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][0] ),
    .S1(net540),
    .X(_06540_));
 sg13g2_mux4_1 _14904_ (.S0(net541),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[8][0] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][0] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][0] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[11][0] ),
    .S1(net540),
    .X(_06541_));
 sg13g2_mux4_1 _14905_ (.S0(net541),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[12][0] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][0] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][0] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[15][0] ),
    .S1(net540),
    .X(_06542_));
 sg13g2_buf_8 _14906_ (.A(_00002_),
    .X(_06543_));
 sg13g2_buf_4 _14907_ (.X(_06544_),
    .A(_00003_));
 sg13g2_mux4_1 _14908_ (.S0(_06543_),
    .A0(_06539_),
    .A1(_06540_),
    .A2(_06541_),
    .A3(_06542_),
    .S1(_06544_),
    .X(_06545_));
 sg13g2_inv_1 _14909_ (.Y(_06546_),
    .A(_06545_));
 sg13g2_buf_1 _14910_ (.A(net617),
    .X(_06547_));
 sg13g2_buf_1 _14911_ (.A(net618),
    .X(_06548_));
 sg13g2_buf_1 _14912_ (.A(net538),
    .X(_06549_));
 sg13g2_inv_1 _14913_ (.Y(_06550_),
    .A(_00061_));
 sg13g2_and2_1 _14914_ (.A(\soc_I.cycle_cnt_ready ),
    .B(_04101_),
    .X(_06551_));
 sg13g2_buf_1 _14915_ (.A(_06551_),
    .X(_06552_));
 sg13g2_buf_1 _14916_ (.A(_06552_),
    .X(_06553_));
 sg13g2_buf_1 _14917_ (.A(_06553_),
    .X(_06554_));
 sg13g2_a221oi_1 _14918_ (.B2(_05814_),
    .C1(net506),
    .B1(net350),
    .A1(_06549_),
    .Y(_06555_),
    .A2(_06550_));
 sg13g2_a21o_1 _14919_ (.A2(_03851_),
    .A1(net414),
    .B1(_03852_),
    .X(_06556_));
 sg13g2_buf_1 _14920_ (.A(_06556_),
    .X(_06557_));
 sg13g2_mux2_1 _14921_ (.A0(_00062_),
    .A1(_00063_),
    .S(_06557_),
    .X(_06558_));
 sg13g2_or3_1 _14922_ (.A(net472),
    .B(_04190_),
    .C(_06558_),
    .X(_06559_));
 sg13g2_buf_1 _14923_ (.A(_04103_),
    .X(_06560_));
 sg13g2_a221oi_1 _14924_ (.B2(_06559_),
    .C1(net537),
    .B1(_06555_),
    .A1(net436),
    .Y(_06561_),
    .A2(_00060_));
 sg13g2_nor2_1 _14925_ (.A(_06547_),
    .B(_06561_),
    .Y(_06562_));
 sg13g2_a21oi_1 _14926_ (.A1(net330),
    .A2(_06546_),
    .Y(_06563_),
    .B1(_06562_));
 sg13g2_nor2_1 _14927_ (.A(_04226_),
    .B(\soc_I.qqspi_I.ready ),
    .Y(_06564_));
 sg13g2_and2_1 _14928_ (.A(_04271_),
    .B(_06564_),
    .X(_06565_));
 sg13g2_buf_8 _14929_ (.A(_06565_),
    .X(_06566_));
 sg13g2_o21ai_1 _14930_ (.B1(net410),
    .Y(_06567_),
    .A1(_04269_),
    .A2(_04271_));
 sg13g2_buf_1 _14931_ (.A(_06567_),
    .X(_06568_));
 sg13g2_a221oi_1 _14932_ (.B2(_06566_),
    .C1(net46),
    .B1(_06563_),
    .A1(net432),
    .Y(_06569_),
    .A2(\soc_I.qqspi_I.rdata[0] ));
 sg13g2_nor3_1 _14933_ (.A(net392),
    .B(_06528_),
    .C(_06569_),
    .Y(_00259_));
 sg13g2_buf_8 _14934_ (.A(_04260_),
    .X(_06570_));
 sg13g2_buf_1 _14935_ (.A(_06570_),
    .X(_06571_));
 sg13g2_buf_1 _14936_ (.A(_06529_),
    .X(_06572_));
 sg13g2_nor2_1 _14937_ (.A(_03807_),
    .B(_04045_),
    .Y(_06573_));
 sg13g2_and2_1 _14938_ (.A(_04190_),
    .B(_04210_),
    .X(_06574_));
 sg13g2_nand4_1 _14939_ (.B(_06573_),
    .C(_04319_),
    .A(_03788_),
    .Y(_06575_),
    .D(_06574_));
 sg13g2_a21oi_1 _14940_ (.A1(_04116_),
    .A2(_04188_),
    .Y(_06576_),
    .B1(_06575_));
 sg13g2_nand3_1 _14941_ (.B(_04218_),
    .C(_06564_),
    .A(_04199_),
    .Y(_06577_));
 sg13g2_a221oi_1 _14942_ (.B2(_06576_),
    .C1(_06577_),
    .B1(_04112_),
    .A1(_03672_),
    .Y(_06578_),
    .A2(_04098_));
 sg13g2_buf_8 _14943_ (.A(_06578_),
    .X(_06579_));
 sg13g2_buf_1 _14944_ (.A(_06579_),
    .X(_06580_));
 sg13g2_buf_1 _14945_ (.A(net578),
    .X(_06581_));
 sg13g2_nor2b_1 _14946_ (.A(_05516_),
    .B_N(net470),
    .Y(_06582_));
 sg13g2_a221oi_1 _14947_ (.B2(net350),
    .C1(net470),
    .B1(\soc_I.cycle_cnt[10] ),
    .A1(net472),
    .Y(_06583_),
    .A2(_05674_));
 sg13g2_nor3_1 _14948_ (.A(net537),
    .B(_06582_),
    .C(_06583_),
    .Y(_06584_));
 sg13g2_nor2_1 _14949_ (.A(net539),
    .B(_06584_),
    .Y(_06585_));
 sg13g2_nor2_1 _14950_ (.A(net330),
    .B(_06585_),
    .Y(_06586_));
 sg13g2_a22oi_1 _14951_ (.Y(_06587_),
    .B1(_06580_),
    .B2(_06586_),
    .A2(\soc_I.qqspi_I.rdata[10] ),
    .A1(net471));
 sg13g2_o21ai_1 _14952_ (.B1(net433),
    .Y(_06588_),
    .A1(_02289_),
    .A2(net47));
 sg13g2_a21oi_1 _14953_ (.A1(net40),
    .A2(_06587_),
    .Y(_00260_),
    .B1(_06588_));
 sg13g2_nor2b_1 _14954_ (.A(net608),
    .B_N(net507),
    .Y(_06589_));
 sg13g2_a221oi_1 _14955_ (.B2(net350),
    .C1(net470),
    .B1(_05825_),
    .A1(net472),
    .Y(_06590_),
    .A2(_05713_));
 sg13g2_nor3_1 _14956_ (.A(net537),
    .B(_06589_),
    .C(_06590_),
    .Y(_06591_));
 sg13g2_nor2_1 _14957_ (.A(net539),
    .B(_06591_),
    .Y(_06592_));
 sg13g2_nor2_1 _14958_ (.A(net330),
    .B(_06592_),
    .Y(_06593_));
 sg13g2_a22oi_1 _14959_ (.Y(_06594_),
    .B1(net67),
    .B2(_06593_),
    .A2(\soc_I.qqspi_I.rdata[11] ),
    .A1(net471));
 sg13g2_o21ai_1 _14960_ (.B1(net433),
    .Y(_06595_),
    .A1(\soc_I.kianv_I.Instr[11] ),
    .A2(net47));
 sg13g2_a21oi_1 _14961_ (.A1(net40),
    .A2(_06594_),
    .Y(_00261_),
    .B1(_06595_));
 sg13g2_nor2b_1 _14962_ (.A(_05544_),
    .B_N(_05903_),
    .Y(_06596_));
 sg13g2_a221oi_1 _14963_ (.B2(net350),
    .C1(_06581_),
    .B1(\soc_I.cycle_cnt[12] ),
    .A1(net472),
    .Y(_06597_),
    .A2(_05714_));
 sg13g2_nor3_1 _14964_ (.A(_06560_),
    .B(_06596_),
    .C(_06597_),
    .Y(_06598_));
 sg13g2_nor2_1 _14965_ (.A(net539),
    .B(_06598_),
    .Y(_06599_));
 sg13g2_nor2_1 _14966_ (.A(net330),
    .B(_06599_),
    .Y(_06600_));
 sg13g2_a22oi_1 _14967_ (.Y(_06601_),
    .B1(net67),
    .B2(_06600_),
    .A2(\soc_I.qqspi_I.rdata[12] ),
    .A1(net471));
 sg13g2_o21ai_1 _14968_ (.B1(net433),
    .Y(_06602_),
    .A1(_05996_),
    .A2(net47));
 sg13g2_a21oi_1 _14969_ (.A1(_06571_),
    .A2(_06601_),
    .Y(_00262_),
    .B1(_06602_));
 sg13g2_nand2_1 _14970_ (.Y(_06603_),
    .A(_06530_),
    .B(\soc_I.qqspi_I.rdata[13] ));
 sg13g2_buf_1 _14971_ (.A(_05911_),
    .X(_06604_));
 sg13g2_a22oi_1 _14972_ (.Y(_06605_),
    .B1(\soc_I.cycle_cnt[13] ),
    .B2(_06554_),
    .A2(_05718_),
    .A1(net472));
 sg13g2_nor2_1 _14973_ (.A(net436),
    .B(_06605_),
    .Y(_06606_));
 sg13g2_a21oi_1 _14974_ (.A1(net431),
    .A2(_05560_),
    .Y(_06607_),
    .B1(_06606_));
 sg13g2_a21oi_1 _14975_ (.A1(net539),
    .A2(_05795_),
    .Y(_06608_),
    .B1(_04226_));
 sg13g2_o21ai_1 _14976_ (.B1(_06608_),
    .Y(_06609_),
    .A1(_04107_),
    .A2(_06607_));
 sg13g2_nor2b_1 _14977_ (.A(_05448_),
    .B_N(_04226_),
    .Y(_06610_));
 sg13g2_nor2_1 _14978_ (.A(net542),
    .B(_06610_),
    .Y(_06611_));
 sg13g2_nand3_1 _14979_ (.B(_06609_),
    .C(_06611_),
    .A(_04271_),
    .Y(_06612_));
 sg13g2_and2_1 _14980_ (.A(_06603_),
    .B(_06612_),
    .X(_06613_));
 sg13g2_o21ai_1 _14981_ (.B1(net433),
    .Y(_06614_),
    .A1(net434),
    .A2(net47));
 sg13g2_a21oi_1 _14982_ (.A1(net40),
    .A2(_06613_),
    .Y(_00263_),
    .B1(_06614_));
 sg13g2_nand2_1 _14983_ (.Y(_06615_),
    .A(net471),
    .B(\soc_I.qqspi_I.rdata[14] ));
 sg13g2_a22oi_1 _14984_ (.Y(_06616_),
    .B1(_05834_),
    .B2(_06554_),
    .A2(_05734_),
    .A1(net472));
 sg13g2_nor2_1 _14985_ (.A(net436),
    .B(_06616_),
    .Y(_06617_));
 sg13g2_a21oi_1 _14986_ (.A1(_06604_),
    .A2(_05568_),
    .Y(_06618_),
    .B1(_06617_));
 sg13g2_o21ai_1 _14987_ (.B1(_06608_),
    .Y(_06619_),
    .A1(_04107_),
    .A2(_06618_));
 sg13g2_nand3_1 _14988_ (.B(_06611_),
    .C(_06619_),
    .A(_04271_),
    .Y(_06620_));
 sg13g2_and2_1 _14989_ (.A(_06615_),
    .B(_06620_),
    .X(_06621_));
 sg13g2_o21ai_1 _14990_ (.B1(net433),
    .Y(_06622_),
    .A1(net602),
    .A2(_06527_));
 sg13g2_a21oi_1 _14991_ (.A1(_06571_),
    .A2(_06621_),
    .Y(_00264_),
    .B1(_06622_));
 sg13g2_a22oi_1 _14992_ (.Y(_06623_),
    .B1(_05837_),
    .B2(_06552_),
    .A2(_05731_),
    .A1(net618));
 sg13g2_nor2_1 _14993_ (.A(_05902_),
    .B(_06623_),
    .Y(_06624_));
 sg13g2_a21oi_1 _14994_ (.A1(_05902_),
    .A2(_05581_),
    .Y(_06625_),
    .B1(_06624_));
 sg13g2_buf_1 _14995_ (.A(_04106_),
    .X(_06626_));
 sg13g2_o21ai_1 _14996_ (.B1(net469),
    .Y(_06627_),
    .A1(_04103_),
    .A2(_06625_));
 sg13g2_inv_1 _14997_ (.Y(_06628_),
    .A(_05795_));
 sg13g2_nand2_1 _14998_ (.Y(_06629_),
    .A(net617),
    .B(_06628_));
 sg13g2_and4_1 _14999_ (.A(_04238_),
    .B(_04256_),
    .C(_06629_),
    .D(_06579_),
    .X(_06630_));
 sg13g2_buf_2 _15000_ (.A(_06630_),
    .X(_06631_));
 sg13g2_buf_8 _15001_ (.A(_06631_),
    .X(_06632_));
 sg13g2_a22oi_1 _15002_ (.Y(_06633_),
    .B1(_06627_),
    .B2(net57),
    .A2(\soc_I.qqspi_I.rdata[15] ),
    .A1(net432));
 sg13g2_buf_1 _15003_ (.A(net523),
    .X(_06634_));
 sg13g2_o21ai_1 _15004_ (.B1(net430),
    .Y(_06635_),
    .A1(_06053_),
    .A2(_06527_));
 sg13g2_a21oi_1 _15005_ (.A1(net40),
    .A2(_06633_),
    .Y(_00265_),
    .B1(_06635_));
 sg13g2_a22oi_1 _15006_ (.Y(_06636_),
    .B1(net350),
    .B2(\soc_I.cycle_cnt[16] ),
    .A2(\soc_I.spi_div_reg[16] ),
    .A1(_06549_));
 sg13g2_nand2_1 _15007_ (.Y(_06637_),
    .A(_05911_),
    .B(\soc_I.div_reg[16] ));
 sg13g2_o21ai_1 _15008_ (.B1(_06637_),
    .Y(_06638_),
    .A1(net431),
    .A2(_06636_));
 sg13g2_a21oi_1 _15009_ (.A1(_04104_),
    .A2(_06638_),
    .Y(_06639_),
    .B1(net539));
 sg13g2_inv_1 _15010_ (.Y(_06640_),
    .A(_06639_));
 sg13g2_a22oi_1 _15011_ (.Y(_06641_),
    .B1(net57),
    .B2(_06640_),
    .A2(\soc_I.qqspi_I.rdata[16] ),
    .A1(_06530_));
 sg13g2_buf_1 _15012_ (.A(_04260_),
    .X(_06642_));
 sg13g2_o21ai_1 _15013_ (.B1(net430),
    .Y(_06643_),
    .A1(net500),
    .A2(net45));
 sg13g2_a21oi_1 _15014_ (.A1(net40),
    .A2(_06641_),
    .Y(_00266_),
    .B1(_06643_));
 sg13g2_buf_1 _15015_ (.A(net537),
    .X(_06644_));
 sg13g2_buf_1 _15016_ (.A(net538),
    .X(_06645_));
 sg13g2_buf_1 _15017_ (.A(_06553_),
    .X(_06646_));
 sg13g2_a22oi_1 _15018_ (.Y(_06647_),
    .B1(net349),
    .B2(\soc_I.cycle_cnt[17] ),
    .A2(\soc_I.spi_div_reg[17] ),
    .A1(net467));
 sg13g2_nor2_1 _15019_ (.A(net431),
    .B(_06647_),
    .Y(_06648_));
 sg13g2_a21oi_1 _15020_ (.A1(net399),
    .A2(\soc_I.div_reg[17] ),
    .Y(_06649_),
    .B1(_06648_));
 sg13g2_o21ai_1 _15021_ (.B1(net469),
    .Y(_06650_),
    .A1(net468),
    .A2(_06649_));
 sg13g2_a22oi_1 _15022_ (.Y(_06651_),
    .B1(_06631_),
    .B2(_06650_),
    .A2(\soc_I.qqspi_I.rdata[17] ),
    .A1(net471));
 sg13g2_o21ai_1 _15023_ (.B1(net430),
    .Y(_06652_),
    .A1(_06071_),
    .A2(net45));
 sg13g2_a21oi_1 _15024_ (.A1(net40),
    .A2(_06651_),
    .Y(_00267_),
    .B1(_06652_));
 sg13g2_a22oi_1 _15025_ (.Y(_06653_),
    .B1(net349),
    .B2(_05846_),
    .A2(\soc_I.spi_div_reg[18] ),
    .A1(net467));
 sg13g2_nor2_1 _15026_ (.A(net431),
    .B(_06653_),
    .Y(_06654_));
 sg13g2_a21oi_1 _15027_ (.A1(net399),
    .A2(\soc_I.div_reg[18] ),
    .Y(_06655_),
    .B1(_06654_));
 sg13g2_o21ai_1 _15028_ (.B1(net469),
    .Y(_06656_),
    .A1(net468),
    .A2(_06655_));
 sg13g2_a22oi_1 _15029_ (.Y(_06657_),
    .B1(_06631_),
    .B2(_06656_),
    .A2(\soc_I.qqspi_I.rdata[18] ),
    .A1(net471));
 sg13g2_o21ai_1 _15030_ (.B1(_06634_),
    .Y(_06658_),
    .A1(net572),
    .A2(_06642_));
 sg13g2_a21oi_1 _15031_ (.A1(net40),
    .A2(_06657_),
    .Y(_00268_),
    .B1(_06658_));
 sg13g2_a22oi_1 _15032_ (.Y(_06659_),
    .B1(net349),
    .B2(\soc_I.cycle_cnt[19] ),
    .A2(\soc_I.spi_div_reg[19] ),
    .A1(net467));
 sg13g2_nor2_1 _15033_ (.A(net431),
    .B(_06659_),
    .Y(_06660_));
 sg13g2_a21oi_1 _15034_ (.A1(net399),
    .A2(\soc_I.div_reg[19] ),
    .Y(_06661_),
    .B1(_06660_));
 sg13g2_o21ai_1 _15035_ (.B1(_06626_),
    .Y(_06662_),
    .A1(net468),
    .A2(_06661_));
 sg13g2_a22oi_1 _15036_ (.Y(_06663_),
    .B1(_06631_),
    .B2(_06662_),
    .A2(\soc_I.qqspi_I.rdata[19] ),
    .A1(net471));
 sg13g2_o21ai_1 _15037_ (.B1(_06634_),
    .Y(_06664_),
    .A1(\soc_I.kianv_I.Instr[19] ),
    .A2(_06642_));
 sg13g2_a21oi_1 _15038_ (.A1(net40),
    .A2(_06663_),
    .Y(_00269_),
    .B1(_06664_));
 sg13g2_buf_1 _15039_ (.A(_06570_),
    .X(_06665_));
 sg13g2_buf_1 _15040_ (.A(_06547_),
    .X(_06666_));
 sg13g2_inv_1 _15041_ (.Y(_06667_),
    .A(_00065_));
 sg13g2_a221oi_1 _15042_ (.B2(_05815_),
    .C1(net436),
    .B1(net349),
    .A1(net467),
    .Y(_06668_),
    .A2(_06667_));
 sg13g2_nor3_1 _15043_ (.A(_04100_),
    .B(_03854_),
    .C(_04190_),
    .Y(_06669_));
 sg13g2_buf_2 _15044_ (.A(_06669_),
    .X(_06670_));
 sg13g2_nand2_1 _15045_ (.Y(_06671_),
    .A(\soc_I.spi0_I.rx_data[1] ),
    .B(_06670_));
 sg13g2_a221oi_1 _15046_ (.B2(_06671_),
    .C1(net468),
    .B1(_06668_),
    .A1(net399),
    .Y(_06672_),
    .A2(_00064_));
 sg13g2_buf_2 _15047_ (.A(net541),
    .X(_06673_));
 sg13g2_buf_1 _15048_ (.A(net540),
    .X(_06674_));
 sg13g2_mux4_1 _15049_ (.S0(net465),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][1] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][1] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][1] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][1] ),
    .S1(net464),
    .X(_06675_));
 sg13g2_mux4_1 _15050_ (.S0(net465),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][1] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][1] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][1] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][1] ),
    .S1(net464),
    .X(_06676_));
 sg13g2_buf_2 _15051_ (.A(net541),
    .X(_06677_));
 sg13g2_buf_1 _15052_ (.A(net540),
    .X(_06678_));
 sg13g2_mux4_1 _15053_ (.S0(net463),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[8][1] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][1] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][1] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[11][1] ),
    .S1(net462),
    .X(_06679_));
 sg13g2_mux4_1 _15054_ (.S0(net463),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[12][1] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][1] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][1] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[15][1] ),
    .S1(net462),
    .X(_06680_));
 sg13g2_mux4_1 _15055_ (.S0(_06543_),
    .A0(_06675_),
    .A1(_06676_),
    .A2(_06679_),
    .A3(_06680_),
    .S1(_06544_),
    .X(_06681_));
 sg13g2_nand2b_1 _15056_ (.Y(_06682_),
    .B(_06534_),
    .A_N(_06681_));
 sg13g2_o21ai_1 _15057_ (.B1(_06682_),
    .Y(_06683_),
    .A1(net466),
    .A2(_06672_));
 sg13g2_inv_1 _15058_ (.Y(_06684_),
    .A(_06683_));
 sg13g2_a22oi_1 _15059_ (.Y(_06685_),
    .B1(_06566_),
    .B2(_06684_),
    .A2(\soc_I.qqspi_I.rdata[1] ),
    .A1(net473));
 sg13g2_o21ai_1 _15060_ (.B1(net430),
    .Y(_06686_),
    .A1(\soc_I.kianv_I.Instr[1] ),
    .A2(net45));
 sg13g2_a21oi_1 _15061_ (.A1(net39),
    .A2(_06685_),
    .Y(_00270_),
    .B1(_06686_));
 sg13g2_a22oi_1 _15062_ (.Y(_06687_),
    .B1(net349),
    .B2(\soc_I.cycle_cnt[20] ),
    .A2(\soc_I.spi_div_reg[20] ),
    .A1(net467));
 sg13g2_nor2_1 _15063_ (.A(net431),
    .B(_06687_),
    .Y(_06688_));
 sg13g2_a21oi_1 _15064_ (.A1(net399),
    .A2(\soc_I.div_reg[20] ),
    .Y(_06689_),
    .B1(_06688_));
 sg13g2_o21ai_1 _15065_ (.B1(_06626_),
    .Y(_06690_),
    .A1(net468),
    .A2(_06689_));
 sg13g2_a22oi_1 _15066_ (.Y(_06691_),
    .B1(_06631_),
    .B2(_06690_),
    .A2(\soc_I.qqspi_I.rdata[20] ),
    .A1(_06572_));
 sg13g2_o21ai_1 _15067_ (.B1(net430),
    .Y(_06692_),
    .A1(net486),
    .A2(net45));
 sg13g2_a21oi_1 _15068_ (.A1(net39),
    .A2(_06691_),
    .Y(_00271_),
    .B1(_06692_));
 sg13g2_buf_1 _15069_ (.A(_06570_),
    .X(_06693_));
 sg13g2_a22oi_1 _15070_ (.Y(_06694_),
    .B1(net350),
    .B2(_05855_),
    .A2(\soc_I.spi_div_reg[21] ),
    .A1(net472));
 sg13g2_nor2_1 _15071_ (.A(net506),
    .B(_06694_),
    .Y(_06695_));
 sg13g2_a21oi_1 _15072_ (.A1(net431),
    .A2(\soc_I.div_reg[21] ),
    .Y(_06696_),
    .B1(_06695_));
 sg13g2_o21ai_1 _15073_ (.B1(net469),
    .Y(_06697_),
    .A1(net537),
    .A2(_06696_));
 sg13g2_and2_1 _15074_ (.A(_06529_),
    .B(\soc_I.qqspi_I.rdata[21] ),
    .X(_06698_));
 sg13g2_a21o_1 _15075_ (.A2(_06697_),
    .A1(net57),
    .B1(_06698_),
    .X(_06699_));
 sg13g2_nand2_1 _15076_ (.Y(_06700_),
    .A(net38),
    .B(_06699_));
 sg13g2_buf_8 _15077_ (.A(net46),
    .X(_06701_));
 sg13g2_nand2_1 _15078_ (.Y(_06702_),
    .A(net485),
    .B(_06701_));
 sg13g2_buf_1 _15079_ (.A(_06002_),
    .X(_06703_));
 sg13g2_a21oi_1 _15080_ (.A1(_06700_),
    .A2(_06702_),
    .Y(_00272_),
    .B1(_06703_));
 sg13g2_a22oi_1 _15081_ (.Y(_06704_),
    .B1(net350),
    .B2(\soc_I.cycle_cnt[22] ),
    .A2(\soc_I.spi_div_reg[22] ),
    .A1(_06548_));
 sg13g2_nor2_1 _15082_ (.A(net506),
    .B(_06704_),
    .Y(_06705_));
 sg13g2_a21oi_1 _15083_ (.A1(net431),
    .A2(\soc_I.div_reg[22] ),
    .Y(_06706_),
    .B1(_06705_));
 sg13g2_o21ai_1 _15084_ (.B1(net469),
    .Y(_06707_),
    .A1(net537),
    .A2(_06706_));
 sg13g2_and2_1 _15085_ (.A(net542),
    .B(\soc_I.qqspi_I.rdata[22] ),
    .X(_06708_));
 sg13g2_a21o_1 _15086_ (.A2(_06707_),
    .A1(net57),
    .B1(_06708_),
    .X(_06709_));
 sg13g2_nand2_1 _15087_ (.Y(_06710_),
    .A(net38),
    .B(_06709_));
 sg13g2_nand2_1 _15088_ (.Y(_06711_),
    .A(net555),
    .B(_06701_));
 sg13g2_a21oi_1 _15089_ (.A1(_06710_),
    .A2(_06711_),
    .Y(_00273_),
    .B1(_06703_));
 sg13g2_a22oi_1 _15090_ (.Y(_06712_),
    .B1(_06552_),
    .B2(\soc_I.cycle_cnt[23] ),
    .A2(\soc_I.spi_div_reg[23] ),
    .A1(net618));
 sg13g2_nor2_1 _15091_ (.A(net578),
    .B(_06712_),
    .Y(_06713_));
 sg13g2_a21oi_1 _15092_ (.A1(net578),
    .A2(\soc_I.div_reg[23] ),
    .Y(_06714_),
    .B1(_06713_));
 sg13g2_o21ai_1 _15093_ (.B1(net469),
    .Y(_06715_),
    .A1(_04103_),
    .A2(_06714_));
 sg13g2_and2_1 _15094_ (.A(_06629_),
    .B(_06715_),
    .X(_06716_));
 sg13g2_a22oi_1 _15095_ (.Y(_06717_),
    .B1(_06579_),
    .B2(_06716_),
    .A2(\soc_I.qqspi_I.rdata[23] ),
    .A1(net542));
 sg13g2_o21ai_1 _15096_ (.B1(net430),
    .Y(_06718_),
    .A1(net554),
    .A2(net45));
 sg13g2_a21oi_1 _15097_ (.A1(net39),
    .A2(_06717_),
    .Y(_00274_),
    .B1(_06718_));
 sg13g2_a22oi_1 _15098_ (.Y(_06719_),
    .B1(net390),
    .B2(_05863_),
    .A2(\soc_I.spi_div_reg[24] ),
    .A1(net618));
 sg13g2_nor2_1 _15099_ (.A(net578),
    .B(_06719_),
    .Y(_06720_));
 sg13g2_a21oi_1 _15100_ (.A1(net507),
    .A2(\soc_I.div_reg[24] ),
    .Y(_06721_),
    .B1(_06720_));
 sg13g2_o21ai_1 _15101_ (.B1(net469),
    .Y(_06722_),
    .A1(net537),
    .A2(_06721_));
 sg13g2_and2_1 _15102_ (.A(_06629_),
    .B(_06722_),
    .X(_06723_));
 sg13g2_and2_1 _15103_ (.A(net615),
    .B(\soc_I.qqspi_I.rdata[24] ),
    .X(_06724_));
 sg13g2_a21o_1 _15104_ (.A2(_06723_),
    .A1(_06579_),
    .B1(_06724_),
    .X(_06725_));
 sg13g2_buf_1 _15105_ (.A(_06725_),
    .X(_06726_));
 sg13g2_inv_1 _15106_ (.Y(_06727_),
    .A(_06726_));
 sg13g2_o21ai_1 _15107_ (.B1(net430),
    .Y(_06728_),
    .A1(\soc_I.kianv_I.Instr[24] ),
    .A2(net45));
 sg13g2_a21oi_1 _15108_ (.A1(net39),
    .A2(_06727_),
    .Y(_00275_),
    .B1(_06728_));
 sg13g2_a22oi_1 _15109_ (.Y(_06729_),
    .B1(net390),
    .B2(\soc_I.cycle_cnt[25] ),
    .A2(\soc_I.spi_div_reg[25] ),
    .A1(net538));
 sg13g2_nand2_1 _15110_ (.Y(_06730_),
    .A(net507),
    .B(\soc_I.div_reg[25] ));
 sg13g2_o21ai_1 _15111_ (.B1(_06730_),
    .Y(_06731_),
    .A1(net506),
    .A2(_06729_));
 sg13g2_a21oi_1 _15112_ (.A1(net594),
    .A2(_06731_),
    .Y(_06732_),
    .B1(net617));
 sg13g2_nor2_1 _15113_ (.A(net351),
    .B(_06732_),
    .Y(_06733_));
 sg13g2_and2_1 _15114_ (.A(net542),
    .B(\soc_I.qqspi_I.rdata[25] ),
    .X(_06734_));
 sg13g2_a21o_1 _15115_ (.A2(_06733_),
    .A1(_06580_),
    .B1(_06734_),
    .X(_06735_));
 sg13g2_buf_1 _15116_ (.A(_06735_),
    .X(_06736_));
 sg13g2_inv_1 _15117_ (.Y(_06737_),
    .A(_06736_));
 sg13g2_o21ai_1 _15118_ (.B1(net430),
    .Y(_06738_),
    .A1(\soc_I.kianv_I.Instr[25] ),
    .A2(net45));
 sg13g2_a21oi_1 _15119_ (.A1(net39),
    .A2(_06737_),
    .Y(_00276_),
    .B1(_06738_));
 sg13g2_a22oi_1 _15120_ (.Y(_06739_),
    .B1(net390),
    .B2(\soc_I.cycle_cnt[26] ),
    .A2(\soc_I.spi_div_reg[26] ),
    .A1(net538));
 sg13g2_nand2_1 _15121_ (.Y(_06740_),
    .A(net507),
    .B(\soc_I.div_reg[26] ));
 sg13g2_o21ai_1 _15122_ (.B1(_06740_),
    .Y(_06741_),
    .A1(net506),
    .A2(_06739_));
 sg13g2_a21oi_1 _15123_ (.A1(net594),
    .A2(_06741_),
    .Y(_06742_),
    .B1(net617));
 sg13g2_nor2_1 _15124_ (.A(net351),
    .B(_06742_),
    .Y(_06743_));
 sg13g2_and2_1 _15125_ (.A(net615),
    .B(\soc_I.qqspi_I.rdata[26] ),
    .X(_06744_));
 sg13g2_a21o_1 _15126_ (.A2(_06743_),
    .A1(net67),
    .B1(_06744_),
    .X(_06745_));
 sg13g2_buf_1 _15127_ (.A(_06745_),
    .X(_06746_));
 sg13g2_inv_1 _15128_ (.Y(_06747_),
    .A(_06746_));
 sg13g2_buf_1 _15129_ (.A(net523),
    .X(_06748_));
 sg13g2_o21ai_1 _15130_ (.B1(net429),
    .Y(_06749_),
    .A1(\soc_I.kianv_I.Instr[26] ),
    .A2(net45));
 sg13g2_a21oi_1 _15131_ (.A1(_06665_),
    .A2(_06747_),
    .Y(_00277_),
    .B1(_06749_));
 sg13g2_a22oi_1 _15132_ (.Y(_06750_),
    .B1(net390),
    .B2(_05872_),
    .A2(\soc_I.spi_div_reg[27] ),
    .A1(net538));
 sg13g2_nand2_1 _15133_ (.Y(_06751_),
    .A(net507),
    .B(\soc_I.div_reg[27] ));
 sg13g2_o21ai_1 _15134_ (.B1(_06751_),
    .Y(_06752_),
    .A1(net470),
    .A2(_06750_));
 sg13g2_a21oi_1 _15135_ (.A1(net594),
    .A2(_06752_),
    .Y(_06753_),
    .B1(net617));
 sg13g2_nor2_1 _15136_ (.A(net351),
    .B(_06753_),
    .Y(_06754_));
 sg13g2_and2_1 _15137_ (.A(net615),
    .B(\soc_I.qqspi_I.rdata[27] ),
    .X(_06755_));
 sg13g2_a21o_1 _15138_ (.A2(_06754_),
    .A1(net67),
    .B1(_06755_),
    .X(_06756_));
 sg13g2_buf_1 _15139_ (.A(_06756_),
    .X(_06757_));
 sg13g2_inv_1 _15140_ (.Y(_06758_),
    .A(_06757_));
 sg13g2_buf_1 _15141_ (.A(_04260_),
    .X(_06759_));
 sg13g2_o21ai_1 _15142_ (.B1(net429),
    .Y(_06760_),
    .A1(_02322_),
    .A2(net44));
 sg13g2_a21oi_1 _15143_ (.A1(_06665_),
    .A2(_06758_),
    .Y(_00278_),
    .B1(_06760_));
 sg13g2_a22oi_1 _15144_ (.Y(_06761_),
    .B1(net390),
    .B2(_05875_),
    .A2(\soc_I.spi_div_reg[28] ),
    .A1(net538));
 sg13g2_nand2_1 _15145_ (.Y(_06762_),
    .A(net507),
    .B(\soc_I.div_reg[28] ));
 sg13g2_o21ai_1 _15146_ (.B1(_06762_),
    .Y(_06763_),
    .A1(net470),
    .A2(_06761_));
 sg13g2_a21oi_1 _15147_ (.A1(net594),
    .A2(_06763_),
    .Y(_06764_),
    .B1(net617));
 sg13g2_nor2_1 _15148_ (.A(net351),
    .B(_06764_),
    .Y(_06765_));
 sg13g2_and2_1 _15149_ (.A(net615),
    .B(\soc_I.qqspi_I.rdata[28] ),
    .X(_06766_));
 sg13g2_a21o_1 _15150_ (.A2(_06765_),
    .A1(_06579_),
    .B1(_06766_),
    .X(_06767_));
 sg13g2_buf_1 _15151_ (.A(_06767_),
    .X(_06768_));
 sg13g2_inv_1 _15152_ (.Y(_06769_),
    .A(_06768_));
 sg13g2_o21ai_1 _15153_ (.B1(_06748_),
    .Y(_06770_),
    .A1(_01934_),
    .A2(_06759_));
 sg13g2_a21oi_1 _15154_ (.A1(net39),
    .A2(_06769_),
    .Y(_00279_),
    .B1(_06770_));
 sg13g2_a22oi_1 _15155_ (.Y(_06771_),
    .B1(net390),
    .B2(\soc_I.cycle_cnt[29] ),
    .A2(\soc_I.spi_div_reg[29] ),
    .A1(net538));
 sg13g2_nand2_1 _15156_ (.Y(_06772_),
    .A(net470),
    .B(\soc_I.div_reg[29] ));
 sg13g2_o21ai_1 _15157_ (.B1(_06772_),
    .Y(_06773_),
    .A1(net506),
    .A2(_06771_));
 sg13g2_a21oi_1 _15158_ (.A1(net594),
    .A2(_06773_),
    .Y(_06774_),
    .B1(net539));
 sg13g2_nor2_1 _15159_ (.A(net330),
    .B(_06774_),
    .Y(_06775_));
 sg13g2_a22oi_1 _15160_ (.Y(_06776_),
    .B1(net67),
    .B2(_06775_),
    .A2(\soc_I.qqspi_I.rdata[29] ),
    .A1(_06572_));
 sg13g2_o21ai_1 _15161_ (.B1(_06748_),
    .Y(_06777_),
    .A1(_01950_),
    .A2(_06759_));
 sg13g2_a21oi_1 _15162_ (.A1(net39),
    .A2(_06776_),
    .Y(_00280_),
    .B1(_06777_));
 sg13g2_inv_1 _15163_ (.Y(_06778_),
    .A(_00067_));
 sg13g2_a221oi_1 _15164_ (.B2(_05816_),
    .C1(net436),
    .B1(net349),
    .A1(net467),
    .Y(_06779_),
    .A2(_06778_));
 sg13g2_nand2_1 _15165_ (.Y(_06780_),
    .A(\soc_I.spi0_I.rx_data[2] ),
    .B(_06670_));
 sg13g2_a221oi_1 _15166_ (.B2(_06780_),
    .C1(net468),
    .B1(_06779_),
    .A1(net399),
    .Y(_06781_),
    .A2(_00066_));
 sg13g2_mux4_1 _15167_ (.S0(_06677_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][2] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][2] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][2] ),
    .S1(_06678_),
    .X(_06782_));
 sg13g2_mux4_1 _15168_ (.S0(net465),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][2] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][2] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][2] ),
    .S1(net464),
    .X(_06783_));
 sg13g2_mux4_1 _15169_ (.S0(net541),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[8][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][2] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][2] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[11][2] ),
    .S1(net540),
    .X(_06784_));
 sg13g2_mux4_1 _15170_ (.S0(net463),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[12][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][2] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][2] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[15][2] ),
    .S1(net462),
    .X(_06785_));
 sg13g2_mux4_1 _15171_ (.S0(_06543_),
    .A0(_06782_),
    .A1(_06783_),
    .A2(_06784_),
    .A3(_06785_),
    .S1(_06544_),
    .X(_06786_));
 sg13g2_nand2b_1 _15172_ (.Y(_06787_),
    .B(net351),
    .A_N(_06786_));
 sg13g2_o21ai_1 _15173_ (.B1(_06787_),
    .Y(_06788_),
    .A1(net466),
    .A2(_06781_));
 sg13g2_inv_1 _15174_ (.Y(_06789_),
    .A(_06788_));
 sg13g2_a22oi_1 _15175_ (.Y(_06790_),
    .B1(_06566_),
    .B2(_06789_),
    .A2(\soc_I.qqspi_I.rdata[2] ),
    .A1(net473));
 sg13g2_o21ai_1 _15176_ (.B1(net429),
    .Y(_06791_),
    .A1(_01652_),
    .A2(net44));
 sg13g2_a21oi_1 _15177_ (.A1(net39),
    .A2(_06790_),
    .Y(_00281_),
    .B1(_06791_));
 sg13g2_a22oi_1 _15178_ (.Y(_06792_),
    .B1(net390),
    .B2(\soc_I.cycle_cnt[30] ),
    .A2(\soc_I.spi_div_reg[30] ),
    .A1(net538));
 sg13g2_nand2_1 _15179_ (.Y(_06793_),
    .A(net470),
    .B(\soc_I.div_reg[30] ));
 sg13g2_o21ai_1 _15180_ (.B1(_06793_),
    .Y(_06794_),
    .A1(net506),
    .A2(_06792_));
 sg13g2_a21oi_1 _15181_ (.A1(net594),
    .A2(_06794_),
    .Y(_06795_),
    .B1(net539));
 sg13g2_nor2_1 _15182_ (.A(net330),
    .B(_06795_),
    .Y(_06796_));
 sg13g2_a22oi_1 _15183_ (.Y(_06797_),
    .B1(net67),
    .B2(_06796_),
    .A2(\soc_I.qqspi_I.rdata[30] ),
    .A1(net542));
 sg13g2_o21ai_1 _15184_ (.B1(net429),
    .Y(_06798_),
    .A1(\soc_I.kianv_I.Instr[30] ),
    .A2(net44));
 sg13g2_a21oi_1 _15185_ (.A1(net38),
    .A2(_06797_),
    .Y(_00282_),
    .B1(_06798_));
 sg13g2_inv_1 _15186_ (.Y(_06799_),
    .A(_00079_));
 sg13g2_a221oi_1 _15187_ (.B2(\soc_I.cycle_cnt[31] ),
    .C1(net578),
    .B1(_06552_),
    .A1(net618),
    .Y(_06800_),
    .A2(_06799_));
 sg13g2_nor4_1 _15188_ (.A(_05745_),
    .B(\soc_I.spi0_I.xfer_cycles[5] ),
    .C(_05746_),
    .D(_05749_),
    .Y(_06801_));
 sg13g2_buf_1 _15189_ (.A(_06801_),
    .X(_06802_));
 sg13g2_or4_1 _15190_ (.A(net618),
    .B(_06557_),
    .C(_04190_),
    .D(_06802_),
    .X(_06803_));
 sg13g2_a221oi_1 _15191_ (.B2(_06803_),
    .C1(_04103_),
    .B1(_06800_),
    .A1(net578),
    .Y(_06804_),
    .A2(_00078_));
 sg13g2_nor2_1 _15192_ (.A(net617),
    .B(_06804_),
    .Y(_06805_));
 sg13g2_inv_1 _15193_ (.Y(_06806_),
    .A(_06805_));
 sg13g2_a22oi_1 _15194_ (.Y(_06807_),
    .B1(_06631_),
    .B2(_06806_),
    .A2(\soc_I.qqspi_I.rdata[31] ),
    .A1(net473));
 sg13g2_o21ai_1 _15195_ (.B1(net429),
    .Y(_06808_),
    .A1(_01819_),
    .A2(net44));
 sg13g2_a21oi_1 _15196_ (.A1(net38),
    .A2(_06807_),
    .Y(_00283_),
    .B1(_06808_));
 sg13g2_inv_1 _15197_ (.Y(_06809_),
    .A(_00069_));
 sg13g2_a221oi_1 _15198_ (.B2(\soc_I.cycle_cnt[3] ),
    .C1(net436),
    .B1(net349),
    .A1(net467),
    .Y(_06810_),
    .A2(_06809_));
 sg13g2_nand2_1 _15199_ (.Y(_06811_),
    .A(\soc_I.spi0_I.rx_data[3] ),
    .B(_06670_));
 sg13g2_a221oi_1 _15200_ (.B2(_06811_),
    .C1(net468),
    .B1(_06810_),
    .A1(net399),
    .Y(_06812_),
    .A2(_00068_));
 sg13g2_mux4_1 _15201_ (.S0(net463),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][3] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][3] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][3] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][3] ),
    .S1(net462),
    .X(_06813_));
 sg13g2_mux4_1 _15202_ (.S0(_06673_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][3] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][3] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][3] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][3] ),
    .S1(_06674_),
    .X(_06814_));
 sg13g2_mux4_1 _15203_ (.S0(_06536_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[8][3] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][3] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][3] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[11][3] ),
    .S1(_06538_),
    .X(_06815_));
 sg13g2_mux4_1 _15204_ (.S0(net463),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[12][3] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][3] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][3] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[15][3] ),
    .S1(net462),
    .X(_06816_));
 sg13g2_mux4_1 _15205_ (.S0(_06543_),
    .A0(_06813_),
    .A1(_06814_),
    .A2(_06815_),
    .A3(_06816_),
    .S1(_06544_),
    .X(_06817_));
 sg13g2_nand2b_1 _15206_ (.Y(_06818_),
    .B(net351),
    .A_N(_06817_));
 sg13g2_o21ai_1 _15207_ (.B1(_06818_),
    .Y(_06819_),
    .A1(net466),
    .A2(_06812_));
 sg13g2_inv_1 _15208_ (.Y(_06820_),
    .A(_06819_));
 sg13g2_a22oi_1 _15209_ (.Y(_06821_),
    .B1(_06566_),
    .B2(_06820_),
    .A2(\soc_I.qqspi_I.rdata[3] ),
    .A1(net473));
 sg13g2_o21ai_1 _15210_ (.B1(net429),
    .Y(_06822_),
    .A1(_01642_),
    .A2(net44));
 sg13g2_a21oi_1 _15211_ (.A1(_06693_),
    .A2(_06821_),
    .Y(_00284_),
    .B1(_06822_));
 sg13g2_inv_1 _15212_ (.Y(_06823_),
    .A(_00071_));
 sg13g2_a221oi_1 _15213_ (.B2(\soc_I.cycle_cnt[4] ),
    .C1(_05904_),
    .B1(net349),
    .A1(net467),
    .Y(_06824_),
    .A2(_06823_));
 sg13g2_nand2_1 _15214_ (.Y(_06825_),
    .A(\soc_I.spi0_I.rx_data[4] ),
    .B(_06670_));
 sg13g2_a221oi_1 _15215_ (.B2(_06825_),
    .C1(net468),
    .B1(_06824_),
    .A1(_05905_),
    .Y(_06826_),
    .A2(_00070_));
 sg13g2_mux4_1 _15216_ (.S0(_06677_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][4] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][4] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][4] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][4] ),
    .S1(_06678_),
    .X(_06827_));
 sg13g2_mux4_1 _15217_ (.S0(_06673_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][4] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][4] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][4] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][4] ),
    .S1(_06674_),
    .X(_06828_));
 sg13g2_mux4_1 _15218_ (.S0(_06536_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[8][4] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][4] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][4] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[11][4] ),
    .S1(_06538_),
    .X(_06829_));
 sg13g2_mux4_1 _15219_ (.S0(net463),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[12][4] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][4] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][4] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[15][4] ),
    .S1(net462),
    .X(_06830_));
 sg13g2_mux4_1 _15220_ (.S0(_06543_),
    .A0(_06827_),
    .A1(_06828_),
    .A2(_06829_),
    .A3(_06830_),
    .S1(_06544_),
    .X(_06831_));
 sg13g2_nand2b_1 _15221_ (.Y(_06832_),
    .B(_06533_),
    .A_N(_06831_));
 sg13g2_o21ai_1 _15222_ (.B1(_06832_),
    .Y(_06833_),
    .A1(net466),
    .A2(_06826_));
 sg13g2_inv_1 _15223_ (.Y(_06834_),
    .A(_06833_));
 sg13g2_a22oi_1 _15224_ (.Y(_06835_),
    .B1(_06566_),
    .B2(_06834_),
    .A2(\soc_I.qqspi_I.rdata[4] ),
    .A1(net473));
 sg13g2_o21ai_1 _15225_ (.B1(net429),
    .Y(_06836_),
    .A1(_01641_),
    .A2(net44));
 sg13g2_a21oi_1 _15226_ (.A1(net38),
    .A2(_06835_),
    .Y(_00285_),
    .B1(_06836_));
 sg13g2_inv_1 _15227_ (.Y(_06837_),
    .A(_00073_));
 sg13g2_a221oi_1 _15228_ (.B2(\soc_I.cycle_cnt[5] ),
    .C1(net436),
    .B1(_06646_),
    .A1(_06645_),
    .Y(_06838_),
    .A2(_06837_));
 sg13g2_nand2_1 _15229_ (.Y(_06839_),
    .A(\soc_I.spi0_I.rx_data[5] ),
    .B(_06670_));
 sg13g2_a221oi_1 _15230_ (.B2(_06839_),
    .C1(_06644_),
    .B1(_06838_),
    .A1(_06604_),
    .Y(_06840_),
    .A2(_00072_));
 sg13g2_mux4_1 _15231_ (.S0(net463),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][5] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][5] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][5] ),
    .S1(net462),
    .X(_06841_));
 sg13g2_mux4_1 _15232_ (.S0(net465),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][5] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][5] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][5] ),
    .S1(net464),
    .X(_06842_));
 sg13g2_mux4_1 _15233_ (.S0(net541),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[8][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][5] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][5] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[11][5] ),
    .S1(net540),
    .X(_06843_));
 sg13g2_mux4_1 _15234_ (.S0(net463),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[12][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][5] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][5] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[15][5] ),
    .S1(net462),
    .X(_06844_));
 sg13g2_mux4_1 _15235_ (.S0(_06543_),
    .A0(_06841_),
    .A1(_06842_),
    .A2(_06843_),
    .A3(_06844_),
    .S1(_06544_),
    .X(_06845_));
 sg13g2_nand2b_1 _15236_ (.Y(_06846_),
    .B(_06533_),
    .A_N(_06845_));
 sg13g2_o21ai_1 _15237_ (.B1(_06846_),
    .Y(_06847_),
    .A1(_06666_),
    .A2(_06840_));
 sg13g2_inv_1 _15238_ (.Y(_06848_),
    .A(_06847_));
 sg13g2_a22oi_1 _15239_ (.Y(_06849_),
    .B1(_06566_),
    .B2(_06848_),
    .A2(\soc_I.qqspi_I.rdata[5] ),
    .A1(net473));
 sg13g2_o21ai_1 _15240_ (.B1(net429),
    .Y(_06850_),
    .A1(_01650_),
    .A2(net44));
 sg13g2_a21oi_1 _15241_ (.A1(net38),
    .A2(_06849_),
    .Y(_00286_),
    .B1(_06850_));
 sg13g2_mux4_1 _15242_ (.S0(net465),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][6] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][6] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][6] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][6] ),
    .S1(net464),
    .X(_06851_));
 sg13g2_mux4_1 _15243_ (.S0(net465),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][6] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][6] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][6] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][6] ),
    .S1(net464),
    .X(_06852_));
 sg13g2_mux4_1 _15244_ (.S0(net465),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[8][6] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][6] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][6] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[11][6] ),
    .S1(net464),
    .X(_06853_));
 sg13g2_mux4_1 _15245_ (.S0(net465),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[12][6] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][6] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][6] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[15][6] ),
    .S1(net464),
    .X(_06854_));
 sg13g2_mux4_1 _15246_ (.S0(_06543_),
    .A0(_06851_),
    .A1(_06852_),
    .A2(_06853_),
    .A3(_06854_),
    .S1(_06544_),
    .X(_06855_));
 sg13g2_inv_1 _15247_ (.Y(_06856_),
    .A(_06855_));
 sg13g2_inv_1 _15248_ (.Y(_06857_),
    .A(_00075_));
 sg13g2_a221oi_1 _15249_ (.B2(_05813_),
    .C1(net436),
    .B1(_06646_),
    .A1(_06645_),
    .Y(_06858_),
    .A2(_06857_));
 sg13g2_nand2_1 _15250_ (.Y(_06859_),
    .A(\soc_I.spi0_I.rx_data[6] ),
    .B(_06670_));
 sg13g2_a221oi_1 _15251_ (.B2(_06859_),
    .C1(_06644_),
    .B1(_06858_),
    .A1(_05905_),
    .Y(_06860_),
    .A2(_00074_));
 sg13g2_nor2_1 _15252_ (.A(_06666_),
    .B(_06860_),
    .Y(_06861_));
 sg13g2_a21oi_1 _15253_ (.A1(_06534_),
    .A2(_06856_),
    .Y(_06862_),
    .B1(_06861_));
 sg13g2_a22oi_1 _15254_ (.Y(_06863_),
    .B1(_06566_),
    .B2(_06862_),
    .A2(\soc_I.qqspi_I.rdata[6] ),
    .A1(net473));
 sg13g2_o21ai_1 _15255_ (.B1(net518),
    .Y(_06864_),
    .A1(net629),
    .A2(net44));
 sg13g2_a21oi_1 _15256_ (.A1(net38),
    .A2(_06863_),
    .Y(_00287_),
    .B1(_06864_));
 sg13g2_nor2_1 _15257_ (.A(_01702_),
    .B(net47),
    .Y(_06865_));
 sg13g2_a22oi_1 _15258_ (.Y(_06866_),
    .B1(_04097_),
    .B2(net76),
    .A2(_03671_),
    .A1(_03655_));
 sg13g2_inv_1 _15259_ (.Y(_06867_),
    .A(_00077_));
 sg13g2_a221oi_1 _15260_ (.B2(\soc_I.cycle_cnt[7] ),
    .C1(_04102_),
    .B1(_06552_),
    .A1(net618),
    .Y(_06868_),
    .A2(_06867_));
 sg13g2_nand2_1 _15261_ (.Y(_06869_),
    .A(\soc_I.spi0_I.rx_data[7] ),
    .B(_06670_));
 sg13g2_a221oi_1 _15262_ (.B2(_06869_),
    .C1(_04103_),
    .B1(_06868_),
    .A1(_04102_),
    .Y(_06870_),
    .A2(_00076_));
 sg13g2_mux4_1 _15263_ (.S0(_06535_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][7] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][7] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][7] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][7] ),
    .S1(_06537_),
    .X(_06871_));
 sg13g2_mux4_1 _15264_ (.S0(_06535_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][7] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][7] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][7] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][7] ),
    .S1(_06537_),
    .X(_06872_));
 sg13g2_mux4_1 _15265_ (.S0(_06535_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[8][7] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][7] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][7] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[11][7] ),
    .S1(_06537_),
    .X(_06873_));
 sg13g2_mux4_1 _15266_ (.S0(_06535_),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[12][7] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][7] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][7] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[15][7] ),
    .S1(_06537_),
    .X(_06874_));
 sg13g2_mux4_1 _15267_ (.S0(_06543_),
    .A0(_06871_),
    .A1(_06872_),
    .A2(_06873_),
    .A3(_06874_),
    .S1(_06544_),
    .X(_06875_));
 sg13g2_nand2b_1 _15268_ (.Y(_06876_),
    .B(_06532_),
    .A_N(_06875_));
 sg13g2_o21ai_1 _15269_ (.B1(_06876_),
    .Y(_06877_),
    .A1(_04105_),
    .A2(_06870_));
 sg13g2_or4_1 _15270_ (.A(_04226_),
    .B(net615),
    .C(_04219_),
    .D(_06877_),
    .X(_06878_));
 sg13g2_nand2_1 _15271_ (.Y(_06879_),
    .A(_04325_),
    .B(\soc_I.qqspi_I.rdata[7] ));
 sg13g2_o21ai_1 _15272_ (.B1(_06879_),
    .Y(_06880_),
    .A1(_06866_),
    .A2(_06878_));
 sg13g2_nor2_1 _15273_ (.A(_06568_),
    .B(_06880_),
    .Y(_06881_));
 sg13g2_nor3_1 _15274_ (.A(net392),
    .B(_06865_),
    .C(_06881_),
    .Y(_00288_));
 sg13g2_a22oi_1 _15275_ (.Y(_06882_),
    .B1(\soc_I.cycle_cnt[8] ),
    .B2(net390),
    .A2(_05659_),
    .A1(_06548_));
 sg13g2_nor2_1 _15276_ (.A(net507),
    .B(_06882_),
    .Y(_06883_));
 sg13g2_a21oi_1 _15277_ (.A1(net470),
    .A2(net609),
    .Y(_06884_),
    .B1(_06883_));
 sg13g2_o21ai_1 _15278_ (.B1(net469),
    .Y(_06885_),
    .A1(net537),
    .A2(_06884_));
 sg13g2_nor2_1 _15279_ (.A(_04226_),
    .B(net351),
    .Y(_06886_));
 sg13g2_a22oi_1 _15280_ (.Y(_06887_),
    .B1(_06885_),
    .B2(_06886_),
    .A2(_06628_),
    .A1(_04226_));
 sg13g2_nor2_1 _15281_ (.A(net542),
    .B(_06887_),
    .Y(_06888_));
 sg13g2_a22oi_1 _15282_ (.Y(_06889_),
    .B1(_04271_),
    .B2(_06888_),
    .A2(\soc_I.qqspi_I.rdata[8] ),
    .A1(net542));
 sg13g2_o21ai_1 _15283_ (.B1(net518),
    .Y(_06890_),
    .A1(_01667_),
    .A2(_06570_));
 sg13g2_a21oi_1 _15284_ (.A1(net38),
    .A2(_06889_),
    .Y(_00289_),
    .B1(_06890_));
 sg13g2_nor2b_1 _15285_ (.A(_05480_),
    .B_N(_05903_),
    .Y(_06891_));
 sg13g2_a221oi_1 _15286_ (.B2(net350),
    .C1(_06581_),
    .B1(_05811_),
    .A1(net472),
    .Y(_06892_),
    .A2(_05657_));
 sg13g2_nor3_1 _15287_ (.A(_06560_),
    .B(_06891_),
    .C(_06892_),
    .Y(_06893_));
 sg13g2_nor2_1 _15288_ (.A(net539),
    .B(_06893_),
    .Y(_06894_));
 sg13g2_nor2_1 _15289_ (.A(net330),
    .B(_06894_),
    .Y(_06895_));
 sg13g2_a22oi_1 _15290_ (.Y(_06896_),
    .B1(net67),
    .B2(_06895_),
    .A2(\soc_I.qqspi_I.rdata[9] ),
    .A1(net471));
 sg13g2_o21ai_1 _15291_ (.B1(_04305_),
    .Y(_06897_),
    .A1(_02273_),
    .A2(_06570_));
 sg13g2_a21oi_1 _15292_ (.A1(_06693_),
    .A2(_06896_),
    .Y(_00290_),
    .B1(_06897_));
 sg13g2_buf_1 _15293_ (.A(_06570_),
    .X(_06898_));
 sg13g2_nand2_1 _15294_ (.Y(_06899_),
    .A(_01712_),
    .B(net36));
 sg13g2_nand2_1 _15295_ (.Y(_06900_),
    .A(\soc_I.PC[0] ),
    .B(net37));
 sg13g2_a21oi_1 _15296_ (.A1(_06899_),
    .A2(_06900_),
    .Y(_00291_),
    .B1(net389));
 sg13g2_nand2_1 _15297_ (.Y(_06901_),
    .A(_01959_),
    .B(net36));
 sg13g2_nand2_1 _15298_ (.Y(_06902_),
    .A(\soc_I.PC[10] ),
    .B(net37));
 sg13g2_a21oi_1 _15299_ (.A1(_06901_),
    .A2(_06902_),
    .Y(_00292_),
    .B1(net389));
 sg13g2_nand2_1 _15300_ (.Y(_06903_),
    .A(_01979_),
    .B(net36));
 sg13g2_nand2_1 _15301_ (.Y(_06904_),
    .A(\soc_I.PC[11] ),
    .B(net37));
 sg13g2_a21oi_1 _15302_ (.A1(_06903_),
    .A2(_06904_),
    .Y(_00293_),
    .B1(net389));
 sg13g2_nand2_1 _15303_ (.Y(_06905_),
    .A(_01864_),
    .B(net36));
 sg13g2_nand2_1 _15304_ (.Y(_06906_),
    .A(\soc_I.PC[12] ),
    .B(net37));
 sg13g2_a21oi_1 _15305_ (.A1(_06905_),
    .A2(_06906_),
    .Y(_00294_),
    .B1(net389));
 sg13g2_nand2_1 _15306_ (.Y(_06907_),
    .A(_01903_),
    .B(net36));
 sg13g2_nand2_1 _15307_ (.Y(_06908_),
    .A(\soc_I.PC[13] ),
    .B(net37));
 sg13g2_a21oi_1 _15308_ (.A1(_06907_),
    .A2(_06908_),
    .Y(_00295_),
    .B1(net389));
 sg13g2_nand2_1 _15309_ (.Y(_06909_),
    .A(_01883_),
    .B(_06898_));
 sg13g2_nand2_1 _15310_ (.Y(_06910_),
    .A(\soc_I.PC[14] ),
    .B(net37));
 sg13g2_a21oi_1 _15311_ (.A1(_06909_),
    .A2(_06910_),
    .Y(_00296_),
    .B1(net389));
 sg13g2_nand2_1 _15312_ (.Y(_06911_),
    .A(_01826_),
    .B(_06898_));
 sg13g2_nand2_1 _15313_ (.Y(_06912_),
    .A(\soc_I.PC[15] ),
    .B(net37));
 sg13g2_a21oi_1 _15314_ (.A1(_06911_),
    .A2(_06912_),
    .Y(_00297_),
    .B1(net389));
 sg13g2_nand2_1 _15315_ (.Y(_06913_),
    .A(_02150_),
    .B(net36));
 sg13g2_nand2_1 _15316_ (.Y(_06914_),
    .A(\soc_I.PC[16] ),
    .B(net37));
 sg13g2_a21oi_1 _15317_ (.A1(_06913_),
    .A2(_06914_),
    .Y(_00298_),
    .B1(net389));
 sg13g2_nand2_1 _15318_ (.Y(_06915_),
    .A(_02134_),
    .B(net36));
 sg13g2_buf_8 _15319_ (.A(net46),
    .X(_06916_));
 sg13g2_nand2_1 _15320_ (.Y(_06917_),
    .A(\soc_I.PC[17] ),
    .B(net35));
 sg13g2_buf_1 _15321_ (.A(_04267_),
    .X(_06918_));
 sg13g2_a21oi_1 _15322_ (.A1(_06915_),
    .A2(_06917_),
    .Y(_00299_),
    .B1(net387));
 sg13g2_nand2_1 _15323_ (.Y(_06919_),
    .A(_02117_),
    .B(net36));
 sg13g2_nand2_1 _15324_ (.Y(_06920_),
    .A(\soc_I.PC[18] ),
    .B(net35));
 sg13g2_a21oi_1 _15325_ (.A1(_06919_),
    .A2(_06920_),
    .Y(_00300_),
    .B1(net387));
 sg13g2_buf_1 _15326_ (.A(_06570_),
    .X(_06921_));
 sg13g2_nand2_1 _15327_ (.Y(_06922_),
    .A(_02099_),
    .B(_06921_));
 sg13g2_nand2_1 _15328_ (.Y(_06923_),
    .A(\soc_I.PC[19] ),
    .B(_06916_));
 sg13g2_a21oi_1 _15329_ (.A1(_06922_),
    .A2(_06923_),
    .Y(_00301_),
    .B1(_06918_));
 sg13g2_nand2_1 _15330_ (.Y(_06924_),
    .A(_01573_),
    .B(net34));
 sg13g2_nand2_1 _15331_ (.Y(_06925_),
    .A(\soc_I.PC[1] ),
    .B(net35));
 sg13g2_a21oi_1 _15332_ (.A1(_06924_),
    .A2(_06925_),
    .Y(_00302_),
    .B1(net387));
 sg13g2_nand2_1 _15333_ (.Y(_06926_),
    .A(_02049_),
    .B(_06921_));
 sg13g2_nand2_1 _15334_ (.Y(_06927_),
    .A(\soc_I.PC[20] ),
    .B(net35));
 sg13g2_a21oi_1 _15335_ (.A1(_06926_),
    .A2(_06927_),
    .Y(_00303_),
    .B1(net387));
 sg13g2_nand2_1 _15336_ (.Y(_06928_),
    .A(_02039_),
    .B(net34));
 sg13g2_nand2_1 _15337_ (.Y(_06929_),
    .A(\soc_I.PC[21] ),
    .B(net35));
 sg13g2_a21oi_1 _15338_ (.A1(_06928_),
    .A2(_06929_),
    .Y(_00304_),
    .B1(net387));
 sg13g2_nand2_1 _15339_ (.Y(_06930_),
    .A(_02064_),
    .B(net34));
 sg13g2_nand2_1 _15340_ (.Y(_06931_),
    .A(\soc_I.PC[22] ),
    .B(net35));
 sg13g2_a21oi_1 _15341_ (.A1(_06930_),
    .A2(_06931_),
    .Y(_00305_),
    .B1(net387));
 sg13g2_nand2_1 _15342_ (.Y(_06932_),
    .A(_02074_),
    .B(net34));
 sg13g2_nand2_1 _15343_ (.Y(_06933_),
    .A(\soc_I.PC[23] ),
    .B(_06916_));
 sg13g2_a21oi_1 _15344_ (.A1(_06932_),
    .A2(_06933_),
    .Y(_00306_),
    .B1(_06918_));
 sg13g2_nand2_1 _15345_ (.Y(_06934_),
    .A(_02489_),
    .B(net34));
 sg13g2_nand2_1 _15346_ (.Y(_06935_),
    .A(\soc_I.PC[24] ),
    .B(net35));
 sg13g2_a21oi_1 _15347_ (.A1(_06934_),
    .A2(_06935_),
    .Y(_00307_),
    .B1(net387));
 sg13g2_nand2_1 _15348_ (.Y(_06936_),
    .A(_02479_),
    .B(net34));
 sg13g2_nand2_1 _15349_ (.Y(_06937_),
    .A(\soc_I.PC[25] ),
    .B(net35));
 sg13g2_a21oi_1 _15350_ (.A1(_06936_),
    .A2(_06937_),
    .Y(_00308_),
    .B1(net387));
 sg13g2_nand2_1 _15351_ (.Y(_06938_),
    .A(_02551_),
    .B(net34));
 sg13g2_buf_8 _15352_ (.A(net46),
    .X(_06939_));
 sg13g2_nand2_1 _15353_ (.Y(_06940_),
    .A(\soc_I.PC[26] ),
    .B(net33));
 sg13g2_buf_1 _15354_ (.A(_04267_),
    .X(_06941_));
 sg13g2_a21oi_1 _15355_ (.A1(_06938_),
    .A2(_06940_),
    .Y(_00309_),
    .B1(net386));
 sg13g2_nand2_1 _15356_ (.Y(_06942_),
    .A(_02544_),
    .B(net34));
 sg13g2_nand2_1 _15357_ (.Y(_06943_),
    .A(\soc_I.PC[27] ),
    .B(net33));
 sg13g2_a21oi_1 _15358_ (.A1(_06942_),
    .A2(_06943_),
    .Y(_00310_),
    .B1(net386));
 sg13g2_buf_8 _15359_ (.A(_06570_),
    .X(_06944_));
 sg13g2_nand2_1 _15360_ (.Y(_06945_),
    .A(_02514_),
    .B(net32));
 sg13g2_nand2_1 _15361_ (.Y(_06946_),
    .A(\soc_I.PC[28] ),
    .B(net33));
 sg13g2_a21oi_1 _15362_ (.A1(_06945_),
    .A2(_06946_),
    .Y(_00311_),
    .B1(net386));
 sg13g2_nand2_1 _15363_ (.Y(_06947_),
    .A(_02527_),
    .B(net32));
 sg13g2_nand2_1 _15364_ (.Y(_06948_),
    .A(\soc_I.PC[29] ),
    .B(_06939_));
 sg13g2_a21oi_1 _15365_ (.A1(_06947_),
    .A2(_06948_),
    .Y(_00312_),
    .B1(net386));
 sg13g2_nand2_1 _15366_ (.Y(_06949_),
    .A(_02268_),
    .B(net32));
 sg13g2_nand2_1 _15367_ (.Y(_06950_),
    .A(\soc_I.PC[2] ),
    .B(net33));
 sg13g2_a21oi_1 _15368_ (.A1(_06949_),
    .A2(_06950_),
    .Y(_00313_),
    .B1(net386));
 sg13g2_nand2_1 _15369_ (.Y(_06951_),
    .A(_02665_),
    .B(net32));
 sg13g2_nand2_1 _15370_ (.Y(_06952_),
    .A(\soc_I.PC[30] ),
    .B(net33));
 sg13g2_a21oi_1 _15371_ (.A1(_06951_),
    .A2(_06952_),
    .Y(_00314_),
    .B1(net386));
 sg13g2_nand2_1 _15372_ (.Y(_06953_),
    .A(_02658_),
    .B(net32));
 sg13g2_nand2_1 _15373_ (.Y(_06954_),
    .A(\soc_I.PC[31] ),
    .B(net33));
 sg13g2_a21oi_1 _15374_ (.A1(_06953_),
    .A2(_06954_),
    .Y(_00315_),
    .B1(net386));
 sg13g2_nand2_1 _15375_ (.Y(_06955_),
    .A(_02282_),
    .B(_06944_));
 sg13g2_nand2_1 _15376_ (.Y(_06956_),
    .A(\soc_I.PC[3] ),
    .B(net33));
 sg13g2_a21oi_1 _15377_ (.A1(_06955_),
    .A2(_06956_),
    .Y(_00316_),
    .B1(_06941_));
 sg13g2_nand2_1 _15378_ (.Y(_06957_),
    .A(_02397_),
    .B(net32));
 sg13g2_nand2_1 _15379_ (.Y(_06958_),
    .A(\soc_I.PC[4] ),
    .B(net33));
 sg13g2_a21oi_1 _15380_ (.A1(_06957_),
    .A2(_06958_),
    .Y(_00317_),
    .B1(net386));
 sg13g2_nand2_1 _15381_ (.Y(_06959_),
    .A(_02425_),
    .B(net32));
 sg13g2_nand2_1 _15382_ (.Y(_06960_),
    .A(\soc_I.PC[5] ),
    .B(_06939_));
 sg13g2_a21oi_1 _15383_ (.A1(_06959_),
    .A2(_06960_),
    .Y(_00318_),
    .B1(_06941_));
 sg13g2_nand2_1 _15384_ (.Y(_06961_),
    .A(_02337_),
    .B(net32));
 sg13g2_nand2_1 _15385_ (.Y(_06962_),
    .A(\soc_I.PC[6] ),
    .B(net46));
 sg13g2_buf_1 _15386_ (.A(_04267_),
    .X(_06963_));
 sg13g2_a21oi_1 _15387_ (.A1(_06961_),
    .A2(_06962_),
    .Y(_00319_),
    .B1(net385));
 sg13g2_nand2_1 _15388_ (.Y(_06964_),
    .A(_02330_),
    .B(_06944_));
 sg13g2_nand2_1 _15389_ (.Y(_06965_),
    .A(\soc_I.PC[7] ),
    .B(net46));
 sg13g2_a21oi_1 _15390_ (.A1(_06964_),
    .A2(_06965_),
    .Y(_00320_),
    .B1(net385));
 sg13g2_nand2_1 _15391_ (.Y(_06966_),
    .A(_01929_),
    .B(net47));
 sg13g2_nand2_1 _15392_ (.Y(_06967_),
    .A(\soc_I.PC[8] ),
    .B(net46));
 sg13g2_a21oi_1 _15393_ (.A1(_06966_),
    .A2(_06967_),
    .Y(_00321_),
    .B1(net385));
 sg13g2_nand2_1 _15394_ (.Y(_06968_),
    .A(_01943_),
    .B(net47));
 sg13g2_nand2_1 _15395_ (.Y(_06969_),
    .A(\soc_I.PC[9] ),
    .B(net46));
 sg13g2_a21oi_1 _15396_ (.A1(_06968_),
    .A2(_06969_),
    .Y(_00322_),
    .B1(net385));
 sg13g2_inv_1 _15397_ (.Y(_06970_),
    .A(_01712_));
 sg13g2_inv_1 _15398_ (.Y(_06971_),
    .A(_01594_));
 sg13g2_nor3_1 _15399_ (.A(_04134_),
    .B(_04152_),
    .C(_04185_),
    .Y(_06972_));
 sg13g2_nand3b_1 _15400_ (.B(_04118_),
    .C(_06972_),
    .Y(_06973_),
    .A_N(_03529_));
 sg13g2_a21o_1 _15401_ (.A2(_06973_),
    .A1(_06971_),
    .B1(_01577_),
    .X(_06974_));
 sg13g2_or3_1 _15402_ (.A(_04269_),
    .B(_03580_),
    .C(_06974_),
    .X(_06975_));
 sg13g2_a21oi_1 _15403_ (.A1(_04238_),
    .A2(_04256_),
    .Y(_06976_),
    .B1(_06975_));
 sg13g2_buf_2 _15404_ (.A(_06976_),
    .X(_06977_));
 sg13g2_a21o_1 _15405_ (.A2(_04261_),
    .A1(net447),
    .B1(_06974_),
    .X(_06978_));
 sg13g2_o21ai_1 _15406_ (.B1(_06978_),
    .Y(_06979_),
    .A1(_04221_),
    .A2(_06975_));
 sg13g2_buf_2 _15407_ (.A(_06979_),
    .X(_06980_));
 sg13g2_nor2_1 _15408_ (.A(_06977_),
    .B(_06980_),
    .Y(_06981_));
 sg13g2_buf_4 _15409_ (.X(_06982_),
    .A(_06981_));
 sg13g2_buf_8 _15410_ (.A(_06982_),
    .X(_06983_));
 sg13g2_mux2_1 _15411_ (.A0(_06970_),
    .A1(_04549_),
    .S(_06983_),
    .X(_06984_));
 sg13g2_nor2_1 _15412_ (.A(net391),
    .B(_06984_),
    .Y(_00323_));
 sg13g2_inv_1 _15413_ (.Y(_06985_),
    .A(_01959_));
 sg13g2_buf_8 _15414_ (.A(_06982_),
    .X(_06986_));
 sg13g2_mux2_1 _15415_ (.A0(_06985_),
    .A1(net117),
    .S(net30),
    .X(_06987_));
 sg13g2_nor2_1 _15416_ (.A(net391),
    .B(_06987_),
    .Y(_00324_));
 sg13g2_buf_8 _15417_ (.A(_06982_),
    .X(_06988_));
 sg13g2_mux2_1 _15418_ (.A0(_01979_),
    .A1(net129),
    .S(net29),
    .X(_06989_));
 sg13g2_and2_1 _15419_ (.A(net435),
    .B(_06989_),
    .X(_00325_));
 sg13g2_mux2_1 _15420_ (.A0(_01865_),
    .A1(net131),
    .S(net30),
    .X(_06990_));
 sg13g2_nor2_1 _15421_ (.A(net391),
    .B(_06990_),
    .Y(_00326_));
 sg13g2_mux2_1 _15422_ (.A0(_01903_),
    .A1(net99),
    .S(net29),
    .X(_06991_));
 sg13g2_and2_1 _15423_ (.A(net435),
    .B(_06991_),
    .X(_00327_));
 sg13g2_mux2_1 _15424_ (.A0(_03995_),
    .A1(net98),
    .S(net30),
    .X(_06992_));
 sg13g2_nor2_1 _15425_ (.A(net391),
    .B(_06992_),
    .Y(_00328_));
 sg13g2_or2_1 _15426_ (.X(_06993_),
    .B(_06988_),
    .A(_01826_));
 sg13g2_nand2_1 _15427_ (.Y(_06994_),
    .A(_03933_),
    .B(net31));
 sg13g2_and3_1 _15428_ (.X(_00329_),
    .A(net433),
    .B(_06993_),
    .C(_06994_));
 sg13g2_inv_1 _15429_ (.Y(_06995_),
    .A(_02150_));
 sg13g2_mux2_1 _15430_ (.A0(_06995_),
    .A1(net85),
    .S(_06986_),
    .X(_06996_));
 sg13g2_nor2_1 _15431_ (.A(net391),
    .B(_06996_),
    .Y(_00330_));
 sg13g2_mux2_1 _15432_ (.A0(_02753_),
    .A1(net121),
    .S(net30),
    .X(_06997_));
 sg13g2_nor2_1 _15433_ (.A(net391),
    .B(_06997_),
    .Y(_00331_));
 sg13g2_mux2_1 _15434_ (.A0(_02754_),
    .A1(net97),
    .S(net30),
    .X(_06998_));
 sg13g2_nor2_1 _15435_ (.A(net391),
    .B(_06998_),
    .Y(_00332_));
 sg13g2_inv_1 _15436_ (.Y(_06999_),
    .A(_02099_));
 sg13g2_mux2_1 _15437_ (.A0(_06999_),
    .A1(net120),
    .S(net30),
    .X(_07000_));
 sg13g2_nor2_1 _15438_ (.A(net391),
    .B(_07000_),
    .Y(_00333_));
 sg13g2_inv_1 _15439_ (.Y(_07001_),
    .A(_01573_));
 sg13g2_mux2_1 _15440_ (.A0(_07001_),
    .A1(net124),
    .S(_06986_),
    .X(_07002_));
 sg13g2_nor2_1 _15441_ (.A(_06522_),
    .B(_07002_),
    .Y(_00334_));
 sg13g2_nor2_1 _15442_ (.A(_02049_),
    .B(_06983_),
    .Y(_07003_));
 sg13g2_nor3_1 _15443_ (.A(net96),
    .B(_06977_),
    .C(_06980_),
    .Y(_07004_));
 sg13g2_o21ai_1 _15444_ (.B1(net437),
    .Y(_00335_),
    .A1(_07003_),
    .A2(_07004_));
 sg13g2_nor2_1 _15445_ (.A(_02039_),
    .B(net31),
    .Y(_07005_));
 sg13g2_and2_1 _15446_ (.A(_04609_),
    .B(net31),
    .X(_07006_));
 sg13g2_nor3_1 _15447_ (.A(net392),
    .B(_07005_),
    .C(_07006_),
    .Y(_00336_));
 sg13g2_o21ai_1 _15448_ (.B1(_02064_),
    .Y(_07007_),
    .A1(_06977_),
    .A2(_06980_));
 sg13g2_nand2b_1 _15449_ (.Y(_07008_),
    .B(net31),
    .A_N(_04207_));
 sg13g2_a21oi_1 _15450_ (.A1(_07007_),
    .A2(_07008_),
    .Y(_00337_),
    .B1(_06963_));
 sg13g2_buf_1 _15451_ (.A(net438),
    .X(_07009_));
 sg13g2_inv_1 _15452_ (.Y(_07010_),
    .A(_02074_));
 sg13g2_mux2_1 _15453_ (.A0(_07010_),
    .A1(_03714_),
    .S(net30),
    .X(_07011_));
 sg13g2_nor2_1 _15454_ (.A(net384),
    .B(_07011_),
    .Y(_00338_));
 sg13g2_nor2_1 _15455_ (.A(_02489_),
    .B(net31),
    .Y(_07012_));
 sg13g2_nor3_1 _15456_ (.A(_04203_),
    .B(_06977_),
    .C(_06980_),
    .Y(_07013_));
 sg13g2_nor3_1 _15457_ (.A(_06509_),
    .B(_07012_),
    .C(_07013_),
    .Y(_00339_));
 sg13g2_nor2_1 _15458_ (.A(_02479_),
    .B(net31),
    .Y(_07014_));
 sg13g2_nor3_1 _15459_ (.A(_04619_),
    .B(_06977_),
    .C(_06980_),
    .Y(_07015_));
 sg13g2_nor3_1 _15460_ (.A(_06509_),
    .B(_07014_),
    .C(_07015_),
    .Y(_00340_));
 sg13g2_inv_1 _15461_ (.Y(_07016_),
    .A(_02551_));
 sg13g2_mux2_1 _15462_ (.A0(_07016_),
    .A1(_04626_),
    .S(net30),
    .X(_07017_));
 sg13g2_nor2_1 _15463_ (.A(net384),
    .B(_07017_),
    .Y(_00341_));
 sg13g2_inv_1 _15464_ (.Y(_07018_),
    .A(_02544_));
 sg13g2_mux2_1 _15465_ (.A0(_07018_),
    .A1(_04632_),
    .S(net29),
    .X(_07019_));
 sg13g2_nor2_1 _15466_ (.A(net384),
    .B(_07019_),
    .Y(_00342_));
 sg13g2_mux2_1 _15467_ (.A0(_03783_),
    .A1(_04215_),
    .S(net29),
    .X(_07020_));
 sg13g2_nor2_1 _15468_ (.A(net384),
    .B(_07020_),
    .Y(_00343_));
 sg13g2_mux2_1 _15469_ (.A0(_04328_),
    .A1(_04330_),
    .S(net31),
    .X(_07021_));
 sg13g2_nand2_1 _15470_ (.Y(_00344_),
    .A(net437),
    .B(_07021_));
 sg13g2_mux2_1 _15471_ (.A0(_02268_),
    .A1(_03851_),
    .S(_06982_),
    .X(_07022_));
 sg13g2_and2_1 _15472_ (.A(net435),
    .B(_07022_),
    .X(_00345_));
 sg13g2_mux2_1 _15473_ (.A0(_04320_),
    .A1(_03650_),
    .S(_06988_),
    .X(_07023_));
 sg13g2_nor2_1 _15474_ (.A(_07009_),
    .B(_07023_),
    .Y(_00346_));
 sg13g2_buf_1 _15475_ (.A(_05918_),
    .X(_07024_));
 sg13g2_nor2_1 _15476_ (.A(_02658_),
    .B(net31),
    .Y(_07025_));
 sg13g2_nor3_1 _15477_ (.A(_04332_),
    .B(_06977_),
    .C(_06980_),
    .Y(_07026_));
 sg13g2_nor3_1 _15478_ (.A(net383),
    .B(_07025_),
    .C(_07026_),
    .Y(_00347_));
 sg13g2_inv_1 _15479_ (.Y(_07027_),
    .A(_02282_));
 sg13g2_mux2_1 _15480_ (.A0(_07027_),
    .A1(_03832_),
    .S(net29),
    .X(_07028_));
 sg13g2_nor2_1 _15481_ (.A(net384),
    .B(_07028_),
    .Y(_00348_));
 sg13g2_inv_1 _15482_ (.Y(_07029_),
    .A(_02397_));
 sg13g2_mux2_1 _15483_ (.A0(_07029_),
    .A1(_03804_),
    .S(net29),
    .X(_07030_));
 sg13g2_nor2_1 _15484_ (.A(net384),
    .B(_07030_),
    .Y(_00349_));
 sg13g2_mux2_1 _15485_ (.A0(_02426_),
    .A1(net123),
    .S(net29),
    .X(_07031_));
 sg13g2_nor2_1 _15486_ (.A(net384),
    .B(_07031_),
    .Y(_00350_));
 sg13g2_buf_1 _15487_ (.A(net515),
    .X(_07032_));
 sg13g2_mux2_1 _15488_ (.A0(_02337_),
    .A1(_03902_),
    .S(_06982_),
    .X(_07033_));
 sg13g2_and2_1 _15489_ (.A(net428),
    .B(_07033_),
    .X(_00351_));
 sg13g2_inv_1 _15490_ (.Y(_07034_),
    .A(_02330_));
 sg13g2_mux2_1 _15491_ (.A0(_07034_),
    .A1(net101),
    .S(net29),
    .X(_07035_));
 sg13g2_nor2_1 _15492_ (.A(net384),
    .B(_07035_),
    .Y(_00352_));
 sg13g2_mux2_1 _15493_ (.A0(_01929_),
    .A1(net100),
    .S(_06982_),
    .X(_07036_));
 sg13g2_and2_1 _15494_ (.A(net428),
    .B(_07036_),
    .X(_00353_));
 sg13g2_mux2_1 _15495_ (.A0(_01943_),
    .A1(net128),
    .S(_06982_),
    .X(_07037_));
 sg13g2_and2_1 _15496_ (.A(net428),
    .B(_07037_),
    .X(_00354_));
 sg13g2_nor2_1 _15497_ (.A(_01711_),
    .B(_02281_),
    .Y(_07038_));
 sg13g2_nand4_1 _15498_ (.B(_02853_),
    .C(_02891_),
    .A(_01686_),
    .Y(_07039_),
    .D(_07038_));
 sg13g2_buf_1 _15499_ (.A(_07039_),
    .X(_07040_));
 sg13g2_nor3_1 _15500_ (.A(_04390_),
    .B(_04386_),
    .C(_07040_),
    .Y(_07041_));
 sg13g2_a21oi_1 _15501_ (.A1(_04384_),
    .A2(_04386_),
    .Y(_07042_),
    .B1(_07041_));
 sg13g2_buf_1 _15502_ (.A(_07042_),
    .X(_07043_));
 sg13g2_buf_1 _15503_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[0] ),
    .X(_07044_));
 sg13g2_nand2b_1 _15504_ (.Y(_07045_),
    .B(_07044_),
    .A_N(net132));
 sg13g2_nand2_1 _15505_ (.Y(_07046_),
    .A(net589),
    .B(_00086_));
 sg13g2_o21ai_1 _15506_ (.B1(_07046_),
    .Y(_07047_),
    .A1(net590),
    .A2(_01718_));
 sg13g2_nand2_1 _15507_ (.Y(_07048_),
    .A(net132),
    .B(_07047_));
 sg13g2_a21oi_1 _15508_ (.A1(_07045_),
    .A2(_07048_),
    .Y(_00355_),
    .B1(net385));
 sg13g2_buf_1 _15509_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[1] ),
    .X(_07049_));
 sg13g2_nor2_1 _15510_ (.A(_07044_),
    .B(_07049_),
    .Y(_07050_));
 sg13g2_nand2_1 _15511_ (.Y(_07051_),
    .A(net589),
    .B(_07050_));
 sg13g2_o21ai_1 _15512_ (.B1(_07051_),
    .Y(_07052_),
    .A1(_04395_),
    .A2(_01686_));
 sg13g2_inv_1 _15513_ (.Y(_07053_),
    .A(_07044_));
 sg13g2_o21ai_1 _15514_ (.B1(_07043_),
    .Y(_07054_),
    .A1(_07053_),
    .A2(_04391_));
 sg13g2_a22oi_1 _15515_ (.Y(_07055_),
    .B1(_07054_),
    .B2(_07049_),
    .A2(_07052_),
    .A1(net132));
 sg13g2_nor2_1 _15516_ (.A(_07009_),
    .B(_07055_),
    .Y(_00356_));
 sg13g2_buf_1 _15517_ (.A(_06002_),
    .X(_07056_));
 sg13g2_nor3_1 _15518_ (.A(_07044_),
    .B(_07049_),
    .C(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[2] ),
    .Y(_07057_));
 sg13g2_mux2_1 _15519_ (.A0(_02281_),
    .A1(_07057_),
    .S(_04402_),
    .X(_07058_));
 sg13g2_o21ai_1 _15520_ (.B1(net132),
    .Y(_07059_),
    .A1(_04391_),
    .A2(_07050_));
 sg13g2_a22oi_1 _15521_ (.Y(_07060_),
    .B1(_07059_),
    .B2(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[2] ),
    .A2(_07058_),
    .A1(_07043_));
 sg13g2_nor2_1 _15522_ (.A(net382),
    .B(_07060_),
    .Y(_00357_));
 sg13g2_o21ai_1 _15523_ (.B1(net132),
    .Y(_07061_),
    .A1(_04391_),
    .A2(_07057_));
 sg13g2_nor2b_1 _15524_ (.A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[3] ),
    .B_N(_07057_),
    .Y(_07062_));
 sg13g2_nand2_1 _15525_ (.Y(_07063_),
    .A(_04402_),
    .B(_07062_));
 sg13g2_o21ai_1 _15526_ (.B1(_07063_),
    .Y(_07064_),
    .A1(net590),
    .A2(_02891_));
 sg13g2_a22oi_1 _15527_ (.Y(_07065_),
    .B1(_07064_),
    .B2(net132),
    .A2(_07061_),
    .A1(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[3] ));
 sg13g2_nor2_1 _15528_ (.A(net382),
    .B(_07065_),
    .Y(_00358_));
 sg13g2_nand3_1 _15529_ (.B(net589),
    .C(_07062_),
    .A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[4] ),
    .Y(_07066_));
 sg13g2_o21ai_1 _15530_ (.B1(_07066_),
    .Y(_07067_),
    .A1(_04403_),
    .A2(_03793_));
 sg13g2_o21ai_1 _15531_ (.B1(net132),
    .Y(_07068_),
    .A1(_04391_),
    .A2(_07062_));
 sg13g2_inv_1 _15532_ (.Y(_07069_),
    .A(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[4] ));
 sg13g2_a221oi_1 _15533_ (.B2(_07069_),
    .C1(net398),
    .B1(_07068_),
    .A1(net132),
    .Y(_00359_),
    .A2(_07067_));
 sg13g2_nor4_1 _15534_ (.A(_07049_),
    .B(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[3] ),
    .C(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[2] ),
    .D(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[4] ),
    .Y(_07070_));
 sg13g2_nand2_1 _15535_ (.Y(_07071_),
    .A(_07044_),
    .B(_07070_));
 sg13g2_nand2b_1 _15536_ (.Y(_07072_),
    .B(_07071_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_ready ));
 sg13g2_o21ai_1 _15537_ (.B1(_04384_),
    .Y(_07073_),
    .A1(_04386_),
    .A2(_07040_));
 sg13g2_o21ai_1 _15538_ (.B1(_07073_),
    .Y(_07074_),
    .A1(_04384_),
    .A2(_07072_));
 sg13g2_nor2_1 _15539_ (.A(net382),
    .B(_07074_),
    .Y(_00360_));
 sg13g2_inv_1 _15540_ (.Y(_07075_),
    .A(_07040_));
 sg13g2_nor3_1 _15541_ (.A(_04403_),
    .B(_04386_),
    .C(_07075_),
    .Y(_07076_));
 sg13g2_a21oi_1 _15542_ (.A1(_04400_),
    .A2(_07071_),
    .Y(_07077_),
    .B1(_07076_));
 sg13g2_nor2_1 _15543_ (.A(net382),
    .B(_07077_),
    .Y(_00393_));
 sg13g2_or4_1 _15544_ (.A(\soc_I.pwm_ready ),
    .B(net106),
    .C(_05907_),
    .D(_05913_),
    .X(_07078_));
 sg13g2_buf_4 _15545_ (.X(_07079_),
    .A(_07078_));
 sg13g2_mux2_1 _15546_ (.A0(net607),
    .A1(\soc_I.pwm_I.pcm[0] ),
    .S(_07079_),
    .X(_07080_));
 sg13g2_and2_1 _15547_ (.A(net428),
    .B(_07080_),
    .X(_00906_));
 sg13g2_buf_1 _15548_ (.A(\soc_I.pwm_I.pcm[1] ),
    .X(_07081_));
 sg13g2_mux2_1 _15549_ (.A0(net604),
    .A1(_07081_),
    .S(_07079_),
    .X(_07082_));
 sg13g2_and2_1 _15550_ (.A(net428),
    .B(_07082_),
    .X(_00907_));
 sg13g2_mux2_1 _15551_ (.A0(net619),
    .A1(\soc_I.pwm_I.pcm[2] ),
    .S(_07079_),
    .X(_07083_));
 sg13g2_and2_1 _15552_ (.A(net428),
    .B(_07083_),
    .X(_00908_));
 sg13g2_mux2_1 _15553_ (.A0(_05929_),
    .A1(\soc_I.pwm_I.pcm[3] ),
    .S(_07079_),
    .X(_07084_));
 sg13g2_and2_1 _15554_ (.A(net428),
    .B(_07084_),
    .X(_00909_));
 sg13g2_mux2_1 _15555_ (.A0(net606),
    .A1(\soc_I.pwm_I.pcm[4] ),
    .S(_07079_),
    .X(_07085_));
 sg13g2_and2_1 _15556_ (.A(net428),
    .B(_07085_),
    .X(_00910_));
 sg13g2_mux2_1 _15557_ (.A0(_05941_),
    .A1(\soc_I.pwm_I.pcm[5] ),
    .S(_07079_),
    .X(_07086_));
 sg13g2_and2_1 _15558_ (.A(_07032_),
    .B(_07086_),
    .X(_00911_));
 sg13g2_mux2_1 _15559_ (.A0(_05946_),
    .A1(\soc_I.pwm_I.pcm[6] ),
    .S(_07079_),
    .X(_07087_));
 sg13g2_and2_1 _15560_ (.A(_07032_),
    .B(_07087_),
    .X(_00912_));
 sg13g2_buf_1 _15561_ (.A(net515),
    .X(_07088_));
 sg13g2_buf_1 _15562_ (.A(\soc_I.pwm_I.pcm[7] ),
    .X(_07089_));
 sg13g2_mux2_1 _15563_ (.A0(net605),
    .A1(_07089_),
    .S(_07079_),
    .X(_07090_));
 sg13g2_and2_1 _15564_ (.A(net427),
    .B(_07090_),
    .X(_00913_));
 sg13g2_xnor2_1 _15565_ (.Y(_07091_),
    .A(\soc_I.pwm_I.pcm[0] ),
    .B(\soc_I.pwm_I.pwm_accumulator[0] ));
 sg13g2_nor2_1 _15566_ (.A(net382),
    .B(_07091_),
    .Y(_00914_));
 sg13g2_nand2_1 _15567_ (.Y(_07092_),
    .A(\soc_I.pwm_I.pcm[0] ),
    .B(\soc_I.pwm_I.pwm_accumulator[0] ));
 sg13g2_xnor2_1 _15568_ (.Y(_07093_),
    .A(_07081_),
    .B(\soc_I.pwm_I.pwm_accumulator[1] ));
 sg13g2_xnor2_1 _15569_ (.Y(_07094_),
    .A(_07092_),
    .B(_07093_));
 sg13g2_nor2_1 _15570_ (.A(net382),
    .B(_07094_),
    .Y(_00915_));
 sg13g2_nor2_1 _15571_ (.A(_07081_),
    .B(\soc_I.pwm_I.pwm_accumulator[1] ),
    .Y(_07095_));
 sg13g2_nand2_1 _15572_ (.Y(_07096_),
    .A(_07081_),
    .B(\soc_I.pwm_I.pwm_accumulator[1] ));
 sg13g2_o21ai_1 _15573_ (.B1(_07096_),
    .Y(_07097_),
    .A1(_07092_),
    .A2(_07095_));
 sg13g2_buf_1 _15574_ (.A(_07097_),
    .X(_07098_));
 sg13g2_xor2_1 _15575_ (.B(\soc_I.pwm_I.pwm_accumulator[2] ),
    .A(\soc_I.pwm_I.pcm[2] ),
    .X(_07099_));
 sg13g2_xnor2_1 _15576_ (.Y(_07100_),
    .A(_07098_),
    .B(_07099_));
 sg13g2_nor2_1 _15577_ (.A(net382),
    .B(_07100_),
    .Y(_00916_));
 sg13g2_nor2_1 _15578_ (.A(\soc_I.pwm_I.pwm_accumulator[2] ),
    .B(_07098_),
    .Y(_07101_));
 sg13g2_a21oi_1 _15579_ (.A1(\soc_I.pwm_I.pwm_accumulator[2] ),
    .A2(_07098_),
    .Y(_07102_),
    .B1(\soc_I.pwm_I.pcm[2] ));
 sg13g2_nor2_1 _15580_ (.A(_07101_),
    .B(_07102_),
    .Y(_07103_));
 sg13g2_xor2_1 _15581_ (.B(\soc_I.pwm_I.pwm_accumulator[3] ),
    .A(\soc_I.pwm_I.pcm[3] ),
    .X(_07104_));
 sg13g2_xnor2_1 _15582_ (.Y(_07105_),
    .A(_07103_),
    .B(_07104_));
 sg13g2_nor2_1 _15583_ (.A(net382),
    .B(_07105_),
    .Y(_00917_));
 sg13g2_nor2_1 _15584_ (.A(\soc_I.pwm_I.pwm_accumulator[3] ),
    .B(_07103_),
    .Y(_07106_));
 sg13g2_a21oi_1 _15585_ (.A1(\soc_I.pwm_I.pwm_accumulator[3] ),
    .A2(_07103_),
    .Y(_07107_),
    .B1(\soc_I.pwm_I.pcm[3] ));
 sg13g2_nor2_1 _15586_ (.A(_07106_),
    .B(_07107_),
    .Y(_07108_));
 sg13g2_xor2_1 _15587_ (.B(\soc_I.pwm_I.pwm_accumulator[4] ),
    .A(\soc_I.pwm_I.pcm[4] ),
    .X(_07109_));
 sg13g2_xnor2_1 _15588_ (.Y(_07110_),
    .A(_07108_),
    .B(_07109_));
 sg13g2_nor2_1 _15589_ (.A(_07056_),
    .B(_07110_),
    .Y(_00918_));
 sg13g2_a21o_1 _15590_ (.A2(_07108_),
    .A1(\soc_I.pwm_I.pwm_accumulator[4] ),
    .B1(\soc_I.pwm_I.pcm[4] ),
    .X(_07111_));
 sg13g2_o21ai_1 _15591_ (.B1(_07111_),
    .Y(_07112_),
    .A1(\soc_I.pwm_I.pwm_accumulator[4] ),
    .A2(_07108_));
 sg13g2_buf_1 _15592_ (.A(_07112_),
    .X(_07113_));
 sg13g2_xnor2_1 _15593_ (.Y(_07114_),
    .A(\soc_I.pwm_I.pcm[5] ),
    .B(\soc_I.pwm_I.pwm_accumulator[5] ));
 sg13g2_xnor2_1 _15594_ (.Y(_07115_),
    .A(_07113_),
    .B(_07114_));
 sg13g2_nor2_1 _15595_ (.A(_07056_),
    .B(_07115_),
    .Y(_00919_));
 sg13g2_buf_1 _15596_ (.A(_06002_),
    .X(_07116_));
 sg13g2_inv_1 _15597_ (.Y(_07117_),
    .A(\soc_I.pwm_I.pwm_accumulator[5] ));
 sg13g2_inv_1 _15598_ (.Y(_07118_),
    .A(_07113_));
 sg13g2_a21oi_1 _15599_ (.A1(\soc_I.pwm_I.pwm_accumulator[5] ),
    .A2(_07118_),
    .Y(_07119_),
    .B1(\soc_I.pwm_I.pcm[5] ));
 sg13g2_a21oi_2 _15600_ (.B1(_07119_),
    .Y(_07120_),
    .A2(_07113_),
    .A1(_07117_));
 sg13g2_xor2_1 _15601_ (.B(\soc_I.pwm_I.pwm_accumulator[6] ),
    .A(\soc_I.pwm_I.pcm[6] ),
    .X(_07121_));
 sg13g2_xnor2_1 _15602_ (.Y(_07122_),
    .A(_07120_),
    .B(_07121_));
 sg13g2_nor2_1 _15603_ (.A(_07116_),
    .B(_07122_),
    .Y(_00920_));
 sg13g2_a21o_1 _15604_ (.A2(_07120_),
    .A1(\soc_I.pwm_I.pwm_accumulator[6] ),
    .B1(\soc_I.pwm_I.pcm[6] ),
    .X(_07123_));
 sg13g2_o21ai_1 _15605_ (.B1(_07123_),
    .Y(_07124_),
    .A1(\soc_I.pwm_I.pwm_accumulator[6] ),
    .A2(_07120_));
 sg13g2_xnor2_1 _15606_ (.Y(_07125_),
    .A(_07089_),
    .B(\soc_I.pwm_I.pwm_accumulator[7] ));
 sg13g2_xnor2_1 _15607_ (.Y(_07126_),
    .A(_07124_),
    .B(_07125_));
 sg13g2_nor2_1 _15608_ (.A(net381),
    .B(_07126_),
    .Y(_00921_));
 sg13g2_nor2_1 _15609_ (.A(_07089_),
    .B(\soc_I.pwm_I.pwm_accumulator[7] ),
    .Y(_07127_));
 sg13g2_nor2_1 _15610_ (.A(_07124_),
    .B(_07127_),
    .Y(_07128_));
 sg13g2_a21oi_1 _15611_ (.A1(_07089_),
    .A2(\soc_I.pwm_I.pwm_accumulator[7] ),
    .Y(_07129_),
    .B1(_07128_));
 sg13g2_nor2_1 _15612_ (.A(net381),
    .B(_07129_),
    .Y(_00922_));
 sg13g2_nor3_1 _15613_ (.A(\soc_I.pwm_ready ),
    .B(net520),
    .C(_03854_),
    .Y(_07130_));
 sg13g2_nand2_1 _15614_ (.Y(_07131_),
    .A(_05912_),
    .B(_07130_));
 sg13g2_nor2_1 _15615_ (.A(_05907_),
    .B(_07131_),
    .Y(_00923_));
 sg13g2_nor4_1 _15616_ (.A(_00055_),
    .B(_04356_),
    .C(_04327_),
    .D(_04341_),
    .Y(_07132_));
 sg13g2_nor2_1 _15617_ (.A(_04311_),
    .B(_07132_),
    .Y(_07133_));
 sg13g2_and2_1 _15618_ (.A(_04307_),
    .B(_07133_),
    .X(_07134_));
 sg13g2_nor3_1 _15619_ (.A(net74),
    .B(_04327_),
    .C(_04339_),
    .Y(_07135_));
 sg13g2_o21ai_1 _15620_ (.B1(_07133_),
    .Y(_07136_),
    .A1(_04315_),
    .A2(_04307_));
 sg13g2_inv_1 _15621_ (.Y(_07137_),
    .A(net12));
 sg13g2_a22oi_1 _15622_ (.Y(_07138_),
    .B1(_07136_),
    .B2(_07137_),
    .A2(_07135_),
    .A1(_07134_));
 sg13g2_nand2b_1 _15623_ (.Y(_00924_),
    .B(net437),
    .A_N(_07138_));
 sg13g2_nor2b_1 _15624_ (.A(net18),
    .B_N(_07136_),
    .Y(_07139_));
 sg13g2_and2_1 _15625_ (.A(_05199_),
    .B(_07134_),
    .X(_07140_));
 sg13g2_o21ai_1 _15626_ (.B1(net437),
    .Y(_00925_),
    .A1(_07139_),
    .A2(_07140_));
 sg13g2_buf_2 _15627_ (.A(\soc_I.qqspi_I.is_quad ),
    .X(_07141_));
 sg13g2_buf_1 _15628_ (.A(_07141_),
    .X(_07142_));
 sg13g2_buf_1 _15629_ (.A(net536),
    .X(_07143_));
 sg13g2_buf_1 _15630_ (.A(net461),
    .X(_07144_));
 sg13g2_inv_1 _15631_ (.Y(_07145_),
    .A(_04347_));
 sg13g2_nor2_1 _15632_ (.A(_04344_),
    .B(_04302_),
    .Y(_07146_));
 sg13g2_buf_1 _15633_ (.A(_07146_),
    .X(_07147_));
 sg13g2_nand2_1 _15634_ (.Y(_07148_),
    .A(_07145_),
    .B(_07147_));
 sg13g2_o21ai_1 _15635_ (.B1(net412),
    .Y(_07149_),
    .A1(_04315_),
    .A2(_07148_));
 sg13g2_buf_1 _15636_ (.A(_07149_),
    .X(_07150_));
 sg13g2_nor2_1 _15637_ (.A(net334),
    .B(_07147_),
    .Y(_07151_));
 sg13g2_a21oi_1 _15638_ (.A1(net426),
    .A2(_07150_),
    .Y(_07152_),
    .B1(_07151_));
 sg13g2_nor2_1 _15639_ (.A(_07116_),
    .B(_07152_),
    .Y(_00926_));
 sg13g2_nor2_1 _15640_ (.A(_04315_),
    .B(_00056_),
    .Y(_07153_));
 sg13g2_nor4_1 _15641_ (.A(_00048_),
    .B(_04316_),
    .C(_05196_),
    .D(_07135_),
    .Y(_07154_));
 sg13g2_buf_1 _15642_ (.A(_04297_),
    .X(_07155_));
 sg13g2_o21ai_1 _15643_ (.B1(_07155_),
    .Y(_07156_),
    .A1(_07153_),
    .A2(_07154_));
 sg13g2_mux2_1 _15644_ (.A0(\soc_I.qqspi_I.state[3] ),
    .A1(net432),
    .S(_07156_),
    .X(_07157_));
 sg13g2_and2_1 _15645_ (.A(net427),
    .B(_07157_),
    .X(_00959_));
 sg13g2_nand2_1 _15646_ (.Y(_07158_),
    .A(sclk),
    .B(_04300_));
 sg13g2_nand2_1 _15647_ (.Y(_07159_),
    .A(_00025_),
    .B(net335));
 sg13g2_nand3_1 _15648_ (.B(_07158_),
    .C(_07159_),
    .A(net437),
    .Y(_00960_));
 sg13g2_inv_1 _15649_ (.Y(_07160_),
    .A(net8));
 sg13g2_nor2_1 _15650_ (.A(_04347_),
    .B(net519),
    .Y(_07161_));
 sg13g2_buf_1 _15651_ (.A(_00081_),
    .X(_07162_));
 sg13g2_nand2b_1 _15652_ (.Y(_07163_),
    .B(net593),
    .A_N(_00082_));
 sg13g2_nand3b_1 _15653_ (.B(_07162_),
    .C(_07163_),
    .Y(_07164_),
    .A_N(_07161_));
 sg13g2_o21ai_1 _15654_ (.B1(net518),
    .Y(_07165_),
    .A1(net335),
    .A2(_07164_));
 sg13g2_a21oi_1 _15655_ (.A1(_07160_),
    .A2(_07150_),
    .Y(_00961_),
    .B1(_07165_));
 sg13g2_nor2b_1 _15656_ (.A(net11),
    .B_N(_07150_),
    .Y(_07166_));
 sg13g2_o21ai_1 _15657_ (.B1(_07162_),
    .Y(_07167_),
    .A1(_07163_),
    .A2(_07161_));
 sg13g2_nor2_1 _15658_ (.A(_07150_),
    .B(_07167_),
    .Y(_07168_));
 sg13g2_nor3_1 _15659_ (.A(net383),
    .B(_07166_),
    .C(_07168_),
    .Y(_00962_));
 sg13g2_nor2_1 _15660_ (.A(sio0_si_mosi_o),
    .B(net335),
    .Y(_07169_));
 sg13g2_nor2b_1 _15661_ (.A(net426),
    .B_N(_05310_),
    .Y(_07170_));
 sg13g2_a221oi_1 _15662_ (.B2(net516),
    .C1(_07170_),
    .B1(net517),
    .A1(_05291_),
    .Y(_07171_),
    .A2(net426));
 sg13g2_nor3_1 _15663_ (.A(net383),
    .B(_07169_),
    .C(_07171_),
    .Y(_00963_));
 sg13g2_nand2_1 _15664_ (.Y(_07172_),
    .A(sio1_so_miso_o),
    .B(net336));
 sg13g2_nand3_1 _15665_ (.B(_05297_),
    .C(net335),
    .A(net426),
    .Y(_07173_));
 sg13g2_a21oi_1 _15666_ (.A1(_07172_),
    .A2(_07173_),
    .Y(_00964_),
    .B1(net385));
 sg13g2_nand2_1 _15667_ (.Y(_07174_),
    .A(sio2_o),
    .B(net336));
 sg13g2_nand3_1 _15668_ (.B(_05305_),
    .C(_04313_),
    .A(net426),
    .Y(_07175_));
 sg13g2_a21oi_1 _15669_ (.A1(_07174_),
    .A2(_07175_),
    .Y(_00965_),
    .B1(net385));
 sg13g2_nand2_1 _15670_ (.Y(_07176_),
    .A(sio3_o),
    .B(net336));
 sg13g2_nand3_1 _15671_ (.B(net426),
    .C(_04313_),
    .A(_05310_),
    .Y(_07177_));
 sg13g2_a21oi_1 _15672_ (.A1(_07176_),
    .A2(_07177_),
    .Y(_00966_),
    .B1(net385));
 sg13g2_inv_1 _15673_ (.Y(_07178_),
    .A(_07141_));
 sg13g2_buf_1 _15674_ (.A(_07178_),
    .X(_07179_));
 sg13g2_buf_1 _15675_ (.A(_07141_),
    .X(_07180_));
 sg13g2_and2_1 _15676_ (.A(net535),
    .B(net4),
    .X(_07181_));
 sg13g2_a21oi_1 _15677_ (.A1(net460),
    .A2(net5),
    .Y(_07182_),
    .B1(_07181_));
 sg13g2_nand2_1 _15678_ (.Y(_07183_),
    .A(net607),
    .B(net380));
 sg13g2_o21ai_1 _15679_ (.B1(_07183_),
    .Y(_07184_),
    .A1(net361),
    .A2(_07182_));
 sg13g2_nor2_2 _15680_ (.A(sclk),
    .B(net443),
    .Y(_07185_));
 sg13g2_nand3_1 _15681_ (.B(_04302_),
    .C(net443),
    .A(net593),
    .Y(_07186_));
 sg13g2_nand2b_1 _15682_ (.Y(_07187_),
    .B(_07186_),
    .A_N(_07185_));
 sg13g2_buf_4 _15683_ (.X(_07188_),
    .A(_07187_));
 sg13g2_mux2_1 _15684_ (.A0(_05194_),
    .A1(_07184_),
    .S(_07188_),
    .X(_07189_));
 sg13g2_and2_1 _15685_ (.A(net427),
    .B(_07189_),
    .X(_00967_));
 sg13g2_nor2b_1 _15686_ (.A(net593),
    .B_N(_04302_),
    .Y(_07190_));
 sg13g2_nor3_1 _15687_ (.A(_04311_),
    .B(_07147_),
    .C(_07190_),
    .Y(_07191_));
 sg13g2_nor2_1 _15688_ (.A(_07185_),
    .B(_07191_),
    .Y(_07192_));
 sg13g2_buf_1 _15689_ (.A(_07192_),
    .X(_07193_));
 sg13g2_buf_1 _15690_ (.A(_07193_),
    .X(_07194_));
 sg13g2_buf_1 _15691_ (.A(_07193_),
    .X(_07195_));
 sg13g2_buf_1 _15692_ (.A(net412),
    .X(_07196_));
 sg13g2_buf_1 _15693_ (.A(_04302_),
    .X(_07197_));
 sg13g2_mux2_1 _15694_ (.A0(_06557_),
    .A1(_05926_),
    .S(_07197_),
    .X(_07198_));
 sg13g2_and2_1 _15695_ (.A(net536),
    .B(_05306_),
    .X(_07199_));
 sg13g2_a21oi_1 _15696_ (.A1(net460),
    .A2(_05242_),
    .Y(_07200_),
    .B1(_07199_));
 sg13g2_nor2_1 _15697_ (.A(net380),
    .B(_07200_),
    .Y(_07201_));
 sg13g2_a21oi_1 _15698_ (.A1(net348),
    .A2(_07198_),
    .Y(_07202_),
    .B1(_07201_));
 sg13g2_nor2_1 _15699_ (.A(_07195_),
    .B(_07202_),
    .Y(_07203_));
 sg13g2_a21oi_1 _15700_ (.A1(_05205_),
    .A2(_07194_),
    .Y(_07204_),
    .B1(_07203_));
 sg13g2_nor2_1 _15701_ (.A(net381),
    .B(_07204_),
    .Y(_00968_));
 sg13g2_mux2_1 _15702_ (.A0(_04245_),
    .A1(_05931_),
    .S(_07197_),
    .X(_07205_));
 sg13g2_and2_1 _15703_ (.A(net536),
    .B(_05311_),
    .X(_07206_));
 sg13g2_a21oi_1 _15704_ (.A1(_07178_),
    .A2(_05205_),
    .Y(_07207_),
    .B1(_07206_));
 sg13g2_nor2_1 _15705_ (.A(net412),
    .B(_07207_),
    .Y(_07208_));
 sg13g2_a21oi_1 _15706_ (.A1(net348),
    .A2(_07205_),
    .Y(_07209_),
    .B1(_07208_));
 sg13g2_nor2_1 _15707_ (.A(net312),
    .B(_07209_),
    .Y(_07210_));
 sg13g2_a21oi_1 _15708_ (.A1(_05210_),
    .A2(net313),
    .Y(_07211_),
    .B1(_07210_));
 sg13g2_nor2_1 _15709_ (.A(net381),
    .B(_07211_),
    .Y(_00969_));
 sg13g2_mux2_1 _15710_ (.A0(_03807_),
    .A1(_05937_),
    .S(net534),
    .X(_07212_));
 sg13g2_and2_1 _15711_ (.A(net536),
    .B(_05237_),
    .X(_07213_));
 sg13g2_a21oi_1 _15712_ (.A1(_07178_),
    .A2(_05210_),
    .Y(_07214_),
    .B1(_07213_));
 sg13g2_nor2_1 _15713_ (.A(net412),
    .B(_07214_),
    .Y(_07215_));
 sg13g2_a21oi_1 _15714_ (.A1(net348),
    .A2(_07212_),
    .Y(_07216_),
    .B1(_07215_));
 sg13g2_nor2_1 _15715_ (.A(_07195_),
    .B(_07216_),
    .Y(_07217_));
 sg13g2_a21oi_1 _15716_ (.A1(_05215_),
    .A2(_07194_),
    .Y(_07218_),
    .B1(_07217_));
 sg13g2_nor2_1 _15717_ (.A(net381),
    .B(_07218_),
    .Y(_00970_));
 sg13g2_buf_1 _15718_ (.A(_07193_),
    .X(_07219_));
 sg13g2_buf_1 _15719_ (.A(_04302_),
    .X(_07220_));
 sg13g2_buf_1 _15720_ (.A(net411),
    .X(_07221_));
 sg13g2_buf_1 _15721_ (.A(_04321_),
    .X(_07222_));
 sg13g2_nor2_1 _15722_ (.A(net346),
    .B(_04656_),
    .Y(_07223_));
 sg13g2_a21oi_1 _15723_ (.A1(_02425_),
    .A2(net347),
    .Y(_07224_),
    .B1(_07223_));
 sg13g2_nand2_1 _15724_ (.Y(_07225_),
    .A(net591),
    .B(_05943_));
 sg13g2_o21ai_1 _15725_ (.B1(_07225_),
    .Y(_07226_),
    .A1(net533),
    .A2(_07224_));
 sg13g2_nor2_1 _15726_ (.A(net360),
    .B(_07226_),
    .Y(_07227_));
 sg13g2_buf_1 _15727_ (.A(net535),
    .X(_07228_));
 sg13g2_nor2b_1 _15728_ (.A(net461),
    .B_N(_05215_),
    .Y(_07229_));
 sg13g2_a221oi_1 _15729_ (.B2(net516),
    .C1(_07229_),
    .B1(net517),
    .A1(net459),
    .Y(_07230_),
    .A2(_05242_));
 sg13g2_nor3_1 _15730_ (.A(_07219_),
    .B(_07227_),
    .C(_07230_),
    .Y(_07231_));
 sg13g2_a21oi_1 _15731_ (.A1(_05220_),
    .A2(net313),
    .Y(_07232_),
    .B1(_07231_));
 sg13g2_nor2_1 _15732_ (.A(net381),
    .B(_07232_),
    .Y(_00971_));
 sg13g2_mux2_1 _15733_ (.A0(_05220_),
    .A1(_05205_),
    .S(net535),
    .X(_07233_));
 sg13g2_nand2_1 _15734_ (.Y(_07234_),
    .A(_02337_),
    .B(net411));
 sg13g2_o21ai_1 _15735_ (.B1(_07234_),
    .Y(_07235_),
    .A1(net346),
    .A2(_04660_));
 sg13g2_a21oi_1 _15736_ (.A1(_05946_),
    .A2(net397),
    .Y(_07236_),
    .B1(_05947_));
 sg13g2_nand2_1 _15737_ (.Y(_07237_),
    .A(net591),
    .B(_07236_));
 sg13g2_o21ai_1 _15738_ (.B1(_07237_),
    .Y(_07238_),
    .A1(net591),
    .A2(_07235_));
 sg13g2_nor2_1 _15739_ (.A(_04357_),
    .B(_07238_),
    .Y(_07239_));
 sg13g2_a21oi_1 _15740_ (.A1(net334),
    .A2(_07233_),
    .Y(_07240_),
    .B1(_07239_));
 sg13g2_nor2_1 _15741_ (.A(net312),
    .B(_07240_),
    .Y(_07241_));
 sg13g2_a21oi_1 _15742_ (.A1(_05225_),
    .A2(net313),
    .Y(_07242_),
    .B1(_07241_));
 sg13g2_nor2_1 _15743_ (.A(net381),
    .B(_07242_),
    .Y(_00972_));
 sg13g2_nor2_1 _15744_ (.A(net346),
    .B(_04668_),
    .Y(_07243_));
 sg13g2_a21oi_1 _15745_ (.A1(_02330_),
    .A2(net347),
    .Y(_07244_),
    .B1(_07243_));
 sg13g2_nand2_1 _15746_ (.Y(_07245_),
    .A(net591),
    .B(_05953_));
 sg13g2_o21ai_1 _15747_ (.B1(_07245_),
    .Y(_07246_),
    .A1(net533),
    .A2(_07244_));
 sg13g2_nor2_1 _15748_ (.A(net360),
    .B(_07246_),
    .Y(_07247_));
 sg13g2_nor2b_1 _15749_ (.A(net461),
    .B_N(_05225_),
    .Y(_07248_));
 sg13g2_a221oi_1 _15750_ (.B2(net516),
    .C1(_07248_),
    .B1(net517),
    .A1(net459),
    .Y(_07249_),
    .A2(_05210_));
 sg13g2_nor3_1 _15751_ (.A(net311),
    .B(_07247_),
    .C(_07249_),
    .Y(_07250_));
 sg13g2_a21oi_1 _15752_ (.A1(_05230_),
    .A2(net313),
    .Y(_07251_),
    .B1(_07250_));
 sg13g2_nor2_1 _15753_ (.A(net381),
    .B(_07251_),
    .Y(_00973_));
 sg13g2_buf_1 _15754_ (.A(_06002_),
    .X(_07252_));
 sg13g2_and2_1 _15755_ (.A(_01929_),
    .B(net346),
    .X(_07253_));
 sg13g2_a21oi_1 _15756_ (.A1(_04323_),
    .A2(_04673_),
    .Y(_07254_),
    .B1(_07253_));
 sg13g2_nand2_1 _15757_ (.Y(_07255_),
    .A(net534),
    .B(_05958_));
 sg13g2_o21ai_1 _15758_ (.B1(_07255_),
    .Y(_07256_),
    .A1(net533),
    .A2(_07254_));
 sg13g2_and2_1 _15759_ (.A(_07141_),
    .B(_05215_),
    .X(_07257_));
 sg13g2_a21oi_1 _15760_ (.A1(_07178_),
    .A2(_05230_),
    .Y(_07258_),
    .B1(_07257_));
 sg13g2_nor2_1 _15761_ (.A(net412),
    .B(_07258_),
    .Y(_07259_));
 sg13g2_a21oi_1 _15762_ (.A1(net348),
    .A2(_07256_),
    .Y(_07260_),
    .B1(_07259_));
 sg13g2_nor2_1 _15763_ (.A(net311),
    .B(_07260_),
    .Y(_07261_));
 sg13g2_a21oi_1 _15764_ (.A1(_05235_),
    .A2(net313),
    .Y(_07262_),
    .B1(_07261_));
 sg13g2_nor2_1 _15765_ (.A(_07252_),
    .B(_07262_),
    .Y(_00974_));
 sg13g2_and2_1 _15766_ (.A(_01943_),
    .B(net346),
    .X(_07263_));
 sg13g2_a21oi_1 _15767_ (.A1(net359),
    .A2(_03888_),
    .Y(_07264_),
    .B1(_07263_));
 sg13g2_nand2_1 _15768_ (.Y(_07265_),
    .A(net591),
    .B(_05962_));
 sg13g2_o21ai_1 _15769_ (.B1(_07265_),
    .Y(_07266_),
    .A1(net533),
    .A2(_07264_));
 sg13g2_and2_1 _15770_ (.A(_07141_),
    .B(_05220_),
    .X(_07267_));
 sg13g2_a21oi_1 _15771_ (.A1(_07178_),
    .A2(_05235_),
    .Y(_07268_),
    .B1(_07267_));
 sg13g2_nor2_1 _15772_ (.A(net412),
    .B(_07268_),
    .Y(_07269_));
 sg13g2_a21oi_1 _15773_ (.A1(_07196_),
    .A2(_07266_),
    .Y(_07270_),
    .B1(_07269_));
 sg13g2_nor2_1 _15774_ (.A(_07219_),
    .B(_07270_),
    .Y(_07271_));
 sg13g2_a21oi_1 _15775_ (.A1(_05241_),
    .A2(net313),
    .Y(_07272_),
    .B1(_07271_));
 sg13g2_nor2_1 _15776_ (.A(net379),
    .B(_07272_),
    .Y(_00975_));
 sg13g2_nor2_1 _15777_ (.A(net346),
    .B(net117),
    .Y(_07273_));
 sg13g2_a21oi_1 _15778_ (.A1(_01959_),
    .A2(net346),
    .Y(_07274_),
    .B1(_07273_));
 sg13g2_nand2_1 _15779_ (.Y(_07275_),
    .A(_04303_),
    .B(_05966_));
 sg13g2_o21ai_1 _15780_ (.B1(_07275_),
    .Y(_07276_),
    .A1(net533),
    .A2(_07274_));
 sg13g2_nor2_1 _15781_ (.A(net360),
    .B(_07276_),
    .Y(_07277_));
 sg13g2_nor2b_1 _15782_ (.A(net461),
    .B_N(_05241_),
    .Y(_07278_));
 sg13g2_a221oi_1 _15783_ (.B2(net516),
    .C1(_07278_),
    .B1(net517),
    .A1(net459),
    .Y(_07279_),
    .A2(_05225_));
 sg13g2_nor3_1 _15784_ (.A(net311),
    .B(_07277_),
    .C(_07279_),
    .Y(_07280_));
 sg13g2_a21oi_1 _15785_ (.A1(_05206_),
    .A2(net313),
    .Y(_07281_),
    .B1(_07280_));
 sg13g2_nor2_1 _15786_ (.A(net379),
    .B(_07281_),
    .Y(_00976_));
 sg13g2_mux2_1 _15787_ (.A0(_05206_),
    .A1(_05230_),
    .S(net535),
    .X(_07282_));
 sg13g2_nand2_1 _15788_ (.Y(_07283_),
    .A(net359),
    .B(_04014_));
 sg13g2_nand2_1 _15789_ (.Y(_07284_),
    .A(_01979_),
    .B(net411));
 sg13g2_a21oi_1 _15790_ (.A1(_07283_),
    .A2(_07284_),
    .Y(_07285_),
    .B1(net591));
 sg13g2_a21oi_1 _15791_ (.A1(net534),
    .A2(_05970_),
    .Y(_07286_),
    .B1(_07285_));
 sg13g2_nor2_1 _15792_ (.A(net358),
    .B(_07286_),
    .Y(_07287_));
 sg13g2_a21oi_1 _15793_ (.A1(net360),
    .A2(_07282_),
    .Y(_07288_),
    .B1(_07287_));
 sg13g2_nor2_1 _15794_ (.A(net311),
    .B(_07288_),
    .Y(_07289_));
 sg13g2_a21oi_1 _15795_ (.A1(_05211_),
    .A2(net313),
    .Y(_07290_),
    .B1(_07289_));
 sg13g2_nor2_1 _15796_ (.A(net379),
    .B(_07290_),
    .Y(_00977_));
 sg13g2_and2_1 _15797_ (.A(net535),
    .B(net5),
    .X(_07291_));
 sg13g2_a21oi_1 _15798_ (.A1(net460),
    .A2(_05194_),
    .Y(_07292_),
    .B1(_07291_));
 sg13g2_nand2_1 _15799_ (.Y(_07293_),
    .A(net604),
    .B(net380));
 sg13g2_o21ai_1 _15800_ (.B1(_07293_),
    .Y(_07294_),
    .A1(_04299_),
    .A2(_07292_));
 sg13g2_mux2_1 _15801_ (.A0(_05255_),
    .A1(_07294_),
    .S(_07188_),
    .X(_07295_));
 sg13g2_and2_1 _15802_ (.A(net427),
    .B(_07295_),
    .X(_00978_));
 sg13g2_mux2_1 _15803_ (.A0(_05211_),
    .A1(_05235_),
    .S(net535),
    .X(_07296_));
 sg13g2_nor2_1 _15804_ (.A(_01864_),
    .B(net359),
    .Y(_07297_));
 sg13g2_nor3_1 _15805_ (.A(_04302_),
    .B(_03918_),
    .C(_07297_),
    .Y(_07298_));
 sg13g2_a21oi_1 _15806_ (.A1(net534),
    .A2(_05974_),
    .Y(_07299_),
    .B1(_07298_));
 sg13g2_nor2_1 _15807_ (.A(net358),
    .B(_07299_),
    .Y(_07300_));
 sg13g2_a21oi_1 _15808_ (.A1(net360),
    .A2(_07296_),
    .Y(_07301_),
    .B1(_07300_));
 sg13g2_nor2_1 _15809_ (.A(net311),
    .B(_07301_),
    .Y(_07302_));
 sg13g2_a21oi_1 _15810_ (.A1(_05216_),
    .A2(net312),
    .Y(_07303_),
    .B1(_07302_));
 sg13g2_nor2_1 _15811_ (.A(net379),
    .B(_07303_),
    .Y(_00979_));
 sg13g2_mux2_1 _15812_ (.A0(_05216_),
    .A1(_05241_),
    .S(_07180_),
    .X(_07304_));
 sg13g2_nand2_1 _15813_ (.Y(_07305_),
    .A(_01903_),
    .B(_04321_));
 sg13g2_nand2_1 _15814_ (.Y(_07306_),
    .A(net359),
    .B(_04575_));
 sg13g2_a21oi_1 _15815_ (.A1(_07305_),
    .A2(_07306_),
    .Y(_07307_),
    .B1(_04302_));
 sg13g2_a21oi_1 _15816_ (.A1(net534),
    .A2(_05978_),
    .Y(_07308_),
    .B1(_07307_));
 sg13g2_nor2_1 _15817_ (.A(net358),
    .B(_07308_),
    .Y(_07309_));
 sg13g2_a21oi_1 _15818_ (.A1(net360),
    .A2(_07304_),
    .Y(_07310_),
    .B1(_07309_));
 sg13g2_nor2_1 _15819_ (.A(net311),
    .B(_07310_),
    .Y(_07311_));
 sg13g2_a21oi_1 _15820_ (.A1(_05221_),
    .A2(net312),
    .Y(_07312_),
    .B1(_07311_));
 sg13g2_nor2_1 _15821_ (.A(net379),
    .B(_07312_),
    .Y(_00980_));
 sg13g2_nor2_1 _15822_ (.A(_07222_),
    .B(net98),
    .Y(_07313_));
 sg13g2_a21oi_1 _15823_ (.A1(_01883_),
    .A2(_07222_),
    .Y(_07314_),
    .B1(_07313_));
 sg13g2_nand2_1 _15824_ (.Y(_07315_),
    .A(_04303_),
    .B(_05984_));
 sg13g2_o21ai_1 _15825_ (.B1(_07315_),
    .Y(_07316_),
    .A1(net533),
    .A2(_07314_));
 sg13g2_nor2_1 _15826_ (.A(net358),
    .B(_07316_),
    .Y(_07317_));
 sg13g2_nor2b_1 _15827_ (.A(_07143_),
    .B_N(_05221_),
    .Y(_07318_));
 sg13g2_a221oi_1 _15828_ (.B2(_04309_),
    .C1(_07318_),
    .B1(_04308_),
    .A1(_07228_),
    .Y(_07319_),
    .A2(_05206_));
 sg13g2_nor3_1 _15829_ (.A(_07193_),
    .B(_07317_),
    .C(_07319_),
    .Y(_07320_));
 sg13g2_a21oi_1 _15830_ (.A1(_05226_),
    .A2(net312),
    .Y(_07321_),
    .B1(_07320_));
 sg13g2_nor2_1 _15831_ (.A(net379),
    .B(_07321_),
    .Y(_00981_));
 sg13g2_mux2_1 _15832_ (.A0(_05226_),
    .A1(_05211_),
    .S(_07180_),
    .X(_07322_));
 sg13g2_nand2_1 _15833_ (.Y(_07323_),
    .A(net359),
    .B(net130));
 sg13g2_o21ai_1 _15834_ (.B1(_07323_),
    .Y(_07324_),
    .A1(_01826_),
    .A2(net359));
 sg13g2_nor2_1 _15835_ (.A(net591),
    .B(_07324_),
    .Y(_07325_));
 sg13g2_a21oi_1 _15836_ (.A1(net534),
    .A2(_05988_),
    .Y(_07326_),
    .B1(_07325_));
 sg13g2_nor2_1 _15837_ (.A(net358),
    .B(_07326_),
    .Y(_07327_));
 sg13g2_a21oi_1 _15838_ (.A1(_04312_),
    .A2(_07322_),
    .Y(_07328_),
    .B1(_07327_));
 sg13g2_nor2_1 _15839_ (.A(net311),
    .B(_07328_),
    .Y(_07329_));
 sg13g2_a21oi_1 _15840_ (.A1(_05231_),
    .A2(net312),
    .Y(_07330_),
    .B1(_07329_));
 sg13g2_nor2_1 _15841_ (.A(net379),
    .B(_07330_),
    .Y(_00982_));
 sg13g2_inv_1 _15842_ (.Y(_07331_),
    .A(_04350_));
 sg13g2_a21oi_1 _15843_ (.A1(_07331_),
    .A2(_07147_),
    .Y(_07332_),
    .B1(_07190_));
 sg13g2_a21oi_2 _15844_ (.B1(_07185_),
    .Y(_07333_),
    .A2(_07332_),
    .A1(net443));
 sg13g2_inv_1 _15845_ (.Y(_07334_),
    .A(_07333_));
 sg13g2_nor2_2 _15846_ (.A(net520),
    .B(_07334_),
    .Y(_07335_));
 sg13g2_nand2b_1 _15847_ (.Y(_07336_),
    .B(net461),
    .A_N(_05216_));
 sg13g2_o21ai_1 _15848_ (.B1(_07336_),
    .Y(_07337_),
    .A1(_07144_),
    .A2(_05231_));
 sg13g2_nor2_1 _15849_ (.A(_07162_),
    .B(_07147_),
    .Y(_07338_));
 sg13g2_nand2_1 _15850_ (.Y(_07339_),
    .A(_02150_),
    .B(net347));
 sg13g2_o21ai_1 _15851_ (.B1(_07339_),
    .Y(_07340_),
    .A1(net347),
    .A2(_04589_));
 sg13g2_a21o_1 _15852_ (.A2(_07147_),
    .A1(net521),
    .B1(_04311_),
    .X(_07341_));
 sg13g2_buf_1 _15853_ (.A(_07341_),
    .X(_07342_));
 sg13g2_a21oi_1 _15854_ (.A1(_07338_),
    .A2(_07340_),
    .Y(_07343_),
    .B1(_07342_));
 sg13g2_nor2_1 _15855_ (.A(net521),
    .B(net505),
    .Y(_07344_));
 sg13g2_buf_1 _15856_ (.A(_07344_),
    .X(_07345_));
 sg13g2_nand2_1 _15857_ (.Y(_07346_),
    .A(_04603_),
    .B(_07345_));
 sg13g2_a21oi_2 _15858_ (.B1(_07346_),
    .Y(_07347_),
    .A2(net397),
    .A1(net76));
 sg13g2_nand2b_1 _15859_ (.Y(_07348_),
    .B(_07347_),
    .A_N(_06046_));
 sg13g2_and3_1 _15860_ (.X(_07349_),
    .A(_03574_),
    .B(_05924_),
    .C(_07345_));
 sg13g2_buf_2 _15861_ (.A(_07349_),
    .X(_07350_));
 sg13g2_nand2b_1 _15862_ (.Y(_07351_),
    .B(_07350_),
    .A_N(net607));
 sg13g2_and2_1 _15863_ (.A(_04603_),
    .B(_07345_),
    .X(_07352_));
 sg13g2_buf_1 _15864_ (.A(_07352_),
    .X(_07353_));
 sg13g2_a21oi_1 _15865_ (.A1(\soc_I.cpu_mem_addr[1] ),
    .A2(_07350_),
    .Y(_07354_),
    .B1(_07353_));
 sg13g2_nand2b_1 _15866_ (.Y(_07355_),
    .B(_07354_),
    .A_N(_05993_));
 sg13g2_nand4_1 _15867_ (.B(_07348_),
    .C(_07351_),
    .A(net519),
    .Y(_07356_),
    .D(_07355_));
 sg13g2_nand2_1 _15868_ (.Y(_07357_),
    .A(_03576_),
    .B(_07334_));
 sg13g2_a221oi_1 _15869_ (.B2(_07356_),
    .C1(_07357_),
    .B1(_07343_),
    .A1(net334),
    .Y(_07358_),
    .A2(_07337_));
 sg13g2_a21o_1 _15870_ (.A2(_07335_),
    .A1(_05200_),
    .B1(_07358_),
    .X(_00983_));
 sg13g2_inv_1 _15871_ (.Y(_07359_),
    .A(_07162_));
 sg13g2_nand2_1 _15872_ (.Y(_07360_),
    .A(_02134_),
    .B(net411));
 sg13g2_o21ai_1 _15873_ (.B1(_07360_),
    .Y(_07361_),
    .A1(net411),
    .A2(_03730_));
 sg13g2_nand2_1 _15874_ (.Y(_07362_),
    .A(_07359_),
    .B(_07361_));
 sg13g2_nor2_1 _15875_ (.A(_03765_),
    .B(_04344_),
    .Y(_07363_));
 sg13g2_a21oi_1 _15876_ (.A1(_04344_),
    .A2(_07362_),
    .Y(_07364_),
    .B1(_07363_));
 sg13g2_nor3_1 _15877_ (.A(net519),
    .B(net334),
    .C(_07364_),
    .Y(_07365_));
 sg13g2_nor2b_1 _15878_ (.A(net459),
    .B_N(_05200_),
    .Y(_07366_));
 sg13g2_a221oi_1 _15879_ (.B2(net516),
    .C1(_07366_),
    .B1(net517),
    .A1(net459),
    .Y(_07367_),
    .A2(_05221_));
 sg13g2_a21o_1 _15880_ (.A2(_07347_),
    .A1(net397),
    .B1(_07350_),
    .X(_07368_));
 sg13g2_nand3b_1 _15881_ (.B(_07353_),
    .C(_01952_),
    .Y(_07369_),
    .A_N(net397));
 sg13g2_nand4_1 _15882_ (.B(_04298_),
    .C(_07362_),
    .A(net519),
    .Y(_07370_),
    .D(_07369_));
 sg13g2_a221oi_1 _15883_ (.B2(net604),
    .C1(_07370_),
    .B1(_07368_),
    .A1(_05999_),
    .Y(_07371_),
    .A2(_07354_));
 sg13g2_nor4_1 _15884_ (.A(_07357_),
    .B(_07365_),
    .C(_07367_),
    .D(_07371_),
    .Y(_07372_));
 sg13g2_a21o_1 _15885_ (.A2(_07335_),
    .A1(_05256_),
    .B1(_07372_),
    .X(_00984_));
 sg13g2_nand2_1 _15886_ (.Y(_07373_),
    .A(_06009_),
    .B(_07354_));
 sg13g2_nand2_1 _15887_ (.Y(_07374_),
    .A(_02117_),
    .B(net346));
 sg13g2_o21ai_1 _15888_ (.B1(_07374_),
    .Y(_07375_),
    .A1(net347),
    .A2(_04597_));
 sg13g2_and2_1 _15889_ (.A(_07141_),
    .B(_05226_),
    .X(_07376_));
 sg13g2_a21oi_1 _15890_ (.A1(_07178_),
    .A2(_05256_),
    .Y(_07377_),
    .B1(_07376_));
 sg13g2_o21ai_1 _15891_ (.B1(_07334_),
    .Y(_07378_),
    .A1(net443),
    .A2(_07377_));
 sg13g2_a21oi_1 _15892_ (.A1(_07359_),
    .A2(_07375_),
    .Y(_07379_),
    .B1(_07378_));
 sg13g2_a22oi_1 _15893_ (.Y(_07380_),
    .B1(_07350_),
    .B2(net619),
    .A2(_07347_),
    .A1(_05926_));
 sg13g2_and3_1 _15894_ (.X(_07381_),
    .A(_07373_),
    .B(_07379_),
    .C(_07380_));
 sg13g2_o21ai_1 _15895_ (.B1(net515),
    .Y(_07382_),
    .A1(_05279_),
    .A2(_07334_));
 sg13g2_nand2_1 _15896_ (.Y(_07383_),
    .A(_00082_),
    .B(_07379_));
 sg13g2_o21ai_1 _15897_ (.B1(_07383_),
    .Y(_07384_),
    .A1(_07151_),
    .A2(_07378_));
 sg13g2_nor3_1 _15898_ (.A(_07381_),
    .B(_07382_),
    .C(_07384_),
    .Y(_00985_));
 sg13g2_inv_1 _15899_ (.Y(_07385_),
    .A(_06014_));
 sg13g2_and2_1 _15900_ (.A(\soc_I.cpu_mem_addr[1] ),
    .B(_07350_),
    .X(_07386_));
 sg13g2_buf_1 _15901_ (.A(_07386_),
    .X(_07387_));
 sg13g2_or2_1 _15902_ (.X(_07388_),
    .B(_07387_),
    .A(_07353_));
 sg13g2_buf_2 _15903_ (.A(_07388_),
    .X(_07389_));
 sg13g2_a22oi_1 _15904_ (.Y(_07390_),
    .B1(_07387_),
    .B2(_05970_),
    .A2(_07353_),
    .A1(_05931_));
 sg13g2_o21ai_1 _15905_ (.B1(_07390_),
    .Y(_07391_),
    .A1(_07385_),
    .A2(_07389_));
 sg13g2_nor2_1 _15906_ (.A(net347),
    .B(_03749_),
    .Y(_07392_));
 sg13g2_a21oi_1 _15907_ (.A1(_02099_),
    .A2(net347),
    .Y(_07393_),
    .B1(_07392_));
 sg13g2_o21ai_1 _15908_ (.B1(_07191_),
    .Y(_07394_),
    .A1(_07162_),
    .A2(_07393_));
 sg13g2_a21oi_1 _15909_ (.A1(_04304_),
    .A2(_07391_),
    .Y(_07395_),
    .B1(_07394_));
 sg13g2_nand2b_1 _15910_ (.Y(_07396_),
    .B(net461),
    .A_N(_05231_));
 sg13g2_o21ai_1 _15911_ (.B1(_07396_),
    .Y(_07397_),
    .A1(net459),
    .A2(_05279_));
 sg13g2_a21oi_1 _15912_ (.A1(net334),
    .A2(_07397_),
    .Y(_07398_),
    .B1(_07333_));
 sg13g2_a21oi_1 _15913_ (.A1(_05285_),
    .A2(_07333_),
    .Y(_07399_),
    .B1(_07398_));
 sg13g2_nor3_1 _15914_ (.A(net383),
    .B(_07395_),
    .C(_07399_),
    .Y(_00986_));
 sg13g2_or3_1 _15915_ (.A(_01856_),
    .B(net397),
    .C(_07346_),
    .X(_07400_));
 sg13g2_nand2b_1 _15916_ (.Y(_07401_),
    .B(net535),
    .A_N(_05200_));
 sg13g2_o21ai_1 _15917_ (.B1(_07401_),
    .Y(_07402_),
    .A1(net535),
    .A2(_05285_));
 sg13g2_a21oi_1 _15918_ (.A1(net358),
    .A2(_07402_),
    .Y(_07403_),
    .B1(_07357_));
 sg13g2_nand3_1 _15919_ (.B(_07400_),
    .C(_07403_),
    .A(net519),
    .Y(_07404_));
 sg13g2_nand2b_1 _15920_ (.Y(_07405_),
    .B(_07368_),
    .A_N(net606));
 sg13g2_o21ai_1 _15921_ (.B1(_07405_),
    .Y(_07406_),
    .A1(_06019_),
    .A2(_07389_));
 sg13g2_a21oi_1 _15922_ (.A1(_07359_),
    .A2(_04606_),
    .Y(_07407_),
    .B1(_07147_));
 sg13g2_a22oi_1 _15923_ (.Y(_07408_),
    .B1(_04606_),
    .B2(_01556_),
    .A2(net347),
    .A1(_02049_));
 sg13g2_nor2b_1 _15924_ (.A(_07408_),
    .B_N(_07338_),
    .Y(_07409_));
 sg13g2_nor2_1 _15925_ (.A(net360),
    .B(_07409_),
    .Y(_07410_));
 sg13g2_o21ai_1 _15926_ (.B1(_07410_),
    .Y(_07411_),
    .A1(_03765_),
    .A2(_07407_));
 sg13g2_a22oi_1 _15927_ (.Y(_07412_),
    .B1(_07403_),
    .B2(_07411_),
    .A2(_07335_),
    .A1(_05291_));
 sg13g2_o21ai_1 _15928_ (.B1(_07412_),
    .Y(_00987_),
    .A1(_07404_),
    .A2(_07406_));
 sg13g2_inv_1 _15929_ (.Y(_07413_),
    .A(_06024_));
 sg13g2_a22oi_1 _15930_ (.Y(_07414_),
    .B1(_07387_),
    .B2(_05978_),
    .A2(_07353_),
    .A1(_05943_));
 sg13g2_o21ai_1 _15931_ (.B1(_07414_),
    .Y(_07415_),
    .A1(_07413_),
    .A2(_07389_));
 sg13g2_o21ai_1 _15932_ (.B1(_07359_),
    .Y(_07416_),
    .A1(_02039_),
    .A2(_04323_));
 sg13g2_o21ai_1 _15933_ (.B1(_07191_),
    .Y(_07417_),
    .A1(_03782_),
    .A2(_07416_));
 sg13g2_a21oi_1 _15934_ (.A1(net519),
    .A2(_07415_),
    .Y(_07418_),
    .B1(_07417_));
 sg13g2_nand2b_1 _15935_ (.Y(_07419_),
    .B(net461),
    .A_N(_05256_));
 sg13g2_o21ai_1 _15936_ (.B1(_07419_),
    .Y(_07420_),
    .A1(_05291_),
    .A2(net459));
 sg13g2_a21oi_1 _15937_ (.A1(net334),
    .A2(_07420_),
    .Y(_07421_),
    .B1(_07333_));
 sg13g2_a21oi_1 _15938_ (.A1(_05297_),
    .A2(_07333_),
    .Y(_07422_),
    .B1(_07421_));
 sg13g2_nor3_1 _15939_ (.A(net383),
    .B(_07418_),
    .C(_07422_),
    .Y(_00988_));
 sg13g2_and2_1 _15940_ (.A(net536),
    .B(net6),
    .X(_07423_));
 sg13g2_a21oi_1 _15941_ (.A1(net460),
    .A2(_05255_),
    .Y(_07424_),
    .B1(_07423_));
 sg13g2_nand2_1 _15942_ (.Y(_07425_),
    .A(_02277_),
    .B(net380));
 sg13g2_o21ai_1 _15943_ (.B1(_07425_),
    .Y(_07426_),
    .A1(net361),
    .A2(_07424_));
 sg13g2_mux2_1 _15944_ (.A0(_05280_),
    .A1(_07426_),
    .S(_07188_),
    .X(_07427_));
 sg13g2_and2_1 _15945_ (.A(net427),
    .B(_07427_),
    .X(_00989_));
 sg13g2_nand2b_1 _15946_ (.Y(_07428_),
    .B(net461),
    .A_N(_05279_));
 sg13g2_o21ai_1 _15947_ (.B1(_07428_),
    .Y(_07429_),
    .A1(_07144_),
    .A2(_05297_));
 sg13g2_nand2_1 _15948_ (.Y(_07430_),
    .A(_02064_),
    .B(_07221_));
 sg13g2_o21ai_1 _15949_ (.B1(_07430_),
    .Y(_07431_),
    .A1(_07221_),
    .A2(_04207_));
 sg13g2_a21oi_1 _15950_ (.A1(_07338_),
    .A2(_07431_),
    .Y(_07432_),
    .B1(_07342_));
 sg13g2_a22oi_1 _15951_ (.Y(_07433_),
    .B1(_07350_),
    .B2(_05982_),
    .A2(_07347_),
    .A1(_07236_));
 sg13g2_and2_1 _15952_ (.A(net533),
    .B(_07433_),
    .X(_07434_));
 sg13g2_o21ai_1 _15953_ (.B1(_07434_),
    .Y(_07435_),
    .A1(_06030_),
    .A2(_07389_));
 sg13g2_a221oi_1 _15954_ (.B2(_07435_),
    .C1(_07357_),
    .B1(_07432_),
    .A1(_04358_),
    .Y(_07436_),
    .A2(_07429_));
 sg13g2_a21o_1 _15955_ (.A2(_07335_),
    .A1(_05305_),
    .B1(_07436_),
    .X(_00990_));
 sg13g2_nand2b_1 _15956_ (.Y(_07437_),
    .B(net459),
    .A_N(_05285_));
 sg13g2_o21ai_1 _15957_ (.B1(_07437_),
    .Y(_07438_),
    .A1(net426),
    .A2(_05305_));
 sg13g2_a21o_1 _15958_ (.A2(_07438_),
    .A1(net335),
    .B1(_07357_),
    .X(_07439_));
 sg13g2_inv_1 _15959_ (.Y(_07440_),
    .A(_06035_));
 sg13g2_a22oi_1 _15960_ (.Y(_07441_),
    .B1(_07350_),
    .B2(net605),
    .A2(_07347_),
    .A1(_05953_));
 sg13g2_o21ai_1 _15961_ (.B1(_07441_),
    .Y(_07442_),
    .A1(_07440_),
    .A2(_07389_));
 sg13g2_a221oi_1 _15962_ (.B2(net519),
    .C1(_07342_),
    .B1(_07442_),
    .A1(_04344_),
    .Y(_07443_),
    .A2(_04335_));
 sg13g2_nand2_1 _15963_ (.Y(_07444_),
    .A(_05310_),
    .B(_07335_));
 sg13g2_o21ai_1 _15964_ (.B1(_07444_),
    .Y(_00991_),
    .A1(_07439_),
    .A2(_07443_));
 sg13g2_and2_1 _15965_ (.A(net536),
    .B(net7),
    .X(_07445_));
 sg13g2_a21oi_1 _15966_ (.A1(_07179_),
    .A2(_05280_),
    .Y(_07446_),
    .B1(_07445_));
 sg13g2_nand2_1 _15967_ (.Y(_07447_),
    .A(_05929_),
    .B(_07155_));
 sg13g2_o21ai_1 _15968_ (.B1(_07447_),
    .Y(_07448_),
    .A1(net348),
    .A2(_07446_));
 sg13g2_mux2_1 _15969_ (.A0(_05286_),
    .A1(_07448_),
    .S(_07188_),
    .X(_07449_));
 sg13g2_and2_1 _15970_ (.A(net427),
    .B(_07449_),
    .X(_00992_));
 sg13g2_and2_1 _15971_ (.A(_07142_),
    .B(_05194_),
    .X(_07450_));
 sg13g2_a21oi_1 _15972_ (.A1(net460),
    .A2(_05286_),
    .Y(_07451_),
    .B1(_07450_));
 sg13g2_nand2_1 _15973_ (.Y(_07452_),
    .A(net606),
    .B(net380));
 sg13g2_o21ai_1 _15974_ (.B1(_07452_),
    .Y(_07453_),
    .A1(net348),
    .A2(_07451_));
 sg13g2_mux2_1 _15975_ (.A0(_05293_),
    .A1(_07453_),
    .S(_07188_),
    .X(_07454_));
 sg13g2_and2_1 _15976_ (.A(_07088_),
    .B(_07454_),
    .X(_00993_));
 sg13g2_and2_1 _15977_ (.A(_07142_),
    .B(_05255_),
    .X(_07455_));
 sg13g2_a21oi_1 _15978_ (.A1(net460),
    .A2(_05293_),
    .Y(_07456_),
    .B1(_07455_));
 sg13g2_nand2_1 _15979_ (.Y(_07457_),
    .A(_05941_),
    .B(net380));
 sg13g2_o21ai_1 _15980_ (.B1(_07457_),
    .Y(_07458_),
    .A1(_07196_),
    .A2(_07456_));
 sg13g2_mux2_1 _15981_ (.A0(_05298_),
    .A1(_07458_),
    .S(_07188_),
    .X(_07459_));
 sg13g2_and2_1 _15982_ (.A(_07088_),
    .B(_07459_),
    .X(_00994_));
 sg13g2_mux2_1 _15983_ (.A0(_05298_),
    .A1(_05280_),
    .S(net536),
    .X(_07460_));
 sg13g2_nand2_1 _15984_ (.Y(_07461_),
    .A(_04357_),
    .B(_07460_));
 sg13g2_o21ai_1 _15985_ (.B1(_07461_),
    .Y(_07462_),
    .A1(_05982_),
    .A2(_04358_));
 sg13g2_mux2_1 _15986_ (.A0(_05306_),
    .A1(_07462_),
    .S(_07188_),
    .X(_07463_));
 sg13g2_and2_1 _15987_ (.A(net427),
    .B(_07463_),
    .X(_00995_));
 sg13g2_and2_1 _15988_ (.A(net536),
    .B(_05286_),
    .X(_07464_));
 sg13g2_a21oi_1 _15989_ (.A1(_07179_),
    .A2(_05306_),
    .Y(_07465_),
    .B1(_07464_));
 sg13g2_nand2_1 _15990_ (.Y(_07466_),
    .A(net605),
    .B(net380));
 sg13g2_o21ai_1 _15991_ (.B1(_07466_),
    .Y(_07467_),
    .A1(net348),
    .A2(_07465_));
 sg13g2_mux2_1 _15992_ (.A0(_05311_),
    .A1(_07467_),
    .S(_07188_),
    .X(_07468_));
 sg13g2_and2_1 _15993_ (.A(net427),
    .B(_07468_),
    .X(_00996_));
 sg13g2_mux2_1 _15994_ (.A0(_07350_),
    .A1(_06046_),
    .S(net534),
    .X(_07469_));
 sg13g2_and2_1 _15995_ (.A(_07141_),
    .B(_05293_),
    .X(_07470_));
 sg13g2_a21oi_1 _15996_ (.A1(_07178_),
    .A2(_05311_),
    .Y(_07471_),
    .B1(_07470_));
 sg13g2_nor2_1 _15997_ (.A(net412),
    .B(_07471_),
    .Y(_07472_));
 sg13g2_a21oi_1 _15998_ (.A1(net348),
    .A2(_07469_),
    .Y(_07473_),
    .B1(_07472_));
 sg13g2_nor2_1 _15999_ (.A(net311),
    .B(_07473_),
    .Y(_07474_));
 sg13g2_a21oi_1 _16000_ (.A1(_05237_),
    .A2(net312),
    .Y(_07475_),
    .B1(_07474_));
 sg13g2_nor2_1 _16001_ (.A(_07252_),
    .B(_07475_),
    .Y(_00997_));
 sg13g2_nor2b_1 _16002_ (.A(_07143_),
    .B_N(_05237_),
    .Y(_07476_));
 sg13g2_a221oi_1 _16003_ (.B2(_04309_),
    .C1(_07476_),
    .B1(_04308_),
    .A1(_07228_),
    .Y(_07477_),
    .A2(_05298_));
 sg13g2_nand2_1 _16004_ (.Y(_07478_),
    .A(net534),
    .B(_06049_));
 sg13g2_o21ai_1 _16005_ (.B1(_07478_),
    .Y(_07479_),
    .A1(net533),
    .A2(_07346_));
 sg13g2_nor2_1 _16006_ (.A(_04312_),
    .B(_07479_),
    .Y(_07480_));
 sg13g2_nor3_1 _16007_ (.A(_07193_),
    .B(_07477_),
    .C(_07480_),
    .Y(_07481_));
 sg13g2_a21oi_1 _16008_ (.A1(_05242_),
    .A2(net312),
    .Y(_07482_),
    .B1(_07481_));
 sg13g2_nor2_1 _16009_ (.A(net379),
    .B(_07482_),
    .Y(_00998_));
 sg13g2_buf_1 _16010_ (.A(_06002_),
    .X(_07483_));
 sg13g2_nand2b_1 _16011_ (.Y(_07484_),
    .B(_00051_),
    .A_N(sclk));
 sg13g2_nor4_1 _16012_ (.A(_04291_),
    .B(net426),
    .C(_04299_),
    .D(_07484_),
    .Y(_07485_));
 sg13g2_a21oi_1 _16013_ (.A1(_04291_),
    .A2(_07484_),
    .Y(_07486_),
    .B1(_07485_));
 sg13g2_nor2_1 _16014_ (.A(_07483_),
    .B(_07486_),
    .Y(_00999_));
 sg13g2_nor2_1 _16015_ (.A(_04350_),
    .B(_07148_),
    .Y(_07487_));
 sg13g2_nor2_1 _16016_ (.A(_04315_),
    .B(_07487_),
    .Y(_07488_));
 sg13g2_o21ai_1 _16017_ (.B1(net443),
    .Y(_07489_),
    .A1(_04342_),
    .A2(_07488_));
 sg13g2_nor2b_1 _16018_ (.A(_07185_),
    .B_N(_07489_),
    .Y(_07490_));
 sg13g2_buf_2 _16019_ (.A(_07490_),
    .X(_07491_));
 sg13g2_nor2b_1 _16020_ (.A(net516),
    .B_N(_00051_),
    .Y(_07492_));
 sg13g2_a21oi_1 _16021_ (.A1(_04347_),
    .A2(net516),
    .Y(_07493_),
    .B1(_07492_));
 sg13g2_or4_1 _16022_ (.A(_04291_),
    .B(\soc_I.qqspi_I.xfer_cycles[1] ),
    .C(_07491_),
    .D(_07493_),
    .X(_07494_));
 sg13g2_o21ai_1 _16023_ (.B1(\soc_I.qqspi_I.xfer_cycles[1] ),
    .Y(_07495_),
    .A1(_04291_),
    .A2(_07484_));
 sg13g2_a21oi_1 _16024_ (.A1(_07494_),
    .A2(_07495_),
    .Y(_01000_),
    .B1(_06963_));
 sg13g2_buf_1 _16025_ (.A(net515),
    .X(_07496_));
 sg13g2_xnor2_1 _16026_ (.Y(_07497_),
    .A(_04294_),
    .B(net517));
 sg13g2_nor3_1 _16027_ (.A(net460),
    .B(_00085_),
    .C(_04298_),
    .Y(_07498_));
 sg13g2_a221oi_1 _16028_ (.B2(net460),
    .C1(_07498_),
    .B1(_07497_),
    .A1(_07145_),
    .Y(_07499_),
    .A2(net380));
 sg13g2_mux2_1 _16029_ (.A0(_07499_),
    .A1(_04294_),
    .S(_07491_),
    .X(_07500_));
 sg13g2_and2_1 _16030_ (.A(_07496_),
    .B(_07500_),
    .X(_01001_));
 sg13g2_inv_1 _16031_ (.Y(_07501_),
    .A(_04294_));
 sg13g2_o21ai_1 _16032_ (.B1(_07501_),
    .Y(_07502_),
    .A1(_07141_),
    .A2(net517));
 sg13g2_and3_1 _16033_ (.X(_07503_),
    .A(_01840_),
    .B(_07220_),
    .C(_07345_));
 sg13g2_nor4_1 _16034_ (.A(_04350_),
    .B(_04344_),
    .C(net358),
    .D(_07503_),
    .Y(_07504_));
 sg13g2_or4_1 _16035_ (.A(_04293_),
    .B(_07491_),
    .C(_07502_),
    .D(_07504_),
    .X(_07505_));
 sg13g2_o21ai_1 _16036_ (.B1(_04293_),
    .Y(_07506_),
    .A1(_07491_),
    .A2(_07502_));
 sg13g2_buf_1 _16037_ (.A(_04267_),
    .X(_07507_));
 sg13g2_a21oi_1 _16038_ (.A1(_07505_),
    .A2(_07506_),
    .Y(_01002_),
    .B1(net377));
 sg13g2_or2_1 _16039_ (.X(_07508_),
    .B(_07502_),
    .A(_04293_));
 sg13g2_nor2_1 _16040_ (.A(\soc_I.qqspi_I.xfer_cycles[4] ),
    .B(_07508_),
    .Y(_07509_));
 sg13g2_nand3_1 _16041_ (.B(_07220_),
    .C(_07345_),
    .A(_05996_),
    .Y(_07510_));
 sg13g2_o21ai_1 _16042_ (.B1(net443),
    .Y(_07511_),
    .A1(_04350_),
    .A2(_07148_));
 sg13g2_a21oi_1 _16043_ (.A1(_07162_),
    .A2(_07510_),
    .Y(_07512_),
    .B1(_07511_));
 sg13g2_a21o_1 _16044_ (.A2(_07509_),
    .A1(net334),
    .B1(_07512_),
    .X(_07513_));
 sg13g2_nand3b_1 _16045_ (.B(_07513_),
    .C(net518),
    .Y(_07514_),
    .A_N(_07491_));
 sg13g2_and2_1 _16046_ (.A(\soc_I.qqspi_I.xfer_cycles[4] ),
    .B(net596),
    .X(_07515_));
 sg13g2_o21ai_1 _16047_ (.B1(_07515_),
    .Y(_07516_),
    .A1(_07491_),
    .A2(_07508_));
 sg13g2_nand2_1 _16048_ (.Y(_01003_),
    .A(_07514_),
    .B(_07516_));
 sg13g2_inv_1 _16049_ (.Y(_07517_),
    .A(_07509_));
 sg13g2_nor3_1 _16050_ (.A(\soc_I.qqspi_I.xfer_cycles[5] ),
    .B(net361),
    .C(_07517_),
    .Y(_07518_));
 sg13g2_nor3_1 _16051_ (.A(_00082_),
    .B(_07345_),
    .C(_07511_),
    .Y(_07519_));
 sg13g2_o21ai_1 _16052_ (.B1(_04371_),
    .Y(_07520_),
    .A1(_07518_),
    .A2(_07519_));
 sg13g2_and2_1 _16053_ (.A(\soc_I.qqspi_I.xfer_cycles[5] ),
    .B(net596),
    .X(_07521_));
 sg13g2_o21ai_1 _16054_ (.B1(_07521_),
    .Y(_07522_),
    .A1(_07491_),
    .A2(_07517_));
 sg13g2_o21ai_1 _16055_ (.B1(_07522_),
    .Y(_01004_),
    .A1(_07491_),
    .A2(_07520_));
 sg13g2_inv_1 _16056_ (.Y(_07523_),
    .A(net1));
 sg13g2_buf_1 _16057_ (.A(\soc_I.rst_cnt[0] ),
    .X(_07524_));
 sg13g2_nor2b_1 _16058_ (.A(net596),
    .B_N(_07524_),
    .Y(_07525_));
 sg13g2_nor2_1 _16059_ (.A(net438),
    .B(_07524_),
    .Y(_07526_));
 sg13g2_nor3_1 _16060_ (.A(_07523_),
    .B(_07525_),
    .C(_07526_),
    .Y(_01005_));
 sg13g2_xnor2_1 _16061_ (.Y(_07527_),
    .A(\soc_I.rst_cnt[1] ),
    .B(_07525_));
 sg13g2_nor2_1 _16062_ (.A(_07523_),
    .B(_07527_),
    .Y(_01006_));
 sg13g2_nand3_1 _16063_ (.B(_07524_),
    .C(\soc_I.rst_cnt[1] ),
    .A(net520),
    .Y(_07528_));
 sg13g2_xor2_1 _16064_ (.B(_07528_),
    .A(\soc_I.rst_cnt[2] ),
    .X(_07529_));
 sg13g2_nor2_1 _16065_ (.A(_07523_),
    .B(_07529_),
    .Y(_01007_));
 sg13g2_nand3_1 _16066_ (.B(\soc_I.rst_cnt[1] ),
    .C(\soc_I.rst_cnt[2] ),
    .A(_07524_),
    .Y(_07530_));
 sg13g2_a21oi_1 _16067_ (.A1(net398),
    .A2(_07530_),
    .Y(_01008_),
    .B1(_07523_));
 sg13g2_nand2_1 _16068_ (.Y(_07531_),
    .A(_00088_),
    .B(_05416_));
 sg13g2_o21ai_1 _16069_ (.B1(_05419_),
    .Y(_07532_),
    .A1(net580),
    .A2(_05415_));
 sg13g2_a21oi_1 _16070_ (.A1(_07531_),
    .A2(_07532_),
    .Y(_01009_),
    .B1(net377));
 sg13g2_inv_1 _16071_ (.Y(_07533_),
    .A(_05418_));
 sg13g2_nand2_1 _16072_ (.Y(_07534_),
    .A(_05419_),
    .B(_05416_));
 sg13g2_xnor2_1 _16073_ (.Y(_07535_),
    .A(_07533_),
    .B(_07534_));
 sg13g2_nor2_1 _16074_ (.A(net378),
    .B(_07535_),
    .Y(_01010_));
 sg13g2_nor3_1 _16075_ (.A(net580),
    .B(_05415_),
    .C(_05420_),
    .Y(_07536_));
 sg13g2_xnor2_1 _16076_ (.Y(_07537_),
    .A(_05410_),
    .B(_07536_));
 sg13g2_nor2_1 _16077_ (.A(net378),
    .B(_07537_),
    .Y(_01011_));
 sg13g2_xnor2_1 _16078_ (.Y(_07538_),
    .A(_00084_),
    .B(net442));
 sg13g2_and2_1 _16079_ (.A(_05799_),
    .B(_07538_),
    .X(_07539_));
 sg13g2_inv_1 _16080_ (.Y(_07540_),
    .A(_05793_));
 sg13g2_and2_1 _16081_ (.A(_00084_),
    .B(net442),
    .X(_07541_));
 sg13g2_a221oi_1 _16082_ (.B2(_07540_),
    .C1(_07541_),
    .B1(_06628_),
    .A1(_05341_),
    .Y(_07542_),
    .A2(_05345_));
 sg13g2_nor3_1 _16083_ (.A(net383),
    .B(_07539_),
    .C(_07542_),
    .Y(_01012_));
 sg13g2_nor2_1 _16084_ (.A(_05341_),
    .B(_05379_),
    .Y(_07543_));
 sg13g2_and3_1 _16085_ (.X(_07544_),
    .A(_05793_),
    .B(_05341_),
    .C(_05344_));
 sg13g2_a21oi_1 _16086_ (.A1(_05799_),
    .A2(_07543_),
    .Y(_07545_),
    .B1(_07544_));
 sg13g2_xor2_1 _16087_ (.B(_07545_),
    .A(_05340_),
    .X(_07546_));
 sg13g2_nor2_1 _16088_ (.A(_07483_),
    .B(_07546_),
    .Y(_01013_));
 sg13g2_nand3b_1 _16089_ (.B(_05799_),
    .C(_07543_),
    .Y(_07547_),
    .A_N(_05340_));
 sg13g2_buf_1 _16090_ (.A(_07547_),
    .X(_07548_));
 sg13g2_nand4_1 _16091_ (.B(_05340_),
    .C(_05341_),
    .A(_05793_),
    .Y(_07549_),
    .D(_05344_));
 sg13g2_buf_1 _16092_ (.A(_07549_),
    .X(_07550_));
 sg13g2_a21o_1 _16093_ (.A2(_07550_),
    .A1(_07548_),
    .B1(_05342_),
    .X(_07551_));
 sg13g2_nand3_1 _16094_ (.B(_07548_),
    .C(_07550_),
    .A(_05342_),
    .Y(_07552_));
 sg13g2_a21oi_1 _16095_ (.A1(_07551_),
    .A2(_07552_),
    .Y(_01014_),
    .B1(net377));
 sg13g2_inv_1 _16096_ (.Y(_07553_),
    .A(_07550_));
 sg13g2_nand2_1 _16097_ (.Y(_07554_),
    .A(_05342_),
    .B(_07553_));
 sg13g2_o21ai_1 _16098_ (.B1(_07554_),
    .Y(_07555_),
    .A1(_05342_),
    .A2(_07548_));
 sg13g2_xnor2_1 _16099_ (.Y(_07556_),
    .A(\soc_I.rx_uart_i.fifo_i.cnt[3] ),
    .B(_07555_));
 sg13g2_nor2_1 _16100_ (.A(net378),
    .B(_07556_),
    .Y(_01015_));
 sg13g2_nand2_1 _16101_ (.Y(_07557_),
    .A(_07540_),
    .B(_05343_));
 sg13g2_nand3_1 _16102_ (.B(_05342_),
    .C(_07553_),
    .A(\soc_I.rx_uart_i.fifo_i.cnt[3] ),
    .Y(_07558_));
 sg13g2_nand3_1 _16103_ (.B(_07557_),
    .C(_07558_),
    .A(_05339_),
    .Y(_07559_));
 sg13g2_or2_1 _16104_ (.X(_07560_),
    .B(_07558_),
    .A(_05339_));
 sg13g2_a21oi_1 _16105_ (.A1(_07559_),
    .A2(_07560_),
    .Y(_01016_),
    .B1(net377));
 sg13g2_nand2_1 _16106_ (.Y(_07561_),
    .A(_00090_),
    .B(_05799_));
 sg13g2_a21oi_1 _16107_ (.A1(_05797_),
    .A2(_07561_),
    .Y(_01145_),
    .B1(net377));
 sg13g2_nand2_1 _16108_ (.Y(_07562_),
    .A(_00089_),
    .B(net442));
 sg13g2_nand2_1 _16109_ (.Y(_07563_),
    .A(_05350_),
    .B(_05347_));
 sg13g2_a21oi_1 _16110_ (.A1(_07562_),
    .A2(_07563_),
    .Y(_01146_),
    .B1(_07507_));
 sg13g2_nand2_1 _16111_ (.Y(_07564_),
    .A(_05350_),
    .B(net442));
 sg13g2_xor2_1 _16112_ (.B(_07564_),
    .A(_05349_),
    .X(_07565_));
 sg13g2_nor2_1 _16113_ (.A(net378),
    .B(_07565_),
    .Y(_01147_));
 sg13g2_nor2_1 _16114_ (.A(_05347_),
    .B(_05375_),
    .Y(_07566_));
 sg13g2_xnor2_1 _16115_ (.Y(_07567_),
    .A(net613),
    .B(_07566_));
 sg13g2_nor2_1 _16116_ (.A(net378),
    .B(_07567_),
    .Y(_01148_));
 sg13g2_o21ai_1 _16117_ (.B1(net614),
    .Y(_07568_),
    .A1(_05375_),
    .A2(_05396_));
 sg13g2_nor2b_1 _16118_ (.A(net331),
    .B_N(_07568_),
    .Y(_07569_));
 sg13g2_nor2_1 _16119_ (.A(net378),
    .B(_07569_),
    .Y(_01149_));
 sg13g2_buf_2 _16120_ (.A(\soc_I.rx_uart_i.state[2] ),
    .X(_07570_));
 sg13g2_nand2_1 _16121_ (.Y(_07571_),
    .A(net612),
    .B(_05421_));
 sg13g2_o21ai_1 _16122_ (.B1(_05344_),
    .Y(_07572_),
    .A1(_07570_),
    .A2(_07571_));
 sg13g2_nand2_1 _16123_ (.Y(_07573_),
    .A(_07570_),
    .B(_05421_));
 sg13g2_buf_1 _16124_ (.A(_07573_),
    .X(_07574_));
 sg13g2_buf_1 _16125_ (.A(net424),
    .X(_07575_));
 sg13g2_buf_1 _16126_ (.A(\soc_I.rx_uart_i.wait_states[9] ),
    .X(_07576_));
 sg13g2_nor4_1 _16127_ (.A(_07576_),
    .B(\soc_I.rx_uart_i.wait_states[11] ),
    .C(\soc_I.rx_uart_i.wait_states[10] ),
    .D(\soc_I.rx_uart_i.wait_states[13] ),
    .Y(_07577_));
 sg13g2_buf_1 _16128_ (.A(\soc_I.rx_uart_i.wait_states[7] ),
    .X(_07578_));
 sg13g2_buf_1 _16129_ (.A(\soc_I.rx_uart_i.wait_states[6] ),
    .X(_07579_));
 sg13g2_nor4_1 _16130_ (.A(\soc_I.rx_uart_i.wait_states[4] ),
    .B(_07578_),
    .C(_07579_),
    .D(\soc_I.rx_uart_i.wait_states[8] ),
    .Y(_07580_));
 sg13g2_nor2b_1 _16131_ (.A(\soc_I.rx_uart_i.wait_states[5] ),
    .B_N(_07580_),
    .Y(_07581_));
 sg13g2_buf_1 _16132_ (.A(\soc_I.rx_uart_i.wait_states[14] ),
    .X(_07582_));
 sg13g2_inv_1 _16133_ (.Y(_07583_),
    .A(_00054_));
 sg13g2_nor4_1 _16134_ (.A(\soc_I.rx_uart_i.wait_states[12] ),
    .B(\soc_I.rx_uart_i.wait_states[15] ),
    .C(_07582_),
    .D(_07583_),
    .Y(_07584_));
 sg13g2_buf_1 _16135_ (.A(\soc_I.rx_uart_i.wait_states[0] ),
    .X(_07585_));
 sg13g2_inv_1 _16136_ (.Y(_07586_),
    .A(_07585_));
 sg13g2_buf_1 _16137_ (.A(\soc_I.rx_uart_i.wait_states[1] ),
    .X(_07587_));
 sg13g2_buf_1 _16138_ (.A(\soc_I.rx_uart_i.wait_states[3] ),
    .X(_07588_));
 sg13g2_nor4_1 _16139_ (.A(_07586_),
    .B(_07587_),
    .C(_07588_),
    .D(\soc_I.rx_uart_i.wait_states[2] ),
    .Y(_07589_));
 sg13g2_nand4_1 _16140_ (.B(_07581_),
    .C(_07584_),
    .A(_07577_),
    .Y(_07590_),
    .D(_07589_));
 sg13g2_or4_1 _16141_ (.A(\soc_I.rx_uart_i.return_state[1] ),
    .B(\soc_I.rx_uart_i.return_state[0] ),
    .C(net376),
    .D(_07590_),
    .X(_07591_));
 sg13g2_a21oi_1 _16142_ (.A1(_07572_),
    .A2(_07591_),
    .Y(_01150_),
    .B1(_07507_));
 sg13g2_inv_1 _16143_ (.Y(_07592_),
    .A(_05419_));
 sg13g2_nor3_2 _16144_ (.A(net580),
    .B(_05410_),
    .C(_05415_),
    .Y(_07593_));
 sg13g2_and3_1 _16145_ (.X(_07594_),
    .A(_07533_),
    .B(_07592_),
    .C(_07593_));
 sg13g2_nand2_1 _16146_ (.Y(_07595_),
    .A(_00088_),
    .B(_07594_));
 sg13g2_a22oi_1 _16147_ (.Y(_07596_),
    .B1(_07595_),
    .B2(_05336_),
    .A2(_07594_),
    .A1(net611));
 sg13g2_nor2_1 _16148_ (.A(net378),
    .B(_07596_),
    .Y(_01153_));
 sg13g2_nand3_1 _16149_ (.B(_05419_),
    .C(_07593_),
    .A(_07533_),
    .Y(_07597_));
 sg13g2_mux2_1 _16150_ (.A0(net611),
    .A1(_05354_),
    .S(_07597_),
    .X(_07598_));
 sg13g2_and2_1 _16151_ (.A(net425),
    .B(_07598_),
    .X(_01154_));
 sg13g2_nand3_1 _16152_ (.B(_07592_),
    .C(_07593_),
    .A(_05418_),
    .Y(_07599_));
 sg13g2_nand2_1 _16153_ (.Y(_07600_),
    .A(_05355_),
    .B(_07599_));
 sg13g2_o21ai_1 _16154_ (.B1(_07600_),
    .Y(_07601_),
    .A1(_00059_),
    .A2(_07599_));
 sg13g2_and2_1 _16155_ (.A(net425),
    .B(_07601_),
    .X(_01155_));
 sg13g2_nand2b_1 _16156_ (.Y(_07602_),
    .B(_07593_),
    .A_N(_05420_));
 sg13g2_mux2_1 _16157_ (.A0(net611),
    .A1(_05356_),
    .S(_07602_),
    .X(_07603_));
 sg13g2_and2_1 _16158_ (.A(net425),
    .B(_07603_),
    .X(_01156_));
 sg13g2_inv_1 _16159_ (.Y(_07604_),
    .A(_00059_));
 sg13g2_nor3_1 _16160_ (.A(_05418_),
    .B(_05419_),
    .C(_05417_),
    .Y(_07605_));
 sg13g2_mux2_1 _16161_ (.A0(_05357_),
    .A1(_07604_),
    .S(_07605_),
    .X(_07606_));
 sg13g2_and2_1 _16162_ (.A(net425),
    .B(_07606_),
    .X(_01157_));
 sg13g2_nor3_1 _16163_ (.A(_05418_),
    .B(_07592_),
    .C(_05417_),
    .Y(_07607_));
 sg13g2_mux2_1 _16164_ (.A0(_05358_),
    .A1(net611),
    .S(_07607_),
    .X(_07608_));
 sg13g2_and2_1 _16165_ (.A(net425),
    .B(_07608_),
    .X(_01158_));
 sg13g2_nor3_1 _16166_ (.A(_07533_),
    .B(_05419_),
    .C(_05417_),
    .Y(_07609_));
 sg13g2_mux2_1 _16167_ (.A0(_05359_),
    .A1(_07604_),
    .S(_07609_),
    .X(_07610_));
 sg13g2_and2_1 _16168_ (.A(net425),
    .B(_07610_),
    .X(_01159_));
 sg13g2_nor2_1 _16169_ (.A(_05417_),
    .B(_05420_),
    .Y(_07611_));
 sg13g2_mux2_1 _16170_ (.A0(_05360_),
    .A1(net611),
    .S(_07611_),
    .X(_07612_));
 sg13g2_and2_1 _16171_ (.A(net425),
    .B(_07612_),
    .X(_01160_));
 sg13g2_and2_1 _16172_ (.A(_07496_),
    .B(net3),
    .X(_01161_));
 sg13g2_and2_1 _16173_ (.A(net425),
    .B(\soc_I.rx_uart_i.rx_in_sync[0] ),
    .X(_01162_));
 sg13g2_buf_1 _16174_ (.A(net515),
    .X(_07613_));
 sg13g2_and2_1 _16175_ (.A(net423),
    .B(\soc_I.rx_uart_i.rx_in_sync[1] ),
    .X(_01163_));
 sg13g2_nor2_2 _16176_ (.A(_05429_),
    .B(_07571_),
    .Y(_07614_));
 sg13g2_nor4_1 _16177_ (.A(net520),
    .B(net376),
    .C(_07590_),
    .D(_07614_),
    .Y(_07615_));
 sg13g2_and2_1 _16178_ (.A(\soc_I.rx_uart_i.return_state[0] ),
    .B(_07615_),
    .X(_01164_));
 sg13g2_and2_1 _16179_ (.A(\soc_I.rx_uart_i.return_state[1] ),
    .B(_07615_),
    .X(_01165_));
 sg13g2_inv_1 _16180_ (.Y(_07616_),
    .A(_05413_));
 sg13g2_nand2_1 _16181_ (.Y(_07617_),
    .A(net580),
    .B(net612));
 sg13g2_nand2b_1 _16182_ (.Y(_07618_),
    .B(_07590_),
    .A_N(net580));
 sg13g2_o21ai_1 _16183_ (.B1(_07618_),
    .Y(_07619_),
    .A1(_05427_),
    .A2(_07617_));
 sg13g2_nand4_1 _16184_ (.B(net580),
    .C(_05414_),
    .A(_05413_),
    .Y(_07620_),
    .D(_05427_));
 sg13g2_o21ai_1 _16185_ (.B1(_07620_),
    .Y(_07621_),
    .A1(_05412_),
    .A2(_07570_));
 sg13g2_a21oi_1 _16186_ (.A1(_07616_),
    .A2(_07619_),
    .Y(_07622_),
    .B1(_07621_));
 sg13g2_nor2_1 _16187_ (.A(_07614_),
    .B(_07622_),
    .Y(_07623_));
 sg13g2_a21oi_1 _16188_ (.A1(_07570_),
    .A2(_07614_),
    .Y(_07624_),
    .B1(_07623_));
 sg13g2_nor2_1 _16189_ (.A(net378),
    .B(_07624_),
    .Y(_01166_));
 sg13g2_nor2_1 _16190_ (.A(net424),
    .B(_07614_),
    .Y(_07625_));
 sg13g2_nand2_1 _16191_ (.Y(_07626_),
    .A(_07586_),
    .B(_07625_));
 sg13g2_and2_1 _16192_ (.A(_07570_),
    .B(_05421_),
    .X(_07627_));
 sg13g2_buf_1 _16193_ (.A(_07627_),
    .X(_07628_));
 sg13g2_nor2_1 _16194_ (.A(net441),
    .B(_07628_),
    .Y(_07629_));
 sg13g2_buf_2 _16195_ (.A(_07629_),
    .X(_07630_));
 sg13g2_buf_1 _16196_ (.A(_07630_),
    .X(_07631_));
 sg13g2_a22oi_1 _16197_ (.Y(_07632_),
    .B1(net329),
    .B2(_05500_),
    .A2(net408),
    .A1(_05468_));
 sg13g2_and2_1 _16198_ (.A(_05411_),
    .B(net612),
    .X(_07633_));
 sg13g2_a21oi_1 _16199_ (.A1(_00059_),
    .A2(_07633_),
    .Y(_07634_),
    .B1(_07570_));
 sg13g2_nand2_1 _16200_ (.Y(_07635_),
    .A(_05413_),
    .B(_07634_));
 sg13g2_nor3_1 _16201_ (.A(_05411_),
    .B(net612),
    .C(_07570_),
    .Y(_07636_));
 sg13g2_a21oi_1 _16202_ (.A1(_07604_),
    .A2(_07633_),
    .Y(_07637_),
    .B1(_07636_));
 sg13g2_nand2_1 _16203_ (.Y(_07638_),
    .A(_07616_),
    .B(_07637_));
 sg13g2_a221oi_1 _16204_ (.B2(_07638_),
    .C1(_07614_),
    .B1(_07635_),
    .A1(_05411_),
    .Y(_07639_),
    .A2(_07570_));
 sg13g2_buf_1 _16205_ (.A(_07639_),
    .X(_07640_));
 sg13g2_buf_1 _16206_ (.A(_07640_),
    .X(_07641_));
 sg13g2_buf_1 _16207_ (.A(net328),
    .X(_07642_));
 sg13g2_mux2_1 _16208_ (.A0(_07586_),
    .A1(_07632_),
    .S(net317),
    .X(_07643_));
 sg13g2_nand3_1 _16209_ (.B(_07626_),
    .C(_07643_),
    .A(_05810_),
    .Y(_01167_));
 sg13g2_buf_1 _16210_ (.A(_06002_),
    .X(_07644_));
 sg13g2_buf_1 _16211_ (.A(net328),
    .X(_07645_));
 sg13g2_nor3_2 _16212_ (.A(_07585_),
    .B(_07587_),
    .C(\soc_I.rx_uart_i.wait_states[2] ),
    .Y(_07646_));
 sg13g2_nor2b_1 _16213_ (.A(_07588_),
    .B_N(_07646_),
    .Y(_07647_));
 sg13g2_and2_1 _16214_ (.A(_07581_),
    .B(_07647_),
    .X(_07648_));
 sg13g2_buf_1 _16215_ (.A(_07648_),
    .X(_07649_));
 sg13g2_nor2b_1 _16216_ (.A(_07576_),
    .B_N(_07649_),
    .Y(_07650_));
 sg13g2_nand2b_1 _16217_ (.Y(_07651_),
    .B(_07650_),
    .A_N(\soc_I.rx_uart_i.wait_states[10] ));
 sg13g2_a22oi_1 _16218_ (.Y(_07652_),
    .B1(net329),
    .B2(net608),
    .A2(net441),
    .A1(_05516_));
 sg13g2_o21ai_1 _16219_ (.B1(_07652_),
    .Y(_07653_),
    .A1(net376),
    .A2(_07651_));
 sg13g2_o21ai_1 _16220_ (.B1(net317),
    .Y(_07654_),
    .A1(net376),
    .A2(_07650_));
 sg13g2_a22oi_1 _16221_ (.Y(_07655_),
    .B1(_07654_),
    .B2(\soc_I.rx_uart_i.wait_states[10] ),
    .A2(_07653_),
    .A1(net316));
 sg13g2_nor2_1 _16222_ (.A(net375),
    .B(_07655_),
    .Y(_01168_));
 sg13g2_nor2_1 _16223_ (.A(\soc_I.rx_uart_i.wait_states[11] ),
    .B(_07651_),
    .Y(_07656_));
 sg13g2_inv_1 _16224_ (.Y(_07657_),
    .A(_07656_));
 sg13g2_a22oi_1 _16225_ (.Y(_07658_),
    .B1(net329),
    .B2(_05544_),
    .A2(net441),
    .A1(_05535_));
 sg13g2_o21ai_1 _16226_ (.B1(_07658_),
    .Y(_07659_),
    .A1(net424),
    .A2(_07657_));
 sg13g2_buf_1 _16227_ (.A(_07628_),
    .X(_07660_));
 sg13g2_inv_1 _16228_ (.Y(_07661_),
    .A(_07640_));
 sg13g2_a21o_1 _16229_ (.A2(_07651_),
    .A1(net374),
    .B1(_07661_),
    .X(_07662_));
 sg13g2_a22oi_1 _16230_ (.Y(_07663_),
    .B1(_07662_),
    .B2(\soc_I.rx_uart_i.wait_states[11] ),
    .A2(_07659_),
    .A1(net316));
 sg13g2_nor2_1 _16231_ (.A(net375),
    .B(_07663_),
    .Y(_01169_));
 sg13g2_nor2_1 _16232_ (.A(\soc_I.rx_uart_i.wait_states[12] ),
    .B(_07657_),
    .Y(_07664_));
 sg13g2_inv_1 _16233_ (.Y(_07665_),
    .A(_07664_));
 sg13g2_a22oi_1 _16234_ (.Y(_07666_),
    .B1(_07630_),
    .B2(_05560_),
    .A2(net441),
    .A1(_05544_));
 sg13g2_o21ai_1 _16235_ (.B1(_07666_),
    .Y(_07667_),
    .A1(net424),
    .A2(_07665_));
 sg13g2_o21ai_1 _16236_ (.B1(net328),
    .Y(_07668_),
    .A1(net376),
    .A2(_07656_));
 sg13g2_a22oi_1 _16237_ (.Y(_07669_),
    .B1(_07668_),
    .B2(\soc_I.rx_uart_i.wait_states[12] ),
    .A2(_07667_),
    .A1(net316));
 sg13g2_nor2_1 _16238_ (.A(net375),
    .B(_07669_),
    .Y(_01170_));
 sg13g2_nand2b_1 _16239_ (.Y(_07670_),
    .B(_07664_),
    .A_N(\soc_I.rx_uart_i.wait_states[13] ));
 sg13g2_buf_1 _16240_ (.A(_07670_),
    .X(_07671_));
 sg13g2_or2_1 _16241_ (.X(_07672_),
    .B(_07671_),
    .A(net424));
 sg13g2_a22oi_1 _16242_ (.Y(_07673_),
    .B1(net329),
    .B2(_05568_),
    .A2(net408),
    .A1(_05560_));
 sg13g2_nand2_1 _16243_ (.Y(_07674_),
    .A(_07672_),
    .B(_07673_));
 sg13g2_o21ai_1 _16244_ (.B1(net328),
    .Y(_07675_),
    .A1(net376),
    .A2(_07664_));
 sg13g2_a22oi_1 _16245_ (.Y(_07676_),
    .B1(_07675_),
    .B2(\soc_I.rx_uart_i.wait_states[13] ),
    .A2(_07674_),
    .A1(net316));
 sg13g2_nor2_1 _16246_ (.A(net375),
    .B(_07676_),
    .Y(_01171_));
 sg13g2_a21o_1 _16247_ (.A2(_07671_),
    .A1(net374),
    .B1(_07661_),
    .X(_07677_));
 sg13g2_a22oi_1 _16248_ (.Y(_07678_),
    .B1(net329),
    .B2(_05581_),
    .A2(_05424_),
    .A1(_05568_));
 sg13g2_o21ai_1 _16249_ (.B1(_07678_),
    .Y(_07679_),
    .A1(_07582_),
    .A2(_07672_));
 sg13g2_a22oi_1 _16250_ (.Y(_07680_),
    .B1(_07679_),
    .B2(net316),
    .A2(_07677_),
    .A1(_07582_));
 sg13g2_nor2_1 _16251_ (.A(net375),
    .B(_07680_),
    .Y(_01172_));
 sg13g2_nor3_1 _16252_ (.A(\soc_I.rx_uart_i.wait_states[15] ),
    .B(_07582_),
    .C(_07671_),
    .Y(_07681_));
 sg13g2_a22oi_1 _16253_ (.Y(_07682_),
    .B1(net374),
    .B2(_07681_),
    .A2(net408),
    .A1(_05581_));
 sg13g2_inv_1 _16254_ (.Y(_07683_),
    .A(_07682_));
 sg13g2_o21ai_1 _16255_ (.B1(net374),
    .Y(_07684_),
    .A1(_07582_),
    .A2(_07671_));
 sg13g2_nand2_1 _16256_ (.Y(_07685_),
    .A(net317),
    .B(_07684_));
 sg13g2_a22oi_1 _16257_ (.Y(_07686_),
    .B1(_07685_),
    .B2(\soc_I.rx_uart_i.wait_states[15] ),
    .A2(_07683_),
    .A1(net316));
 sg13g2_nor2_1 _16258_ (.A(net375),
    .B(_07686_),
    .Y(_01173_));
 sg13g2_xnor2_1 _16259_ (.Y(_07687_),
    .A(_00054_),
    .B(_07681_));
 sg13g2_a22oi_1 _16260_ (.Y(_07688_),
    .B1(_07687_),
    .B2(_07625_),
    .A2(_07661_),
    .A1(\soc_I.rx_uart_i.wait_states[16] ));
 sg13g2_nor2_1 _16261_ (.A(net375),
    .B(_07688_),
    .Y(_01174_));
 sg13g2_xnor2_1 _16262_ (.Y(_07689_),
    .A(_07585_),
    .B(_07587_));
 sg13g2_a22oi_1 _16263_ (.Y(_07690_),
    .B1(net374),
    .B2(_07689_),
    .A2(net408),
    .A1(_05500_));
 sg13g2_nand2_1 _16264_ (.Y(_07691_),
    .A(_05497_),
    .B(net329));
 sg13g2_nand3_1 _16265_ (.B(_07690_),
    .C(_07691_),
    .A(net317),
    .Y(_07692_));
 sg13g2_o21ai_1 _16266_ (.B1(_07692_),
    .Y(_07693_),
    .A1(_07587_),
    .A2(net317));
 sg13g2_nor2_1 _16267_ (.A(net375),
    .B(_07693_),
    .Y(_01175_));
 sg13g2_and2_1 _16268_ (.A(_07628_),
    .B(_07646_),
    .X(_07694_));
 sg13g2_a221oi_1 _16269_ (.B2(_05498_),
    .C1(_07694_),
    .B1(_07630_),
    .A1(_05497_),
    .Y(_07695_),
    .A2(_05423_));
 sg13g2_inv_1 _16270_ (.Y(_07696_),
    .A(_07695_));
 sg13g2_o21ai_1 _16271_ (.B1(net374),
    .Y(_07697_),
    .A1(_07585_),
    .A2(_07587_));
 sg13g2_nand2_1 _16272_ (.Y(_07698_),
    .A(net317),
    .B(_07697_));
 sg13g2_a22oi_1 _16273_ (.Y(_07699_),
    .B1(_07698_),
    .B2(\soc_I.rx_uart_i.wait_states[2] ),
    .A2(_07696_),
    .A1(net316));
 sg13g2_nor2_1 _16274_ (.A(_07644_),
    .B(_07699_),
    .Y(_01176_));
 sg13g2_o21ai_1 _16275_ (.B1(net328),
    .Y(_07700_),
    .A1(net424),
    .A2(_07646_));
 sg13g2_nand2_1 _16276_ (.Y(_07701_),
    .A(_07660_),
    .B(_07646_));
 sg13g2_a22oi_1 _16277_ (.Y(_07702_),
    .B1(_07631_),
    .B2(_05491_),
    .A2(net408),
    .A1(_05498_));
 sg13g2_o21ai_1 _16278_ (.B1(_07702_),
    .Y(_07703_),
    .A1(_07588_),
    .A2(_07701_));
 sg13g2_a22oi_1 _16279_ (.Y(_07704_),
    .B1(_07703_),
    .B2(_07645_),
    .A2(_07700_),
    .A1(_07588_));
 sg13g2_nor2_1 _16280_ (.A(_07644_),
    .B(_07704_),
    .Y(_01177_));
 sg13g2_nand2b_1 _16281_ (.Y(_07705_),
    .B(_07647_),
    .A_N(\soc_I.rx_uart_i.wait_states[4] ));
 sg13g2_a22oi_1 _16282_ (.Y(_07706_),
    .B1(_07630_),
    .B2(_05492_),
    .A2(net441),
    .A1(_05491_));
 sg13g2_o21ai_1 _16283_ (.B1(_07706_),
    .Y(_07707_),
    .A1(net424),
    .A2(_07705_));
 sg13g2_o21ai_1 _16284_ (.B1(net328),
    .Y(_07708_),
    .A1(net376),
    .A2(_07647_));
 sg13g2_a22oi_1 _16285_ (.Y(_07709_),
    .B1(_07708_),
    .B2(\soc_I.rx_uart_i.wait_states[4] ),
    .A2(_07707_),
    .A1(_07645_));
 sg13g2_nor2_1 _16286_ (.A(net404),
    .B(_07709_),
    .Y(_01178_));
 sg13g2_nor2_1 _16287_ (.A(\soc_I.rx_uart_i.wait_states[5] ),
    .B(_07705_),
    .Y(_07710_));
 sg13g2_inv_1 _16288_ (.Y(_07711_),
    .A(_07710_));
 sg13g2_a22oi_1 _16289_ (.Y(_07712_),
    .B1(_07630_),
    .B2(_05485_),
    .A2(net441),
    .A1(_05492_));
 sg13g2_o21ai_1 _16290_ (.B1(_07712_),
    .Y(_07713_),
    .A1(net424),
    .A2(_07711_));
 sg13g2_a21o_1 _16291_ (.A2(_07705_),
    .A1(net374),
    .B1(_07661_),
    .X(_07714_));
 sg13g2_a22oi_1 _16292_ (.Y(_07715_),
    .B1(_07714_),
    .B2(\soc_I.rx_uart_i.wait_states[5] ),
    .A2(_07713_),
    .A1(net317));
 sg13g2_nor2_1 _16293_ (.A(net404),
    .B(_07715_),
    .Y(_01179_));
 sg13g2_nor2_1 _16294_ (.A(_07579_),
    .B(_07711_),
    .Y(_07716_));
 sg13g2_nand2_1 _16295_ (.Y(_07717_),
    .A(net374),
    .B(_07716_));
 sg13g2_a22oi_1 _16296_ (.Y(_07718_),
    .B1(net329),
    .B2(_05486_),
    .A2(net408),
    .A1(_05485_));
 sg13g2_nand2_1 _16297_ (.Y(_07719_),
    .A(_07717_),
    .B(_07718_));
 sg13g2_o21ai_1 _16298_ (.B1(net328),
    .Y(_07720_),
    .A1(net376),
    .A2(_07710_));
 sg13g2_a22oi_1 _16299_ (.Y(_07721_),
    .B1(_07720_),
    .B2(_07579_),
    .A2(_07719_),
    .A1(net317));
 sg13g2_nor2_1 _16300_ (.A(net404),
    .B(_07721_),
    .Y(_01180_));
 sg13g2_a22oi_1 _16301_ (.Y(_07722_),
    .B1(_07630_),
    .B2(_05479_),
    .A2(net441),
    .A1(_05486_));
 sg13g2_o21ai_1 _16302_ (.B1(_07722_),
    .Y(_07723_),
    .A1(_07578_),
    .A2(_07717_));
 sg13g2_o21ai_1 _16303_ (.B1(_07641_),
    .Y(_07724_),
    .A1(_07575_),
    .A2(_07716_));
 sg13g2_a22oi_1 _16304_ (.Y(_07725_),
    .B1(_07724_),
    .B2(_07578_),
    .A2(_07723_),
    .A1(_07642_));
 sg13g2_nor2_1 _16305_ (.A(net404),
    .B(_07725_),
    .Y(_01181_));
 sg13g2_nand2_1 _16306_ (.Y(_07726_),
    .A(_07660_),
    .B(_07649_));
 sg13g2_a22oi_1 _16307_ (.Y(_07727_),
    .B1(net329),
    .B2(_05480_),
    .A2(_05424_),
    .A1(_05479_));
 sg13g2_nand2_1 _16308_ (.Y(_07728_),
    .A(_07726_),
    .B(_07727_));
 sg13g2_nor3_1 _16309_ (.A(_07578_),
    .B(_07579_),
    .C(_07711_),
    .Y(_07729_));
 sg13g2_o21ai_1 _16310_ (.B1(_07641_),
    .Y(_07730_),
    .A1(_07575_),
    .A2(_07729_));
 sg13g2_a22oi_1 _16311_ (.Y(_07731_),
    .B1(_07730_),
    .B2(\soc_I.rx_uart_i.wait_states[8] ),
    .A2(_07728_),
    .A1(_07642_));
 sg13g2_nor2_1 _16312_ (.A(net404),
    .B(_07731_),
    .Y(_01182_));
 sg13g2_o21ai_1 _16313_ (.B1(net328),
    .Y(_07732_),
    .A1(_07574_),
    .A2(_07649_));
 sg13g2_a22oi_1 _16314_ (.Y(_07733_),
    .B1(_07631_),
    .B2(_05516_),
    .A2(net408),
    .A1(_05480_));
 sg13g2_o21ai_1 _16315_ (.B1(_07733_),
    .Y(_07734_),
    .A1(_07576_),
    .A2(_07726_));
 sg13g2_a22oi_1 _16316_ (.Y(_07735_),
    .B1(_07734_),
    .B2(net316),
    .A2(_07732_),
    .A1(_07576_));
 sg13g2_nor2_1 _16317_ (.A(net404),
    .B(_07735_),
    .Y(_01183_));
 sg13g2_and4_1 _16318_ (.A(net433),
    .B(_03854_),
    .C(_04213_),
    .D(_05912_),
    .X(_01184_));
 sg13g2_buf_1 _16319_ (.A(\soc_I.spi0_I.state ),
    .X(_07736_));
 sg13g2_buf_1 _16320_ (.A(_07736_),
    .X(_07737_));
 sg13g2_buf_1 _16321_ (.A(_05751_),
    .X(_07738_));
 sg13g2_o21ai_1 _16322_ (.B1(\soc_I.spi0_I.ready_xfer ),
    .Y(_07739_),
    .A1(net532),
    .A2(net345));
 sg13g2_nor2_2 _16323_ (.A(_07736_),
    .B(_05751_),
    .Y(_07740_));
 sg13g2_and4_1 _16324_ (.A(net76),
    .B(_04099_),
    .C(_06557_),
    .D(_04213_),
    .X(_07741_));
 sg13g2_buf_1 _16325_ (.A(_07741_),
    .X(_07742_));
 sg13g2_nand2_1 _16326_ (.Y(_07743_),
    .A(_07740_),
    .B(_07742_));
 sg13g2_a21oi_1 _16327_ (.A1(_07739_),
    .A2(_07743_),
    .Y(_01185_),
    .B1(net377));
 sg13g2_buf_1 _16328_ (.A(net388),
    .X(_07744_));
 sg13g2_nand3_1 _16329_ (.B(\soc_I.spi0_I.spi_buf[0] ),
    .C(net344),
    .A(net532),
    .Y(_07745_));
 sg13g2_nand2_1 _16330_ (.Y(_07746_),
    .A(_07736_),
    .B(net388));
 sg13g2_buf_2 _16331_ (.A(_07746_),
    .X(_07747_));
 sg13g2_nand2_1 _16332_ (.Y(_07748_),
    .A(\soc_I.spi0_I.rx_data[0] ),
    .B(_07747_));
 sg13g2_a21oi_1 _16333_ (.A1(_07745_),
    .A2(_07748_),
    .Y(_01186_),
    .B1(net377));
 sg13g2_nand3_1 _16334_ (.B(\soc_I.spi0_I.spi_buf[1] ),
    .C(_07744_),
    .A(net532),
    .Y(_07749_));
 sg13g2_nand2_1 _16335_ (.Y(_07750_),
    .A(\soc_I.spi0_I.rx_data[1] ),
    .B(_07747_));
 sg13g2_a21oi_1 _16336_ (.A1(_07749_),
    .A2(_07750_),
    .Y(_01187_),
    .B1(net377));
 sg13g2_nand3_1 _16337_ (.B(\soc_I.spi0_I.spi_buf[2] ),
    .C(net344),
    .A(net532),
    .Y(_07751_));
 sg13g2_nand2_1 _16338_ (.Y(_07752_),
    .A(\soc_I.spi0_I.rx_data[2] ),
    .B(_07747_));
 sg13g2_buf_1 _16339_ (.A(_04267_),
    .X(_07753_));
 sg13g2_a21oi_1 _16340_ (.A1(_07751_),
    .A2(_07752_),
    .Y(_01188_),
    .B1(net373));
 sg13g2_nand3_1 _16341_ (.B(\soc_I.spi0_I.spi_buf[3] ),
    .C(net344),
    .A(net532),
    .Y(_07754_));
 sg13g2_nand2_1 _16342_ (.Y(_07755_),
    .A(\soc_I.spi0_I.rx_data[3] ),
    .B(_07747_));
 sg13g2_a21oi_1 _16343_ (.A1(_07754_),
    .A2(_07755_),
    .Y(_01189_),
    .B1(net373));
 sg13g2_nand3_1 _16344_ (.B(\soc_I.spi0_I.spi_buf[4] ),
    .C(_07744_),
    .A(_07737_),
    .Y(_07756_));
 sg13g2_nand2_1 _16345_ (.Y(_07757_),
    .A(\soc_I.spi0_I.rx_data[4] ),
    .B(_07747_));
 sg13g2_a21oi_1 _16346_ (.A1(_07756_),
    .A2(_07757_),
    .Y(_01190_),
    .B1(net373));
 sg13g2_nand3_1 _16347_ (.B(\soc_I.spi0_I.spi_buf[5] ),
    .C(net344),
    .A(net532),
    .Y(_07758_));
 sg13g2_nand2_1 _16348_ (.Y(_07759_),
    .A(\soc_I.spi0_I.rx_data[5] ),
    .B(_07747_));
 sg13g2_a21oi_1 _16349_ (.A1(_07758_),
    .A2(_07759_),
    .Y(_01191_),
    .B1(net373));
 sg13g2_nand3_1 _16350_ (.B(\soc_I.spi0_I.spi_buf[6] ),
    .C(net344),
    .A(net532),
    .Y(_07760_));
 sg13g2_nand2_1 _16351_ (.Y(_07761_),
    .A(\soc_I.spi0_I.rx_data[6] ),
    .B(_07747_));
 sg13g2_a21oi_1 _16352_ (.A1(_07760_),
    .A2(_07761_),
    .Y(_01192_),
    .B1(_07753_));
 sg13g2_nand3_1 _16353_ (.B(\soc_I.spi0_I.spi_buf[7] ),
    .C(net344),
    .A(net532),
    .Y(_07762_));
 sg13g2_nand2_1 _16354_ (.Y(_07763_),
    .A(\soc_I.spi0_I.rx_data[7] ),
    .B(_07747_));
 sg13g2_a21oi_1 _16355_ (.A1(_07762_),
    .A2(_07763_),
    .Y(_01193_),
    .B1(net373));
 sg13g2_nor2b_1 _16356_ (.A(_07742_),
    .B_N(_07740_),
    .Y(_07764_));
 sg13g2_nand2b_1 _16357_ (.Y(_07765_),
    .B(_05741_),
    .A_N(_05731_));
 sg13g2_a21oi_2 _16358_ (.B1(net388),
    .Y(_07766_),
    .A2(_07765_),
    .A1(_05744_));
 sg13g2_or2_1 _16359_ (.X(_07767_),
    .B(_07766_),
    .A(\soc_I.spi0_I.sclk ));
 sg13g2_nand3b_1 _16360_ (.B(_07738_),
    .C(_07766_),
    .Y(_07768_),
    .A_N(_00058_));
 sg13g2_o21ai_1 _16361_ (.B1(_07768_),
    .Y(_07769_),
    .A1(_07764_),
    .A2(_07767_));
 sg13g2_nand2_1 _16362_ (.Y(_01194_),
    .A(net437),
    .B(_07769_));
 sg13g2_nand2_1 _16363_ (.Y(_07770_),
    .A(\soc_I.spi0_I.spi_buf[7] ),
    .B(_07766_));
 sg13g2_nand2b_1 _16364_ (.Y(_07771_),
    .B(\soc_I.spi0_I.sio0_si_mosi ),
    .A_N(_07766_));
 sg13g2_a21oi_1 _16365_ (.A1(_07770_),
    .A2(_07771_),
    .Y(_01195_),
    .B1(net373));
 sg13g2_o21ai_1 _16366_ (.B1(_01800_),
    .Y(_07772_),
    .A1(_01610_),
    .A2(net76));
 sg13g2_a21oi_1 _16367_ (.A1(_01605_),
    .A2(_07772_),
    .Y(_07773_),
    .B1(net521));
 sg13g2_nand2_1 _16368_ (.Y(_07774_),
    .A(_07742_),
    .B(_07773_));
 sg13g2_a21oi_2 _16369_ (.B1(_07740_),
    .Y(_07775_),
    .A2(_07766_),
    .A1(_00058_));
 sg13g2_a21oi_1 _16370_ (.A1(_07740_),
    .A2(_07774_),
    .Y(_07776_),
    .B1(_07775_));
 sg13g2_buf_1 _16371_ (.A(_07776_),
    .X(_07777_));
 sg13g2_buf_1 _16372_ (.A(_07777_),
    .X(_07778_));
 sg13g2_nor2_1 _16373_ (.A(\soc_I.spi0_I.spi_buf[0] ),
    .B(net56),
    .Y(_07779_));
 sg13g2_and2_1 _16374_ (.A(net607),
    .B(net344),
    .X(_07780_));
 sg13g2_a21oi_1 _16375_ (.A1(net2),
    .A2(net345),
    .Y(_07781_),
    .B1(_07780_));
 sg13g2_and2_1 _16376_ (.A(net56),
    .B(_07781_),
    .X(_07782_));
 sg13g2_nor3_1 _16377_ (.A(net383),
    .B(_07779_),
    .C(_07782_),
    .Y(_01196_));
 sg13g2_nor2_1 _16378_ (.A(\soc_I.spi0_I.spi_buf[1] ),
    .B(_07778_),
    .Y(_07783_));
 sg13g2_and2_1 _16379_ (.A(net604),
    .B(net388),
    .X(_07784_));
 sg13g2_a21oi_1 _16380_ (.A1(\soc_I.spi0_I.spi_buf[0] ),
    .A2(net345),
    .Y(_07785_),
    .B1(_07784_));
 sg13g2_and2_1 _16381_ (.A(net56),
    .B(_07785_),
    .X(_07786_));
 sg13g2_nor3_1 _16382_ (.A(net383),
    .B(_07783_),
    .C(_07786_),
    .Y(_01197_));
 sg13g2_nor2_1 _16383_ (.A(\soc_I.spi0_I.spi_buf[2] ),
    .B(_07778_),
    .Y(_07787_));
 sg13g2_and2_1 _16384_ (.A(net619),
    .B(net388),
    .X(_07788_));
 sg13g2_a21oi_1 _16385_ (.A1(\soc_I.spi0_I.spi_buf[1] ),
    .A2(net345),
    .Y(_07789_),
    .B1(_07788_));
 sg13g2_and2_1 _16386_ (.A(_07777_),
    .B(_07789_),
    .X(_07790_));
 sg13g2_nor3_1 _16387_ (.A(_07024_),
    .B(_07787_),
    .C(_07790_),
    .Y(_01198_));
 sg13g2_nor2_1 _16388_ (.A(\soc_I.spi0_I.spi_buf[3] ),
    .B(net56),
    .Y(_01299_));
 sg13g2_and2_1 _16389_ (.A(_05929_),
    .B(net388),
    .X(_01300_));
 sg13g2_a21oi_1 _16390_ (.A1(\soc_I.spi0_I.spi_buf[2] ),
    .A2(net345),
    .Y(_01301_),
    .B1(_01300_));
 sg13g2_and2_1 _16391_ (.A(_07777_),
    .B(_01301_),
    .X(_01302_));
 sg13g2_nor3_1 _16392_ (.A(_07024_),
    .B(_01299_),
    .C(_01302_),
    .Y(_01199_));
 sg13g2_buf_1 _16393_ (.A(_05918_),
    .X(_01303_));
 sg13g2_nor2_1 _16394_ (.A(\soc_I.spi0_I.spi_buf[4] ),
    .B(net56),
    .Y(_01304_));
 sg13g2_and2_1 _16395_ (.A(net606),
    .B(net388),
    .X(_01305_));
 sg13g2_a21oi_1 _16396_ (.A1(\soc_I.spi0_I.spi_buf[3] ),
    .A2(net345),
    .Y(_01306_),
    .B1(_01305_));
 sg13g2_and2_1 _16397_ (.A(_07777_),
    .B(_01306_),
    .X(_01307_));
 sg13g2_nor3_1 _16398_ (.A(net372),
    .B(_01304_),
    .C(_01307_),
    .Y(_01200_));
 sg13g2_nor2_1 _16399_ (.A(\soc_I.spi0_I.spi_buf[5] ),
    .B(net56),
    .Y(_01308_));
 sg13g2_and2_1 _16400_ (.A(_05941_),
    .B(_06802_),
    .X(_01309_));
 sg13g2_a21oi_1 _16401_ (.A1(\soc_I.spi0_I.spi_buf[4] ),
    .A2(net345),
    .Y(_01310_),
    .B1(_01309_));
 sg13g2_and2_1 _16402_ (.A(_07777_),
    .B(_01310_),
    .X(_01311_));
 sg13g2_nor3_1 _16403_ (.A(net372),
    .B(_01308_),
    .C(_01311_),
    .Y(_01201_));
 sg13g2_nor2_1 _16404_ (.A(\soc_I.spi0_I.spi_buf[6] ),
    .B(net56),
    .Y(_01312_));
 sg13g2_nor2_1 _16405_ (.A(_05982_),
    .B(_05751_),
    .Y(_01313_));
 sg13g2_a21oi_1 _16406_ (.A1(\soc_I.spi0_I.spi_buf[5] ),
    .A2(_07738_),
    .Y(_01314_),
    .B1(_01313_));
 sg13g2_and2_1 _16407_ (.A(_07777_),
    .B(_01314_),
    .X(_01315_));
 sg13g2_nor3_1 _16408_ (.A(_01303_),
    .B(_01312_),
    .C(_01315_),
    .Y(_01202_));
 sg13g2_nor2_1 _16409_ (.A(\soc_I.spi0_I.spi_buf[7] ),
    .B(net56),
    .Y(_01316_));
 sg13g2_and2_1 _16410_ (.A(net605),
    .B(net388),
    .X(_01317_));
 sg13g2_a21oi_1 _16411_ (.A1(\soc_I.spi0_I.spi_buf[6] ),
    .A2(_05751_),
    .Y(_01318_),
    .B1(_01317_));
 sg13g2_and2_1 _16412_ (.A(_07777_),
    .B(_01318_),
    .X(_01319_));
 sg13g2_nor3_1 _16413_ (.A(_01303_),
    .B(_01316_),
    .C(_01319_),
    .Y(_01203_));
 sg13g2_nand4_1 _16414_ (.B(_04213_),
    .C(_05912_),
    .A(_03854_),
    .Y(_01320_),
    .D(_07773_));
 sg13g2_nor2_1 _16415_ (.A(_01691_),
    .B(_01320_),
    .Y(_01321_));
 sg13g2_nor2b_1 _16416_ (.A(\soc_I.spi0_I.cen ),
    .B_N(_01320_),
    .Y(_01322_));
 sg13g2_o21ai_1 _16417_ (.B1(net437),
    .Y(_01204_),
    .A1(_01321_),
    .A2(_01322_));
 sg13g2_nand2_1 _16418_ (.Y(_01323_),
    .A(_07737_),
    .B(net345));
 sg13g2_a21oi_1 _16419_ (.A1(_07743_),
    .A2(_01323_),
    .Y(_01205_),
    .B1(net373));
 sg13g2_o21ai_1 _16420_ (.B1(net596),
    .Y(_01324_),
    .A1(_07736_),
    .A2(_05751_));
 sg13g2_buf_1 _16421_ (.A(_01324_),
    .X(_01325_));
 sg13g2_xor2_1 _16422_ (.B(_07775_),
    .A(\soc_I.spi0_I.xfer_cycles[0] ),
    .X(_01326_));
 sg13g2_nor2_1 _16423_ (.A(_01325_),
    .B(_01326_),
    .Y(_01224_));
 sg13g2_nor2_1 _16424_ (.A(\soc_I.spi0_I.xfer_cycles[0] ),
    .B(_07775_),
    .Y(_01327_));
 sg13g2_xnor2_1 _16425_ (.Y(_01328_),
    .A(\soc_I.spi0_I.xfer_cycles[1] ),
    .B(_01327_));
 sg13g2_nor2_1 _16426_ (.A(_01325_),
    .B(_01328_),
    .Y(_01225_));
 sg13g2_o21ai_1 _16427_ (.B1(\soc_I.spi0_I.xfer_cycles[2] ),
    .Y(_01329_),
    .A1(_05747_),
    .A2(_07775_));
 sg13g2_or2_1 _16428_ (.X(_01330_),
    .B(_07775_),
    .A(_05749_));
 sg13g2_buf_1 _16429_ (.A(_01330_),
    .X(_01331_));
 sg13g2_a21oi_1 _16430_ (.A1(_01329_),
    .A2(_01331_),
    .Y(_01226_),
    .B1(_01325_));
 sg13g2_nand2_1 _16431_ (.Y(_01332_),
    .A(_05745_),
    .B(_01331_));
 sg13g2_nand2_1 _16432_ (.Y(_01333_),
    .A(net344),
    .B(_07774_));
 sg13g2_nor2_1 _16433_ (.A(_05745_),
    .B(_01331_),
    .Y(_01334_));
 sg13g2_nand2_1 _16434_ (.Y(_01335_),
    .A(_01333_),
    .B(_01334_));
 sg13g2_a21oi_1 _16435_ (.A1(_01332_),
    .A2(_01335_),
    .Y(_01227_),
    .B1(net373));
 sg13g2_xnor2_1 _16436_ (.Y(_01336_),
    .A(_05746_),
    .B(_01334_));
 sg13g2_nor2_1 _16437_ (.A(_01325_),
    .B(_01336_),
    .Y(_01228_));
 sg13g2_inv_1 _16438_ (.Y(_01337_),
    .A(_05746_));
 sg13g2_nand2_1 _16439_ (.Y(_01338_),
    .A(\soc_I.spi0_I.xfer_cycles[5] ),
    .B(_06501_));
 sg13g2_a21oi_1 _16440_ (.A1(_01337_),
    .A2(_01334_),
    .Y(_01229_),
    .B1(_01338_));
 sg13g2_nor3_1 _16441_ (.A(_05899_),
    .B(_04240_),
    .C(_04251_),
    .Y(_01339_));
 sg13g2_nor2b_1 _16442_ (.A(_05908_),
    .B_N(_01339_),
    .Y(_01230_));
 sg13g2_nand4_1 _16443_ (.B(_04640_),
    .C(_05912_),
    .A(net593),
    .Y(_01340_),
    .D(_01339_));
 sg13g2_buf_2 _16444_ (.A(_01340_),
    .X(_01341_));
 sg13g2_buf_1 _16445_ (.A(_01341_),
    .X(_01342_));
 sg13g2_mux2_1 _16446_ (.A0(net607),
    .A1(_05662_),
    .S(net55),
    .X(_01343_));
 sg13g2_and2_1 _16447_ (.A(net423),
    .B(_01343_),
    .X(_01231_));
 sg13g2_buf_1 _16448_ (.A(_01341_),
    .X(_01344_));
 sg13g2_nor2b_1 _16449_ (.A(_05674_),
    .B_N(net54),
    .Y(_01345_));
 sg13g2_buf_1 _16450_ (.A(_01341_),
    .X(_01346_));
 sg13g2_nor2_1 _16451_ (.A(_05926_),
    .B(net53),
    .Y(_01347_));
 sg13g2_nor3_1 _16452_ (.A(net372),
    .B(_01345_),
    .C(_01347_),
    .Y(_01232_));
 sg13g2_nor2b_1 _16453_ (.A(_05713_),
    .B_N(net54),
    .Y(_01348_));
 sg13g2_nor2_1 _16454_ (.A(_05931_),
    .B(net53),
    .Y(_01349_));
 sg13g2_nor3_1 _16455_ (.A(net372),
    .B(_01348_),
    .C(_01349_),
    .Y(_01233_));
 sg13g2_nor2b_1 _16456_ (.A(_05714_),
    .B_N(net54),
    .Y(_01350_));
 sg13g2_nor2_1 _16457_ (.A(_05937_),
    .B(net53),
    .Y(_01351_));
 sg13g2_nor3_1 _16458_ (.A(net372),
    .B(_01350_),
    .C(_01351_),
    .Y(_01234_));
 sg13g2_nor2b_1 _16459_ (.A(_05718_),
    .B_N(net54),
    .Y(_01352_));
 sg13g2_nor2_1 _16460_ (.A(_05943_),
    .B(net53),
    .Y(_01353_));
 sg13g2_nor3_1 _16461_ (.A(net372),
    .B(_01352_),
    .C(_01353_),
    .Y(_01235_));
 sg13g2_nor2b_1 _16462_ (.A(_05734_),
    .B_N(_01344_),
    .Y(_01354_));
 sg13g2_nor2_1 _16463_ (.A(_05948_),
    .B(_01346_),
    .Y(_01355_));
 sg13g2_nor3_1 _16464_ (.A(net372),
    .B(_01354_),
    .C(_01355_),
    .Y(_01236_));
 sg13g2_nor2b_1 _16465_ (.A(_05731_),
    .B_N(net54),
    .Y(_01356_));
 sg13g2_nor2_1 _16466_ (.A(_05953_),
    .B(_01346_),
    .Y(_01357_));
 sg13g2_nor3_1 _16467_ (.A(net372),
    .B(_01356_),
    .C(_01357_),
    .Y(_01237_));
 sg13g2_buf_1 _16468_ (.A(net520),
    .X(_01358_));
 sg13g2_nor2b_1 _16469_ (.A(\soc_I.spi_div_reg[16] ),
    .B_N(net54),
    .Y(_01359_));
 sg13g2_nor2_1 _16470_ (.A(_05958_),
    .B(net53),
    .Y(_01360_));
 sg13g2_nor3_1 _16471_ (.A(net422),
    .B(_01359_),
    .C(_01360_),
    .Y(_01238_));
 sg13g2_nor2b_1 _16472_ (.A(\soc_I.spi_div_reg[17] ),
    .B_N(net54),
    .Y(_01361_));
 sg13g2_nor2_1 _16473_ (.A(_05962_),
    .B(net53),
    .Y(_01362_));
 sg13g2_nor3_1 _16474_ (.A(net422),
    .B(_01361_),
    .C(_01362_),
    .Y(_01239_));
 sg13g2_nor2b_1 _16475_ (.A(\soc_I.spi_div_reg[18] ),
    .B_N(net54),
    .Y(_01363_));
 sg13g2_nor2_1 _16476_ (.A(_05966_),
    .B(net53),
    .Y(_01364_));
 sg13g2_nor3_1 _16477_ (.A(_01358_),
    .B(_01363_),
    .C(_01364_),
    .Y(_01240_));
 sg13g2_buf_1 _16478_ (.A(_01341_),
    .X(_01365_));
 sg13g2_nor2b_1 _16479_ (.A(\soc_I.spi_div_reg[19] ),
    .B_N(net52),
    .Y(_01366_));
 sg13g2_nor2_1 _16480_ (.A(_05970_),
    .B(net53),
    .Y(_01367_));
 sg13g2_nor3_1 _16481_ (.A(_01358_),
    .B(_01366_),
    .C(_01367_),
    .Y(_01241_));
 sg13g2_mux2_1 _16482_ (.A0(net604),
    .A1(_05663_),
    .S(net55),
    .X(_01368_));
 sg13g2_and2_1 _16483_ (.A(net423),
    .B(_01368_),
    .X(_01242_));
 sg13g2_nor2b_1 _16484_ (.A(\soc_I.spi_div_reg[20] ),
    .B_N(net52),
    .Y(_01369_));
 sg13g2_buf_1 _16485_ (.A(_01341_),
    .X(_01370_));
 sg13g2_nor2_1 _16486_ (.A(_05974_),
    .B(net51),
    .Y(_01371_));
 sg13g2_nor3_1 _16487_ (.A(net422),
    .B(_01369_),
    .C(_01371_),
    .Y(_01243_));
 sg13g2_nor2b_1 _16488_ (.A(\soc_I.spi_div_reg[21] ),
    .B_N(net52),
    .Y(_01372_));
 sg13g2_nor2_1 _16489_ (.A(_05978_),
    .B(net51),
    .Y(_01373_));
 sg13g2_nor3_1 _16490_ (.A(net422),
    .B(_01372_),
    .C(_01373_),
    .Y(_01244_));
 sg13g2_nor2b_1 _16491_ (.A(\soc_I.spi_div_reg[22] ),
    .B_N(net52),
    .Y(_01374_));
 sg13g2_nor2_1 _16492_ (.A(_05984_),
    .B(net51),
    .Y(_01375_));
 sg13g2_nor3_1 _16493_ (.A(net422),
    .B(_01374_),
    .C(_01375_),
    .Y(_01245_));
 sg13g2_nor2b_1 _16494_ (.A(\soc_I.spi_div_reg[23] ),
    .B_N(net52),
    .Y(_01376_));
 sg13g2_nor2_1 _16495_ (.A(_05988_),
    .B(net51),
    .Y(_01377_));
 sg13g2_nor3_1 _16496_ (.A(net422),
    .B(_01376_),
    .C(_01377_),
    .Y(_01246_));
 sg13g2_mux2_1 _16497_ (.A0(_05993_),
    .A1(\soc_I.spi_div_reg[24] ),
    .S(net55),
    .X(_01378_));
 sg13g2_and2_1 _16498_ (.A(net423),
    .B(_01378_),
    .X(_01247_));
 sg13g2_mux2_1 _16499_ (.A0(_05999_),
    .A1(\soc_I.spi_div_reg[25] ),
    .S(net55),
    .X(_01379_));
 sg13g2_and2_1 _16500_ (.A(net423),
    .B(_01379_),
    .X(_01248_));
 sg13g2_nor2b_1 _16501_ (.A(\soc_I.spi_div_reg[26] ),
    .B_N(net52),
    .Y(_01380_));
 sg13g2_nor2_1 _16502_ (.A(_06009_),
    .B(net51),
    .Y(_01381_));
 sg13g2_nor3_1 _16503_ (.A(net422),
    .B(_01380_),
    .C(_01381_),
    .Y(_01249_));
 sg13g2_or2_1 _16504_ (.X(_01382_),
    .B(net52),
    .A(_07385_));
 sg13g2_nand2_1 _16505_ (.Y(_01383_),
    .A(\soc_I.spi_div_reg[27] ),
    .B(net51));
 sg13g2_a21oi_1 _16506_ (.A1(_01382_),
    .A2(_01383_),
    .Y(_01250_),
    .B1(_07753_));
 sg13g2_mux2_1 _16507_ (.A0(_06019_),
    .A1(\soc_I.spi_div_reg[28] ),
    .S(net55),
    .X(_01384_));
 sg13g2_and2_1 _16508_ (.A(net423),
    .B(_01384_),
    .X(_01251_));
 sg13g2_or2_1 _16509_ (.X(_01385_),
    .B(net52),
    .A(_07413_));
 sg13g2_nand2_1 _16510_ (.Y(_01386_),
    .A(\soc_I.spi_div_reg[29] ),
    .B(net51));
 sg13g2_a21oi_1 _16511_ (.A1(_01385_),
    .A2(_01386_),
    .Y(_01252_),
    .B1(net398));
 sg13g2_mux2_1 _16512_ (.A0(_02277_),
    .A1(_05664_),
    .S(_01342_),
    .X(_01387_));
 sg13g2_and2_1 _16513_ (.A(net423),
    .B(_01387_),
    .X(_01253_));
 sg13g2_mux2_1 _16514_ (.A0(_06030_),
    .A1(\soc_I.spi_div_reg[30] ),
    .S(net55),
    .X(_01388_));
 sg13g2_and2_1 _16515_ (.A(net423),
    .B(_01388_),
    .X(_01254_));
 sg13g2_or2_1 _16516_ (.X(_01389_),
    .B(net55),
    .A(_07440_));
 sg13g2_nand2_1 _16517_ (.Y(_01390_),
    .A(\soc_I.spi_div_reg[31] ),
    .B(net51));
 sg13g2_a21oi_1 _16518_ (.A1(_01389_),
    .A2(_01390_),
    .Y(_01255_),
    .B1(net398));
 sg13g2_mux2_1 _16519_ (.A0(_05929_),
    .A1(\soc_I.spi0_I.div[3] ),
    .S(net55),
    .X(_01391_));
 sg13g2_and2_1 _16520_ (.A(_07613_),
    .B(_01391_),
    .X(_01256_));
 sg13g2_mux2_1 _16521_ (.A0(net606),
    .A1(_05661_),
    .S(_01341_),
    .X(_01392_));
 sg13g2_and2_1 _16522_ (.A(_07613_),
    .B(_01392_),
    .X(_01257_));
 sg13g2_buf_1 _16523_ (.A(_03578_),
    .X(_01393_));
 sg13g2_mux2_1 _16524_ (.A0(_05941_),
    .A1(\soc_I.spi0_I.div[5] ),
    .S(_01341_),
    .X(_01394_));
 sg13g2_and2_1 _16525_ (.A(net421),
    .B(_01394_),
    .X(_01258_));
 sg13g2_or2_1 _16526_ (.X(_01395_),
    .B(_01342_),
    .A(_05982_));
 sg13g2_nand2_1 _16527_ (.Y(_01396_),
    .A(_05660_),
    .B(_01344_));
 sg13g2_a21oi_1 _16528_ (.A1(_01395_),
    .A2(_01396_),
    .Y(_01259_),
    .B1(net398));
 sg13g2_mux2_1 _16529_ (.A0(net605),
    .A1(\soc_I.spi0_I.div[7] ),
    .S(_01341_),
    .X(_01397_));
 sg13g2_and2_1 _16530_ (.A(net421),
    .B(_01397_),
    .X(_01260_));
 sg13g2_nor2b_1 _16531_ (.A(_05659_),
    .B_N(_01365_),
    .Y(_01398_));
 sg13g2_nor2_1 _16532_ (.A(_06046_),
    .B(_01370_),
    .Y(_01399_));
 sg13g2_nor3_1 _16533_ (.A(net422),
    .B(_01398_),
    .C(_01399_),
    .Y(_01261_));
 sg13g2_nor2b_1 _16534_ (.A(_05657_),
    .B_N(_01365_),
    .Y(_01400_));
 sg13g2_nor2_1 _16535_ (.A(_06049_),
    .B(_01370_),
    .Y(_01401_));
 sg13g2_nor3_1 _16536_ (.A(net438),
    .B(_01400_),
    .C(_01401_),
    .Y(_01262_));
 sg13g2_nand2_1 _16537_ (.Y(_01402_),
    .A(_00092_),
    .B(_05459_));
 sg13g2_o21ai_1 _16538_ (.B1(_05456_),
    .Y(_01403_),
    .A1(net579),
    .A2(_05458_));
 sg13g2_a21oi_1 _16539_ (.A1(_01402_),
    .A2(_01403_),
    .Y(_01263_),
    .B1(_05919_));
 sg13g2_nand2_1 _16540_ (.Y(_01404_),
    .A(_05456_),
    .B(_05459_));
 sg13g2_xor2_1 _16541_ (.B(_01404_),
    .A(_05457_),
    .X(_01405_));
 sg13g2_nor2_1 _16542_ (.A(_05801_),
    .B(_01405_),
    .Y(_01264_));
 sg13g2_buf_1 _16543_ (.A(\soc_I.tx_uart_i.bit_idx[2] ),
    .X(_01406_));
 sg13g2_xor2_1 _16544_ (.B(_05460_),
    .A(_01406_),
    .X(_01407_));
 sg13g2_nor2_1 _16545_ (.A(_05801_),
    .B(_01407_),
    .Y(_01265_));
 sg13g2_nor2_1 _16546_ (.A(\soc_I.tx_uart_i.return_state[0] ),
    .B(net407),
    .Y(_01408_));
 sg13g2_nor4_1 _16547_ (.A(_05502_),
    .B(\soc_I.tx_uart_i.wait_states[10] ),
    .C(\soc_I.tx_uart_i.wait_states[13] ),
    .D(_05573_),
    .Y(_01409_));
 sg13g2_nor4_1 _16548_ (.A(_05464_),
    .B(_05494_),
    .C(_05495_),
    .D(\soc_I.tx_uart_i.wait_states[15] ),
    .Y(_01410_));
 sg13g2_nor4_1 _16549_ (.A(_05476_),
    .B(_05477_),
    .C(_05534_),
    .D(_05543_),
    .Y(_01411_));
 sg13g2_nor4_1 _16550_ (.A(_05488_),
    .B(_05489_),
    .C(_05482_),
    .D(_05483_),
    .Y(_01412_));
 sg13g2_and4_1 _16551_ (.A(_01409_),
    .B(_01410_),
    .C(_01411_),
    .D(_01412_),
    .X(_01413_));
 sg13g2_nand2b_1 _16552_ (.Y(_01414_),
    .B(net439),
    .A_N(_01413_));
 sg13g2_o21ai_1 _16553_ (.B1(_01414_),
    .Y(_01415_),
    .A1(_05455_),
    .A2(_01408_));
 sg13g2_and2_1 _16554_ (.A(net421),
    .B(_01415_),
    .X(_01268_));
 sg13g2_nor2_1 _16555_ (.A(\soc_I.tx_uart_i.return_state[1] ),
    .B(net407),
    .Y(_01416_));
 sg13g2_o21ai_1 _16556_ (.B1(_01414_),
    .Y(_01417_),
    .A1(_05455_),
    .A2(_01416_));
 sg13g2_and2_1 _16557_ (.A(net421),
    .B(_01417_),
    .X(_01269_));
 sg13g2_nand2_1 _16558_ (.Y(_01418_),
    .A(_05448_),
    .B(_05454_));
 sg13g2_buf_2 _16559_ (.A(_01418_),
    .X(_01419_));
 sg13g2_mux2_1 _16560_ (.A0(_05910_),
    .A1(\soc_I.tx_uart_i.tx_data_reg[0] ),
    .S(_01419_),
    .X(_01420_));
 sg13g2_and2_1 _16561_ (.A(net421),
    .B(_01420_),
    .X(_01270_));
 sg13g2_mux2_1 _16562_ (.A0(_05961_),
    .A1(\soc_I.tx_uart_i.tx_data_reg[1] ),
    .S(_01419_),
    .X(_01421_));
 sg13g2_and2_1 _16563_ (.A(net421),
    .B(_01421_),
    .X(_01271_));
 sg13g2_mux2_1 _16564_ (.A0(net619),
    .A1(\soc_I.tx_uart_i.tx_data_reg[2] ),
    .S(_01419_),
    .X(_01422_));
 sg13g2_and2_1 _16565_ (.A(_01393_),
    .B(_01422_),
    .X(_01272_));
 sg13g2_mux2_1 _16566_ (.A0(_05929_),
    .A1(\soc_I.tx_uart_i.tx_data_reg[3] ),
    .S(_01419_),
    .X(_01423_));
 sg13g2_and2_1 _16567_ (.A(_01393_),
    .B(_01423_),
    .X(_01273_));
 sg13g2_mux2_1 _16568_ (.A0(_05935_),
    .A1(\soc_I.tx_uart_i.tx_data_reg[4] ),
    .S(_01419_),
    .X(_01424_));
 sg13g2_and2_1 _16569_ (.A(net421),
    .B(_01424_),
    .X(_01274_));
 sg13g2_mux2_1 _16570_ (.A0(_05941_),
    .A1(\soc_I.tx_uart_i.tx_data_reg[5] ),
    .S(_01419_),
    .X(_01425_));
 sg13g2_and2_1 _16571_ (.A(net421),
    .B(_01425_),
    .X(_01275_));
 sg13g2_nand3_1 _16572_ (.B(_05448_),
    .C(_05454_),
    .A(_05946_),
    .Y(_01426_));
 sg13g2_nand2_1 _16573_ (.Y(_01427_),
    .A(\soc_I.tx_uart_i.tx_data_reg[6] ),
    .B(_01419_));
 sg13g2_a21oi_1 _16574_ (.A1(_01426_),
    .A2(_01427_),
    .Y(_01276_),
    .B1(_05919_));
 sg13g2_mux2_1 _16575_ (.A0(_05951_),
    .A1(\soc_I.tx_uart_i.tx_data_reg[7] ),
    .S(_01419_),
    .X(_01428_));
 sg13g2_and2_1 _16576_ (.A(_06501_),
    .B(_01428_),
    .X(_01277_));
 sg13g2_mux4_1 _16577_ (.S0(_05456_),
    .A0(\soc_I.tx_uart_i.tx_data_reg[2] ),
    .A1(\soc_I.tx_uart_i.tx_data_reg[3] ),
    .A2(\soc_I.tx_uart_i.tx_data_reg[6] ),
    .A3(\soc_I.tx_uart_i.tx_data_reg[7] ),
    .S1(_01406_),
    .X(_01429_));
 sg13g2_nand2_1 _16578_ (.Y(_01430_),
    .A(_05457_),
    .B(_01429_));
 sg13g2_mux4_1 _16579_ (.S0(_05456_),
    .A0(\soc_I.tx_uart_i.tx_data_reg[0] ),
    .A1(\soc_I.tx_uart_i.tx_data_reg[1] ),
    .A2(\soc_I.tx_uart_i.tx_data_reg[4] ),
    .A3(\soc_I.tx_uart_i.tx_data_reg[5] ),
    .S1(_01406_),
    .X(_01431_));
 sg13g2_nand2b_1 _16580_ (.Y(_01432_),
    .B(_01431_),
    .A_N(_05457_));
 sg13g2_nand3_1 _16581_ (.B(_01430_),
    .C(_01432_),
    .A(net610),
    .Y(_01433_));
 sg13g2_nand2_1 _16582_ (.Y(_01434_),
    .A(_05458_),
    .B(_05454_));
 sg13g2_a21oi_1 _16583_ (.A1(_01433_),
    .A2(_01434_),
    .Y(_01435_),
    .B1(net579));
 sg13g2_nor3_1 _16584_ (.A(_05467_),
    .B(_05458_),
    .C(\soc_I.tx_uart_i.tx_out ),
    .Y(_01436_));
 sg13g2_o21ai_1 _16585_ (.B1(_05810_),
    .Y(_01278_),
    .A1(_01435_),
    .A2(_01436_));
 sg13g2_nor3_1 _16586_ (.A(\soc_I.tx_uart_i.return_state[1] ),
    .B(\soc_I.tx_uart_i.return_state[0] ),
    .C(_05442_),
    .Y(_01437_));
 sg13g2_a21oi_1 _16587_ (.A1(_01413_),
    .A2(_01437_),
    .Y(_01438_),
    .B1(\soc_I.tx_uart_i.ready ));
 sg13g2_nor3_1 _16588_ (.A(_05802_),
    .B(_05448_),
    .C(_01438_),
    .Y(_01279_));
 sg13g2_nand3_1 _16589_ (.B(\soc_I.cpu_mem_addr[0] ),
    .C(_04228_),
    .A(net515),
    .Y(_01439_));
 sg13g2_nor3_1 _16590_ (.A(_05899_),
    .B(_04223_),
    .C(_01439_),
    .Y(_01296_));
 sg13g2_or2_1 _16591_ (.X(_01440_),
    .B(_05901_),
    .A(_05444_));
 sg13g2_nor3_1 _16592_ (.A(net593),
    .B(_07540_),
    .C(_01440_),
    .Y(_01297_));
 sg13g2_nor2_1 _16593_ (.A(_05445_),
    .B(_01440_),
    .Y(_01298_));
 sg13g2_buf_1 _16594_ (.A(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[1] ),
    .X(_01441_));
 sg13g2_buf_1 _16595_ (.A(_01441_),
    .X(_01442_));
 sg13g2_nor2b_1 _16596_ (.A(_01610_),
    .B_N(net631),
    .Y(_01443_));
 sg13g2_nand2_1 _16597_ (.Y(_01444_),
    .A(net505),
    .B(_01443_));
 sg13g2_buf_1 _16598_ (.A(_01444_),
    .X(_01445_));
 sg13g2_buf_1 _16599_ (.A(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ),
    .X(_01446_));
 sg13g2_and3_1 _16600_ (.X(_01447_),
    .A(_01840_),
    .B(_01624_),
    .C(_01723_));
 sg13g2_nand2_1 _16601_ (.Y(_01448_),
    .A(_01446_),
    .B(_01447_));
 sg13g2_buf_2 _16602_ (.A(_01448_),
    .X(_01449_));
 sg13g2_inv_1 _16603_ (.Y(_01450_),
    .A(_01449_));
 sg13g2_nand2_1 _16604_ (.Y(_01451_),
    .A(_01445_),
    .B(_01450_));
 sg13g2_buf_1 _16605_ (.A(_01451_),
    .X(_01452_));
 sg13g2_inv_1 _16606_ (.Y(_01453_),
    .A(_01452_));
 sg13g2_nand3_1 _16607_ (.B(_06726_),
    .C(_01453_),
    .A(net531),
    .Y(_01454_));
 sg13g2_o21ai_1 _16608_ (.B1(_01444_),
    .Y(_01455_),
    .A1(net531),
    .A2(_01450_));
 sg13g2_buf_1 _16609_ (.A(_01455_),
    .X(_01456_));
 sg13g2_nand2_1 _16610_ (.Y(_01457_),
    .A(net531),
    .B(_01444_));
 sg13g2_nor2_2 _16611_ (.A(_01450_),
    .B(_01457_),
    .Y(_01458_));
 sg13g2_a22oi_1 _16612_ (.Y(_01459_),
    .B1(_01458_),
    .B2(\soc_I.qqspi_I.rdata[16] ),
    .A2(_01456_),
    .A1(\soc_I.qqspi_I.rdata[0] ));
 sg13g2_inv_1 _16613_ (.Y(_01460_),
    .A(_01459_));
 sg13g2_nor4_1 _16614_ (.A(net330),
    .B(_06639_),
    .C(_01450_),
    .D(_01457_),
    .Y(_01461_));
 sg13g2_a22oi_1 _16615_ (.Y(_01462_),
    .B1(_01461_),
    .B2(net67),
    .A2(_01460_),
    .A1(net432));
 sg13g2_nor2_1 _16616_ (.A(net531),
    .B(_01452_),
    .Y(_01463_));
 sg13g2_nand2b_1 _16617_ (.Y(_01464_),
    .B(_01463_),
    .A_N(_06889_));
 sg13g2_and2_1 _16618_ (.A(_05957_),
    .B(_01443_),
    .X(_01465_));
 sg13g2_buf_1 _16619_ (.A(_01465_),
    .X(_01466_));
 sg13g2_nor2_1 _16620_ (.A(net531),
    .B(_01450_),
    .Y(_01467_));
 sg13g2_and3_1 _16621_ (.X(_01468_),
    .A(_04271_),
    .B(_06563_),
    .C(_06564_));
 sg13g2_o21ai_1 _16622_ (.B1(_01468_),
    .Y(_01469_),
    .A1(_01466_),
    .A2(_01467_));
 sg13g2_nand4_1 _16623_ (.B(_01462_),
    .C(_01464_),
    .A(_01454_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[0] ),
    .D(_01469_));
 sg13g2_inv_1 _16624_ (.Y(_01470_),
    .A(_01441_));
 sg13g2_a221oi_1 _16625_ (.B2(_06716_),
    .C1(_01470_),
    .B1(_06579_),
    .A1(net615),
    .Y(_01471_),
    .A2(\soc_I.qqspi_I.rdata[23] ));
 sg13g2_nor2_1 _16626_ (.A(_01441_),
    .B(_06880_),
    .Y(_01472_));
 sg13g2_or3_1 _16627_ (.A(_01446_),
    .B(_01471_),
    .C(_01472_),
    .X(_01473_));
 sg13g2_nor2_1 _16628_ (.A(_01441_),
    .B(_06627_),
    .Y(_01474_));
 sg13g2_a221oi_1 _16629_ (.B2(_01441_),
    .C1(_01474_),
    .B1(_06805_),
    .A1(net617),
    .Y(_01475_),
    .A2(_06628_));
 sg13g2_mux2_1 _16630_ (.A0(\soc_I.qqspi_I.rdata[15] ),
    .A1(\soc_I.qqspi_I.rdata[31] ),
    .S(_01441_),
    .X(_01476_));
 sg13g2_and2_1 _16631_ (.A(_04325_),
    .B(_01476_),
    .X(_01477_));
 sg13g2_a21o_1 _16632_ (.A2(_01475_),
    .A1(_06579_),
    .B1(_01477_),
    .X(_01478_));
 sg13g2_buf_1 _16633_ (.A(_01478_),
    .X(_01479_));
 sg13g2_nand2_1 _16634_ (.Y(_01480_),
    .A(_01446_),
    .B(_01479_));
 sg13g2_nor2_1 _16635_ (.A(net602),
    .B(net505),
    .Y(_01481_));
 sg13g2_nand2_1 _16636_ (.Y(_01482_),
    .A(_01840_),
    .B(_01481_));
 sg13g2_a21oi_1 _16637_ (.A1(_01473_),
    .A2(_01480_),
    .Y(_01483_),
    .B1(_01482_));
 sg13g2_buf_2 _16638_ (.A(_01483_),
    .X(_01484_));
 sg13g2_buf_1 _16639_ (.A(_01470_),
    .X(_01485_));
 sg13g2_nor2_1 _16640_ (.A(net458),
    .B(_01447_),
    .Y(_01486_));
 sg13g2_buf_2 _16641_ (.A(_01486_),
    .X(_01487_));
 sg13g2_a21oi_1 _16642_ (.A1(net602),
    .A2(net631),
    .Y(_01488_),
    .B1(net504));
 sg13g2_o21ai_1 _16643_ (.B1(_05957_),
    .Y(_01489_),
    .A1(_01470_),
    .A2(_01443_));
 sg13g2_o21ai_1 _16644_ (.B1(_01489_),
    .Y(_01490_),
    .A1(net531),
    .A2(_01488_));
 sg13g2_buf_2 _16645_ (.A(_01490_),
    .X(_01491_));
 sg13g2_inv_1 _16646_ (.Y(_01492_),
    .A(_06587_));
 sg13g2_a22oi_1 _16647_ (.Y(_01493_),
    .B1(_01491_),
    .B2(_01492_),
    .A2(_01487_),
    .A1(_06746_));
 sg13g2_nand2b_1 _16648_ (.Y(\soc_I.kianv_I.datapath_unit_I.Data[10] ),
    .B(_01493_),
    .A_N(_01484_));
 sg13g2_inv_1 _16649_ (.Y(_01494_),
    .A(_06594_));
 sg13g2_a22oi_1 _16650_ (.Y(_01495_),
    .B1(_01491_),
    .B2(_01494_),
    .A2(_01487_),
    .A1(_06757_));
 sg13g2_nand2b_1 _16651_ (.Y(\soc_I.kianv_I.datapath_unit_I.Data[11] ),
    .B(_01495_),
    .A_N(_01484_));
 sg13g2_inv_1 _16652_ (.Y(_01496_),
    .A(_06601_));
 sg13g2_a22oi_1 _16653_ (.Y(_01497_),
    .B1(_01491_),
    .B2(_01496_),
    .A2(_01487_),
    .A1(_06768_));
 sg13g2_nand2b_1 _16654_ (.Y(\soc_I.kianv_I.datapath_unit_I.Data[12] ),
    .B(_01497_),
    .A_N(_01484_));
 sg13g2_nor2b_1 _16655_ (.A(_06776_),
    .B_N(_01487_),
    .Y(_01498_));
 sg13g2_inv_1 _16656_ (.Y(_01499_),
    .A(_01491_));
 sg13g2_a21oi_1 _16657_ (.A1(_06603_),
    .A2(_06612_),
    .Y(_01500_),
    .B1(_01499_));
 sg13g2_or3_1 _16658_ (.A(_01484_),
    .B(_01498_),
    .C(_01500_),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[13] ));
 sg13g2_nor2b_1 _16659_ (.A(_06797_),
    .B_N(_01487_),
    .Y(_01501_));
 sg13g2_a21oi_1 _16660_ (.A1(_06615_),
    .A2(_06620_),
    .Y(_01502_),
    .B1(_01499_));
 sg13g2_or3_1 _16661_ (.A(_01484_),
    .B(_01501_),
    .C(_01502_),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[14] ));
 sg13g2_buf_1 _16662_ (.A(_01466_),
    .X(_01503_));
 sg13g2_nor3_1 _16663_ (.A(_01446_),
    .B(_01471_),
    .C(_01472_),
    .Y(_01504_));
 sg13g2_nand2b_1 _16664_ (.Y(_01505_),
    .B(_01504_),
    .A_N(_01482_));
 sg13g2_nand2_1 _16665_ (.Y(_01506_),
    .A(_01613_),
    .B(_01601_));
 sg13g2_inv_1 _16666_ (.Y(_01507_),
    .A(_01613_));
 sg13g2_nand2_1 _16667_ (.Y(_01508_),
    .A(_01507_),
    .B(_01446_));
 sg13g2_nand3_1 _16668_ (.B(_01506_),
    .C(_01508_),
    .A(net397),
    .Y(_01509_));
 sg13g2_a21oi_1 _16669_ (.A1(_01479_),
    .A2(_01509_),
    .Y(_01510_),
    .B1(_01503_));
 sg13g2_a22oi_1 _16670_ (.Y(\soc_I.kianv_I.datapath_unit_I.Data[15] ),
    .B1(_01505_),
    .B2(_01510_),
    .A2(net327),
    .A1(_06633_));
 sg13g2_o21ai_1 _16671_ (.B1(_01481_),
    .Y(_01511_),
    .A1(_05990_),
    .A2(_01446_));
 sg13g2_nand2b_1 _16672_ (.Y(_01512_),
    .B(_01479_),
    .A_N(_01511_));
 sg13g2_o21ai_1 _16673_ (.B1(_01512_),
    .Y(_01513_),
    .A1(_01482_),
    .A2(_01473_));
 sg13g2_buf_8 _16674_ (.A(_01513_),
    .X(_01514_));
 sg13g2_buf_2 _16675_ (.A(_01514_),
    .X(_01515_));
 sg13g2_nor2_1 _16676_ (.A(_06641_),
    .B(net371),
    .Y(_01516_));
 sg13g2_or2_1 _16677_ (.X(\soc_I.kianv_I.datapath_unit_I.Data[16] ),
    .B(_01516_),
    .A(net28));
 sg13g2_nor2_1 _16678_ (.A(_06651_),
    .B(net371),
    .Y(_01517_));
 sg13g2_or2_1 _16679_ (.X(\soc_I.kianv_I.datapath_unit_I.Data[17] ),
    .B(_01517_),
    .A(_01515_));
 sg13g2_nor2_1 _16680_ (.A(_06657_),
    .B(net371),
    .Y(_01518_));
 sg13g2_or2_1 _16681_ (.X(\soc_I.kianv_I.datapath_unit_I.Data[18] ),
    .B(_01518_),
    .A(_01514_));
 sg13g2_nor2_1 _16682_ (.A(_06663_),
    .B(net371),
    .Y(_01519_));
 sg13g2_or2_1 _16683_ (.X(\soc_I.kianv_I.datapath_unit_I.Data[19] ),
    .B(_01519_),
    .A(_01514_));
 sg13g2_mux2_1 _16684_ (.A0(\soc_I.qqspi_I.rdata[9] ),
    .A1(\soc_I.qqspi_I.rdata[25] ),
    .S(net531),
    .X(_01520_));
 sg13g2_o21ai_1 _16685_ (.B1(net458),
    .Y(_01521_),
    .A1(net466),
    .A2(_06893_));
 sg13g2_o21ai_1 _16686_ (.B1(_01521_),
    .Y(_01522_),
    .A1(net458),
    .A2(_06732_));
 sg13g2_a221oi_1 _16687_ (.B2(net57),
    .C1(_01452_),
    .B1(_01522_),
    .A1(net432),
    .Y(_01523_),
    .A2(_01520_));
 sg13g2_a221oi_1 _16688_ (.B2(_06651_),
    .C1(_01523_),
    .B1(_01458_),
    .A1(_06685_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[1] ),
    .A2(_01456_));
 sg13g2_nor2_1 _16689_ (.A(_06691_),
    .B(net371),
    .Y(_01524_));
 sg13g2_or2_1 _16690_ (.X(\soc_I.kianv_I.datapath_unit_I.Data[20] ),
    .B(_01524_),
    .A(_01514_));
 sg13g2_a21o_1 _16691_ (.A2(net327),
    .A1(_06699_),
    .B1(net28),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[21] ));
 sg13g2_a21o_1 _16692_ (.A2(net327),
    .A1(_06709_),
    .B1(net28),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[22] ));
 sg13g2_inv_1 _16693_ (.Y(_01525_),
    .A(_06717_));
 sg13g2_a21o_1 _16694_ (.A2(_01503_),
    .A1(_01525_),
    .B1(_01515_),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[23] ));
 sg13g2_a21o_1 _16695_ (.A2(net327),
    .A1(_06726_),
    .B1(net28),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[24] ));
 sg13g2_a21o_1 _16696_ (.A2(net327),
    .A1(_06736_),
    .B1(net28),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[25] ));
 sg13g2_a21o_1 _16697_ (.A2(net327),
    .A1(_06746_),
    .B1(net28),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[26] ));
 sg13g2_a21o_1 _16698_ (.A2(net327),
    .A1(_06757_),
    .B1(net28),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[27] ));
 sg13g2_a21o_1 _16699_ (.A2(net327),
    .A1(_06768_),
    .B1(net28),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[28] ));
 sg13g2_nor2_1 _16700_ (.A(_06776_),
    .B(net371),
    .Y(_01526_));
 sg13g2_or2_1 _16701_ (.X(\soc_I.kianv_I.datapath_unit_I.Data[29] ),
    .B(_01526_),
    .A(_01514_));
 sg13g2_mux2_1 _16702_ (.A0(\soc_I.qqspi_I.rdata[10] ),
    .A1(\soc_I.qqspi_I.rdata[26] ),
    .S(net531),
    .X(_01527_));
 sg13g2_o21ai_1 _16703_ (.B1(net458),
    .Y(_01528_),
    .A1(net466),
    .A2(_06584_));
 sg13g2_o21ai_1 _16704_ (.B1(_01528_),
    .Y(_01529_),
    .A1(net458),
    .A2(_06742_));
 sg13g2_a221oi_1 _16705_ (.B2(net57),
    .C1(_01452_),
    .B1(_01529_),
    .A1(net432),
    .Y(_01530_),
    .A2(_01527_));
 sg13g2_a221oi_1 _16706_ (.B2(_06657_),
    .C1(_01530_),
    .B1(_01458_),
    .A1(_06790_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[2] ),
    .A2(_01456_));
 sg13g2_nor2_1 _16707_ (.A(_06797_),
    .B(net371),
    .Y(_01531_));
 sg13g2_or2_1 _16708_ (.X(\soc_I.kianv_I.datapath_unit_I.Data[30] ),
    .B(_01531_),
    .A(_01514_));
 sg13g2_nor2_1 _16709_ (.A(_06807_),
    .B(net371),
    .Y(_01532_));
 sg13g2_or2_1 _16710_ (.X(\soc_I.kianv_I.datapath_unit_I.Data[31] ),
    .B(_01532_),
    .A(_01514_));
 sg13g2_mux2_1 _16711_ (.A0(\soc_I.qqspi_I.rdata[11] ),
    .A1(\soc_I.qqspi_I.rdata[27] ),
    .S(_01442_),
    .X(_01533_));
 sg13g2_o21ai_1 _16712_ (.B1(net458),
    .Y(_01534_),
    .A1(net466),
    .A2(_06591_));
 sg13g2_o21ai_1 _16713_ (.B1(_01534_),
    .Y(_01535_),
    .A1(net458),
    .A2(_06753_));
 sg13g2_a221oi_1 _16714_ (.B2(_06632_),
    .C1(_01452_),
    .B1(_01535_),
    .A1(net432),
    .Y(_01536_),
    .A2(_01533_));
 sg13g2_a221oi_1 _16715_ (.B2(_06663_),
    .C1(_01536_),
    .B1(_01458_),
    .A1(_06821_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[3] ),
    .A2(_01456_));
 sg13g2_mux2_1 _16716_ (.A0(\soc_I.qqspi_I.rdata[12] ),
    .A1(\soc_I.qqspi_I.rdata[28] ),
    .S(_01442_),
    .X(_01537_));
 sg13g2_o21ai_1 _16717_ (.B1(_01485_),
    .Y(_01538_),
    .A1(net466),
    .A2(_06598_));
 sg13g2_o21ai_1 _16718_ (.B1(_01538_),
    .Y(_01539_),
    .A1(_01485_),
    .A2(_06764_));
 sg13g2_a221oi_1 _16719_ (.B2(_06632_),
    .C1(_01452_),
    .B1(_01539_),
    .A1(net432),
    .Y(_01540_),
    .A2(_01537_));
 sg13g2_a221oi_1 _16720_ (.B2(_06691_),
    .C1(_01540_),
    .B1(_01458_),
    .A1(_06835_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[4] ),
    .A2(_01456_));
 sg13g2_mux2_1 _16721_ (.A0(\soc_I.qqspi_I.rdata[29] ),
    .A1(\soc_I.qqspi_I.rdata[21] ),
    .S(_01449_),
    .X(_01541_));
 sg13g2_nand2_1 _16722_ (.Y(_01542_),
    .A(_06697_),
    .B(_01449_));
 sg13g2_o21ai_1 _16723_ (.B1(_01542_),
    .Y(_01543_),
    .A1(_06774_),
    .A2(_01449_));
 sg13g2_a221oi_1 _16724_ (.B2(net57),
    .C1(_01457_),
    .B1(_01543_),
    .A1(_06531_),
    .Y(_01544_),
    .A2(_01541_));
 sg13g2_a221oi_1 _16725_ (.B2(_06613_),
    .C1(_01544_),
    .B1(_01463_),
    .A1(_06849_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[5] ),
    .A2(_01456_));
 sg13g2_mux2_1 _16726_ (.A0(\soc_I.qqspi_I.rdata[30] ),
    .A1(\soc_I.qqspi_I.rdata[22] ),
    .S(_01449_),
    .X(_01545_));
 sg13g2_nand2_1 _16727_ (.Y(_01546_),
    .A(_06707_),
    .B(_01449_));
 sg13g2_o21ai_1 _16728_ (.B1(_01546_),
    .Y(_01547_),
    .A1(_06795_),
    .A2(_01449_));
 sg13g2_a221oi_1 _16729_ (.B2(net57),
    .C1(_01457_),
    .B1(_01547_),
    .A1(_06531_),
    .Y(_01548_),
    .A2(_01545_));
 sg13g2_a221oi_1 _16730_ (.B2(_06621_),
    .C1(_01548_),
    .B1(_01463_),
    .A1(_06863_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[6] ),
    .A2(_01456_));
 sg13g2_nand2_1 _16731_ (.Y(_01549_),
    .A(_01453_),
    .B(_01479_));
 sg13g2_o21ai_1 _16732_ (.B1(_01504_),
    .Y(_01550_),
    .A1(net458),
    .A2(_01445_));
 sg13g2_a22oi_1 _16733_ (.Y(_01551_),
    .B1(_01491_),
    .B2(_06880_),
    .A2(_01487_),
    .A1(_01525_));
 sg13g2_nand3_1 _16734_ (.B(_01550_),
    .C(_01551_),
    .A(_01549_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[7] ));
 sg13g2_nand2_1 _16735_ (.Y(_01552_),
    .A(_06726_),
    .B(_01487_));
 sg13g2_o21ai_1 _16736_ (.B1(_01552_),
    .Y(_01553_),
    .A1(_06889_),
    .A2(_01499_));
 sg13g2_or2_1 _16737_ (.X(\soc_I.kianv_I.datapath_unit_I.Data[8] ),
    .B(_01553_),
    .A(_01484_));
 sg13g2_inv_1 _16738_ (.Y(_01554_),
    .A(_06896_));
 sg13g2_a22oi_1 _16739_ (.Y(_01555_),
    .B1(_01491_),
    .B2(_01554_),
    .A2(_01487_),
    .A1(_06736_));
 sg13g2_nand2b_1 _16740_ (.Y(\soc_I.kianv_I.datapath_unit_I.Data[9] ),
    .B(_01555_),
    .A_N(_01484_));
 sg13g2_dfrbp_1 _16741_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net634),
    .D(_00093_),
    .Q_N(_08936_),
    .Q(_00000_));
 sg13g2_dfrbp_1 _16742_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net635),
    .D(_00094_),
    .Q_N(_08935_),
    .Q(_00001_));
 sg13g2_dfrbp_1 _16743_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net636),
    .D(_00095_),
    .Q_N(_08934_),
    .Q(_00002_));
 sg13g2_dfrbp_1 _16744_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net637),
    .D(_00096_),
    .Q_N(_08933_),
    .Q(_00003_));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _16746_ (.A(net638),
    .X(uio_oe[0]));
 sg13g2_buf_1 _16747_ (.A(net11),
    .X(net9));
 sg13g2_buf_1 _16748_ (.A(net639),
    .X(uio_oe[3]));
 sg13g2_buf_1 _16749_ (.A(net11),
    .X(net10));
 sg13g2_buf_1 _16750_ (.A(net640),
    .X(uio_oe[6]));
 sg13g2_buf_1 _16751_ (.A(net641),
    .X(uio_oe[7]));
 sg13g2_buf_1 _16752_ (.A(sio0_si_mosi_o),
    .X(net13));
 sg13g2_buf_1 _16753_ (.A(sio1_so_miso_o),
    .X(net14));
 sg13g2_buf_1 _16754_ (.A(sclk),
    .X(net15));
 sg13g2_buf_1 _16755_ (.A(sio2_o),
    .X(net16));
 sg13g2_buf_1 _16756_ (.A(sio3_o),
    .X(net17));
 sg13g2_buf_1 _16757_ (.A(net642),
    .X(uio_out[7]));
 sg13g2_buf_1 _16758_ (.A(\soc_I.spi0_I.cen ),
    .X(net19));
 sg13g2_buf_1 _16759_ (.A(\soc_I.spi0_I.sclk ),
    .X(net20));
 sg13g2_buf_1 _16760_ (.A(\soc_I.spi0_I.sio0_si_mosi ),
    .X(net21));
 sg13g2_buf_1 _16761_ (.A(pwm_o),
    .X(net22));
 sg13g2_buf_1 _16762_ (.A(\soc_I.tx_uart_i.tx_out ),
    .X(net23));
 sg13g2_buf_1 _16763_ (.A(\soc_I.PC[16] ),
    .X(net24));
 sg13g2_buf_1 _16764_ (.A(\soc_I.PC[17] ),
    .X(net25));
 sg13g2_buf_1 _16765_ (.A(\soc_I.PC[18] ),
    .X(net26));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[0]$_SDFF_PN0_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net643),
    .D(_00097_),
    .Q_N(_00087_),
    .Q(\soc_I.cycle_cnt[0] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[10]$_SDFF_PN0_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net644),
    .D(_00098_),
    .Q_N(_08932_),
    .Q(\soc_I.cycle_cnt[10] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[11]$_SDFF_PN0_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net645),
    .D(_00099_),
    .Q_N(_08931_),
    .Q(\soc_I.cycle_cnt[11] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[12]$_SDFF_PN0_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net646),
    .D(_00100_),
    .Q_N(_08930_),
    .Q(\soc_I.cycle_cnt[12] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[13]$_SDFF_PN0_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net647),
    .D(_00101_),
    .Q_N(_08929_),
    .Q(\soc_I.cycle_cnt[13] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[14]$_SDFF_PN0_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net648),
    .D(_00102_),
    .Q_N(_08928_),
    .Q(\soc_I.cycle_cnt[14] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[15]$_SDFF_PN0_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net649),
    .D(_00103_),
    .Q_N(_08927_),
    .Q(\soc_I.cycle_cnt[15] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[16]$_SDFF_PN0_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net650),
    .D(_00104_),
    .Q_N(_08926_),
    .Q(\soc_I.cycle_cnt[16] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[17]$_SDFF_PN0_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net651),
    .D(_00105_),
    .Q_N(_08925_),
    .Q(\soc_I.cycle_cnt[17] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[18]$_SDFF_PN0_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net652),
    .D(_00106_),
    .Q_N(_08924_),
    .Q(\soc_I.cycle_cnt[18] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[19]$_SDFF_PN0_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net653),
    .D(_00107_),
    .Q_N(_08923_),
    .Q(\soc_I.cycle_cnt[19] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[1]$_SDFF_PN0_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net654),
    .D(_00108_),
    .Q_N(_08922_),
    .Q(\soc_I.cycle_cnt[1] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[20]$_SDFF_PN0_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net655),
    .D(_00109_),
    .Q_N(_08921_),
    .Q(\soc_I.cycle_cnt[20] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[21]$_SDFF_PN0_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net656),
    .D(_00110_),
    .Q_N(_08920_),
    .Q(\soc_I.cycle_cnt[21] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[22]$_SDFF_PN0_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net657),
    .D(_00111_),
    .Q_N(_08919_),
    .Q(\soc_I.cycle_cnt[22] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[23]$_SDFF_PN0_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net658),
    .D(_00112_),
    .Q_N(_08918_),
    .Q(\soc_I.cycle_cnt[23] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[24]$_SDFF_PN0_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net659),
    .D(_00113_),
    .Q_N(_08917_),
    .Q(\soc_I.cycle_cnt[24] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[25]$_SDFF_PN0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net660),
    .D(_00114_),
    .Q_N(_08916_),
    .Q(\soc_I.cycle_cnt[25] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[26]$_SDFF_PN0_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net661),
    .D(_00115_),
    .Q_N(_08915_),
    .Q(\soc_I.cycle_cnt[26] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[27]$_SDFF_PN0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net662),
    .D(_00116_),
    .Q_N(_08914_),
    .Q(\soc_I.cycle_cnt[27] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[28]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net663),
    .D(_00117_),
    .Q_N(_08913_),
    .Q(\soc_I.cycle_cnt[28] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[29]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net664),
    .D(_00118_),
    .Q_N(_08912_),
    .Q(\soc_I.cycle_cnt[29] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[2]$_SDFF_PN0_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net665),
    .D(_00119_),
    .Q_N(_08911_),
    .Q(\soc_I.cycle_cnt[2] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[30]$_SDFF_PN0_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net666),
    .D(_00120_),
    .Q_N(_08910_),
    .Q(\soc_I.cycle_cnt[30] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[31]$_SDFF_PN0_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net667),
    .D(_00121_),
    .Q_N(_08909_),
    .Q(\soc_I.cycle_cnt[31] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[3]$_SDFF_PN0_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net668),
    .D(_00122_),
    .Q_N(_08908_),
    .Q(\soc_I.cycle_cnt[3] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[4]$_SDFF_PN0_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net669),
    .D(_00123_),
    .Q_N(_08907_),
    .Q(\soc_I.cycle_cnt[4] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[5]$_SDFF_PN0_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net670),
    .D(_00124_),
    .Q_N(_08906_),
    .Q(\soc_I.cycle_cnt[5] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[6]$_SDFF_PN0_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net671),
    .D(_00125_),
    .Q_N(_08905_),
    .Q(\soc_I.cycle_cnt[6] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[7]$_SDFF_PN0_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net672),
    .D(_00126_),
    .Q_N(_08904_),
    .Q(\soc_I.cycle_cnt[7] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[8]$_SDFF_PN0_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net673),
    .D(_00127_),
    .Q_N(_08903_),
    .Q(\soc_I.cycle_cnt[8] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt[9]$_SDFF_PN0_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net674),
    .D(_00128_),
    .Q_N(_08902_),
    .Q(\soc_I.cycle_cnt[9] ));
 sg13g2_dfrbp_1 \soc_I.cycle_cnt_ready$_SDFF_PN0_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net675),
    .D(_00129_),
    .Q_N(_08901_),
    .Q(\soc_I.cycle_cnt_ready ));
 sg13g2_dfrbp_1 \soc_I.div_ready$_SDFF_PN0_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net676),
    .D(_00130_),
    .Q_N(_08900_),
    .Q(\soc_I.div_ready ));
 sg13g2_dfrbp_1 \soc_I.div_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net677),
    .D(_00131_),
    .Q_N(_00060_),
    .Q(\soc_I.div_reg[0] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net678),
    .D(_00132_),
    .Q_N(_08899_),
    .Q(\soc_I.div_reg[10] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net679),
    .D(_00133_),
    .Q_N(_08898_),
    .Q(\soc_I.div_reg[11] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net680),
    .D(_00134_),
    .Q_N(_08897_),
    .Q(\soc_I.div_reg[12] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net681),
    .D(_00135_),
    .Q_N(_08896_),
    .Q(\soc_I.div_reg[13] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net682),
    .D(_00136_),
    .Q_N(_08895_),
    .Q(\soc_I.div_reg[14] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net683),
    .D(_00137_),
    .Q_N(_08894_),
    .Q(\soc_I.div_reg[15] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net684),
    .D(_00138_),
    .Q_N(_08893_),
    .Q(\soc_I.div_reg[16] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net685),
    .D(_00139_),
    .Q_N(_08892_),
    .Q(\soc_I.div_reg[17] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net686),
    .D(_00140_),
    .Q_N(_08891_),
    .Q(\soc_I.div_reg[18] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net687),
    .D(_00141_),
    .Q_N(_08890_),
    .Q(\soc_I.div_reg[19] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net688),
    .D(_00142_),
    .Q_N(_00064_),
    .Q(\soc_I.div_reg[1] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net689),
    .D(_00143_),
    .Q_N(_08889_),
    .Q(\soc_I.div_reg[20] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net690),
    .D(_00144_),
    .Q_N(_08888_),
    .Q(\soc_I.div_reg[21] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net691),
    .D(_00145_),
    .Q_N(_08887_),
    .Q(\soc_I.div_reg[22] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net692),
    .D(_00146_),
    .Q_N(_08886_),
    .Q(\soc_I.div_reg[23] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net693),
    .D(_00147_),
    .Q_N(_08885_),
    .Q(\soc_I.div_reg[24] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net694),
    .D(_00148_),
    .Q_N(_08884_),
    .Q(\soc_I.div_reg[25] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net695),
    .D(_00149_),
    .Q_N(_08883_),
    .Q(\soc_I.div_reg[26] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net696),
    .D(_00150_),
    .Q_N(_08882_),
    .Q(\soc_I.div_reg[27] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net697),
    .D(_00151_),
    .Q_N(_08881_),
    .Q(\soc_I.div_reg[28] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net698),
    .D(_00152_),
    .Q_N(_08880_),
    .Q(\soc_I.div_reg[29] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net699),
    .D(_00153_),
    .Q_N(_00066_),
    .Q(\soc_I.div_reg[2] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net700),
    .D(_00154_),
    .Q_N(_08879_),
    .Q(\soc_I.div_reg[30] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net701),
    .D(_00155_),
    .Q_N(_00078_),
    .Q(\soc_I.div_reg[31] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net702),
    .D(_00156_),
    .Q_N(_00068_),
    .Q(\soc_I.div_reg[3] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net703),
    .D(_00157_),
    .Q_N(_00070_),
    .Q(\soc_I.div_reg[4] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net704),
    .D(_00158_),
    .Q_N(_00072_),
    .Q(\soc_I.div_reg[5] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net705),
    .D(_00159_),
    .Q_N(_00074_),
    .Q(\soc_I.div_reg[6] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net706),
    .D(_00160_),
    .Q_N(_00076_),
    .Q(\soc_I.div_reg[7] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net707),
    .D(_00161_),
    .Q_N(_08878_),
    .Q(\soc_I.div_reg[8] ));
 sg13g2_dfrbp_1 \soc_I.div_reg[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net708),
    .D(_00162_),
    .Q_N(_08937_),
    .Q(\soc_I.div_reg[9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[0]$_DFF_P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net709),
    .D(_00007_),
    .Q_N(_08938_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[10]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net710),
    .D(_00008_),
    .Q_N(_00032_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[11]$_DFF_P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net711),
    .D(_00009_),
    .Q_N(_08939_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[12]$_DFF_P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net712),
    .D(_00010_),
    .Q_N(_08940_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[13]$_DFF_P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net713),
    .D(_00006_),
    .Q_N(_08941_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[1]$_DFF_P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net714),
    .D(_00011_),
    .Q_N(_08942_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[2]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net715),
    .D(_00004_),
    .Q_N(_08943_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[3]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net716),
    .D(_00012_),
    .Q_N(_08944_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[4]$_DFF_P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net717),
    .D(_00005_),
    .Q_N(_08945_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[5]$_DFF_P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net718),
    .D(_00013_),
    .Q_N(_00031_),
    .Q(\soc_I.kianv_I.control_unit_I.Branch ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[6]$_DFF_P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net719),
    .D(_00014_),
    .Q_N(_08946_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[7]$_DFF_P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net720),
    .D(_00015_),
    .Q_N(_08947_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[8]$_DFF_P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net721),
    .D(_00016_),
    .Q_N(_08948_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.control_unit_I.main_fsm_I.state[9]$_DFF_P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net722),
    .D(_00017_),
    .Q_N(_08877_),
    .Q(\soc_I.kianv_I.MemWrite ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[0]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net723),
    .D(_00163_),
    .Q_N(_08876_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[10]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net724),
    .D(_00164_),
    .Q_N(_08875_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[11]$_SDFF_PN0_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net725),
    .D(_00165_),
    .Q_N(_08874_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[12]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net726),
    .D(_00166_),
    .Q_N(_08873_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[13]$_SDFF_PN0_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net727),
    .D(_00167_),
    .Q_N(_08872_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[14]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net728),
    .D(_00168_),
    .Q_N(_08871_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[15]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net729),
    .D(_00169_),
    .Q_N(_08870_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[16]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net730),
    .D(_00170_),
    .Q_N(_08869_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[17]$_SDFF_PN0_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net731),
    .D(_00171_),
    .Q_N(_08868_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[18]$_SDFF_PN0_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net732),
    .D(_00172_),
    .Q_N(_08867_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[19]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net733),
    .D(_00173_),
    .Q_N(_08866_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[1]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net734),
    .D(_00174_),
    .Q_N(_08865_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[20]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net735),
    .D(_00175_),
    .Q_N(_08864_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[21]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net736),
    .D(_00176_),
    .Q_N(_08863_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[22]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net737),
    .D(_00177_),
    .Q_N(_08862_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[23]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net738),
    .D(_00178_),
    .Q_N(_08861_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[24]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net739),
    .D(_00179_),
    .Q_N(_08860_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[25]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net740),
    .D(_00180_),
    .Q_N(_08859_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[26]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net741),
    .D(_00181_),
    .Q_N(_08858_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[27]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net742),
    .D(_00182_),
    .Q_N(_08857_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[28]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net743),
    .D(_00183_),
    .Q_N(_08856_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[29]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net744),
    .D(_00184_),
    .Q_N(_08855_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[2]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net745),
    .D(_00185_),
    .Q_N(_08854_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[30]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net746),
    .D(_00186_),
    .Q_N(_08853_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[31]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net747),
    .D(_00187_),
    .Q_N(_08852_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[3]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net748),
    .D(_00188_),
    .Q_N(_08851_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[4]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net749),
    .D(_00189_),
    .Q_N(_08850_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[5]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net750),
    .D(_00190_),
    .Q_N(_08849_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[6]$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net751),
    .D(_00191_),
    .Q_N(_08848_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[7]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net752),
    .D(_00192_),
    .Q_N(_08847_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[8]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net753),
    .D(_00193_),
    .Q_N(_08846_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A1_I.q[9]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net754),
    .D(_00194_),
    .Q_N(_08845_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[0]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net755),
    .D(_00195_),
    .Q_N(_00026_),
    .Q(\soc_I.cpu_mem_wdata[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[10]$_SDFF_PN0_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net756),
    .D(_00196_),
    .Q_N(_00046_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[11]$_SDFF_PN0_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net757),
    .D(_00197_),
    .Q_N(_08844_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[12]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net758),
    .D(_00198_),
    .Q_N(_08843_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[13]$_SDFF_PN0_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net759),
    .D(_00199_),
    .Q_N(_08842_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[14]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net760),
    .D(_00200_),
    .Q_N(_08841_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[15]$_SDFF_PN0_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net761),
    .D(_00201_),
    .Q_N(_08840_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[16]$_SDFF_PN0_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net762),
    .D(_00202_),
    .Q_N(_08839_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[17]$_SDFF_PN0_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net763),
    .D(_00203_),
    .Q_N(_08838_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[18]$_SDFF_PN0_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net764),
    .D(_00204_),
    .Q_N(_08837_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[19]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net765),
    .D(_00205_),
    .Q_N(_08836_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[1]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net766),
    .D(_00206_),
    .Q_N(_00033_),
    .Q(\soc_I.cpu_mem_wdata[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[20]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net767),
    .D(_00207_),
    .Q_N(_08835_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[21]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net768),
    .D(_00208_),
    .Q_N(_08834_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[22]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net769),
    .D(_00209_),
    .Q_N(_08833_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[23]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net770),
    .D(_00210_),
    .Q_N(_08832_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[24]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net771),
    .D(_00211_),
    .Q_N(_08831_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[25]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net772),
    .D(_00212_),
    .Q_N(_08830_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[26]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net773),
    .D(_00213_),
    .Q_N(_08829_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[27]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net774),
    .D(_00214_),
    .Q_N(_08828_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[28]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net775),
    .D(_00215_),
    .Q_N(_08827_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[29]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net776),
    .D(_00216_),
    .Q_N(_08826_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[2]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net777),
    .D(_00217_),
    .Q_N(_00080_),
    .Q(\soc_I.cpu_mem_wdata[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[30]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net778),
    .D(_00218_),
    .Q_N(_08825_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[31]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net779),
    .D(_00219_),
    .Q_N(_08824_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[3]$_SDFF_PN0_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net780),
    .D(_00220_),
    .Q_N(_00036_),
    .Q(\soc_I.cpu_mem_wdata[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[4]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net781),
    .D(_00221_),
    .Q_N(_00038_),
    .Q(\soc_I.cpu_mem_wdata[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[5]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net782),
    .D(_00222_),
    .Q_N(_00040_),
    .Q(\soc_I.cpu_mem_wdata[5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[6]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net783),
    .D(_00223_),
    .Q_N(_00042_),
    .Q(\soc_I.cpu_mem_wdata[6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[7]$_SDFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net784),
    .D(_00224_),
    .Q_N(_00044_),
    .Q(\soc_I.cpu_mem_wdata[7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[8]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net785),
    .D(_00225_),
    .Q_N(_08823_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.A2_I.q[9]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net786),
    .D(_00226_),
    .Q_N(_08949_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net787),
    .D(\soc_I.cpu_mem_addr[0] ),
    .Q_N(_08950_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ADDR_I.q[1]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net788),
    .D(\soc_I.cpu_mem_addr[1] ),
    .Q_N(_08822_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net789),
    .D(_00227_),
    .Q_N(_08821_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net790),
    .D(_00228_),
    .Q_N(_08820_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net791),
    .D(_00229_),
    .Q_N(_08819_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net792),
    .D(_00230_),
    .Q_N(_08818_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net793),
    .D(_00231_),
    .Q_N(_08817_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net794),
    .D(_00232_),
    .Q_N(_08816_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net795),
    .D(_00233_),
    .Q_N(_08815_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net796),
    .D(_00234_),
    .Q_N(_08814_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net797),
    .D(_00235_),
    .Q_N(_08813_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net798),
    .D(_00236_),
    .Q_N(_08812_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net799),
    .D(_00237_),
    .Q_N(_08811_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net800),
    .D(_00238_),
    .Q_N(_08810_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net801),
    .D(_00239_),
    .Q_N(_08809_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net802),
    .D(_00240_),
    .Q_N(_08808_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net803),
    .D(_00241_),
    .Q_N(_08807_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net804),
    .D(_00242_),
    .Q_N(_08806_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net805),
    .D(_00243_),
    .Q_N(_08805_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net806),
    .D(_00244_),
    .Q_N(_08804_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net807),
    .D(_00245_),
    .Q_N(_08803_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net808),
    .D(_00246_),
    .Q_N(_08802_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net809),
    .D(_00247_),
    .Q_N(_08801_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net810),
    .D(_00248_),
    .Q_N(_08800_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net811),
    .D(_00249_),
    .Q_N(_08799_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net812),
    .D(_00250_),
    .Q_N(_08798_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net813),
    .D(_00251_),
    .Q_N(_08797_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net814),
    .D(_00252_),
    .Q_N(_08796_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net815),
    .D(_00253_),
    .Q_N(_08795_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net816),
    .D(_00254_),
    .Q_N(_08794_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net817),
    .D(_00255_),
    .Q_N(_08793_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net818),
    .D(_00256_),
    .Q_N(_08792_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net819),
    .D(_00257_),
    .Q_N(_08791_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net820),
    .D(_00258_),
    .Q_N(_08951_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[0]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net821),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[0] ),
    .Q_N(_08952_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[10]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net822),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[10] ),
    .Q_N(_08953_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[11]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net823),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[11] ),
    .Q_N(_08954_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[12]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net824),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[12] ),
    .Q_N(_08955_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[13]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net825),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[13] ),
    .Q_N(_08956_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[14]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net826),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[14] ),
    .Q_N(_08957_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[15]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net827),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[15] ),
    .Q_N(_08958_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[16]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net828),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[16] ),
    .Q_N(_08959_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[17]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net829),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[17] ),
    .Q_N(_08960_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[18]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net830),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[18] ),
    .Q_N(_08961_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[19]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net831),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[19] ),
    .Q_N(_08962_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[1]$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net832),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[1] ),
    .Q_N(_08963_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[20]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net833),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[20] ),
    .Q_N(_08964_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[21]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net834),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[21] ),
    .Q_N(_08965_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[22]$_DFF_P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net835),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[22] ),
    .Q_N(_08966_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[23]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net836),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[23] ),
    .Q_N(_08967_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[24]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net837),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[24] ),
    .Q_N(_08968_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[25]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net838),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[25] ),
    .Q_N(_08969_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[26]$_DFF_P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net839),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[26] ),
    .Q_N(_08970_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[27]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net840),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[27] ),
    .Q_N(_08971_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[28]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net841),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[28] ),
    .Q_N(_08972_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[29]$_DFF_P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net842),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[29] ),
    .Q_N(_08973_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[2]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net843),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[2] ),
    .Q_N(_08974_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[30]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net844),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[30] ),
    .Q_N(_08975_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[31]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net845),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[31] ),
    .Q_N(_08976_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[3]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net846),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[3] ),
    .Q_N(_08977_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[4]$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net847),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[4] ),
    .Q_N(_08978_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[5]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net848),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[5] ),
    .Q_N(_08979_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[6]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net849),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[6] ),
    .Q_N(_08980_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[7]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net850),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[7] ),
    .Q_N(_08981_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[8]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net851),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[8] ),
    .Q_N(_08982_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Data_I.q[9]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net852),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[9] ),
    .Q_N(_08790_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net853),
    .D(_00259_),
    .Q_N(_08789_),
    .Q(\soc_I.kianv_I.Instr[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net854),
    .D(_00260_),
    .Q_N(_08788_),
    .Q(\soc_I.kianv_I.Instr[10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net855),
    .D(_00261_),
    .Q_N(_08787_),
    .Q(\soc_I.kianv_I.Instr[11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net856),
    .D(_00262_),
    .Q_N(_00027_),
    .Q(\soc_I.kianv_I.Instr[12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net857),
    .D(_00263_),
    .Q_N(_08786_),
    .Q(\soc_I.kianv_I.Instr[13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net858),
    .D(_00264_),
    .Q_N(_00028_),
    .Q(\soc_I.kianv_I.Instr[14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net859),
    .D(_00265_),
    .Q_N(_08785_),
    .Q(\soc_I.kianv_I.Instr[15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net860),
    .D(_00266_),
    .Q_N(_08784_),
    .Q(\soc_I.kianv_I.Instr[16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net861),
    .D(_00267_),
    .Q_N(_08783_),
    .Q(\soc_I.kianv_I.Instr[17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net862),
    .D(_00268_),
    .Q_N(_08782_),
    .Q(\soc_I.kianv_I.Instr[18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net863),
    .D(_00269_),
    .Q_N(_08781_),
    .Q(\soc_I.kianv_I.Instr[19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net864),
    .D(_00270_),
    .Q_N(_08780_),
    .Q(\soc_I.kianv_I.Instr[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net865),
    .D(_00271_),
    .Q_N(_00035_),
    .Q(\soc_I.kianv_I.Instr[20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net866),
    .D(_00272_),
    .Q_N(_00034_),
    .Q(\soc_I.kianv_I.Instr[21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net867),
    .D(_00273_),
    .Q_N(_08779_),
    .Q(\soc_I.kianv_I.Instr[22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net868),
    .D(_00274_),
    .Q_N(_00037_),
    .Q(\soc_I.kianv_I.Instr[23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net869),
    .D(_00275_),
    .Q_N(_00039_),
    .Q(\soc_I.kianv_I.Instr[24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net870),
    .D(_00276_),
    .Q_N(_00041_),
    .Q(\soc_I.kianv_I.Instr[25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net871),
    .D(_00277_),
    .Q_N(_00043_),
    .Q(\soc_I.kianv_I.Instr[26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net872),
    .D(_00278_),
    .Q_N(_00045_),
    .Q(\soc_I.kianv_I.Instr[27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net873),
    .D(_00279_),
    .Q_N(_08778_),
    .Q(\soc_I.kianv_I.Instr[28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net874),
    .D(_00280_),
    .Q_N(_08777_),
    .Q(\soc_I.kianv_I.Instr[29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net875),
    .D(_00281_),
    .Q_N(_08776_),
    .Q(\soc_I.kianv_I.Instr[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net876),
    .D(_00282_),
    .Q_N(_00029_),
    .Q(\soc_I.kianv_I.Instr[30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net877),
    .D(_00283_),
    .Q_N(_08775_),
    .Q(\soc_I.kianv_I.Instr[31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net878),
    .D(_00284_),
    .Q_N(_08774_),
    .Q(\soc_I.kianv_I.Instr[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net879),
    .D(_00285_),
    .Q_N(_08773_),
    .Q(\soc_I.kianv_I.Instr[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net880),
    .D(_00286_),
    .Q_N(_08772_),
    .Q(\soc_I.kianv_I.Instr[5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net881),
    .D(_00287_),
    .Q_N(_00030_),
    .Q(\soc_I.kianv_I.Instr[6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net882),
    .D(_00288_),
    .Q_N(_08771_),
    .Q(\soc_I.kianv_I.Instr[7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net883),
    .D(_00289_),
    .Q_N(_08770_),
    .Q(\soc_I.kianv_I.Instr[8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.Instr_I.q[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net884),
    .D(_00290_),
    .Q_N(_08769_),
    .Q(\soc_I.kianv_I.Instr[9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net885),
    .D(_00291_),
    .Q_N(_08768_),
    .Q(\soc_I.PC[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net886),
    .D(_00292_),
    .Q_N(_08767_),
    .Q(\soc_I.PC[10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net887),
    .D(_00293_),
    .Q_N(_08766_),
    .Q(\soc_I.PC[11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net888),
    .D(_00294_),
    .Q_N(_08765_),
    .Q(\soc_I.PC[12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net889),
    .D(_00295_),
    .Q_N(_08764_),
    .Q(\soc_I.PC[13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net890),
    .D(_00296_),
    .Q_N(_08763_),
    .Q(\soc_I.PC[14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net891),
    .D(_00297_),
    .Q_N(_08762_),
    .Q(\soc_I.PC[15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net892),
    .D(_00298_),
    .Q_N(_08761_),
    .Q(\soc_I.PC[16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net893),
    .D(_00299_),
    .Q_N(_08760_),
    .Q(\soc_I.PC[17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net894),
    .D(_00300_),
    .Q_N(_08759_),
    .Q(\soc_I.PC[18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net895),
    .D(_00301_),
    .Q_N(_08758_),
    .Q(\soc_I.PC[19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net896),
    .D(_00302_),
    .Q_N(_08757_),
    .Q(\soc_I.PC[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net897),
    .D(_00303_),
    .Q_N(_08756_),
    .Q(\soc_I.PC[20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[21]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net898),
    .D(_00304_),
    .Q_N(_08755_),
    .Q(\soc_I.PC[21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net899),
    .D(_00305_),
    .Q_N(_08754_),
    .Q(\soc_I.PC[22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net900),
    .D(_00306_),
    .Q_N(_08753_),
    .Q(\soc_I.PC[23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net901),
    .D(_00307_),
    .Q_N(_08752_),
    .Q(\soc_I.PC[24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net902),
    .D(_00308_),
    .Q_N(_08751_),
    .Q(\soc_I.PC[25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net903),
    .D(_00309_),
    .Q_N(_08750_),
    .Q(\soc_I.PC[26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net904),
    .D(_00310_),
    .Q_N(_08749_),
    .Q(\soc_I.PC[27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net905),
    .D(_00311_),
    .Q_N(_08748_),
    .Q(\soc_I.PC[28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net906),
    .D(_00312_),
    .Q_N(_08747_),
    .Q(\soc_I.PC[29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net907),
    .D(_00313_),
    .Q_N(_08746_),
    .Q(\soc_I.PC[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net908),
    .D(_00314_),
    .Q_N(_08745_),
    .Q(\soc_I.PC[30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net909),
    .D(_00315_),
    .Q_N(_08744_),
    .Q(\soc_I.PC[31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net910),
    .D(_00316_),
    .Q_N(_08743_),
    .Q(\soc_I.PC[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net911),
    .D(_00317_),
    .Q_N(_08742_),
    .Q(\soc_I.PC[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net912),
    .D(_00318_),
    .Q_N(_08741_),
    .Q(\soc_I.PC[5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net913),
    .D(_00319_),
    .Q_N(_08740_),
    .Q(\soc_I.PC[6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net914),
    .D(_00320_),
    .Q_N(_08739_),
    .Q(\soc_I.PC[7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net915),
    .D(_00321_),
    .Q_N(_08738_),
    .Q(\soc_I.PC[8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net916),
    .D(_00322_),
    .Q_N(_08737_),
    .Q(\soc_I.PC[9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net917),
    .D(_00323_),
    .Q_N(_08736_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net918),
    .D(_00324_),
    .Q_N(_08735_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net919),
    .D(_00325_),
    .Q_N(_08734_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net920),
    .D(_00326_),
    .Q_N(_08733_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net921),
    .D(_00327_),
    .Q_N(_08732_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net922),
    .D(_00328_),
    .Q_N(_08731_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net923),
    .D(_00329_),
    .Q_N(_08730_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net924),
    .D(_00330_),
    .Q_N(_08729_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net925),
    .D(_00331_),
    .Q_N(_08728_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net926),
    .D(_00332_),
    .Q_N(_08727_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net927),
    .D(_00333_),
    .Q_N(_08726_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net928),
    .D(_00334_),
    .Q_N(_08725_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[20]$_SDFFE_PN1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net929),
    .D(_00335_),
    .Q_N(_08724_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net930),
    .D(_00336_),
    .Q_N(_08723_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net931),
    .D(_00337_),
    .Q_N(_08722_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net932),
    .D(_00338_),
    .Q_N(_08721_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net933),
    .D(_00339_),
    .Q_N(_08720_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net934),
    .D(_00340_),
    .Q_N(_08719_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net935),
    .D(_00341_),
    .Q_N(_08718_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net936),
    .D(_00342_),
    .Q_N(_08717_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net937),
    .D(_00343_),
    .Q_N(_08716_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[29]$_SDFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net938),
    .D(_00344_),
    .Q_N(_08715_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net939),
    .D(_00345_),
    .Q_N(_08714_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net940),
    .D(_00346_),
    .Q_N(_08713_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net941),
    .D(_00347_),
    .Q_N(_08712_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net942),
    .D(_00348_),
    .Q_N(_08711_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net943),
    .D(_00349_),
    .Q_N(_08710_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net944),
    .D(_00350_),
    .Q_N(_08709_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net945),
    .D(_00351_),
    .Q_N(_08708_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net946),
    .D(_00352_),
    .Q_N(_08707_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net947),
    .D(_00353_),
    .Q_N(_08706_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.PC_I.q[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net948),
    .D(_00354_),
    .Q_N(_08705_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Addr_I.d0[9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net949),
    .D(_00355_),
    .Q_N(_00086_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net950),
    .D(_00356_),
    .Q_N(_08704_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net951),
    .D(_00357_),
    .Q_N(_08703_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net952),
    .D(_00358_),
    .Q_N(_08702_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net953),
    .D(_00359_),
    .Q_N(_08701_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_ready$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net954),
    .D(_00360_),
    .Q_N(_00053_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_ready ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[0]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net955),
    .D(_00361_),
    .Q_N(_08700_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net956),
    .D(_00362_),
    .Q_N(_08699_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[11]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net957),
    .D(_00363_),
    .Q_N(_08698_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[12]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net958),
    .D(_00364_),
    .Q_N(_08697_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net959),
    .D(_00365_),
    .Q_N(_08696_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[14]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net960),
    .D(_00366_),
    .Q_N(_08695_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[15]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net961),
    .D(_00367_),
    .Q_N(_08694_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[16]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net962),
    .D(_00368_),
    .Q_N(_08693_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[17]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net963),
    .D(_00369_),
    .Q_N(_08692_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[18]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net964),
    .D(_00370_),
    .Q_N(_08691_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[19]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net965),
    .D(_00371_),
    .Q_N(_08690_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net966),
    .D(_00372_),
    .Q_N(_08689_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[20]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net967),
    .D(_00373_),
    .Q_N(_08688_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[21]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net968),
    .D(_00374_),
    .Q_N(_08687_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[22]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net969),
    .D(_00375_),
    .Q_N(_08686_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[23]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net970),
    .D(_00376_),
    .Q_N(_08685_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[24]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net971),
    .D(_00377_),
    .Q_N(_08684_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[25]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net972),
    .D(_00378_),
    .Q_N(_08683_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[26]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net973),
    .D(_00379_),
    .Q_N(_08682_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[27]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net974),
    .D(_00380_),
    .Q_N(_08681_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[28]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net975),
    .D(_00381_),
    .Q_N(_08680_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[29]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net976),
    .D(_00382_),
    .Q_N(_08679_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net977),
    .D(_00383_),
    .Q_N(_08678_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[30]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net978),
    .D(_00384_),
    .Q_N(_08677_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[31]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net979),
    .D(_00385_),
    .Q_N(_08676_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net980),
    .D(_00386_),
    .Q_N(_08675_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net981),
    .D(_00387_),
    .Q_N(_08674_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net982),
    .D(_00388_),
    .Q_N(_08673_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net983),
    .D(_00389_),
    .Q_N(_08672_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net984),
    .D(_00390_),
    .Q_N(_08671_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net985),
    .D(_00391_),
    .Q_N(_08670_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[9]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net986),
    .D(_00392_),
    .Q_N(_08669_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.alu_I.shift_state$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net987),
    .D(_00393_),
    .Q_N(_00052_),
    .Q(\soc_I.kianv_I.datapath_unit_I.alu_I.shift_state ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net988),
    .D(_00394_),
    .Q_N(_08668_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net989),
    .D(_00395_),
    .Q_N(_08667_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net990),
    .D(_00396_),
    .Q_N(_08666_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net991),
    .D(_00397_),
    .Q_N(_08665_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net992),
    .D(_00398_),
    .Q_N(_08664_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net993),
    .D(_00399_),
    .Q_N(_08663_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net994),
    .D(_00400_),
    .Q_N(_08662_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net995),
    .D(_00401_),
    .Q_N(_08661_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net996),
    .D(_00402_),
    .Q_N(_08660_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net997),
    .D(_00403_),
    .Q_N(_08659_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net998),
    .D(_00404_),
    .Q_N(_08658_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net999),
    .D(_00405_),
    .Q_N(_08657_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1000),
    .D(_00406_),
    .Q_N(_08656_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1001),
    .D(_00407_),
    .Q_N(_08655_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1002),
    .D(_00408_),
    .Q_N(_08654_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1003),
    .D(_00409_),
    .Q_N(_08653_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1004),
    .D(_00410_),
    .Q_N(_08652_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1005),
    .D(_00411_),
    .Q_N(_08651_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1006),
    .D(_00412_),
    .Q_N(_08650_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1007),
    .D(_00413_),
    .Q_N(_08649_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1008),
    .D(_00414_),
    .Q_N(_08648_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1009),
    .D(_00415_),
    .Q_N(_08647_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1010),
    .D(_00416_),
    .Q_N(_08646_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1011),
    .D(_00417_),
    .Q_N(_08645_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1012),
    .D(_00418_),
    .Q_N(_08644_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1013),
    .D(_00419_),
    .Q_N(_08643_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1014),
    .D(_00420_),
    .Q_N(_08642_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1015),
    .D(_00421_),
    .Q_N(_08641_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1016),
    .D(_00422_),
    .Q_N(_08640_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1017),
    .D(_00423_),
    .Q_N(_08639_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1018),
    .D(_00424_),
    .Q_N(_08638_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1019),
    .D(_00425_),
    .Q_N(_08637_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1020),
    .D(_00426_),
    .Q_N(_08636_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1021),
    .D(_00427_),
    .Q_N(_08635_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1022),
    .D(_00428_),
    .Q_N(_08634_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1023),
    .D(_00429_),
    .Q_N(_08633_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1024),
    .D(_00430_),
    .Q_N(_08632_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1025),
    .D(_00431_),
    .Q_N(_08631_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1026),
    .D(_00432_),
    .Q_N(_08630_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1027),
    .D(_00433_),
    .Q_N(_08629_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1028),
    .D(_00434_),
    .Q_N(_08628_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1029),
    .D(_00435_),
    .Q_N(_08627_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1030),
    .D(_00436_),
    .Q_N(_08626_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1031),
    .D(_00437_),
    .Q_N(_08625_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1032),
    .D(_00438_),
    .Q_N(_08624_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1033),
    .D(_00439_),
    .Q_N(_08623_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1034),
    .D(_00440_),
    .Q_N(_08622_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1035),
    .D(_00441_),
    .Q_N(_08621_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1036),
    .D(_00442_),
    .Q_N(_08620_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1037),
    .D(_00443_),
    .Q_N(_08619_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1038),
    .D(_00444_),
    .Q_N(_08618_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1039),
    .D(_00445_),
    .Q_N(_08617_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1040),
    .D(_00446_),
    .Q_N(_08616_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1041),
    .D(_00447_),
    .Q_N(_08615_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1042),
    .D(_00448_),
    .Q_N(_08614_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1043),
    .D(_00449_),
    .Q_N(_08613_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1044),
    .D(_00450_),
    .Q_N(_08612_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1045),
    .D(_00451_),
    .Q_N(_08611_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1046),
    .D(_00452_),
    .Q_N(_08610_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1047),
    .D(_00453_),
    .Q_N(_08609_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1048),
    .D(_00454_),
    .Q_N(_08608_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1049),
    .D(_00455_),
    .Q_N(_08607_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1050),
    .D(_00456_),
    .Q_N(_08606_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1051),
    .D(_00457_),
    .Q_N(_08605_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1052),
    .D(_00458_),
    .Q_N(_08604_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1053),
    .D(_00459_),
    .Q_N(_08603_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1054),
    .D(_00460_),
    .Q_N(_08602_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1055),
    .D(_00461_),
    .Q_N(_08601_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1056),
    .D(_00462_),
    .Q_N(_08600_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1057),
    .D(_00463_),
    .Q_N(_08599_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1058),
    .D(_00464_),
    .Q_N(_08598_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1059),
    .D(_00465_),
    .Q_N(_08597_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1060),
    .D(_00466_),
    .Q_N(_08596_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1061),
    .D(_00467_),
    .Q_N(_08595_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1062),
    .D(_00468_),
    .Q_N(_08594_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1063),
    .D(_00469_),
    .Q_N(_08593_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1064),
    .D(_00470_),
    .Q_N(_08592_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1065),
    .D(_00471_),
    .Q_N(_08591_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1066),
    .D(_00472_),
    .Q_N(_08590_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1067),
    .D(_00473_),
    .Q_N(_08589_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1068),
    .D(_00474_),
    .Q_N(_08588_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1069),
    .D(_00475_),
    .Q_N(_08587_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1070),
    .D(_00476_),
    .Q_N(_08586_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1071),
    .D(_00477_),
    .Q_N(_08585_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1072),
    .D(_00478_),
    .Q_N(_08584_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1073),
    .D(_00479_),
    .Q_N(_08583_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1074),
    .D(_00480_),
    .Q_N(_08582_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1075),
    .D(_00481_),
    .Q_N(_08581_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1076),
    .D(_00482_),
    .Q_N(_08580_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1077),
    .D(_00483_),
    .Q_N(_08579_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1078),
    .D(_00484_),
    .Q_N(_08578_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1079),
    .D(_00485_),
    .Q_N(_08577_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1080),
    .D(_00486_),
    .Q_N(_08576_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1081),
    .D(_00487_),
    .Q_N(_08575_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1082),
    .D(_00488_),
    .Q_N(_08574_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1083),
    .D(_00489_),
    .Q_N(_08573_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1084),
    .D(_00490_),
    .Q_N(_08572_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1085),
    .D(_00491_),
    .Q_N(_08571_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1086),
    .D(_00492_),
    .Q_N(_08570_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1087),
    .D(_00493_),
    .Q_N(_08569_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1088),
    .D(_00494_),
    .Q_N(_08568_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1089),
    .D(_00495_),
    .Q_N(_08567_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1090),
    .D(_00496_),
    .Q_N(_08566_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1091),
    .D(_00497_),
    .Q_N(_08565_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1092),
    .D(_00498_),
    .Q_N(_08564_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1093),
    .D(_00499_),
    .Q_N(_08563_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1094),
    .D(_00500_),
    .Q_N(_08562_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1095),
    .D(_00501_),
    .Q_N(_08561_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1096),
    .D(_00502_),
    .Q_N(_08560_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1097),
    .D(_00503_),
    .Q_N(_08559_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1098),
    .D(_00504_),
    .Q_N(_08558_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1099),
    .D(_00505_),
    .Q_N(_08557_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1100),
    .D(_00506_),
    .Q_N(_08556_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1101),
    .D(_00507_),
    .Q_N(_08555_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1102),
    .D(_00508_),
    .Q_N(_08554_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1103),
    .D(_00509_),
    .Q_N(_08553_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1104),
    .D(_00510_),
    .Q_N(_08552_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1105),
    .D(_00511_),
    .Q_N(_08551_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1106),
    .D(_00512_),
    .Q_N(_08550_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1107),
    .D(_00513_),
    .Q_N(_08549_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1108),
    .D(_00514_),
    .Q_N(_08548_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1109),
    .D(_00515_),
    .Q_N(_08547_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1110),
    .D(_00516_),
    .Q_N(_08546_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1111),
    .D(_00517_),
    .Q_N(_08545_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1112),
    .D(_00518_),
    .Q_N(_08544_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1113),
    .D(_00519_),
    .Q_N(_08543_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1114),
    .D(_00520_),
    .Q_N(_08542_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1115),
    .D(_00521_),
    .Q_N(_08541_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1116),
    .D(_00522_),
    .Q_N(_08540_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1117),
    .D(_00523_),
    .Q_N(_08539_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1118),
    .D(_00524_),
    .Q_N(_08538_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1119),
    .D(_00525_),
    .Q_N(_08537_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1120),
    .D(_00526_),
    .Q_N(_08536_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1121),
    .D(_00527_),
    .Q_N(_08535_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1122),
    .D(_00528_),
    .Q_N(_08534_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1123),
    .D(_00529_),
    .Q_N(_08533_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1124),
    .D(_00530_),
    .Q_N(_08532_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1125),
    .D(_00531_),
    .Q_N(_08531_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1126),
    .D(_00532_),
    .Q_N(_08530_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1127),
    .D(_00533_),
    .Q_N(_08529_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1128),
    .D(_00534_),
    .Q_N(_08528_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1129),
    .D(_00535_),
    .Q_N(_08527_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1130),
    .D(_00536_),
    .Q_N(_08526_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1131),
    .D(_00537_),
    .Q_N(_08525_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1132),
    .D(_00538_),
    .Q_N(_08524_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1133),
    .D(_00539_),
    .Q_N(_08523_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1134),
    .D(_00540_),
    .Q_N(_08522_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1135),
    .D(_00541_),
    .Q_N(_08521_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1136),
    .D(_00542_),
    .Q_N(_08520_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1137),
    .D(_00543_),
    .Q_N(_08519_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1138),
    .D(_00544_),
    .Q_N(_08518_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1139),
    .D(_00545_),
    .Q_N(_08517_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1140),
    .D(_00546_),
    .Q_N(_08516_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1141),
    .D(_00547_),
    .Q_N(_08515_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1142),
    .D(_00548_),
    .Q_N(_08514_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1143),
    .D(_00549_),
    .Q_N(_08513_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1144),
    .D(_00550_),
    .Q_N(_08512_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1145),
    .D(_00551_),
    .Q_N(_08511_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1146),
    .D(_00552_),
    .Q_N(_08510_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1147),
    .D(_00553_),
    .Q_N(_08509_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1148),
    .D(_00554_),
    .Q_N(_08508_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1149),
    .D(_00555_),
    .Q_N(_08507_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1150),
    .D(_00556_),
    .Q_N(_08506_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1151),
    .D(_00557_),
    .Q_N(_08505_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1152),
    .D(_00558_),
    .Q_N(_08504_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1153),
    .D(_00559_),
    .Q_N(_08503_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1154),
    .D(_00560_),
    .Q_N(_08502_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1155),
    .D(_00561_),
    .Q_N(_08501_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1156),
    .D(_00562_),
    .Q_N(_08500_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1157),
    .D(_00563_),
    .Q_N(_08499_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1158),
    .D(_00564_),
    .Q_N(_08498_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1159),
    .D(_00565_),
    .Q_N(_08497_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1160),
    .D(_00566_),
    .Q_N(_08496_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1161),
    .D(_00567_),
    .Q_N(_08495_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1162),
    .D(_00568_),
    .Q_N(_08494_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1163),
    .D(_00569_),
    .Q_N(_08493_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1164),
    .D(_00570_),
    .Q_N(_08492_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1165),
    .D(_00571_),
    .Q_N(_08491_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1166),
    .D(_00572_),
    .Q_N(_08490_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1167),
    .D(_00573_),
    .Q_N(_08489_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1168),
    .D(_00574_),
    .Q_N(_08488_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1169),
    .D(_00575_),
    .Q_N(_08487_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1170),
    .D(_00576_),
    .Q_N(_08486_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1171),
    .D(_00577_),
    .Q_N(_08485_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1172),
    .D(_00578_),
    .Q_N(_08484_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1173),
    .D(_00579_),
    .Q_N(_08483_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1174),
    .D(_00580_),
    .Q_N(_08482_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1175),
    .D(_00581_),
    .Q_N(_08481_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1176),
    .D(_00582_),
    .Q_N(_08480_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1177),
    .D(_00583_),
    .Q_N(_08479_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1178),
    .D(_00584_),
    .Q_N(_08478_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1179),
    .D(_00585_),
    .Q_N(_08477_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1180),
    .D(_00586_),
    .Q_N(_08476_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1181),
    .D(_00587_),
    .Q_N(_08475_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1182),
    .D(_00588_),
    .Q_N(_08474_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1183),
    .D(_00589_),
    .Q_N(_08473_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1184),
    .D(_00590_),
    .Q_N(_08472_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1185),
    .D(_00591_),
    .Q_N(_08471_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1186),
    .D(_00592_),
    .Q_N(_08470_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1187),
    .D(_00593_),
    .Q_N(_08469_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1188),
    .D(_00594_),
    .Q_N(_08468_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1189),
    .D(_00595_),
    .Q_N(_08467_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1190),
    .D(_00596_),
    .Q_N(_08466_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1191),
    .D(_00597_),
    .Q_N(_08465_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1192),
    .D(_00598_),
    .Q_N(_08464_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1193),
    .D(_00599_),
    .Q_N(_08463_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1194),
    .D(_00600_),
    .Q_N(_08462_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1195),
    .D(_00601_),
    .Q_N(_08461_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1196),
    .D(_00602_),
    .Q_N(_08460_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1197),
    .D(_00603_),
    .Q_N(_08459_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1198),
    .D(_00604_),
    .Q_N(_08458_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1199),
    .D(_00605_),
    .Q_N(_08457_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1200),
    .D(_00606_),
    .Q_N(_08456_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1201),
    .D(_00607_),
    .Q_N(_08455_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1202),
    .D(_00608_),
    .Q_N(_08454_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1203),
    .D(_00609_),
    .Q_N(_08453_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1204),
    .D(_00610_),
    .Q_N(_08452_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1205),
    .D(_00611_),
    .Q_N(_08451_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1206),
    .D(_00612_),
    .Q_N(_08450_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1207),
    .D(_00613_),
    .Q_N(_08449_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1208),
    .D(_00614_),
    .Q_N(_08448_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1209),
    .D(_00615_),
    .Q_N(_08447_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1210),
    .D(_00616_),
    .Q_N(_08446_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1211),
    .D(_00617_),
    .Q_N(_08445_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1212),
    .D(_00618_),
    .Q_N(_08444_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1213),
    .D(_00619_),
    .Q_N(_08443_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1214),
    .D(_00620_),
    .Q_N(_08442_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1215),
    .D(_00621_),
    .Q_N(_08441_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1216),
    .D(_00622_),
    .Q_N(_08440_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1217),
    .D(_00623_),
    .Q_N(_08439_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1218),
    .D(_00624_),
    .Q_N(_08438_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1219),
    .D(_00625_),
    .Q_N(_08437_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1220),
    .D(_00626_),
    .Q_N(_08436_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1221),
    .D(_00627_),
    .Q_N(_08435_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1222),
    .D(_00628_),
    .Q_N(_08434_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1223),
    .D(_00629_),
    .Q_N(_08433_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1224),
    .D(_00630_),
    .Q_N(_08432_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1225),
    .D(_00631_),
    .Q_N(_08431_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1226),
    .D(_00632_),
    .Q_N(_08430_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1227),
    .D(_00633_),
    .Q_N(_08429_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1228),
    .D(_00634_),
    .Q_N(_08428_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1229),
    .D(_00635_),
    .Q_N(_08427_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1230),
    .D(_00636_),
    .Q_N(_08426_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1231),
    .D(_00637_),
    .Q_N(_08425_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1232),
    .D(_00638_),
    .Q_N(_08424_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1233),
    .D(_00639_),
    .Q_N(_08423_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1234),
    .D(_00640_),
    .Q_N(_08422_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1235),
    .D(_00641_),
    .Q_N(_08421_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1236),
    .D(_00642_),
    .Q_N(_08420_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1237),
    .D(_00643_),
    .Q_N(_08419_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1238),
    .D(_00644_),
    .Q_N(_08418_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1239),
    .D(_00645_),
    .Q_N(_08417_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1240),
    .D(_00646_),
    .Q_N(_08416_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1241),
    .D(_00647_),
    .Q_N(_08415_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1242),
    .D(_00648_),
    .Q_N(_08414_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1243),
    .D(_00649_),
    .Q_N(_08413_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1244),
    .D(_00650_),
    .Q_N(_08412_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1245),
    .D(_00651_),
    .Q_N(_08411_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1246),
    .D(_00652_),
    .Q_N(_08410_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1247),
    .D(_00653_),
    .Q_N(_08409_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1248),
    .D(_00654_),
    .Q_N(_08408_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1249),
    .D(_00655_),
    .Q_N(_08407_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1250),
    .D(_00656_),
    .Q_N(_08406_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1251),
    .D(_00657_),
    .Q_N(_08405_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1252),
    .D(_00658_),
    .Q_N(_08404_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1253),
    .D(_00659_),
    .Q_N(_08403_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1254),
    .D(_00660_),
    .Q_N(_08402_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1255),
    .D(_00661_),
    .Q_N(_08401_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1256),
    .D(_00662_),
    .Q_N(_08400_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1257),
    .D(_00663_),
    .Q_N(_08399_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1258),
    .D(_00664_),
    .Q_N(_08398_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1259),
    .D(_00665_),
    .Q_N(_08397_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1260),
    .D(_00666_),
    .Q_N(_08396_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1261),
    .D(_00667_),
    .Q_N(_08395_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1262),
    .D(_00668_),
    .Q_N(_08394_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1263),
    .D(_00669_),
    .Q_N(_08393_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1264),
    .D(_00670_),
    .Q_N(_08392_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1265),
    .D(_00671_),
    .Q_N(_08391_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1266),
    .D(_00672_),
    .Q_N(_08390_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1267),
    .D(_00673_),
    .Q_N(_08389_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1268),
    .D(_00674_),
    .Q_N(_08388_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1269),
    .D(_00675_),
    .Q_N(_08387_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1270),
    .D(_00676_),
    .Q_N(_08386_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1271),
    .D(_00677_),
    .Q_N(_08385_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1272),
    .D(_00678_),
    .Q_N(_08384_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1273),
    .D(_00679_),
    .Q_N(_08383_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1274),
    .D(_00680_),
    .Q_N(_08382_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1275),
    .D(_00681_),
    .Q_N(_08381_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1276),
    .D(_00682_),
    .Q_N(_08380_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1277),
    .D(_00683_),
    .Q_N(_08379_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1278),
    .D(_00684_),
    .Q_N(_08378_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1279),
    .D(_00685_),
    .Q_N(_08377_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1280),
    .D(_00686_),
    .Q_N(_08376_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1281),
    .D(_00687_),
    .Q_N(_08375_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1282),
    .D(_00688_),
    .Q_N(_08374_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1283),
    .D(_00689_),
    .Q_N(_08373_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1284),
    .D(_00690_),
    .Q_N(_08372_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1285),
    .D(_00691_),
    .Q_N(_08371_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1286),
    .D(_00692_),
    .Q_N(_08370_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1287),
    .D(_00693_),
    .Q_N(_08369_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1288),
    .D(_00694_),
    .Q_N(_08368_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1289),
    .D(_00695_),
    .Q_N(_08367_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1290),
    .D(_00696_),
    .Q_N(_08366_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1291),
    .D(_00697_),
    .Q_N(_08365_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1292),
    .D(_00698_),
    .Q_N(_08364_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1293),
    .D(_00699_),
    .Q_N(_08363_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1294),
    .D(_00700_),
    .Q_N(_08362_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1295),
    .D(_00701_),
    .Q_N(_08361_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1296),
    .D(_00702_),
    .Q_N(_08360_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1297),
    .D(_00703_),
    .Q_N(_08359_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1298),
    .D(_00704_),
    .Q_N(_08358_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1299),
    .D(_00705_),
    .Q_N(_08357_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1300),
    .D(_00706_),
    .Q_N(_08356_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1301),
    .D(_00707_),
    .Q_N(_08355_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1302),
    .D(_00708_),
    .Q_N(_08354_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1303),
    .D(_00709_),
    .Q_N(_08353_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1304),
    .D(_00710_),
    .Q_N(_08352_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1305),
    .D(_00711_),
    .Q_N(_08351_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1306),
    .D(_00712_),
    .Q_N(_08350_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1307),
    .D(_00713_),
    .Q_N(_08349_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1308),
    .D(_00714_),
    .Q_N(_08348_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1309),
    .D(_00715_),
    .Q_N(_08347_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1310),
    .D(_00716_),
    .Q_N(_08346_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1311),
    .D(_00717_),
    .Q_N(_08345_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1312),
    .D(_00718_),
    .Q_N(_08344_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1313),
    .D(_00719_),
    .Q_N(_08343_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1314),
    .D(_00720_),
    .Q_N(_08342_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1315),
    .D(_00721_),
    .Q_N(_08341_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1316),
    .D(_00722_),
    .Q_N(_08340_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1317),
    .D(_00723_),
    .Q_N(_08339_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1318),
    .D(_00724_),
    .Q_N(_08338_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1319),
    .D(_00725_),
    .Q_N(_08337_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1320),
    .D(_00726_),
    .Q_N(_08336_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1321),
    .D(_00727_),
    .Q_N(_08335_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1322),
    .D(_00728_),
    .Q_N(_08334_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1323),
    .D(_00729_),
    .Q_N(_08333_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1324),
    .D(_00730_),
    .Q_N(_08332_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1325),
    .D(_00731_),
    .Q_N(_08331_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1326),
    .D(_00732_),
    .Q_N(_08330_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1327),
    .D(_00733_),
    .Q_N(_08329_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1328),
    .D(_00734_),
    .Q_N(_08328_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1329),
    .D(_00735_),
    .Q_N(_08327_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1330),
    .D(_00736_),
    .Q_N(_08326_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1331),
    .D(_00737_),
    .Q_N(_08325_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1332),
    .D(_00738_),
    .Q_N(_08324_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1333),
    .D(_00739_),
    .Q_N(_08323_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1334),
    .D(_00740_),
    .Q_N(_08322_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1335),
    .D(_00741_),
    .Q_N(_08321_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1336),
    .D(_00742_),
    .Q_N(_08320_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1337),
    .D(_00743_),
    .Q_N(_08319_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1338),
    .D(_00744_),
    .Q_N(_08318_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1339),
    .D(_00745_),
    .Q_N(_08317_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1340),
    .D(_00746_),
    .Q_N(_08316_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1341),
    .D(_00747_),
    .Q_N(_08315_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1342),
    .D(_00748_),
    .Q_N(_08314_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1343),
    .D(_00749_),
    .Q_N(_08313_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1344),
    .D(_00750_),
    .Q_N(_08312_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1345),
    .D(_00751_),
    .Q_N(_08311_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1346),
    .D(_00752_),
    .Q_N(_08310_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1347),
    .D(_00753_),
    .Q_N(_08309_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1348),
    .D(_00754_),
    .Q_N(_08308_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1349),
    .D(_00755_),
    .Q_N(_08307_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1350),
    .D(_00756_),
    .Q_N(_08306_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1351),
    .D(_00757_),
    .Q_N(_08305_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1352),
    .D(_00758_),
    .Q_N(_08304_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1353),
    .D(_00759_),
    .Q_N(_08303_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1354),
    .D(_00760_),
    .Q_N(_08302_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1355),
    .D(_00761_),
    .Q_N(_08301_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1356),
    .D(_00762_),
    .Q_N(_08300_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1357),
    .D(_00763_),
    .Q_N(_08299_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1358),
    .D(_00764_),
    .Q_N(_08298_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1359),
    .D(_00765_),
    .Q_N(_08297_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1360),
    .D(_00766_),
    .Q_N(_08296_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1361),
    .D(_00767_),
    .Q_N(_08295_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1362),
    .D(_00768_),
    .Q_N(_08294_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1363),
    .D(_00769_),
    .Q_N(_08293_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1364),
    .D(_00770_),
    .Q_N(_08292_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1365),
    .D(_00771_),
    .Q_N(_08291_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1366),
    .D(_00772_),
    .Q_N(_08290_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1367),
    .D(_00773_),
    .Q_N(_08289_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1368),
    .D(_00774_),
    .Q_N(_08288_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1369),
    .D(_00775_),
    .Q_N(_08287_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1370),
    .D(_00776_),
    .Q_N(_08286_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1371),
    .D(_00777_),
    .Q_N(_08285_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1372),
    .D(_00778_),
    .Q_N(_08284_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1373),
    .D(_00779_),
    .Q_N(_08283_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1374),
    .D(_00780_),
    .Q_N(_08282_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1375),
    .D(_00781_),
    .Q_N(_08281_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1376),
    .D(_00782_),
    .Q_N(_08280_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1377),
    .D(_00783_),
    .Q_N(_08279_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1378),
    .D(_00784_),
    .Q_N(_08278_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1379),
    .D(_00785_),
    .Q_N(_08277_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1380),
    .D(_00786_),
    .Q_N(_08276_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1381),
    .D(_00787_),
    .Q_N(_08275_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1382),
    .D(_00788_),
    .Q_N(_08274_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1383),
    .D(_00789_),
    .Q_N(_08273_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1384),
    .D(_00790_),
    .Q_N(_08272_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1385),
    .D(_00791_),
    .Q_N(_08271_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1386),
    .D(_00792_),
    .Q_N(_08270_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1387),
    .D(_00793_),
    .Q_N(_08269_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1388),
    .D(_00794_),
    .Q_N(_08268_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1389),
    .D(_00795_),
    .Q_N(_08267_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1390),
    .D(_00796_),
    .Q_N(_08266_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1391),
    .D(_00797_),
    .Q_N(_08265_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1392),
    .D(_00798_),
    .Q_N(_08264_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1393),
    .D(_00799_),
    .Q_N(_08263_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1394),
    .D(_00800_),
    .Q_N(_08262_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1395),
    .D(_00801_),
    .Q_N(_08261_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1396),
    .D(_00802_),
    .Q_N(_08260_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1397),
    .D(_00803_),
    .Q_N(_08259_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1398),
    .D(_00804_),
    .Q_N(_08258_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1399),
    .D(_00805_),
    .Q_N(_08257_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1400),
    .D(_00806_),
    .Q_N(_08256_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1401),
    .D(_00807_),
    .Q_N(_08255_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1402),
    .D(_00808_),
    .Q_N(_08254_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1403),
    .D(_00809_),
    .Q_N(_08253_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1404),
    .D(_00810_),
    .Q_N(_08252_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1405),
    .D(_00811_),
    .Q_N(_08251_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1406),
    .D(_00812_),
    .Q_N(_08250_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1407),
    .D(_00813_),
    .Q_N(_08249_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1408),
    .D(_00814_),
    .Q_N(_08248_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1409),
    .D(_00815_),
    .Q_N(_08247_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1410),
    .D(_00816_),
    .Q_N(_08246_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1411),
    .D(_00817_),
    .Q_N(_08245_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1412),
    .D(_00818_),
    .Q_N(_08244_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1413),
    .D(_00819_),
    .Q_N(_08243_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1414),
    .D(_00820_),
    .Q_N(_08242_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1415),
    .D(_00821_),
    .Q_N(_08241_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1416),
    .D(_00822_),
    .Q_N(_08240_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1417),
    .D(_00823_),
    .Q_N(_08239_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1418),
    .D(_00824_),
    .Q_N(_08238_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1419),
    .D(_00825_),
    .Q_N(_08237_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1420),
    .D(_00826_),
    .Q_N(_08236_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1421),
    .D(_00827_),
    .Q_N(_08235_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1422),
    .D(_00828_),
    .Q_N(_08234_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1423),
    .D(_00829_),
    .Q_N(_08233_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1424),
    .D(_00830_),
    .Q_N(_08232_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1425),
    .D(_00831_),
    .Q_N(_08231_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1426),
    .D(_00832_),
    .Q_N(_08230_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1427),
    .D(_00833_),
    .Q_N(_08229_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1428),
    .D(_00834_),
    .Q_N(_08228_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1429),
    .D(_00835_),
    .Q_N(_08227_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1430),
    .D(_00836_),
    .Q_N(_08226_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1431),
    .D(_00837_),
    .Q_N(_08225_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1432),
    .D(_00838_),
    .Q_N(_08224_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1433),
    .D(_00839_),
    .Q_N(_08223_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1434),
    .D(_00840_),
    .Q_N(_08222_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1435),
    .D(_00841_),
    .Q_N(_08221_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1436),
    .D(_00842_),
    .Q_N(_08220_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1437),
    .D(_00843_),
    .Q_N(_08219_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1438),
    .D(_00844_),
    .Q_N(_08218_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1439),
    .D(_00845_),
    .Q_N(_08217_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1440),
    .D(_00846_),
    .Q_N(_08216_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1441),
    .D(_00847_),
    .Q_N(_08215_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1442),
    .D(_00848_),
    .Q_N(_08214_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1443),
    .D(_00849_),
    .Q_N(_08213_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1444),
    .D(_00850_),
    .Q_N(_08212_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1445),
    .D(_00851_),
    .Q_N(_08211_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1446),
    .D(_00852_),
    .Q_N(_08210_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1447),
    .D(_00853_),
    .Q_N(_08209_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1448),
    .D(_00854_),
    .Q_N(_08208_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1449),
    .D(_00855_),
    .Q_N(_08207_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1450),
    .D(_00856_),
    .Q_N(_08206_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1451),
    .D(_00857_),
    .Q_N(_08205_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1452),
    .D(_00858_),
    .Q_N(_08204_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1453),
    .D(_00859_),
    .Q_N(_08203_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1454),
    .D(_00860_),
    .Q_N(_08202_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1455),
    .D(_00861_),
    .Q_N(_08201_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1456),
    .D(_00862_),
    .Q_N(_08200_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1457),
    .D(_00863_),
    .Q_N(_08199_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1458),
    .D(_00864_),
    .Q_N(_08198_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1459),
    .D(_00865_),
    .Q_N(_08197_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1460),
    .D(_00866_),
    .Q_N(_08196_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1461),
    .D(_00867_),
    .Q_N(_08195_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1462),
    .D(_00868_),
    .Q_N(_08194_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1463),
    .D(_00869_),
    .Q_N(_08193_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1464),
    .D(_00870_),
    .Q_N(_08192_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1465),
    .D(_00871_),
    .Q_N(_08191_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1466),
    .D(_00872_),
    .Q_N(_08190_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1467),
    .D(_00873_),
    .Q_N(_08189_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1468),
    .D(_00874_),
    .Q_N(_08188_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1469),
    .D(_00875_),
    .Q_N(_08187_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1470),
    .D(_00876_),
    .Q_N(_08186_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1471),
    .D(_00877_),
    .Q_N(_08185_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1472),
    .D(_00878_),
    .Q_N(_08184_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1473),
    .D(_00879_),
    .Q_N(_08183_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1474),
    .D(_00880_),
    .Q_N(_08182_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1475),
    .D(_00881_),
    .Q_N(_08181_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1476),
    .D(_00882_),
    .Q_N(_08180_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1477),
    .D(_00883_),
    .Q_N(_08179_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1478),
    .D(_00884_),
    .Q_N(_08178_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1479),
    .D(_00885_),
    .Q_N(_08177_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1480),
    .D(_00886_),
    .Q_N(_08176_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1481),
    .D(_00887_),
    .Q_N(_08175_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1482),
    .D(_00888_),
    .Q_N(_08174_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1483),
    .D(_00889_),
    .Q_N(_08173_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1484),
    .D(_00890_),
    .Q_N(_08172_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1485),
    .D(_00891_),
    .Q_N(_08171_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1486),
    .D(_00892_),
    .Q_N(_08170_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1487),
    .D(_00893_),
    .Q_N(_08169_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1488),
    .D(_00894_),
    .Q_N(_08168_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1489),
    .D(_00895_),
    .Q_N(_08167_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1490),
    .D(_00896_),
    .Q_N(_08166_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1491),
    .D(_00897_),
    .Q_N(_08165_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1492),
    .D(_00898_),
    .Q_N(_08164_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1493),
    .D(_00899_),
    .Q_N(_08163_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1494),
    .D(_00900_),
    .Q_N(_08162_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1495),
    .D(_00901_),
    .Q_N(_08161_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1496),
    .D(_00902_),
    .Q_N(_08160_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1497),
    .D(_00903_),
    .Q_N(_08159_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1498),
    .D(_00904_),
    .Q_N(_08158_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ));
 sg13g2_dfrbp_1 \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1499),
    .D(_00905_),
    .Q_N(_08157_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pcm[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1500),
    .D(_00906_),
    .Q_N(_08156_),
    .Q(\soc_I.pwm_I.pcm[0] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pcm[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1501),
    .D(_00907_),
    .Q_N(_08155_),
    .Q(\soc_I.pwm_I.pcm[1] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pcm[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1502),
    .D(_00908_),
    .Q_N(_08154_),
    .Q(\soc_I.pwm_I.pcm[2] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pcm[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1503),
    .D(_00909_),
    .Q_N(_08153_),
    .Q(\soc_I.pwm_I.pcm[3] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pcm[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1504),
    .D(_00910_),
    .Q_N(_08152_),
    .Q(\soc_I.pwm_I.pcm[4] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pcm[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1505),
    .D(_00911_),
    .Q_N(_08151_),
    .Q(\soc_I.pwm_I.pcm[5] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pcm[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1506),
    .D(_00912_),
    .Q_N(_08150_),
    .Q(\soc_I.pwm_I.pcm[6] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pcm[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1507),
    .D(_00913_),
    .Q_N(_08149_),
    .Q(\soc_I.pwm_I.pcm[7] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pwm_accumulator[0]$_SDFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1508),
    .D(_00914_),
    .Q_N(_08148_),
    .Q(\soc_I.pwm_I.pwm_accumulator[0] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pwm_accumulator[1]$_SDFF_PN0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1509),
    .D(_00915_),
    .Q_N(_08147_),
    .Q(\soc_I.pwm_I.pwm_accumulator[1] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pwm_accumulator[2]$_SDFF_PN0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1510),
    .D(_00916_),
    .Q_N(_08146_),
    .Q(\soc_I.pwm_I.pwm_accumulator[2] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pwm_accumulator[3]$_SDFF_PN0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1511),
    .D(_00917_),
    .Q_N(_08145_),
    .Q(\soc_I.pwm_I.pwm_accumulator[3] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pwm_accumulator[4]$_SDFF_PN0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1512),
    .D(_00918_),
    .Q_N(_08144_),
    .Q(\soc_I.pwm_I.pwm_accumulator[4] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pwm_accumulator[5]$_SDFF_PN0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1513),
    .D(_00919_),
    .Q_N(_08143_),
    .Q(\soc_I.pwm_I.pwm_accumulator[5] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pwm_accumulator[6]$_SDFF_PN0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1514),
    .D(_00920_),
    .Q_N(_08142_),
    .Q(\soc_I.pwm_I.pwm_accumulator[6] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pwm_accumulator[7]$_SDFF_PN0_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1515),
    .D(_00921_),
    .Q_N(_08141_),
    .Q(\soc_I.pwm_I.pwm_accumulator[7] ));
 sg13g2_dfrbp_1 \soc_I.pwm_I.pwm_accumulator[8]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1516),
    .D(_00922_),
    .Q_N(_08140_),
    .Q(pwm_o));
 sg13g2_dfrbp_1 \soc_I.pwm_ready$_SDFF_PN0_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1517),
    .D(_00923_),
    .Q_N(_08139_),
    .Q(\soc_I.pwm_ready ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.ce[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1518),
    .D(_00924_),
    .Q_N(_08138_),
    .Q(net12));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.ce[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1519),
    .D(_00925_),
    .Q_N(_08137_),
    .Q(net18));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.is_quad$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1520),
    .D(_00926_),
    .Q_N(_00051_),
    .Q(\soc_I.qqspi_I.is_quad ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1521),
    .D(_00927_),
    .Q_N(_08136_),
    .Q(\soc_I.qqspi_I.rdata[0] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1522),
    .D(_00928_),
    .Q_N(_08135_),
    .Q(\soc_I.qqspi_I.rdata[10] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1523),
    .D(_00929_),
    .Q_N(_08134_),
    .Q(\soc_I.qqspi_I.rdata[11] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1524),
    .D(_00930_),
    .Q_N(_08133_),
    .Q(\soc_I.qqspi_I.rdata[12] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1525),
    .D(_00931_),
    .Q_N(_08132_),
    .Q(\soc_I.qqspi_I.rdata[13] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1526),
    .D(_00932_),
    .Q_N(_08131_),
    .Q(\soc_I.qqspi_I.rdata[14] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1527),
    .D(_00933_),
    .Q_N(_08130_),
    .Q(\soc_I.qqspi_I.rdata[15] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[16]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1528),
    .D(_00934_),
    .Q_N(_08129_),
    .Q(\soc_I.qqspi_I.rdata[16] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[17]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1529),
    .D(_00935_),
    .Q_N(_08128_),
    .Q(\soc_I.qqspi_I.rdata[17] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[18]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1530),
    .D(_00936_),
    .Q_N(_08127_),
    .Q(\soc_I.qqspi_I.rdata[18] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[19]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1531),
    .D(_00937_),
    .Q_N(_08126_),
    .Q(\soc_I.qqspi_I.rdata[19] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1532),
    .D(_00938_),
    .Q_N(_08125_),
    .Q(\soc_I.qqspi_I.rdata[1] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[20]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1533),
    .D(_00939_),
    .Q_N(_08124_),
    .Q(\soc_I.qqspi_I.rdata[20] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[21]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1534),
    .D(_00940_),
    .Q_N(_08123_),
    .Q(\soc_I.qqspi_I.rdata[21] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[22]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1535),
    .D(_00941_),
    .Q_N(_08122_),
    .Q(\soc_I.qqspi_I.rdata[22] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[23]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1536),
    .D(_00942_),
    .Q_N(_08121_),
    .Q(\soc_I.qqspi_I.rdata[23] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[24]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1537),
    .D(_00943_),
    .Q_N(_08120_),
    .Q(\soc_I.qqspi_I.rdata[24] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[25]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1538),
    .D(_00944_),
    .Q_N(_08119_),
    .Q(\soc_I.qqspi_I.rdata[25] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[26]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1539),
    .D(_00945_),
    .Q_N(_08118_),
    .Q(\soc_I.qqspi_I.rdata[26] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[27]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1540),
    .D(_00946_),
    .Q_N(_08117_),
    .Q(\soc_I.qqspi_I.rdata[27] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[28]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1541),
    .D(_00947_),
    .Q_N(_08116_),
    .Q(\soc_I.qqspi_I.rdata[28] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[29]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1542),
    .D(_00948_),
    .Q_N(_08115_),
    .Q(\soc_I.qqspi_I.rdata[29] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1543),
    .D(_00949_),
    .Q_N(_08114_),
    .Q(\soc_I.qqspi_I.rdata[2] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[30]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1544),
    .D(_00950_),
    .Q_N(_08113_),
    .Q(\soc_I.qqspi_I.rdata[30] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[31]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1545),
    .D(_00951_),
    .Q_N(_08112_),
    .Q(\soc_I.qqspi_I.rdata[31] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1546),
    .D(_00952_),
    .Q_N(_08111_),
    .Q(\soc_I.qqspi_I.rdata[3] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1547),
    .D(_00953_),
    .Q_N(_08110_),
    .Q(\soc_I.qqspi_I.rdata[4] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1548),
    .D(_00954_),
    .Q_N(_08109_),
    .Q(\soc_I.qqspi_I.rdata[5] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1549),
    .D(_00955_),
    .Q_N(_08108_),
    .Q(\soc_I.qqspi_I.rdata[6] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1550),
    .D(_00956_),
    .Q_N(_08107_),
    .Q(\soc_I.qqspi_I.rdata[7] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1551),
    .D(_00957_),
    .Q_N(_08106_),
    .Q(\soc_I.qqspi_I.rdata[8] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.rdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1552),
    .D(_00958_),
    .Q_N(_08105_),
    .Q(\soc_I.qqspi_I.rdata[9] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.ready$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1553),
    .D(_00959_),
    .Q_N(_00048_),
    .Q(\soc_I.qqspi_I.ready ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.sclk$_SDFFE_PN1N_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1554),
    .D(_00960_),
    .Q_N(_00025_),
    .Q(sclk));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.sio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1555),
    .D(_00961_),
    .Q_N(_08104_),
    .Q(net8));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.sio_oe[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1556),
    .D(_00962_),
    .Q_N(_08103_),
    .Q(net11));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.sio_out[0]$_SDFFE_PN0N_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1557),
    .D(_00963_),
    .Q_N(_08102_),
    .Q(sio0_si_mosi_o));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.sio_out[1]$_SDFFE_PN0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1558),
    .D(_00964_),
    .Q_N(_08101_),
    .Q(sio1_so_miso_o));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.sio_out[2]$_SDFFE_PN0N_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1559),
    .D(_00965_),
    .Q_N(_08100_),
    .Q(sio2_o));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.sio_out[3]$_SDFFE_PN0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1560),
    .D(_00966_),
    .Q_N(_08099_),
    .Q(sio3_o));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1561),
    .D(_00967_),
    .Q_N(_08098_),
    .Q(\soc_I.qqspi_I.spi_buf[0] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1562),
    .D(_00968_),
    .Q_N(_08097_),
    .Q(\soc_I.qqspi_I.spi_buf[10] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1563),
    .D(_00969_),
    .Q_N(_08096_),
    .Q(\soc_I.qqspi_I.spi_buf[11] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1564),
    .D(_00970_),
    .Q_N(_08095_),
    .Q(\soc_I.qqspi_I.spi_buf[12] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1565),
    .D(_00971_),
    .Q_N(_08094_),
    .Q(\soc_I.qqspi_I.spi_buf[13] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1566),
    .D(_00972_),
    .Q_N(_08093_),
    .Q(\soc_I.qqspi_I.spi_buf[14] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1567),
    .D(_00973_),
    .Q_N(_08092_),
    .Q(\soc_I.qqspi_I.spi_buf[15] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1568),
    .D(_00974_),
    .Q_N(_08091_),
    .Q(\soc_I.qqspi_I.spi_buf[16] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1569),
    .D(_00975_),
    .Q_N(_08090_),
    .Q(\soc_I.qqspi_I.spi_buf[17] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1570),
    .D(_00976_),
    .Q_N(_08089_),
    .Q(\soc_I.qqspi_I.spi_buf[18] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1571),
    .D(_00977_),
    .Q_N(_08088_),
    .Q(\soc_I.qqspi_I.spi_buf[19] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1572),
    .D(_00978_),
    .Q_N(_08087_),
    .Q(\soc_I.qqspi_I.spi_buf[1] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1573),
    .D(_00979_),
    .Q_N(_08086_),
    .Q(\soc_I.qqspi_I.spi_buf[20] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1574),
    .D(_00980_),
    .Q_N(_08085_),
    .Q(\soc_I.qqspi_I.spi_buf[21] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1575),
    .D(_00981_),
    .Q_N(_08084_),
    .Q(\soc_I.qqspi_I.spi_buf[22] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1576),
    .D(_00982_),
    .Q_N(_08083_),
    .Q(\soc_I.qqspi_I.spi_buf[23] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1577),
    .D(_00983_),
    .Q_N(_08082_),
    .Q(\soc_I.qqspi_I.spi_buf[24] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1578),
    .D(_00984_),
    .Q_N(_08081_),
    .Q(\soc_I.qqspi_I.spi_buf[25] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1579),
    .D(_00985_),
    .Q_N(_08080_),
    .Q(\soc_I.qqspi_I.spi_buf[26] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1580),
    .D(_00986_),
    .Q_N(_08079_),
    .Q(\soc_I.qqspi_I.spi_buf[27] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1581),
    .D(_00987_),
    .Q_N(_08078_),
    .Q(\soc_I.qqspi_I.spi_buf[28] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1582),
    .D(_00988_),
    .Q_N(_08077_),
    .Q(\soc_I.qqspi_I.spi_buf[29] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1583),
    .D(_00989_),
    .Q_N(_08076_),
    .Q(\soc_I.qqspi_I.spi_buf[2] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1584),
    .D(_00990_),
    .Q_N(_08075_),
    .Q(\soc_I.qqspi_I.spi_buf[30] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1585),
    .D(_00991_),
    .Q_N(_08074_),
    .Q(\soc_I.qqspi_I.spi_buf[31] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1586),
    .D(_00992_),
    .Q_N(_08073_),
    .Q(\soc_I.qqspi_I.spi_buf[3] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1587),
    .D(_00993_),
    .Q_N(_08072_),
    .Q(\soc_I.qqspi_I.spi_buf[4] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1588),
    .D(_00994_),
    .Q_N(_08071_),
    .Q(\soc_I.qqspi_I.spi_buf[5] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1589),
    .D(_00995_),
    .Q_N(_08070_),
    .Q(\soc_I.qqspi_I.spi_buf[6] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1590),
    .D(_00996_),
    .Q_N(_08069_),
    .Q(\soc_I.qqspi_I.spi_buf[7] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1591),
    .D(_00997_),
    .Q_N(_08068_),
    .Q(\soc_I.qqspi_I.spi_buf[8] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.spi_buf[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1592),
    .D(_00998_),
    .Q_N(_08983_),
    .Q(\soc_I.qqspi_I.spi_buf[9] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.state[0]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1593),
    .D(_00018_),
    .Q_N(_00055_),
    .Q(\soc_I.qqspi_I.state[0] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.state[1]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1594),
    .D(_00019_),
    .Q_N(_08984_),
    .Q(\soc_I.qqspi_I.state[1] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.state[2]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1595),
    .D(_00020_),
    .Q_N(_08985_),
    .Q(\soc_I.qqspi_I.state[2] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.state[3]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1596),
    .D(_00021_),
    .Q_N(_00056_),
    .Q(\soc_I.qqspi_I.state[3] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.state[4]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1597),
    .D(_00022_),
    .Q_N(_08986_),
    .Q(\soc_I.qqspi_I.state[4] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.state[5]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1598),
    .D(_00023_),
    .Q_N(_00082_),
    .Q(\soc_I.qqspi_I.state[5] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.state[6]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1599),
    .D(_00024_),
    .Q_N(_00081_),
    .Q(\soc_I.qqspi_I.state[6] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.xfer_cycles[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1600),
    .D(_00999_),
    .Q_N(_08067_),
    .Q(\soc_I.qqspi_I.xfer_cycles[0] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.xfer_cycles[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1601),
    .D(_01000_),
    .Q_N(_08066_),
    .Q(\soc_I.qqspi_I.xfer_cycles[1] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.xfer_cycles[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1602),
    .D(_01001_),
    .Q_N(_00085_),
    .Q(\soc_I.qqspi_I.xfer_cycles[2] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.xfer_cycles[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1603),
    .D(_01002_),
    .Q_N(_08065_),
    .Q(\soc_I.qqspi_I.xfer_cycles[3] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.xfer_cycles[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1604),
    .D(_01003_),
    .Q_N(_08064_),
    .Q(\soc_I.qqspi_I.xfer_cycles[4] ));
 sg13g2_dfrbp_1 \soc_I.qqspi_I.xfer_cycles[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1605),
    .D(_01004_),
    .Q_N(_08063_),
    .Q(\soc_I.qqspi_I.xfer_cycles[5] ));
 sg13g2_dfrbp_1 \soc_I.rst_cnt[0]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1606),
    .D(_01005_),
    .Q_N(_08062_),
    .Q(\soc_I.rst_cnt[0] ));
 sg13g2_dfrbp_1 \soc_I.rst_cnt[1]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1607),
    .D(_01006_),
    .Q_N(_08061_),
    .Q(\soc_I.rst_cnt[1] ));
 sg13g2_dfrbp_1 \soc_I.rst_cnt[2]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1608),
    .D(_01007_),
    .Q_N(_08060_),
    .Q(\soc_I.rst_cnt[2] ));
 sg13g2_dfrbp_1 \soc_I.rst_cnt[3]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1609),
    .D(_01008_),
    .Q_N(_00057_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.resetn ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.bit_idx[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1610),
    .D(_01009_),
    .Q_N(_00088_),
    .Q(\soc_I.rx_uart_i.bit_idx[0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.bit_idx[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1611),
    .D(_01010_),
    .Q_N(_08059_),
    .Q(\soc_I.rx_uart_i.bit_idx[1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.bit_idx[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1612),
    .D(_01011_),
    .Q_N(_08058_),
    .Q(\soc_I.rx_uart_i.bit_idx[2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.cnt[0]$_SDFF_PN0_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1613),
    .D(_01012_),
    .Q_N(_00084_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.cnt[1]$_SDFF_PN0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1614),
    .D(_01013_),
    .Q_N(_08057_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.cnt[2]$_SDFF_PN0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1615),
    .D(_01014_),
    .Q_N(_08056_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.cnt[3]$_SDFF_PN0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1616),
    .D(_01015_),
    .Q_N(_08055_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.cnt[4]$_SDFF_PN0_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1617),
    .D(_01016_),
    .Q_N(_08054_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1618),
    .D(_01017_),
    .Q_N(_08053_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1619),
    .D(_01018_),
    .Q_N(_08052_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1620),
    .D(_01019_),
    .Q_N(_08051_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1621),
    .D(_01020_),
    .Q_N(_08050_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1622),
    .D(_01021_),
    .Q_N(_08049_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1623),
    .D(_01022_),
    .Q_N(_08048_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1624),
    .D(_01023_),
    .Q_N(_08047_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1625),
    .D(_01024_),
    .Q_N(_08046_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1626),
    .D(_01025_),
    .Q_N(_08045_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1627),
    .D(_01026_),
    .Q_N(_08044_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1628),
    .D(_01027_),
    .Q_N(_08043_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1629),
    .D(_01028_),
    .Q_N(_08042_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1630),
    .D(_01029_),
    .Q_N(_08041_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1631),
    .D(_01030_),
    .Q_N(_08040_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1632),
    .D(_01031_),
    .Q_N(_08039_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1633),
    .D(_01032_),
    .Q_N(_08038_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1634),
    .D(_01033_),
    .Q_N(_08037_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1635),
    .D(_01034_),
    .Q_N(_08036_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1636),
    .D(_01035_),
    .Q_N(_08035_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1637),
    .D(_01036_),
    .Q_N(_08034_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1638),
    .D(_01037_),
    .Q_N(_08033_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1639),
    .D(_01038_),
    .Q_N(_08032_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1640),
    .D(_01039_),
    .Q_N(_08031_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1641),
    .D(_01040_),
    .Q_N(_08030_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1642),
    .D(_01041_),
    .Q_N(_08029_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1643),
    .D(_01042_),
    .Q_N(_08028_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1644),
    .D(_01043_),
    .Q_N(_08027_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1645),
    .D(_01044_),
    .Q_N(_08026_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1646),
    .D(_01045_),
    .Q_N(_08025_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1647),
    .D(_01046_),
    .Q_N(_08024_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1648),
    .D(_01047_),
    .Q_N(_08023_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1649),
    .D(_01048_),
    .Q_N(_08022_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1650),
    .D(_01049_),
    .Q_N(_08021_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1651),
    .D(_01050_),
    .Q_N(_08020_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1652),
    .D(_01051_),
    .Q_N(_08019_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1653),
    .D(_01052_),
    .Q_N(_08018_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1654),
    .D(_01053_),
    .Q_N(_08017_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1655),
    .D(_01054_),
    .Q_N(_08016_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1656),
    .D(_01055_),
    .Q_N(_08015_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1657),
    .D(_01056_),
    .Q_N(_08014_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1658),
    .D(_01057_),
    .Q_N(_08013_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1659),
    .D(_01058_),
    .Q_N(_08012_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1660),
    .D(_01059_),
    .Q_N(_08011_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1661),
    .D(_01060_),
    .Q_N(_08010_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1662),
    .D(_01061_),
    .Q_N(_08009_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1663),
    .D(_01062_),
    .Q_N(_08008_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1664),
    .D(_01063_),
    .Q_N(_08007_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1665),
    .D(_01064_),
    .Q_N(_08006_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1666),
    .D(_01065_),
    .Q_N(_08005_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1667),
    .D(_01066_),
    .Q_N(_08004_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1668),
    .D(_01067_),
    .Q_N(_08003_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1669),
    .D(_01068_),
    .Q_N(_08002_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1670),
    .D(_01069_),
    .Q_N(_08001_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1671),
    .D(_01070_),
    .Q_N(_08000_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1672),
    .D(_01071_),
    .Q_N(_07999_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1673),
    .D(_01072_),
    .Q_N(_07998_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1674),
    .D(_01073_),
    .Q_N(_07997_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1675),
    .D(_01074_),
    .Q_N(_07996_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1676),
    .D(_01075_),
    .Q_N(_07995_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1677),
    .D(_01076_),
    .Q_N(_07994_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1678),
    .D(_01077_),
    .Q_N(_07993_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1679),
    .D(_01078_),
    .Q_N(_07992_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1680),
    .D(_01079_),
    .Q_N(_07991_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1681),
    .D(_01080_),
    .Q_N(_07990_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1682),
    .D(_01081_),
    .Q_N(_07989_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1683),
    .D(_01082_),
    .Q_N(_07988_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1684),
    .D(_01083_),
    .Q_N(_07987_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1685),
    .D(_01084_),
    .Q_N(_07986_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1686),
    .D(_01085_),
    .Q_N(_07985_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1687),
    .D(_01086_),
    .Q_N(_07984_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1688),
    .D(_01087_),
    .Q_N(_07983_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1689),
    .D(_01088_),
    .Q_N(_07982_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1690),
    .D(_01089_),
    .Q_N(_07981_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1691),
    .D(_01090_),
    .Q_N(_07980_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1692),
    .D(_01091_),
    .Q_N(_07979_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1693),
    .D(_01092_),
    .Q_N(_07978_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1694),
    .D(_01093_),
    .Q_N(_07977_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1695),
    .D(_01094_),
    .Q_N(_07976_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1696),
    .D(_01095_),
    .Q_N(_07975_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1697),
    .D(_01096_),
    .Q_N(_07974_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1698),
    .D(_01097_),
    .Q_N(_07973_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1699),
    .D(_01098_),
    .Q_N(_07972_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1700),
    .D(_01099_),
    .Q_N(_07971_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1701),
    .D(_01100_),
    .Q_N(_07970_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1702),
    .D(_01101_),
    .Q_N(_07969_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1703),
    .D(_01102_),
    .Q_N(_07968_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1704),
    .D(_01103_),
    .Q_N(_07967_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1705),
    .D(_01104_),
    .Q_N(_07966_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1706),
    .D(_01105_),
    .Q_N(_07965_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1707),
    .D(_01106_),
    .Q_N(_07964_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1708),
    .D(_01107_),
    .Q_N(_07963_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1709),
    .D(_01108_),
    .Q_N(_07962_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1710),
    .D(_01109_),
    .Q_N(_07961_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1711),
    .D(_01110_),
    .Q_N(_07960_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1712),
    .D(_01111_),
    .Q_N(_07959_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1713),
    .D(_01112_),
    .Q_N(_07958_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1714),
    .D(_01113_),
    .Q_N(_07957_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1715),
    .D(_01114_),
    .Q_N(_07956_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1716),
    .D(_01115_),
    .Q_N(_07955_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1717),
    .D(_01116_),
    .Q_N(_07954_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1718),
    .D(_01117_),
    .Q_N(_07953_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1719),
    .D(_01118_),
    .Q_N(_07952_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1720),
    .D(_01119_),
    .Q_N(_07951_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1721),
    .D(_01120_),
    .Q_N(_07950_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1722),
    .D(_01121_),
    .Q_N(_07949_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1723),
    .D(_01122_),
    .Q_N(_07948_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1724),
    .D(_01123_),
    .Q_N(_07947_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1725),
    .D(_01124_),
    .Q_N(_07946_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1726),
    .D(_01125_),
    .Q_N(_07945_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1727),
    .D(_01126_),
    .Q_N(_07944_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1728),
    .D(_01127_),
    .Q_N(_07943_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1729),
    .D(_01128_),
    .Q_N(_07942_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1730),
    .D(_01129_),
    .Q_N(_07941_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1731),
    .D(_01130_),
    .Q_N(_07940_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1732),
    .D(_01131_),
    .Q_N(_07939_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1733),
    .D(_01132_),
    .Q_N(_07938_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1734),
    .D(_01133_),
    .Q_N(_07937_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1735),
    .D(_01134_),
    .Q_N(_07936_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1736),
    .D(_01135_),
    .Q_N(_07935_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1737),
    .D(_01136_),
    .Q_N(_07934_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1738),
    .D(_01137_),
    .Q_N(_07933_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1739),
    .D(_01138_),
    .Q_N(_07932_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1740),
    .D(_01139_),
    .Q_N(_07931_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1741),
    .D(_01140_),
    .Q_N(_07930_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1742),
    .D(_01141_),
    .Q_N(_07929_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1743),
    .D(_01142_),
    .Q_N(_07928_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1744),
    .D(_01143_),
    .Q_N(_07927_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.ram[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1745),
    .D(_01144_),
    .Q_N(_07926_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.rd_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1746),
    .D(_01145_),
    .Q_N(_00090_),
    .Q(\soc_I.rx_uart_i.fifo_i.rd_ptr[0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.rd_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1747),
    .D(_00094_),
    .Q_N(_07925_),
    .Q(\soc_I.rx_uart_i.fifo_i.rd_ptr[1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.rd_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1748),
    .D(_00095_),
    .Q_N(_07924_),
    .Q(\soc_I.rx_uart_i.fifo_i.rd_ptr[2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.rd_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1749),
    .D(_00096_),
    .Q_N(_07923_),
    .Q(\soc_I.rx_uart_i.fifo_i.rd_ptr[3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.wr_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1750),
    .D(_01146_),
    .Q_N(_00089_),
    .Q(\soc_I.rx_uart_i.fifo_i.wr_ptr[0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.wr_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1751),
    .D(_01147_),
    .Q_N(_07922_),
    .Q(\soc_I.rx_uart_i.fifo_i.wr_ptr[1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.wr_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1752),
    .D(_01148_),
    .Q_N(_07921_),
    .Q(\soc_I.rx_uart_i.fifo_i.wr_ptr[2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.fifo_i.wr_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1753),
    .D(_01149_),
    .Q_N(_07920_),
    .Q(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.ready$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1754),
    .D(_01150_),
    .Q_N(_07919_),
    .Q(\soc_I.rx_uart_i.ready ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.return_state[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1755),
    .D(_01151_),
    .Q_N(_07918_),
    .Q(\soc_I.rx_uart_i.return_state[0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.return_state[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1756),
    .D(_01152_),
    .Q_N(_07917_),
    .Q(\soc_I.rx_uart_i.return_state[1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_data[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1757),
    .D(_01153_),
    .Q_N(_07916_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_data[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1758),
    .D(_01154_),
    .Q_N(_07915_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_data[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1759),
    .D(_01155_),
    .Q_N(_07914_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_data[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1760),
    .D(_01156_),
    .Q_N(_07913_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_data[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1761),
    .D(_01157_),
    .Q_N(_07912_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_data[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1762),
    .D(_01158_),
    .Q_N(_07911_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_data[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1763),
    .D(_01159_),
    .Q_N(_07910_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_data[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1764),
    .D(_01160_),
    .Q_N(_07909_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_in_sync[0]$_SDFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1765),
    .D(_01161_),
    .Q_N(_07908_),
    .Q(\soc_I.rx_uart_i.rx_in_sync[0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_in_sync[1]$_SDFF_PN0_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1766),
    .D(_01162_),
    .Q_N(_07907_),
    .Q(\soc_I.rx_uart_i.rx_in_sync[1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.rx_in_sync[2]$_SDFF_PN0_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1767),
    .D(_01163_),
    .Q_N(_00059_),
    .Q(\soc_I.rx_uart_i.rx_in_sync[2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1768),
    .D(_01164_),
    .Q_N(_07906_),
    .Q(\soc_I.rx_uart_i.state[0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1769),
    .D(_01165_),
    .Q_N(_07905_),
    .Q(\soc_I.rx_uart_i.state[1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1770),
    .D(_01166_),
    .Q_N(_00047_),
    .Q(\soc_I.rx_uart_i.state[2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1771),
    .D(_01167_),
    .Q_N(_07904_),
    .Q(\soc_I.rx_uart_i.wait_states[0] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1772),
    .D(_01168_),
    .Q_N(_07903_),
    .Q(\soc_I.rx_uart_i.wait_states[10] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1773),
    .D(_01169_),
    .Q_N(_07902_),
    .Q(\soc_I.rx_uart_i.wait_states[11] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1774),
    .D(_01170_),
    .Q_N(_07901_),
    .Q(\soc_I.rx_uart_i.wait_states[12] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1775),
    .D(_01171_),
    .Q_N(_07900_),
    .Q(\soc_I.rx_uart_i.wait_states[13] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1776),
    .D(_01172_),
    .Q_N(_07899_),
    .Q(\soc_I.rx_uart_i.wait_states[14] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1777),
    .D(_01173_),
    .Q_N(_07898_),
    .Q(\soc_I.rx_uart_i.wait_states[15] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1778),
    .D(_01174_),
    .Q_N(_00054_),
    .Q(\soc_I.rx_uart_i.wait_states[16] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1779),
    .D(_01175_),
    .Q_N(_07897_),
    .Q(\soc_I.rx_uart_i.wait_states[1] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1780),
    .D(_01176_),
    .Q_N(_07896_),
    .Q(\soc_I.rx_uart_i.wait_states[2] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1781),
    .D(_01177_),
    .Q_N(_07895_),
    .Q(\soc_I.rx_uart_i.wait_states[3] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1782),
    .D(_01178_),
    .Q_N(_07894_),
    .Q(\soc_I.rx_uart_i.wait_states[4] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1783),
    .D(_01179_),
    .Q_N(_07893_),
    .Q(\soc_I.rx_uart_i.wait_states[5] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1784),
    .D(_01180_),
    .Q_N(_07892_),
    .Q(\soc_I.rx_uart_i.wait_states[6] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1785),
    .D(_01181_),
    .Q_N(_07891_),
    .Q(\soc_I.rx_uart_i.wait_states[7] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1786),
    .D(_01182_),
    .Q_N(_07890_),
    .Q(\soc_I.rx_uart_i.wait_states[8] ));
 sg13g2_dfrbp_1 \soc_I.rx_uart_i.wait_states[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1787),
    .D(_01183_),
    .Q_N(_07889_),
    .Q(\soc_I.rx_uart_i.wait_states[9] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.ready_ctrl$_SDFF_PN0_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1788),
    .D(_01184_),
    .Q_N(_07888_),
    .Q(\soc_I.spi0_I.ready_ctrl ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.ready_xfer$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1789),
    .D(_01185_),
    .Q_N(_07887_),
    .Q(\soc_I.spi0_I.ready_xfer ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.rx_data[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1790),
    .D(_01186_),
    .Q_N(_00063_),
    .Q(\soc_I.spi0_I.rx_data[0] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.rx_data[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1791),
    .D(_01187_),
    .Q_N(_07886_),
    .Q(\soc_I.spi0_I.rx_data[1] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.rx_data[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1792),
    .D(_01188_),
    .Q_N(_07885_),
    .Q(\soc_I.spi0_I.rx_data[2] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.rx_data[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1793),
    .D(_01189_),
    .Q_N(_07884_),
    .Q(\soc_I.spi0_I.rx_data[3] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.rx_data[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1794),
    .D(_01190_),
    .Q_N(_07883_),
    .Q(\soc_I.spi0_I.rx_data[4] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.rx_data[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1795),
    .D(_01191_),
    .Q_N(_07882_),
    .Q(\soc_I.spi0_I.rx_data[5] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.rx_data[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1796),
    .D(_01192_),
    .Q_N(_07881_),
    .Q(\soc_I.spi0_I.rx_data[6] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.rx_data[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1797),
    .D(_01193_),
    .Q_N(_07880_),
    .Q(\soc_I.spi0_I.rx_data[7] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.sclk$_SDFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1798),
    .D(_01194_),
    .Q_N(_00058_),
    .Q(\soc_I.spi0_I.sclk ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.sio_out$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1799),
    .D(_01195_),
    .Q_N(_07879_),
    .Q(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.spi_buf[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1800),
    .D(_01196_),
    .Q_N(_07878_),
    .Q(\soc_I.spi0_I.spi_buf[0] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.spi_buf[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1801),
    .D(_01197_),
    .Q_N(_07877_),
    .Q(\soc_I.spi0_I.spi_buf[1] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.spi_buf[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1802),
    .D(_01198_),
    .Q_N(_07876_),
    .Q(\soc_I.spi0_I.spi_buf[2] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.spi_buf[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1803),
    .D(_01199_),
    .Q_N(_07875_),
    .Q(\soc_I.spi0_I.spi_buf[3] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.spi_buf[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1804),
    .D(_01200_),
    .Q_N(_07874_),
    .Q(\soc_I.spi0_I.spi_buf[4] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.spi_buf[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1805),
    .D(_01201_),
    .Q_N(_07873_),
    .Q(\soc_I.spi0_I.spi_buf[5] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.spi_buf[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1806),
    .D(_01202_),
    .Q_N(_07872_),
    .Q(\soc_I.spi0_I.spi_buf[6] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.spi_buf[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1807),
    .D(_01203_),
    .Q_N(_07871_),
    .Q(\soc_I.spi0_I.spi_buf[7] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.spi_cen$_SDFFE_PN1P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1808),
    .D(_01204_),
    .Q_N(_00062_),
    .Q(\soc_I.spi0_I.cen ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.state$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1809),
    .D(_01205_),
    .Q_N(_07870_),
    .Q(\soc_I.spi0_I.state ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1810),
    .D(_01206_),
    .Q_N(_00091_),
    .Q(\soc_I.spi0_I.tick_cnt[0] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1811),
    .D(_01207_),
    .Q_N(_07869_),
    .Q(\soc_I.spi0_I.tick_cnt[10] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[11]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1812),
    .D(_01208_),
    .Q_N(_07868_),
    .Q(\soc_I.spi0_I.tick_cnt[11] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[12]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1813),
    .D(_01209_),
    .Q_N(_07867_),
    .Q(\soc_I.spi0_I.tick_cnt[12] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[13]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1814),
    .D(_01210_),
    .Q_N(_07866_),
    .Q(\soc_I.spi0_I.tick_cnt[13] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[14]$_SDFFE_PP0N_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1815),
    .D(_01211_),
    .Q_N(_07865_),
    .Q(\soc_I.spi0_I.tick_cnt[14] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[15]$_SDFFE_PP0N_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1816),
    .D(_01212_),
    .Q_N(_07864_),
    .Q(\soc_I.spi0_I.tick_cnt[15] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[16]$_SDFFE_PP0N_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1817),
    .D(_01213_),
    .Q_N(_07863_),
    .Q(\soc_I.spi0_I.tick_cnt[16] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[17]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1818),
    .D(_01214_),
    .Q_N(_07862_),
    .Q(\soc_I.spi0_I.tick_cnt[17] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1819),
    .D(_01215_),
    .Q_N(_07861_),
    .Q(\soc_I.spi0_I.tick_cnt[1] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1820),
    .D(_01216_),
    .Q_N(_07860_),
    .Q(\soc_I.spi0_I.tick_cnt[2] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1821),
    .D(_01217_),
    .Q_N(_07859_),
    .Q(\soc_I.spi0_I.tick_cnt[3] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1822),
    .D(_01218_),
    .Q_N(_07858_),
    .Q(\soc_I.spi0_I.tick_cnt[4] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1823),
    .D(_01219_),
    .Q_N(_07857_),
    .Q(\soc_I.spi0_I.tick_cnt[5] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1824),
    .D(_01220_),
    .Q_N(_07856_),
    .Q(\soc_I.spi0_I.tick_cnt[6] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1825),
    .D(_01221_),
    .Q_N(_07855_),
    .Q(\soc_I.spi0_I.tick_cnt[7] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1826),
    .D(_01222_),
    .Q_N(_07854_),
    .Q(\soc_I.spi0_I.tick_cnt[8] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.tick_cnt[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1827),
    .D(_01223_),
    .Q_N(_07853_),
    .Q(\soc_I.spi0_I.tick_cnt[9] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.xfer_cycles[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1828),
    .D(_01224_),
    .Q_N(_07852_),
    .Q(\soc_I.spi0_I.xfer_cycles[0] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.xfer_cycles[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1829),
    .D(_01225_),
    .Q_N(_07851_),
    .Q(\soc_I.spi0_I.xfer_cycles[1] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.xfer_cycles[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1830),
    .D(_01226_),
    .Q_N(_07850_),
    .Q(\soc_I.spi0_I.xfer_cycles[2] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.xfer_cycles[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1831),
    .D(_01227_),
    .Q_N(_07849_),
    .Q(\soc_I.spi0_I.xfer_cycles[3] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.xfer_cycles[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1832),
    .D(_01228_),
    .Q_N(_07848_),
    .Q(\soc_I.spi0_I.xfer_cycles[4] ));
 sg13g2_dfrbp_1 \soc_I.spi0_I.xfer_cycles[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1833),
    .D(_01229_),
    .Q_N(_07847_),
    .Q(\soc_I.spi0_I.xfer_cycles[5] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_ready$_SDFF_PN0_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1834),
    .D(_01230_),
    .Q_N(_07846_),
    .Q(\soc_I.spi_div_ready ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1835),
    .D(_01231_),
    .Q_N(_00061_),
    .Q(\soc_I.spi0_I.div[0] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1836),
    .D(_01232_),
    .Q_N(_07845_),
    .Q(\soc_I.spi0_I.div[10] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1837),
    .D(_01233_),
    .Q_N(_07844_),
    .Q(\soc_I.spi0_I.div[11] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1838),
    .D(_01234_),
    .Q_N(_07843_),
    .Q(\soc_I.spi0_I.div[12] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1839),
    .D(_01235_),
    .Q_N(_07842_),
    .Q(\soc_I.spi0_I.div[13] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1840),
    .D(_01236_),
    .Q_N(_07841_),
    .Q(\soc_I.spi0_I.div[14] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1841),
    .D(_01237_),
    .Q_N(_07840_),
    .Q(\soc_I.spi0_I.div[15] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1842),
    .D(_01238_),
    .Q_N(_07839_),
    .Q(\soc_I.spi_div_reg[16] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1843),
    .D(_01239_),
    .Q_N(_07838_),
    .Q(\soc_I.spi_div_reg[17] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1844),
    .D(_01240_),
    .Q_N(_07837_),
    .Q(\soc_I.spi_div_reg[18] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1845),
    .D(_01241_),
    .Q_N(_07836_),
    .Q(\soc_I.spi_div_reg[19] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1846),
    .D(_01242_),
    .Q_N(_00065_),
    .Q(\soc_I.spi0_I.div[1] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1847),
    .D(_01243_),
    .Q_N(_07835_),
    .Q(\soc_I.spi_div_reg[20] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1848),
    .D(_01244_),
    .Q_N(_07834_),
    .Q(\soc_I.spi_div_reg[21] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1849),
    .D(_01245_),
    .Q_N(_07833_),
    .Q(\soc_I.spi_div_reg[22] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1850),
    .D(_01246_),
    .Q_N(_07832_),
    .Q(\soc_I.spi_div_reg[23] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1851),
    .D(_01247_),
    .Q_N(_07831_),
    .Q(\soc_I.spi_div_reg[24] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1852),
    .D(_01248_),
    .Q_N(_07830_),
    .Q(\soc_I.spi_div_reg[25] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1853),
    .D(_01249_),
    .Q_N(_07829_),
    .Q(\soc_I.spi_div_reg[26] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1854),
    .D(_01250_),
    .Q_N(_07828_),
    .Q(\soc_I.spi_div_reg[27] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1855),
    .D(_01251_),
    .Q_N(_07827_),
    .Q(\soc_I.spi_div_reg[28] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1856),
    .D(_01252_),
    .Q_N(_07826_),
    .Q(\soc_I.spi_div_reg[29] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1857),
    .D(_01253_),
    .Q_N(_00067_),
    .Q(\soc_I.spi0_I.div[2] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1858),
    .D(_01254_),
    .Q_N(_07825_),
    .Q(\soc_I.spi_div_reg[30] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1859),
    .D(_01255_),
    .Q_N(_00079_),
    .Q(\soc_I.spi_div_reg[31] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1860),
    .D(_01256_),
    .Q_N(_00069_),
    .Q(\soc_I.spi0_I.div[3] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1861),
    .D(_01257_),
    .Q_N(_00071_),
    .Q(\soc_I.spi0_I.div[4] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1862),
    .D(_01258_),
    .Q_N(_00073_),
    .Q(\soc_I.spi0_I.div[5] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1863),
    .D(_01259_),
    .Q_N(_00075_),
    .Q(\soc_I.spi0_I.div[6] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1864),
    .D(_01260_),
    .Q_N(_00077_),
    .Q(\soc_I.spi0_I.div[7] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1865),
    .D(_01261_),
    .Q_N(_07824_),
    .Q(\soc_I.spi0_I.div[8] ));
 sg13g2_dfrbp_1 \soc_I.spi_div_reg[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1866),
    .D(_01262_),
    .Q_N(_07823_),
    .Q(\soc_I.spi0_I.div[9] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.bit_idx[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1867),
    .D(_01263_),
    .Q_N(_00092_),
    .Q(\soc_I.tx_uart_i.bit_idx[0] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.bit_idx[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1868),
    .D(_01264_),
    .Q_N(_07822_),
    .Q(\soc_I.tx_uart_i.bit_idx[1] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.bit_idx[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1869),
    .D(_01265_),
    .Q_N(_00083_),
    .Q(\soc_I.tx_uart_i.bit_idx[2] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.return_state[0]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1870),
    .D(_01266_),
    .Q_N(_07821_),
    .Q(\soc_I.tx_uart_i.return_state[0] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.return_state[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1871),
    .D(_01267_),
    .Q_N(_07820_),
    .Q(\soc_I.tx_uart_i.return_state[1] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1872),
    .D(_01268_),
    .Q_N(_07819_),
    .Q(\soc_I.tx_uart_i.state[0] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1873),
    .D(_01269_),
    .Q_N(_07818_),
    .Q(\soc_I.tx_uart_i.state[1] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.tx_data_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1874),
    .D(_01270_),
    .Q_N(_07817_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[0] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.tx_data_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1875),
    .D(_01271_),
    .Q_N(_07816_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[1] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.tx_data_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1876),
    .D(_01272_),
    .Q_N(_07815_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[2] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.tx_data_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1877),
    .D(_01273_),
    .Q_N(_07814_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[3] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.tx_data_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1878),
    .D(_01274_),
    .Q_N(_07813_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[4] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.tx_data_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1879),
    .D(_01275_),
    .Q_N(_07812_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[5] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.tx_data_reg[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1880),
    .D(_01276_),
    .Q_N(_07811_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[6] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.tx_data_reg[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1881),
    .D(_01277_),
    .Q_N(_07810_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[7] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.tx_out$_SDFFE_PN1N_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1882),
    .D(_01278_),
    .Q_N(_07809_),
    .Q(\soc_I.tx_uart_i.tx_out ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.txfer_done$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1883),
    .D(_01279_),
    .Q_N(_07808_),
    .Q(\soc_I.tx_uart_i.ready ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1884),
    .D(_01280_),
    .Q_N(_07807_),
    .Q(\soc_I.tx_uart_i.wait_states[0] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[10]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1885),
    .D(_01281_),
    .Q_N(_07806_),
    .Q(\soc_I.tx_uart_i.wait_states[10] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[11]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1886),
    .D(_01282_),
    .Q_N(_07805_),
    .Q(\soc_I.tx_uart_i.wait_states[11] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[12]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1887),
    .D(_01283_),
    .Q_N(_07804_),
    .Q(\soc_I.tx_uart_i.wait_states[12] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[13]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1888),
    .D(_01284_),
    .Q_N(_07803_),
    .Q(\soc_I.tx_uart_i.wait_states[13] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[14]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1889),
    .D(_01285_),
    .Q_N(_07802_),
    .Q(\soc_I.tx_uart_i.wait_states[14] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[15]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1890),
    .D(_01286_),
    .Q_N(_07801_),
    .Q(\soc_I.tx_uart_i.wait_states[15] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[1]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1891),
    .D(_01287_),
    .Q_N(_07800_),
    .Q(\soc_I.tx_uart_i.wait_states[1] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[2]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1892),
    .D(_01288_),
    .Q_N(_07799_),
    .Q(\soc_I.tx_uart_i.wait_states[2] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1893),
    .D(_01289_),
    .Q_N(_07798_),
    .Q(\soc_I.tx_uart_i.wait_states[3] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[4]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1894),
    .D(_01290_),
    .Q_N(_07797_),
    .Q(\soc_I.tx_uart_i.wait_states[4] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[5]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1895),
    .D(_01291_),
    .Q_N(_07796_),
    .Q(\soc_I.tx_uart_i.wait_states[5] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[6]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1896),
    .D(_01292_),
    .Q_N(_07795_),
    .Q(\soc_I.tx_uart_i.wait_states[6] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[7]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1897),
    .D(_01293_),
    .Q_N(_07794_),
    .Q(\soc_I.tx_uart_i.wait_states[7] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[8]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1898),
    .D(_01294_),
    .Q_N(_07793_),
    .Q(\soc_I.tx_uart_i.wait_states[8] ));
 sg13g2_dfrbp_1 \soc_I.tx_uart_i.wait_states[9]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1899),
    .D(_01295_),
    .Q_N(_07792_),
    .Q(\soc_I.tx_uart_i.wait_states[9] ));
 sg13g2_dfrbp_1 \soc_I.uart_lsr_rdy$_SDFF_PN0_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1900),
    .D(_01296_),
    .Q_N(_00049_),
    .Q(\soc_I.uart_lsr_rdy ));
 sg13g2_dfrbp_1 \soc_I.uart_rx_ready$_SDFF_PN0_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1901),
    .D(_01297_),
    .Q_N(_00050_),
    .Q(\soc_I.rx_uart_i.data_rd ));
 sg13g2_dfrbp_1 \soc_I.uart_tx_ready$_SDFF_PN0_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1902),
    .D(_01298_),
    .Q_N(_07791_),
    .Q(\soc_I.uart_tx_ready ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[2]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[5]),
    .X(net7));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[1]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[2]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[5]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[0]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[1]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[2]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[4]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[5]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[6]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout27 (.A(_04264_),
    .X(net27));
 sg13g2_buf_1 fanout28 (.A(_01515_),
    .X(net28));
 sg13g2_buf_4 fanout29 (.X(net29),
    .A(_06988_));
 sg13g2_buf_4 fanout30 (.X(net30),
    .A(_06986_));
 sg13g2_buf_2 fanout31 (.A(_06983_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_06944_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_06939_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_06921_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_06916_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_06898_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_06701_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_06693_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_06665_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_06571_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_05981_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_05934_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_05922_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_06759_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_06642_),
    .X(net45));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(_06568_));
 sg13g2_buf_2 fanout47 (.A(_06527_),
    .X(net47));
 sg13g2_buf_1 fanout48 (.A(_05964_),
    .X(net48));
 sg13g2_buf_1 fanout49 (.A(_05920_),
    .X(net49));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(_05916_));
 sg13g2_buf_2 fanout51 (.A(_01370_),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(_01365_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_01346_),
    .X(net53));
 sg13g2_buf_1 fanout54 (.A(_01344_),
    .X(net54));
 sg13g2_buf_4 fanout55 (.X(net55),
    .A(_01342_));
 sg13g2_buf_2 fanout56 (.A(_07778_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_06632_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_05466_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_05465_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_05292_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_05251_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_05236_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_05199_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_05198_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_05275_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_05197_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_06580_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_06492_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_06462_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_06455_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_06453_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_06467_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_06458_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_04356_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_04550_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_03574_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_04635_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_04590_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_04633_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_04627_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_04620_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_04616_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_04607_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_04598_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_04589_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_04581_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_04576_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_04215_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_04674_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_04669_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_04643_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_04641_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_04637_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_04612_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_04610_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_04606_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_04597_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_04580_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_04575_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_04673_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_04668_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_04661_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_04649_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_04647_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_04645_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_04640_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_04614_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_04600_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_04592_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_04565_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_04330_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_04207_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_03650_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_04675_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_04657_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_04604_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_04564_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_03832_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_03804_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_03749_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_03730_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_03714_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_04656_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_04603_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_04583_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_04569_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_04567_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_03888_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_04014_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_03933_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_03917_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_07043_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_04491_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_04489_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_04441_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_04439_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_04398_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_04389_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_03234_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_03231_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_03127_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_03007_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_05754_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_03217_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_03000_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_02914_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_02701_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_02652_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_05753_),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(_03014_));
 sg13g2_buf_2 fanout151 (.A(_02700_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_02685_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_02651_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_03013_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_02684_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_02176_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_01926_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_01758_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_03546_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_02439_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_02180_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_01920_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_01757_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03612_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03545_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_03536_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_02712_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_02030_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_01919_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_01804_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_01756_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_03944_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_03772_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_03549_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_03544_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_03535_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_02623_),
    .X(net177));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(_01918_));
 sg13g2_buf_2 fanout179 (.A(_01803_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_01755_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_03610_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_03548_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_02903_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_02622_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_01786_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_01782_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_01639_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_05176_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_05162_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_05142_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_05128_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_04869_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_04855_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_04835_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_04821_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_04801_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_04787_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_04766_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_04752_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_04730_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_04716_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_04696_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_04682_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_04473_),
    .X(net204));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(_04443_));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(_04394_));
 sg13g2_buf_2 fanout207 (.A(_03541_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_02670_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_02639_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_02621_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_02591_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_01785_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_01771_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_05173_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_05166_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_05163_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_05161_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_05139_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_05132_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_05129_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_05127_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_05108_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_05094_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_05074_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_05060_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_05040_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_05026_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_05006_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_04992_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_04971_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_04957_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_04937_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_04923_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_04903_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_04889_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_04866_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_04859_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_04856_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_04854_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_04832_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_04825_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_04822_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_04820_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_04798_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_04791_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_04788_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_04786_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_04763_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_04756_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_04753_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_04751_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_04727_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_04720_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_04717_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_04715_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_04693_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_04686_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_04683_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_04681_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_04561_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_04558_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_03540_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_03005_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_02625_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_02604_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_02286_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_02243_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_02213_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_02156_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_02140_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_02110_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_02044_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_05105_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_05098_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_05095_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_05093_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_05071_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_05064_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_05061_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_05059_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_05037_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_05030_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_05027_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_05025_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_05003_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_04996_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_04993_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_04991_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_04968_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_04961_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_04958_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_04956_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_04934_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_04927_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_04924_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_04922_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_04900_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_04893_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_04890_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_04888_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_04601_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_04568_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_04559_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_04557_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_02693_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_02493_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_02487_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_02281_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_02085_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_01768_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_07219_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_07195_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_07194_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_02007_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_01623_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_07645_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_07642_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_05290_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_05283_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_05250_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_05245_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_05193_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_02080_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_01978_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_01746_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_01572_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_01503_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_07641_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_07631_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_06534_),
    .X(net330));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(_05405_));
 sg13g2_buf_2 fanout332 (.A(_05203_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_04362_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_04358_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_04313_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_04300_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_01977_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_01941_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_01818_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_01708_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_01680_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_01666_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_01571_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_07744_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_07738_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_07222_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_07221_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_07196_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_06646_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_06554_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_06533_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_06392_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_06331_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_06257_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_06190_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_06129_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_06057_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_04357_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_04323_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_04312_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_04299_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_03538_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_01927_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_01850_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_01828_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_01707_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_01677_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_01586_),
    .X(net368));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(_01582_));
 sg13g2_buf_2 fanout370 (.A(_01570_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_01445_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_01303_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_07753_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_07660_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_07644_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_07575_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_07507_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_07483_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_07252_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_07155_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_07116_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_07056_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_07024_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_07009_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_06963_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_06941_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_06918_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_06802_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_06703_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_06553_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_06522_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_06509_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_06477_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_06003_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_05986_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_05939_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_05936_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_05919_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_05905_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_05891_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_05868_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_05842_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_05803_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_05801_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_05528_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_05475_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_05442_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_05424_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_04551_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_04546_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_04321_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_04298_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_04258_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_03752_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_03537_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_01846_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_01808_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_01672_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_01585_),
    .X(net419));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(_01581_));
 sg13g2_buf_2 fanout421 (.A(_01393_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_01358_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_07613_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_07574_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_07496_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_07144_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_07088_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_07032_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_06748_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_06634_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_06604_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_06531_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_06501_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_05957_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_05909_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_05904_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_05810_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_05802_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_05470_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_05441_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_05423_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_05379_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_04297_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_03657_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_03584_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_03567_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_03565_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_02035_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_01904_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_01866_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_01807_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_01787_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_01700_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_01697_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_01692_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_01683_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_01560_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_01485_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_07228_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_07179_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_07143_),
    .X(net461));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(_06678_));
 sg13g2_buf_8 fanout463 (.A(_06677_),
    .X(net463));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(_06674_));
 sg13g2_buf_8 fanout465 (.A(_06673_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_06666_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_06645_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_06644_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_06626_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_06581_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_06572_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_06549_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_06530_),
    .X(net473));
 sg13g2_buf_4 fanout474 (.X(net474),
    .A(_06385_));
 sg13g2_buf_8 fanout475 (.A(_06384_),
    .X(net475));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(_06372_));
 sg13g2_buf_8 fanout477 (.A(_06371_),
    .X(net477));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(_06324_));
 sg13g2_buf_8 fanout479 (.A(_06323_),
    .X(net479));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(_06311_));
 sg13g2_buf_8 fanout481 (.A(_06310_),
    .X(net481));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(_06302_));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(_06271_));
 sg13g2_buf_8 fanout484 (.A(_06270_),
    .X(net484));
 sg13g2_buf_4 fanout485 (.X(net485),
    .A(_06265_));
 sg13g2_buf_4 fanout486 (.X(net486),
    .A(_06263_));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(_06261_));
 sg13g2_buf_8 fanout488 (.A(_06259_),
    .X(net488));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(_06183_));
 sg13g2_buf_8 fanout490 (.A(_06177_),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(_06170_));
 sg13g2_buf_8 fanout492 (.A(_06164_),
    .X(net492));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(_06122_));
 sg13g2_buf_8 fanout494 (.A(_06116_),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(_06109_));
 sg13g2_buf_8 fanout496 (.A(_06103_),
    .X(net496));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(_06100_));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(_06069_));
 sg13g2_buf_8 fanout499 (.A(_06068_),
    .X(net499));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(_06063_));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(_06060_));
 sg13g2_buf_8 fanout502 (.A(_06058_),
    .X(net502));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(_06053_));
 sg13g2_buf_2 fanout504 (.A(_05996_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_05956_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_05911_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_05903_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_05440_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_04469_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_04468_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_04442_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_04432_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_04403_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_04400_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_04371_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_04309_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_04308_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_04305_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_04304_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_04266_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_03765_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_03602_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_03578_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_03566_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_03564_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_01863_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_01798_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_01644_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_01605_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_01559_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_01442_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_07737_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_07220_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_07197_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_07180_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_07142_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_06560_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_06548_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_06547_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_06538_),
    .X(net540));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(_06536_));
 sg13g2_buf_2 fanout542 (.A(_06529_),
    .X(net542));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(_06390_));
 sg13g2_buf_8 fanout544 (.A(_06389_),
    .X(net544));
 sg13g2_buf_4 fanout545 (.X(net545),
    .A(_06363_));
 sg13g2_buf_8 fanout546 (.A(_06362_),
    .X(net546));
 sg13g2_buf_4 fanout547 (.X(net547),
    .A(_06350_));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(_06349_));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(_06329_));
 sg13g2_buf_8 fanout550 (.A(_06328_),
    .X(net550));
 sg13g2_buf_8 fanout551 (.A(_06301_),
    .X(net551));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(_06289_));
 sg13g2_buf_8 fanout553 (.A(_06288_),
    .X(net553));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_06274_));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(_06273_));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(_06268_));
 sg13g2_buf_8 fanout557 (.A(_06267_),
    .X(net557));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(_06264_));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(_06253_));
 sg13g2_buf_8 fanout560 (.A(_06203_),
    .X(net560));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(_06188_));
 sg13g2_buf_8 fanout562 (.A(_06187_),
    .X(net562));
 sg13g2_buf_4 fanout563 (.X(net563),
    .A(_06161_));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(_06155_));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(_06148_));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(_06142_));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(_06127_));
 sg13g2_buf_8 fanout568 (.A(_06126_),
    .X(net568));
 sg13g2_buf_8 fanout569 (.A(_06094_),
    .X(net569));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_06087_));
 sg13g2_buf_8 fanout571 (.A(_06081_),
    .X(net571));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(_06072_));
 sg13g2_buf_8 fanout573 (.A(_06071_),
    .X(net573));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(_06066_));
 sg13g2_buf_8 fanout575 (.A(_06065_),
    .X(net575));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(_06062_));
 sg13g2_buf_2 fanout577 (.A(_05990_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_05902_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_05453_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_05412_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_05373_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_05372_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_05371_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_05370_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_05369_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_05368_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_05367_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_05361_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_04402_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_04395_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_04303_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_04285_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_04225_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_04104_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_03603_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_03577_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_03563_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_01902_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_01793_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_01650_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_01641_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_01613_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_01609_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_05961_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_05951_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_05935_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_05910_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_05535_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_05479_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_05438_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_05427_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_05414_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_05338_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_05337_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_04325_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_04273_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_04105_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_04100_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_02277_),
    .X(net619));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(_02131_));
 sg13g2_buf_2 fanout621 (.A(_02114_),
    .X(net621));
 sg13g2_buf_4 fanout622 (.X(net622),
    .A(_02058_));
 sg13g2_buf_2 fanout623 (.A(_01819_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_01796_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_01702_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_01667_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_01654_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_01652_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_01645_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_01610_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_01601_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_01576_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_01561_),
    .X(net633));
 sg13g2_tiehi _16741__634 (.L_HI(net634));
 sg13g2_tiehi _16742__635 (.L_HI(net635));
 sg13g2_tiehi _16743__636 (.L_HI(net636));
 sg13g2_tiehi _16744__637 (.L_HI(net637));
 sg13g2_tiehi _16746__638 (.L_HI(net638));
 sg13g2_tiehi _16748__639 (.L_HI(net639));
 sg13g2_tiehi _16750__640 (.L_HI(net640));
 sg13g2_tiehi _16751__641 (.L_HI(net641));
 sg13g2_tiehi _16757__642 (.L_HI(net642));
 sg13g2_tiehi \soc_I.cycle_cnt[0]$_SDFF_PN0__643  (.L_HI(net643));
 sg13g2_tiehi \soc_I.cycle_cnt[10]$_SDFF_PN0__644  (.L_HI(net644));
 sg13g2_tiehi \soc_I.cycle_cnt[11]$_SDFF_PN0__645  (.L_HI(net645));
 sg13g2_tiehi \soc_I.cycle_cnt[12]$_SDFF_PN0__646  (.L_HI(net646));
 sg13g2_tiehi \soc_I.cycle_cnt[13]$_SDFF_PN0__647  (.L_HI(net647));
 sg13g2_tiehi \soc_I.cycle_cnt[14]$_SDFF_PN0__648  (.L_HI(net648));
 sg13g2_tiehi \soc_I.cycle_cnt[15]$_SDFF_PN0__649  (.L_HI(net649));
 sg13g2_tiehi \soc_I.cycle_cnt[16]$_SDFF_PN0__650  (.L_HI(net650));
 sg13g2_tiehi \soc_I.cycle_cnt[17]$_SDFF_PN0__651  (.L_HI(net651));
 sg13g2_tiehi \soc_I.cycle_cnt[18]$_SDFF_PN0__652  (.L_HI(net652));
 sg13g2_tiehi \soc_I.cycle_cnt[19]$_SDFF_PN0__653  (.L_HI(net653));
 sg13g2_tiehi \soc_I.cycle_cnt[1]$_SDFF_PN0__654  (.L_HI(net654));
 sg13g2_tiehi \soc_I.cycle_cnt[20]$_SDFF_PN0__655  (.L_HI(net655));
 sg13g2_tiehi \soc_I.cycle_cnt[21]$_SDFF_PN0__656  (.L_HI(net656));
 sg13g2_tiehi \soc_I.cycle_cnt[22]$_SDFF_PN0__657  (.L_HI(net657));
 sg13g2_tiehi \soc_I.cycle_cnt[23]$_SDFF_PN0__658  (.L_HI(net658));
 sg13g2_tiehi \soc_I.cycle_cnt[24]$_SDFF_PN0__659  (.L_HI(net659));
 sg13g2_tiehi \soc_I.cycle_cnt[25]$_SDFF_PN0__660  (.L_HI(net660));
 sg13g2_tiehi \soc_I.cycle_cnt[26]$_SDFF_PN0__661  (.L_HI(net661));
 sg13g2_tiehi \soc_I.cycle_cnt[27]$_SDFF_PN0__662  (.L_HI(net662));
 sg13g2_tiehi \soc_I.cycle_cnt[28]$_SDFF_PN0__663  (.L_HI(net663));
 sg13g2_tiehi \soc_I.cycle_cnt[29]$_SDFF_PN0__664  (.L_HI(net664));
 sg13g2_tiehi \soc_I.cycle_cnt[2]$_SDFF_PN0__665  (.L_HI(net665));
 sg13g2_tiehi \soc_I.cycle_cnt[30]$_SDFF_PN0__666  (.L_HI(net666));
 sg13g2_tiehi \soc_I.cycle_cnt[31]$_SDFF_PN0__667  (.L_HI(net667));
 sg13g2_tiehi \soc_I.cycle_cnt[3]$_SDFF_PN0__668  (.L_HI(net668));
 sg13g2_tiehi \soc_I.cycle_cnt[4]$_SDFF_PN0__669  (.L_HI(net669));
 sg13g2_tiehi \soc_I.cycle_cnt[5]$_SDFF_PN0__670  (.L_HI(net670));
 sg13g2_tiehi \soc_I.cycle_cnt[6]$_SDFF_PN0__671  (.L_HI(net671));
 sg13g2_tiehi \soc_I.cycle_cnt[7]$_SDFF_PN0__672  (.L_HI(net672));
 sg13g2_tiehi \soc_I.cycle_cnt[8]$_SDFF_PN0__673  (.L_HI(net673));
 sg13g2_tiehi \soc_I.cycle_cnt[9]$_SDFF_PN0__674  (.L_HI(net674));
 sg13g2_tiehi \soc_I.cycle_cnt_ready$_SDFF_PN0__675  (.L_HI(net675));
 sg13g2_tiehi \soc_I.div_ready$_SDFF_PN0__676  (.L_HI(net676));
 sg13g2_tiehi \soc_I.div_reg[0]$_SDFFE_PN0P__677  (.L_HI(net677));
 sg13g2_tiehi \soc_I.div_reg[10]$_SDFFE_PN0P__678  (.L_HI(net678));
 sg13g2_tiehi \soc_I.div_reg[11]$_SDFFE_PN0P__679  (.L_HI(net679));
 sg13g2_tiehi \soc_I.div_reg[12]$_SDFFE_PN0P__680  (.L_HI(net680));
 sg13g2_tiehi \soc_I.div_reg[13]$_SDFFE_PN0P__681  (.L_HI(net681));
 sg13g2_tiehi \soc_I.div_reg[14]$_SDFFE_PN0P__682  (.L_HI(net682));
 sg13g2_tiehi \soc_I.div_reg[15]$_SDFFE_PN0P__683  (.L_HI(net683));
 sg13g2_tiehi \soc_I.div_reg[16]$_SDFFE_PN0P__684  (.L_HI(net684));
 sg13g2_tiehi \soc_I.div_reg[17]$_SDFFE_PN0P__685  (.L_HI(net685));
 sg13g2_tiehi \soc_I.div_reg[18]$_SDFFE_PN0P__686  (.L_HI(net686));
 sg13g2_tiehi \soc_I.div_reg[19]$_SDFFE_PN0P__687  (.L_HI(net687));
 sg13g2_tiehi \soc_I.div_reg[1]$_SDFFE_PN0P__688  (.L_HI(net688));
 sg13g2_tiehi \soc_I.div_reg[20]$_SDFFE_PN0P__689  (.L_HI(net689));
 sg13g2_tiehi \soc_I.div_reg[21]$_SDFFE_PN0P__690  (.L_HI(net690));
 sg13g2_tiehi \soc_I.div_reg[22]$_SDFFE_PN0P__691  (.L_HI(net691));
 sg13g2_tiehi \soc_I.div_reg[23]$_SDFFE_PN0P__692  (.L_HI(net692));
 sg13g2_tiehi \soc_I.div_reg[24]$_SDFFE_PN0P__693  (.L_HI(net693));
 sg13g2_tiehi \soc_I.div_reg[25]$_SDFFE_PN0P__694  (.L_HI(net694));
 sg13g2_tiehi \soc_I.div_reg[26]$_SDFFE_PN0P__695  (.L_HI(net695));
 sg13g2_tiehi \soc_I.div_reg[27]$_SDFFE_PN0P__696  (.L_HI(net696));
 sg13g2_tiehi \soc_I.div_reg[28]$_SDFFE_PN0P__697  (.L_HI(net697));
 sg13g2_tiehi \soc_I.div_reg[29]$_SDFFE_PN0P__698  (.L_HI(net698));
 sg13g2_tiehi \soc_I.div_reg[2]$_SDFFE_PN0P__699  (.L_HI(net699));
 sg13g2_tiehi \soc_I.div_reg[30]$_SDFFE_PN0P__700  (.L_HI(net700));
 sg13g2_tiehi \soc_I.div_reg[31]$_SDFFE_PN0P__701  (.L_HI(net701));
 sg13g2_tiehi \soc_I.div_reg[3]$_SDFFE_PN0P__702  (.L_HI(net702));
 sg13g2_tiehi \soc_I.div_reg[4]$_SDFFE_PN0P__703  (.L_HI(net703));
 sg13g2_tiehi \soc_I.div_reg[5]$_SDFFE_PN0P__704  (.L_HI(net704));
 sg13g2_tiehi \soc_I.div_reg[6]$_SDFFE_PN0P__705  (.L_HI(net705));
 sg13g2_tiehi \soc_I.div_reg[7]$_SDFFE_PN0P__706  (.L_HI(net706));
 sg13g2_tiehi \soc_I.div_reg[8]$_SDFFE_PN0P__707  (.L_HI(net707));
 sg13g2_tiehi \soc_I.div_reg[9]$_SDFFE_PN0P__708  (.L_HI(net708));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[0]$_DFF_P__709  (.L_HI(net709));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[10]$_DFF_P__710  (.L_HI(net710));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[11]$_DFF_P__711  (.L_HI(net711));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[12]$_DFF_P__712  (.L_HI(net712));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[13]$_DFF_P__713  (.L_HI(net713));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[1]$_DFF_P__714  (.L_HI(net714));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[2]$_DFF_P__715  (.L_HI(net715));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[3]$_DFF_P__716  (.L_HI(net716));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[4]$_DFF_P__717  (.L_HI(net717));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[5]$_DFF_P__718  (.L_HI(net718));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[6]$_DFF_P__719  (.L_HI(net719));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[7]$_DFF_P__720  (.L_HI(net720));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[8]$_DFF_P__721  (.L_HI(net721));
 sg13g2_tiehi \soc_I.kianv_I.control_unit_I.main_fsm_I.state[9]$_DFF_P__722  (.L_HI(net722));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[0]$_SDFF_PN0__723  (.L_HI(net723));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[10]$_SDFF_PN0__724  (.L_HI(net724));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[11]$_SDFF_PN0__725  (.L_HI(net725));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[12]$_SDFF_PN0__726  (.L_HI(net726));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[13]$_SDFF_PN0__727  (.L_HI(net727));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[14]$_SDFF_PN0__728  (.L_HI(net728));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[15]$_SDFF_PN0__729  (.L_HI(net729));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[16]$_SDFF_PN0__730  (.L_HI(net730));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[17]$_SDFF_PN0__731  (.L_HI(net731));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[18]$_SDFF_PN0__732  (.L_HI(net732));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[19]$_SDFF_PN0__733  (.L_HI(net733));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[1]$_SDFF_PN0__734  (.L_HI(net734));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[20]$_SDFF_PN0__735  (.L_HI(net735));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[21]$_SDFF_PN0__736  (.L_HI(net736));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[22]$_SDFF_PN0__737  (.L_HI(net737));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[23]$_SDFF_PN0__738  (.L_HI(net738));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[24]$_SDFF_PN0__739  (.L_HI(net739));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[25]$_SDFF_PN0__740  (.L_HI(net740));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[26]$_SDFF_PN0__741  (.L_HI(net741));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[27]$_SDFF_PN0__742  (.L_HI(net742));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[28]$_SDFF_PN0__743  (.L_HI(net743));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[29]$_SDFF_PN0__744  (.L_HI(net744));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[2]$_SDFF_PN0__745  (.L_HI(net745));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[30]$_SDFF_PN0__746  (.L_HI(net746));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[31]$_SDFF_PN0__747  (.L_HI(net747));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[3]$_SDFF_PN0__748  (.L_HI(net748));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[4]$_SDFF_PN0__749  (.L_HI(net749));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[5]$_SDFF_PN0__750  (.L_HI(net750));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[6]$_SDFF_PN0__751  (.L_HI(net751));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[7]$_SDFF_PN0__752  (.L_HI(net752));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[8]$_SDFF_PN0__753  (.L_HI(net753));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A1_I.q[9]$_SDFF_PN0__754  (.L_HI(net754));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[0]$_SDFF_PN0__755  (.L_HI(net755));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[10]$_SDFF_PN0__756  (.L_HI(net756));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[11]$_SDFF_PN0__757  (.L_HI(net757));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[12]$_SDFF_PN0__758  (.L_HI(net758));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[13]$_SDFF_PN0__759  (.L_HI(net759));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[14]$_SDFF_PN0__760  (.L_HI(net760));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[15]$_SDFF_PN0__761  (.L_HI(net761));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[16]$_SDFF_PN0__762  (.L_HI(net762));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[17]$_SDFF_PN0__763  (.L_HI(net763));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[18]$_SDFF_PN0__764  (.L_HI(net764));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[19]$_SDFF_PN0__765  (.L_HI(net765));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[1]$_SDFF_PN0__766  (.L_HI(net766));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[20]$_SDFF_PN0__767  (.L_HI(net767));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[21]$_SDFF_PN0__768  (.L_HI(net768));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[22]$_SDFF_PN0__769  (.L_HI(net769));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[23]$_SDFF_PN0__770  (.L_HI(net770));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[24]$_SDFF_PN0__771  (.L_HI(net771));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[25]$_SDFF_PN0__772  (.L_HI(net772));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[26]$_SDFF_PN0__773  (.L_HI(net773));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[27]$_SDFF_PN0__774  (.L_HI(net774));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[28]$_SDFF_PN0__775  (.L_HI(net775));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[29]$_SDFF_PN0__776  (.L_HI(net776));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[2]$_SDFF_PN0__777  (.L_HI(net777));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[30]$_SDFF_PN0__778  (.L_HI(net778));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[31]$_SDFF_PN0__779  (.L_HI(net779));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[3]$_SDFF_PN0__780  (.L_HI(net780));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[4]$_SDFF_PN0__781  (.L_HI(net781));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[5]$_SDFF_PN0__782  (.L_HI(net782));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[6]$_SDFF_PN0__783  (.L_HI(net783));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[7]$_SDFF_PN0__784  (.L_HI(net784));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[8]$_SDFF_PN0__785  (.L_HI(net785));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.A2_I.q[9]$_SDFF_PN0__786  (.L_HI(net786));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0]$_DFF_P__787  (.L_HI(net787));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ADDR_I.q[1]$_DFF_P__788  (.L_HI(net788));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[0]$_SDFFE_PN0P__789  (.L_HI(net789));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[10]$_SDFFE_PN0P__790  (.L_HI(net790));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[11]$_SDFFE_PN0P__791  (.L_HI(net791));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[12]$_SDFFE_PN0P__792  (.L_HI(net792));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[13]$_SDFFE_PN0P__793  (.L_HI(net793));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[14]$_SDFFE_PN0P__794  (.L_HI(net794));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[15]$_SDFFE_PN0P__795  (.L_HI(net795));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[16]$_SDFFE_PN0P__796  (.L_HI(net796));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[17]$_SDFFE_PN0P__797  (.L_HI(net797));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[18]$_SDFFE_PN0P__798  (.L_HI(net798));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[19]$_SDFFE_PN0P__799  (.L_HI(net799));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[1]$_SDFFE_PN0P__800  (.L_HI(net800));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[20]$_SDFFE_PN0P__801  (.L_HI(net801));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[21]$_SDFFE_PN0P__802  (.L_HI(net802));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[22]$_SDFFE_PN0P__803  (.L_HI(net803));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[23]$_SDFFE_PN0P__804  (.L_HI(net804));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[24]$_SDFFE_PN0P__805  (.L_HI(net805));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[25]$_SDFFE_PN0P__806  (.L_HI(net806));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[26]$_SDFFE_PN0P__807  (.L_HI(net807));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[27]$_SDFFE_PN0P__808  (.L_HI(net808));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[28]$_SDFFE_PN0P__809  (.L_HI(net809));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[29]$_SDFFE_PN0P__810  (.L_HI(net810));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[2]$_SDFFE_PN0P__811  (.L_HI(net811));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[30]$_SDFFE_PN0P__812  (.L_HI(net812));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[31]$_SDFFE_PN0P__813  (.L_HI(net813));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[3]$_SDFFE_PN0P__814  (.L_HI(net814));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[4]$_SDFFE_PN0P__815  (.L_HI(net815));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[5]$_SDFFE_PN0P__816  (.L_HI(net816));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[6]$_SDFFE_PN0P__817  (.L_HI(net817));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[7]$_SDFFE_PN0P__818  (.L_HI(net818));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[8]$_SDFFE_PN0P__819  (.L_HI(net819));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.ALUOut_I.q[9]$_SDFFE_PN0P__820  (.L_HI(net820));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[0]$_DFF_P__821  (.L_HI(net821));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[10]$_DFF_P__822  (.L_HI(net822));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[11]$_DFF_P__823  (.L_HI(net823));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[12]$_DFF_P__824  (.L_HI(net824));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[13]$_DFF_P__825  (.L_HI(net825));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[14]$_DFF_P__826  (.L_HI(net826));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[15]$_DFF_P__827  (.L_HI(net827));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[16]$_DFF_P__828  (.L_HI(net828));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[17]$_DFF_P__829  (.L_HI(net829));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[18]$_DFF_P__830  (.L_HI(net830));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[19]$_DFF_P__831  (.L_HI(net831));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[1]$_DFF_P__832  (.L_HI(net832));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[20]$_DFF_P__833  (.L_HI(net833));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[21]$_DFF_P__834  (.L_HI(net834));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[22]$_DFF_P__835  (.L_HI(net835));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[23]$_DFF_P__836  (.L_HI(net836));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[24]$_DFF_P__837  (.L_HI(net837));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[25]$_DFF_P__838  (.L_HI(net838));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[26]$_DFF_P__839  (.L_HI(net839));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[27]$_DFF_P__840  (.L_HI(net840));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[28]$_DFF_P__841  (.L_HI(net841));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[29]$_DFF_P__842  (.L_HI(net842));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[2]$_DFF_P__843  (.L_HI(net843));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[30]$_DFF_P__844  (.L_HI(net844));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[31]$_DFF_P__845  (.L_HI(net845));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[3]$_DFF_P__846  (.L_HI(net846));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[4]$_DFF_P__847  (.L_HI(net847));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[5]$_DFF_P__848  (.L_HI(net848));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[6]$_DFF_P__849  (.L_HI(net849));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[7]$_DFF_P__850  (.L_HI(net850));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[8]$_DFF_P__851  (.L_HI(net851));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Data_I.q[9]$_DFF_P__852  (.L_HI(net852));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[0]$_SDFFE_PN0P__853  (.L_HI(net853));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[10]$_SDFFE_PN0P__854  (.L_HI(net854));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[11]$_SDFFE_PN0P__855  (.L_HI(net855));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[12]$_SDFFE_PN0P__856  (.L_HI(net856));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[13]$_SDFFE_PN0P__857  (.L_HI(net857));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[14]$_SDFFE_PN0P__858  (.L_HI(net858));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[15]$_SDFFE_PN0P__859  (.L_HI(net859));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[16]$_SDFFE_PN0P__860  (.L_HI(net860));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[17]$_SDFFE_PN0P__861  (.L_HI(net861));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[18]$_SDFFE_PN0P__862  (.L_HI(net862));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[19]$_SDFFE_PN0P__863  (.L_HI(net863));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[1]$_SDFFE_PN0P__864  (.L_HI(net864));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[20]$_SDFFE_PN0P__865  (.L_HI(net865));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[21]$_SDFFE_PN0P__866  (.L_HI(net866));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[22]$_SDFFE_PN0P__867  (.L_HI(net867));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[23]$_SDFFE_PN0P__868  (.L_HI(net868));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[24]$_SDFFE_PN0P__869  (.L_HI(net869));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[25]$_SDFFE_PN0P__870  (.L_HI(net870));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[26]$_SDFFE_PN0P__871  (.L_HI(net871));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[27]$_SDFFE_PN0P__872  (.L_HI(net872));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[28]$_SDFFE_PN0P__873  (.L_HI(net873));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[29]$_SDFFE_PN0P__874  (.L_HI(net874));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[2]$_SDFFE_PN0P__875  (.L_HI(net875));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[30]$_SDFFE_PN0P__876  (.L_HI(net876));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[31]$_SDFFE_PN0P__877  (.L_HI(net877));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[3]$_SDFFE_PN0P__878  (.L_HI(net878));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[4]$_SDFFE_PN0P__879  (.L_HI(net879));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[5]$_SDFFE_PN0P__880  (.L_HI(net880));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[6]$_SDFFE_PN0P__881  (.L_HI(net881));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[7]$_SDFFE_PN0P__882  (.L_HI(net882));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[8]$_SDFFE_PN0P__883  (.L_HI(net883));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.Instr_I.q[9]$_SDFFE_PN0P__884  (.L_HI(net884));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[0]$_SDFFE_PN0P__885  (.L_HI(net885));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[10]$_SDFFE_PN0P__886  (.L_HI(net886));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[11]$_SDFFE_PN0P__887  (.L_HI(net887));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[12]$_SDFFE_PN0P__888  (.L_HI(net888));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[13]$_SDFFE_PN0P__889  (.L_HI(net889));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[14]$_SDFFE_PN0P__890  (.L_HI(net890));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[15]$_SDFFE_PN0P__891  (.L_HI(net891));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[16]$_SDFFE_PN0P__892  (.L_HI(net892));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[17]$_SDFFE_PN0P__893  (.L_HI(net893));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[18]$_SDFFE_PN0P__894  (.L_HI(net894));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[19]$_SDFFE_PN0P__895  (.L_HI(net895));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[1]$_SDFFE_PN0P__896  (.L_HI(net896));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[20]$_SDFFE_PN0P__897  (.L_HI(net897));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[21]$_SDFFE_PN0P__898  (.L_HI(net898));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[22]$_SDFFE_PN0P__899  (.L_HI(net899));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[23]$_SDFFE_PN0P__900  (.L_HI(net900));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[24]$_SDFFE_PN0P__901  (.L_HI(net901));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[25]$_SDFFE_PN0P__902  (.L_HI(net902));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[26]$_SDFFE_PN0P__903  (.L_HI(net903));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[27]$_SDFFE_PN0P__904  (.L_HI(net904));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[28]$_SDFFE_PN0P__905  (.L_HI(net905));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[29]$_SDFFE_PN0P__906  (.L_HI(net906));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[2]$_SDFFE_PN0P__907  (.L_HI(net907));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[30]$_SDFFE_PN0P__908  (.L_HI(net908));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[31]$_SDFFE_PN0P__909  (.L_HI(net909));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[3]$_SDFFE_PN0P__910  (.L_HI(net910));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[4]$_SDFFE_PN0P__911  (.L_HI(net911));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[5]$_SDFFE_PN0P__912  (.L_HI(net912));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[6]$_SDFFE_PN0P__913  (.L_HI(net913));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[7]$_SDFFE_PN0P__914  (.L_HI(net914));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[8]$_SDFFE_PN0P__915  (.L_HI(net915));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.OldPC_I.q[9]$_SDFFE_PN0P__916  (.L_HI(net916));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[0]$_SDFFE_PN0P__917  (.L_HI(net917));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[10]$_SDFFE_PN0P__918  (.L_HI(net918));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[11]$_SDFFE_PN0P__919  (.L_HI(net919));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[12]$_SDFFE_PN0P__920  (.L_HI(net920));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[13]$_SDFFE_PN0P__921  (.L_HI(net921));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[14]$_SDFFE_PN0P__922  (.L_HI(net922));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[15]$_SDFFE_PN0P__923  (.L_HI(net923));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[16]$_SDFFE_PN0P__924  (.L_HI(net924));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[17]$_SDFFE_PN0P__925  (.L_HI(net925));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[18]$_SDFFE_PN0P__926  (.L_HI(net926));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[19]$_SDFFE_PN0P__927  (.L_HI(net927));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[1]$_SDFFE_PN0P__928  (.L_HI(net928));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[20]$_SDFFE_PN1P__929  (.L_HI(net929));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[21]$_SDFFE_PN0P__930  (.L_HI(net930));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[22]$_SDFFE_PN0P__931  (.L_HI(net931));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[23]$_SDFFE_PN0P__932  (.L_HI(net932));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[24]$_SDFFE_PN0P__933  (.L_HI(net933));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[25]$_SDFFE_PN0P__934  (.L_HI(net934));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[26]$_SDFFE_PN0P__935  (.L_HI(net935));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[27]$_SDFFE_PN0P__936  (.L_HI(net936));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[28]$_SDFFE_PN0P__937  (.L_HI(net937));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[29]$_SDFFE_PN1P__938  (.L_HI(net938));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[2]$_SDFFE_PN0P__939  (.L_HI(net939));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[30]$_SDFFE_PN0P__940  (.L_HI(net940));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[31]$_SDFFE_PN0P__941  (.L_HI(net941));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[3]$_SDFFE_PN0P__942  (.L_HI(net942));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[4]$_SDFFE_PN0P__943  (.L_HI(net943));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[5]$_SDFFE_PN0P__944  (.L_HI(net944));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[6]$_SDFFE_PN0P__945  (.L_HI(net945));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[7]$_SDFFE_PN0P__946  (.L_HI(net946));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[8]$_SDFFE_PN0P__947  (.L_HI(net947));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.PC_I.q[9]$_SDFFE_PN0P__948  (.L_HI(net948));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[0]$_SDFFE_PN0P__949  (.L_HI(net949));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[1]$_SDFFE_PN0P__950  (.L_HI(net950));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[2]$_SDFFE_PN0P__951  (.L_HI(net951));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[3]$_SDFFE_PN0P__952  (.L_HI(net952));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_cnt[4]$_SDFFE_PN0P__953  (.L_HI(net953));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_ready$_SDFFE_PN0P__954  (.L_HI(net954));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[0]$_DFFE_PP__955  (.L_HI(net955));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[10]$_DFFE_PP__956  (.L_HI(net956));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[11]$_DFFE_PP__957  (.L_HI(net957));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[12]$_DFFE_PP__958  (.L_HI(net958));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[13]$_DFFE_PP__959  (.L_HI(net959));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[14]$_DFFE_PP__960  (.L_HI(net960));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[15]$_DFFE_PP__961  (.L_HI(net961));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[16]$_DFFE_PP__962  (.L_HI(net962));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[17]$_DFFE_PP__963  (.L_HI(net963));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[18]$_DFFE_PP__964  (.L_HI(net964));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[19]$_DFFE_PP__965  (.L_HI(net965));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[1]$_DFFE_PP__966  (.L_HI(net966));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[20]$_DFFE_PP__967  (.L_HI(net967));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[21]$_DFFE_PP__968  (.L_HI(net968));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[22]$_DFFE_PP__969  (.L_HI(net969));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[23]$_DFFE_PP__970  (.L_HI(net970));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[24]$_DFFE_PP__971  (.L_HI(net971));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[25]$_DFFE_PP__972  (.L_HI(net972));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[26]$_DFFE_PP__973  (.L_HI(net973));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[27]$_DFFE_PP__974  (.L_HI(net974));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[28]$_DFFE_PP__975  (.L_HI(net975));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[29]$_DFFE_PP__976  (.L_HI(net976));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[2]$_DFFE_PP__977  (.L_HI(net977));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[30]$_DFFE_PP__978  (.L_HI(net978));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[31]$_DFFE_PP__979  (.L_HI(net979));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[3]$_DFFE_PP__980  (.L_HI(net980));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[4]$_DFFE_PP__981  (.L_HI(net981));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[5]$_DFFE_PP__982  (.L_HI(net982));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[6]$_DFFE_PP__983  (.L_HI(net983));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[7]$_DFFE_PP__984  (.L_HI(net984));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[8]$_DFFE_PP__985  (.L_HI(net985));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_result[9]$_DFFE_PP__986  (.L_HI(net986));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.alu_I.shift_state$_SDFF_PN0__987  (.L_HI(net987));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0]$_DFFE_PP__988  (.L_HI(net988));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10]$_DFFE_PP__989  (.L_HI(net989));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11]$_DFFE_PP__990  (.L_HI(net990));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12]$_DFFE_PP__991  (.L_HI(net991));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13]$_DFFE_PP__992  (.L_HI(net992));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14]$_DFFE_PP__993  (.L_HI(net993));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15]$_DFFE_PP__994  (.L_HI(net994));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16]$_DFFE_PP__995  (.L_HI(net995));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17]$_DFFE_PP__996  (.L_HI(net996));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18]$_DFFE_PP__997  (.L_HI(net997));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19]$_DFFE_PP__998  (.L_HI(net998));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1]$_DFFE_PP__999  (.L_HI(net999));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20]$_DFFE_PP__1000  (.L_HI(net1000));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21]$_DFFE_PP__1001  (.L_HI(net1001));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22]$_DFFE_PP__1002  (.L_HI(net1002));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23]$_DFFE_PP__1003  (.L_HI(net1003));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24]$_DFFE_PP__1004  (.L_HI(net1004));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25]$_DFFE_PP__1005  (.L_HI(net1005));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26]$_DFFE_PP__1006  (.L_HI(net1006));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27]$_DFFE_PP__1007  (.L_HI(net1007));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28]$_DFFE_PP__1008  (.L_HI(net1008));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29]$_DFFE_PP__1009  (.L_HI(net1009));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2]$_DFFE_PP__1010  (.L_HI(net1010));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30]$_DFFE_PP__1011  (.L_HI(net1011));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31]$_DFFE_PP__1012  (.L_HI(net1012));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3]$_DFFE_PP__1013  (.L_HI(net1013));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4]$_DFFE_PP__1014  (.L_HI(net1014));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5]$_DFFE_PP__1015  (.L_HI(net1015));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6]$_DFFE_PP__1016  (.L_HI(net1016));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7]$_DFFE_PP__1017  (.L_HI(net1017));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8]$_DFFE_PP__1018  (.L_HI(net1018));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9]$_DFFE_PP__1019  (.L_HI(net1019));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0]$_DFFE_PP__1020  (.L_HI(net1020));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10]$_DFFE_PP__1021  (.L_HI(net1021));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11]$_DFFE_PP__1022  (.L_HI(net1022));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12]$_DFFE_PP__1023  (.L_HI(net1023));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13]$_DFFE_PP__1024  (.L_HI(net1024));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14]$_DFFE_PP__1025  (.L_HI(net1025));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15]$_DFFE_PP__1026  (.L_HI(net1026));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16]$_DFFE_PP__1027  (.L_HI(net1027));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17]$_DFFE_PP__1028  (.L_HI(net1028));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18]$_DFFE_PP__1029  (.L_HI(net1029));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19]$_DFFE_PP__1030  (.L_HI(net1030));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1]$_DFFE_PP__1031  (.L_HI(net1031));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20]$_DFFE_PP__1032  (.L_HI(net1032));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21]$_DFFE_PP__1033  (.L_HI(net1033));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22]$_DFFE_PP__1034  (.L_HI(net1034));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23]$_DFFE_PP__1035  (.L_HI(net1035));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24]$_DFFE_PP__1036  (.L_HI(net1036));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25]$_DFFE_PP__1037  (.L_HI(net1037));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26]$_DFFE_PP__1038  (.L_HI(net1038));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27]$_DFFE_PP__1039  (.L_HI(net1039));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28]$_DFFE_PP__1040  (.L_HI(net1040));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29]$_DFFE_PP__1041  (.L_HI(net1041));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2]$_DFFE_PP__1042  (.L_HI(net1042));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30]$_DFFE_PP__1043  (.L_HI(net1043));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31]$_DFFE_PP__1044  (.L_HI(net1044));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3]$_DFFE_PP__1045  (.L_HI(net1045));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4]$_DFFE_PP__1046  (.L_HI(net1046));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5]$_DFFE_PP__1047  (.L_HI(net1047));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6]$_DFFE_PP__1048  (.L_HI(net1048));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7]$_DFFE_PP__1049  (.L_HI(net1049));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8]$_DFFE_PP__1050  (.L_HI(net1050));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9]$_DFFE_PP__1051  (.L_HI(net1051));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0]$_DFFE_PP__1052  (.L_HI(net1052));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10]$_DFFE_PP__1053  (.L_HI(net1053));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11]$_DFFE_PP__1054  (.L_HI(net1054));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12]$_DFFE_PP__1055  (.L_HI(net1055));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13]$_DFFE_PP__1056  (.L_HI(net1056));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14]$_DFFE_PP__1057  (.L_HI(net1057));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15]$_DFFE_PP__1058  (.L_HI(net1058));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16]$_DFFE_PP__1059  (.L_HI(net1059));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17]$_DFFE_PP__1060  (.L_HI(net1060));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18]$_DFFE_PP__1061  (.L_HI(net1061));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19]$_DFFE_PP__1062  (.L_HI(net1062));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1]$_DFFE_PP__1063  (.L_HI(net1063));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20]$_DFFE_PP__1064  (.L_HI(net1064));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21]$_DFFE_PP__1065  (.L_HI(net1065));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22]$_DFFE_PP__1066  (.L_HI(net1066));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23]$_DFFE_PP__1067  (.L_HI(net1067));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24]$_DFFE_PP__1068  (.L_HI(net1068));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25]$_DFFE_PP__1069  (.L_HI(net1069));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26]$_DFFE_PP__1070  (.L_HI(net1070));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27]$_DFFE_PP__1071  (.L_HI(net1071));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28]$_DFFE_PP__1072  (.L_HI(net1072));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29]$_DFFE_PP__1073  (.L_HI(net1073));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2]$_DFFE_PP__1074  (.L_HI(net1074));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30]$_DFFE_PP__1075  (.L_HI(net1075));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31]$_DFFE_PP__1076  (.L_HI(net1076));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3]$_DFFE_PP__1077  (.L_HI(net1077));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4]$_DFFE_PP__1078  (.L_HI(net1078));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5]$_DFFE_PP__1079  (.L_HI(net1079));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6]$_DFFE_PP__1080  (.L_HI(net1080));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7]$_DFFE_PP__1081  (.L_HI(net1081));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8]$_DFFE_PP__1082  (.L_HI(net1082));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9]$_DFFE_PP__1083  (.L_HI(net1083));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0]$_DFFE_PP__1084  (.L_HI(net1084));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10]$_DFFE_PP__1085  (.L_HI(net1085));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11]$_DFFE_PP__1086  (.L_HI(net1086));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12]$_DFFE_PP__1087  (.L_HI(net1087));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13]$_DFFE_PP__1088  (.L_HI(net1088));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14]$_DFFE_PP__1089  (.L_HI(net1089));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15]$_DFFE_PP__1090  (.L_HI(net1090));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16]$_DFFE_PP__1091  (.L_HI(net1091));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17]$_DFFE_PP__1092  (.L_HI(net1092));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18]$_DFFE_PP__1093  (.L_HI(net1093));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19]$_DFFE_PP__1094  (.L_HI(net1094));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1]$_DFFE_PP__1095  (.L_HI(net1095));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20]$_DFFE_PP__1096  (.L_HI(net1096));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21]$_DFFE_PP__1097  (.L_HI(net1097));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22]$_DFFE_PP__1098  (.L_HI(net1098));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23]$_DFFE_PP__1099  (.L_HI(net1099));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24]$_DFFE_PP__1100  (.L_HI(net1100));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25]$_DFFE_PP__1101  (.L_HI(net1101));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26]$_DFFE_PP__1102  (.L_HI(net1102));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27]$_DFFE_PP__1103  (.L_HI(net1103));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28]$_DFFE_PP__1104  (.L_HI(net1104));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29]$_DFFE_PP__1105  (.L_HI(net1105));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2]$_DFFE_PP__1106  (.L_HI(net1106));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30]$_DFFE_PP__1107  (.L_HI(net1107));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31]$_DFFE_PP__1108  (.L_HI(net1108));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3]$_DFFE_PP__1109  (.L_HI(net1109));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4]$_DFFE_PP__1110  (.L_HI(net1110));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5]$_DFFE_PP__1111  (.L_HI(net1111));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6]$_DFFE_PP__1112  (.L_HI(net1112));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7]$_DFFE_PP__1113  (.L_HI(net1113));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8]$_DFFE_PP__1114  (.L_HI(net1114));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9]$_DFFE_PP__1115  (.L_HI(net1115));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0]$_DFFE_PP__1116  (.L_HI(net1116));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10]$_DFFE_PP__1117  (.L_HI(net1117));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11]$_DFFE_PP__1118  (.L_HI(net1118));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12]$_DFFE_PP__1119  (.L_HI(net1119));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13]$_DFFE_PP__1120  (.L_HI(net1120));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14]$_DFFE_PP__1121  (.L_HI(net1121));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15]$_DFFE_PP__1122  (.L_HI(net1122));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \soc_I.pwm_I.pcm[0]$_SDFFE_PN0P__1500  (.L_HI(net1500));
 sg13g2_tiehi \soc_I.pwm_I.pcm[1]$_SDFFE_PN0P__1501  (.L_HI(net1501));
 sg13g2_tiehi \soc_I.pwm_I.pcm[2]$_SDFFE_PN0P__1502  (.L_HI(net1502));
 sg13g2_tiehi \soc_I.pwm_I.pcm[3]$_SDFFE_PN0P__1503  (.L_HI(net1503));
 sg13g2_tiehi \soc_I.pwm_I.pcm[4]$_SDFFE_PN0P__1504  (.L_HI(net1504));
 sg13g2_tiehi \soc_I.pwm_I.pcm[5]$_SDFFE_PN0P__1505  (.L_HI(net1505));
 sg13g2_tiehi \soc_I.pwm_I.pcm[6]$_SDFFE_PN0P__1506  (.L_HI(net1506));
 sg13g2_tiehi \soc_I.pwm_I.pcm[7]$_SDFFE_PN0P__1507  (.L_HI(net1507));
 sg13g2_tiehi \soc_I.pwm_I.pwm_accumulator[0]$_SDFF_PN0__1508  (.L_HI(net1508));
 sg13g2_tiehi \soc_I.pwm_I.pwm_accumulator[1]$_SDFF_PN0__1509  (.L_HI(net1509));
 sg13g2_tiehi \soc_I.pwm_I.pwm_accumulator[2]$_SDFF_PN0__1510  (.L_HI(net1510));
 sg13g2_tiehi \soc_I.pwm_I.pwm_accumulator[3]$_SDFF_PN0__1511  (.L_HI(net1511));
 sg13g2_tiehi \soc_I.pwm_I.pwm_accumulator[4]$_SDFF_PN0__1512  (.L_HI(net1512));
 sg13g2_tiehi \soc_I.pwm_I.pwm_accumulator[5]$_SDFF_PN0__1513  (.L_HI(net1513));
 sg13g2_tiehi \soc_I.pwm_I.pwm_accumulator[6]$_SDFF_PN0__1514  (.L_HI(net1514));
 sg13g2_tiehi \soc_I.pwm_I.pwm_accumulator[7]$_SDFF_PN0__1515  (.L_HI(net1515));
 sg13g2_tiehi \soc_I.pwm_I.pwm_accumulator[8]$_SDFF_PN0__1516  (.L_HI(net1516));
 sg13g2_tiehi \soc_I.pwm_ready$_SDFF_PN0__1517  (.L_HI(net1517));
 sg13g2_tiehi \soc_I.qqspi_I.ce[0]$_SDFFE_PN1P__1518  (.L_HI(net1518));
 sg13g2_tiehi \soc_I.qqspi_I.ce[1]$_SDFFE_PN1P__1519  (.L_HI(net1519));
 sg13g2_tiehi \soc_I.qqspi_I.is_quad$_SDFFE_PN0P__1520  (.L_HI(net1520));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[0]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[10]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[11]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[12]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[13]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[14]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[15]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[16]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[17]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[18]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[19]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[1]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[20]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[21]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[22]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[23]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[24]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[25]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[26]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[27]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[28]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[29]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[2]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[30]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[31]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[3]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[4]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[5]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[6]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[7]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[8]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \soc_I.qqspi_I.rdata[9]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \soc_I.qqspi_I.ready$_SDFFE_PN0P__1553  (.L_HI(net1553));
 sg13g2_tiehi \soc_I.qqspi_I.sclk$_SDFFE_PN1N__1554  (.L_HI(net1554));
 sg13g2_tiehi \soc_I.qqspi_I.sio_oe[0]$_SDFFE_PN0P__1555  (.L_HI(net1555));
 sg13g2_tiehi \soc_I.qqspi_I.sio_oe[2]$_SDFFE_PN0P__1556  (.L_HI(net1556));
 sg13g2_tiehi \soc_I.qqspi_I.sio_out[0]$_SDFFE_PN0N__1557  (.L_HI(net1557));
 sg13g2_tiehi \soc_I.qqspi_I.sio_out[1]$_SDFFE_PN0N__1558  (.L_HI(net1558));
 sg13g2_tiehi \soc_I.qqspi_I.sio_out[2]$_SDFFE_PN0N__1559  (.L_HI(net1559));
 sg13g2_tiehi \soc_I.qqspi_I.sio_out[3]$_SDFFE_PN0N__1560  (.L_HI(net1560));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[0]$_SDFFE_PN0P__1561  (.L_HI(net1561));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[10]$_SDFFE_PN0P__1562  (.L_HI(net1562));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[11]$_SDFFE_PN0P__1563  (.L_HI(net1563));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[12]$_SDFFE_PN0P__1564  (.L_HI(net1564));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[13]$_SDFFE_PN0P__1565  (.L_HI(net1565));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[14]$_SDFFE_PN0P__1566  (.L_HI(net1566));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[15]$_SDFFE_PN0P__1567  (.L_HI(net1567));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[16]$_SDFFE_PN0P__1568  (.L_HI(net1568));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[17]$_SDFFE_PN0P__1569  (.L_HI(net1569));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[18]$_SDFFE_PN0P__1570  (.L_HI(net1570));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[19]$_SDFFE_PN0P__1571  (.L_HI(net1571));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[1]$_SDFFE_PN0P__1572  (.L_HI(net1572));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[20]$_SDFFE_PN0P__1573  (.L_HI(net1573));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[21]$_SDFFE_PN0P__1574  (.L_HI(net1574));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[22]$_SDFFE_PN0P__1575  (.L_HI(net1575));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[23]$_SDFFE_PN0P__1576  (.L_HI(net1576));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[24]$_SDFFE_PN0P__1577  (.L_HI(net1577));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[25]$_SDFFE_PN0P__1578  (.L_HI(net1578));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[26]$_SDFFE_PN0P__1579  (.L_HI(net1579));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[27]$_SDFFE_PN0P__1580  (.L_HI(net1580));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[28]$_SDFFE_PN0P__1581  (.L_HI(net1581));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[29]$_SDFFE_PN0P__1582  (.L_HI(net1582));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[2]$_SDFFE_PN0P__1583  (.L_HI(net1583));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[30]$_SDFFE_PN0P__1584  (.L_HI(net1584));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[31]$_SDFFE_PN0P__1585  (.L_HI(net1585));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[3]$_SDFFE_PN0P__1586  (.L_HI(net1586));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[4]$_SDFFE_PN0P__1587  (.L_HI(net1587));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[5]$_SDFFE_PN0P__1588  (.L_HI(net1588));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[6]$_SDFFE_PN0P__1589  (.L_HI(net1589));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[7]$_SDFFE_PN0P__1590  (.L_HI(net1590));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[8]$_SDFFE_PN0P__1591  (.L_HI(net1591));
 sg13g2_tiehi \soc_I.qqspi_I.spi_buf[9]$_SDFFE_PN0P__1592  (.L_HI(net1592));
 sg13g2_tiehi \soc_I.qqspi_I.state[0]$_DFF_P__1593  (.L_HI(net1593));
 sg13g2_tiehi \soc_I.qqspi_I.state[1]$_DFF_P__1594  (.L_HI(net1594));
 sg13g2_tiehi \soc_I.qqspi_I.state[2]$_DFF_P__1595  (.L_HI(net1595));
 sg13g2_tiehi \soc_I.qqspi_I.state[3]$_DFF_P__1596  (.L_HI(net1596));
 sg13g2_tiehi \soc_I.qqspi_I.state[4]$_DFF_P__1597  (.L_HI(net1597));
 sg13g2_tiehi \soc_I.qqspi_I.state[5]$_DFF_P__1598  (.L_HI(net1598));
 sg13g2_tiehi \soc_I.qqspi_I.state[6]$_DFF_P__1599  (.L_HI(net1599));
 sg13g2_tiehi \soc_I.qqspi_I.xfer_cycles[0]$_SDFFE_PN0P__1600  (.L_HI(net1600));
 sg13g2_tiehi \soc_I.qqspi_I.xfer_cycles[1]$_SDFFE_PN0P__1601  (.L_HI(net1601));
 sg13g2_tiehi \soc_I.qqspi_I.xfer_cycles[2]$_SDFFE_PN0P__1602  (.L_HI(net1602));
 sg13g2_tiehi \soc_I.qqspi_I.xfer_cycles[3]$_SDFFE_PN0P__1603  (.L_HI(net1603));
 sg13g2_tiehi \soc_I.qqspi_I.xfer_cycles[4]$_SDFFE_PN0P__1604  (.L_HI(net1604));
 sg13g2_tiehi \soc_I.qqspi_I.xfer_cycles[5]$_SDFFE_PN0P__1605  (.L_HI(net1605));
 sg13g2_tiehi \soc_I.rst_cnt[0]$_SDFF_PN0__1606  (.L_HI(net1606));
 sg13g2_tiehi \soc_I.rst_cnt[1]$_SDFF_PN0__1607  (.L_HI(net1607));
 sg13g2_tiehi \soc_I.rst_cnt[2]$_SDFF_PN0__1608  (.L_HI(net1608));
 sg13g2_tiehi \soc_I.rst_cnt[3]$_SDFF_PN0__1609  (.L_HI(net1609));
 sg13g2_tiehi \soc_I.rx_uart_i.bit_idx[0]$_SDFFE_PN0P__1610  (.L_HI(net1610));
 sg13g2_tiehi \soc_I.rx_uart_i.bit_idx[1]$_SDFFE_PN0P__1611  (.L_HI(net1611));
 sg13g2_tiehi \soc_I.rx_uart_i.bit_idx[2]$_SDFFE_PN0P__1612  (.L_HI(net1612));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.cnt[0]$_SDFF_PN0__1613  (.L_HI(net1613));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.cnt[1]$_SDFF_PN0__1614  (.L_HI(net1614));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.cnt[2]$_SDFF_PN0__1615  (.L_HI(net1615));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.cnt[3]$_SDFF_PN0__1616  (.L_HI(net1616));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.cnt[4]$_SDFF_PN0__1617  (.L_HI(net1617));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[0][0]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[0][1]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[0][2]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[0][3]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[0][4]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[0][5]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[0][6]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[0][7]$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[10][0]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[10][1]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[10][2]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[10][3]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[10][4]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[10][5]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[10][6]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[10][7]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[11][0]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[11][1]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[11][2]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[11][3]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[11][4]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[11][5]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[11][6]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[11][7]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[12][0]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[12][1]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[12][2]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[12][3]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[12][4]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[12][5]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[12][6]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[12][7]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[13][0]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[13][1]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[13][2]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[13][3]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[13][4]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[13][5]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[13][6]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[13][7]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[14][0]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[14][1]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[14][2]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[14][3]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[14][4]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[14][5]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[14][6]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[14][7]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[15][0]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[15][1]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[15][2]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[15][3]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[15][4]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[15][5]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[15][6]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[15][7]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[1][0]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[1][1]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[1][2]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[1][3]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[1][4]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[1][5]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[1][6]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[1][7]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[2][0]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[2][1]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[2][2]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[2][3]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[2][4]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[2][5]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[2][6]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[2][7]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[3][0]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[3][1]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[3][2]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[3][3]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[3][4]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[3][5]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[3][6]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[3][7]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[4][0]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[4][1]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[4][2]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[4][3]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[4][4]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[4][5]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[4][6]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[4][7]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[5][0]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[5][1]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[5][2]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[5][3]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[5][4]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[5][5]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[5][6]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[5][7]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[6][0]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[6][1]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[6][2]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[6][3]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[6][4]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[6][5]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[6][6]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[6][7]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[7][0]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[7][1]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[7][2]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[7][3]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[7][4]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[7][5]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[7][6]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[7][7]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[8][0]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[8][1]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[8][2]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[8][3]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[8][4]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[8][5]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[8][6]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[8][7]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[9][0]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[9][1]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[9][2]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[9][3]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[9][4]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[9][5]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[9][6]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.ram[9][7]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.rd_ptr[0]$_SDFFE_PN0P__1746  (.L_HI(net1746));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.rd_ptr[1]$_SDFFE_PN0P__1747  (.L_HI(net1747));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.rd_ptr[2]$_SDFFE_PN0P__1748  (.L_HI(net1748));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.rd_ptr[3]$_SDFFE_PN0P__1749  (.L_HI(net1749));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.wr_ptr[0]$_SDFFE_PN0P__1750  (.L_HI(net1750));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.wr_ptr[1]$_SDFFE_PN0P__1751  (.L_HI(net1751));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.wr_ptr[2]$_SDFFE_PN0P__1752  (.L_HI(net1752));
 sg13g2_tiehi \soc_I.rx_uart_i.fifo_i.wr_ptr[3]$_SDFFE_PN0P__1753  (.L_HI(net1753));
 sg13g2_tiehi \soc_I.rx_uart_i.ready$_SDFFE_PN0P__1754  (.L_HI(net1754));
 sg13g2_tiehi \soc_I.rx_uart_i.return_state[0]$_SDFFCE_PP1P__1755  (.L_HI(net1755));
 sg13g2_tiehi \soc_I.rx_uart_i.return_state[1]$_SDFFCE_PP0P__1756  (.L_HI(net1756));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_data[0]$_SDFFE_PN0P__1757  (.L_HI(net1757));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_data[1]$_SDFFE_PN0P__1758  (.L_HI(net1758));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_data[2]$_SDFFE_PN0P__1759  (.L_HI(net1759));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_data[3]$_SDFFE_PN0P__1760  (.L_HI(net1760));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_data[4]$_SDFFE_PN0P__1761  (.L_HI(net1761));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_data[5]$_SDFFE_PN0P__1762  (.L_HI(net1762));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_data[6]$_SDFFE_PN0P__1763  (.L_HI(net1763));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_data[7]$_SDFFE_PN0P__1764  (.L_HI(net1764));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_in_sync[0]$_SDFF_PN0__1765  (.L_HI(net1765));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_in_sync[1]$_SDFF_PN0__1766  (.L_HI(net1766));
 sg13g2_tiehi \soc_I.rx_uart_i.rx_in_sync[2]$_SDFF_PN0__1767  (.L_HI(net1767));
 sg13g2_tiehi \soc_I.rx_uart_i.state[0]$_SDFFE_PN0P__1768  (.L_HI(net1768));
 sg13g2_tiehi \soc_I.rx_uart_i.state[1]$_SDFFE_PN0P__1769  (.L_HI(net1769));
 sg13g2_tiehi \soc_I.rx_uart_i.state[2]$_SDFFE_PN0P__1770  (.L_HI(net1770));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[0]$_SDFFE_PN1P__1771  (.L_HI(net1771));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[10]$_SDFFE_PN0P__1772  (.L_HI(net1772));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[11]$_SDFFE_PN0P__1773  (.L_HI(net1773));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[12]$_SDFFE_PN0P__1774  (.L_HI(net1774));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[13]$_SDFFE_PN0P__1775  (.L_HI(net1775));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[14]$_SDFFE_PN0P__1776  (.L_HI(net1776));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[15]$_SDFFE_PN0P__1777  (.L_HI(net1777));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[16]$_SDFFE_PN0P__1778  (.L_HI(net1778));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[1]$_SDFFE_PN0P__1779  (.L_HI(net1779));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[2]$_SDFFE_PN0P__1780  (.L_HI(net1780));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[3]$_SDFFE_PN0P__1781  (.L_HI(net1781));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[4]$_SDFFE_PN0P__1782  (.L_HI(net1782));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[5]$_SDFFE_PN0P__1783  (.L_HI(net1783));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[6]$_SDFFE_PN0P__1784  (.L_HI(net1784));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[7]$_SDFFE_PN0P__1785  (.L_HI(net1785));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[8]$_SDFFE_PN0P__1786  (.L_HI(net1786));
 sg13g2_tiehi \soc_I.rx_uart_i.wait_states[9]$_SDFFE_PN0P__1787  (.L_HI(net1787));
 sg13g2_tiehi \soc_I.spi0_I.ready_ctrl$_SDFF_PN0__1788  (.L_HI(net1788));
 sg13g2_tiehi \soc_I.spi0_I.ready_xfer$_SDFFE_PN0P__1789  (.L_HI(net1789));
 sg13g2_tiehi \soc_I.spi0_I.rx_data[0]$_SDFFE_PN0P__1790  (.L_HI(net1790));
 sg13g2_tiehi \soc_I.spi0_I.rx_data[1]$_SDFFE_PN0P__1791  (.L_HI(net1791));
 sg13g2_tiehi \soc_I.spi0_I.rx_data[2]$_SDFFE_PN0P__1792  (.L_HI(net1792));
 sg13g2_tiehi \soc_I.spi0_I.rx_data[3]$_SDFFE_PN0P__1793  (.L_HI(net1793));
 sg13g2_tiehi \soc_I.spi0_I.rx_data[4]$_SDFFE_PN0P__1794  (.L_HI(net1794));
 sg13g2_tiehi \soc_I.spi0_I.rx_data[5]$_SDFFE_PN0P__1795  (.L_HI(net1795));
 sg13g2_tiehi \soc_I.spi0_I.rx_data[6]$_SDFFE_PN0P__1796  (.L_HI(net1796));
 sg13g2_tiehi \soc_I.spi0_I.rx_data[7]$_SDFFE_PN0P__1797  (.L_HI(net1797));
 sg13g2_tiehi \soc_I.spi0_I.sclk$_SDFFE_PN1P__1798  (.L_HI(net1798));
 sg13g2_tiehi \soc_I.spi0_I.sio_out$_SDFFE_PN0P__1799  (.L_HI(net1799));
 sg13g2_tiehi \soc_I.spi0_I.spi_buf[0]$_SDFFE_PN0P__1800  (.L_HI(net1800));
 sg13g2_tiehi \soc_I.spi0_I.spi_buf[1]$_SDFFE_PN0P__1801  (.L_HI(net1801));
 sg13g2_tiehi \soc_I.spi0_I.spi_buf[2]$_SDFFE_PN0P__1802  (.L_HI(net1802));
 sg13g2_tiehi \soc_I.spi0_I.spi_buf[3]$_SDFFE_PN0P__1803  (.L_HI(net1803));
 sg13g2_tiehi \soc_I.spi0_I.spi_buf[4]$_SDFFE_PN0P__1804  (.L_HI(net1804));
 sg13g2_tiehi \soc_I.spi0_I.spi_buf[5]$_SDFFE_PN0P__1805  (.L_HI(net1805));
 sg13g2_tiehi \soc_I.spi0_I.spi_buf[6]$_SDFFE_PN0P__1806  (.L_HI(net1806));
 sg13g2_tiehi \soc_I.spi0_I.spi_buf[7]$_SDFFE_PN0P__1807  (.L_HI(net1807));
 sg13g2_tiehi \soc_I.spi0_I.spi_cen$_SDFFE_PN1P__1808  (.L_HI(net1808));
 sg13g2_tiehi \soc_I.spi0_I.state$_SDFFE_PN0P__1809  (.L_HI(net1809));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[0]$_SDFFE_PP0N__1810  (.L_HI(net1810));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[10]$_SDFFE_PP0N__1811  (.L_HI(net1811));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[11]$_SDFFE_PP0N__1812  (.L_HI(net1812));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[12]$_SDFFE_PP0N__1813  (.L_HI(net1813));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[13]$_SDFFE_PP0N__1814  (.L_HI(net1814));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[14]$_SDFFE_PP0N__1815  (.L_HI(net1815));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[15]$_SDFFE_PP0N__1816  (.L_HI(net1816));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[16]$_SDFFE_PP0N__1817  (.L_HI(net1817));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[17]$_SDFFE_PP0N__1818  (.L_HI(net1818));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[1]$_SDFFE_PP0N__1819  (.L_HI(net1819));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[2]$_SDFFE_PP0N__1820  (.L_HI(net1820));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[3]$_SDFFE_PP0N__1821  (.L_HI(net1821));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[4]$_SDFFE_PP0N__1822  (.L_HI(net1822));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[5]$_SDFFE_PP0N__1823  (.L_HI(net1823));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[6]$_SDFFE_PP0N__1824  (.L_HI(net1824));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[7]$_SDFFE_PP0N__1825  (.L_HI(net1825));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[8]$_SDFFE_PP0N__1826  (.L_HI(net1826));
 sg13g2_tiehi \soc_I.spi0_I.tick_cnt[9]$_SDFFE_PP0N__1827  (.L_HI(net1827));
 sg13g2_tiehi \soc_I.spi0_I.xfer_cycles[0]$_SDFFE_PN0P__1828  (.L_HI(net1828));
 sg13g2_tiehi \soc_I.spi0_I.xfer_cycles[1]$_SDFFE_PN0P__1829  (.L_HI(net1829));
 sg13g2_tiehi \soc_I.spi0_I.xfer_cycles[2]$_SDFFE_PN0P__1830  (.L_HI(net1830));
 sg13g2_tiehi \soc_I.spi0_I.xfer_cycles[3]$_SDFFE_PN0P__1831  (.L_HI(net1831));
 sg13g2_tiehi \soc_I.spi0_I.xfer_cycles[4]$_SDFFE_PN0P__1832  (.L_HI(net1832));
 sg13g2_tiehi \soc_I.spi0_I.xfer_cycles[5]$_SDFFE_PN0P__1833  (.L_HI(net1833));
 sg13g2_tiehi \soc_I.spi_div_ready$_SDFF_PN0__1834  (.L_HI(net1834));
 sg13g2_tiehi \soc_I.spi_div_reg[0]$_SDFFE_PN0P__1835  (.L_HI(net1835));
 sg13g2_tiehi \soc_I.spi_div_reg[10]$_SDFFE_PN0P__1836  (.L_HI(net1836));
 sg13g2_tiehi \soc_I.spi_div_reg[11]$_SDFFE_PN0P__1837  (.L_HI(net1837));
 sg13g2_tiehi \soc_I.spi_div_reg[12]$_SDFFE_PN0P__1838  (.L_HI(net1838));
 sg13g2_tiehi \soc_I.spi_div_reg[13]$_SDFFE_PN0P__1839  (.L_HI(net1839));
 sg13g2_tiehi \soc_I.spi_div_reg[14]$_SDFFE_PN0P__1840  (.L_HI(net1840));
 sg13g2_tiehi \soc_I.spi_div_reg[15]$_SDFFE_PN0P__1841  (.L_HI(net1841));
 sg13g2_tiehi \soc_I.spi_div_reg[16]$_SDFFE_PN0P__1842  (.L_HI(net1842));
 sg13g2_tiehi \soc_I.spi_div_reg[17]$_SDFFE_PN0P__1843  (.L_HI(net1843));
 sg13g2_tiehi \soc_I.spi_div_reg[18]$_SDFFE_PN0P__1844  (.L_HI(net1844));
 sg13g2_tiehi \soc_I.spi_div_reg[19]$_SDFFE_PN0P__1845  (.L_HI(net1845));
 sg13g2_tiehi \soc_I.spi_div_reg[1]$_SDFFE_PN0P__1846  (.L_HI(net1846));
 sg13g2_tiehi \soc_I.spi_div_reg[20]$_SDFFE_PN0P__1847  (.L_HI(net1847));
 sg13g2_tiehi \soc_I.spi_div_reg[21]$_SDFFE_PN0P__1848  (.L_HI(net1848));
 sg13g2_tiehi \soc_I.spi_div_reg[22]$_SDFFE_PN0P__1849  (.L_HI(net1849));
 sg13g2_tiehi \soc_I.spi_div_reg[23]$_SDFFE_PN0P__1850  (.L_HI(net1850));
 sg13g2_tiehi \soc_I.spi_div_reg[24]$_SDFFE_PN0P__1851  (.L_HI(net1851));
 sg13g2_tiehi \soc_I.spi_div_reg[25]$_SDFFE_PN0P__1852  (.L_HI(net1852));
 sg13g2_tiehi \soc_I.spi_div_reg[26]$_SDFFE_PN0P__1853  (.L_HI(net1853));
 sg13g2_tiehi \soc_I.spi_div_reg[27]$_SDFFE_PN0P__1854  (.L_HI(net1854));
 sg13g2_tiehi \soc_I.spi_div_reg[28]$_SDFFE_PN0P__1855  (.L_HI(net1855));
 sg13g2_tiehi \soc_I.spi_div_reg[29]$_SDFFE_PN0P__1856  (.L_HI(net1856));
 sg13g2_tiehi \soc_I.spi_div_reg[2]$_SDFFE_PN0P__1857  (.L_HI(net1857));
 sg13g2_tiehi \soc_I.spi_div_reg[30]$_SDFFE_PN0P__1858  (.L_HI(net1858));
 sg13g2_tiehi \soc_I.spi_div_reg[31]$_SDFFE_PN0P__1859  (.L_HI(net1859));
 sg13g2_tiehi \soc_I.spi_div_reg[3]$_SDFFE_PN0P__1860  (.L_HI(net1860));
 sg13g2_tiehi \soc_I.spi_div_reg[4]$_SDFFE_PN0P__1861  (.L_HI(net1861));
 sg13g2_tiehi \soc_I.spi_div_reg[5]$_SDFFE_PN0P__1862  (.L_HI(net1862));
 sg13g2_tiehi \soc_I.spi_div_reg[6]$_SDFFE_PN0P__1863  (.L_HI(net1863));
 sg13g2_tiehi \soc_I.spi_div_reg[7]$_SDFFE_PN0P__1864  (.L_HI(net1864));
 sg13g2_tiehi \soc_I.spi_div_reg[8]$_SDFFE_PN0P__1865  (.L_HI(net1865));
 sg13g2_tiehi \soc_I.spi_div_reg[9]$_SDFFE_PN0P__1866  (.L_HI(net1866));
 sg13g2_tiehi \soc_I.tx_uart_i.bit_idx[0]$_SDFFE_PN0P__1867  (.L_HI(net1867));
 sg13g2_tiehi \soc_I.tx_uart_i.bit_idx[1]$_SDFFE_PN0P__1868  (.L_HI(net1868));
 sg13g2_tiehi \soc_I.tx_uart_i.bit_idx[2]$_SDFFE_PN0P__1869  (.L_HI(net1869));
 sg13g2_tiehi \soc_I.tx_uart_i.return_state[0]$_SDFFCE_PN1P__1870  (.L_HI(net1870));
 sg13g2_tiehi \soc_I.tx_uart_i.return_state[1]$_SDFFCE_PN0P__1871  (.L_HI(net1871));
 sg13g2_tiehi \soc_I.tx_uart_i.state[0]$_SDFFE_PN0P__1872  (.L_HI(net1872));
 sg13g2_tiehi \soc_I.tx_uart_i.state[1]$_SDFFE_PN0P__1873  (.L_HI(net1873));
 sg13g2_tiehi \soc_I.tx_uart_i.tx_data_reg[0]$_SDFFE_PN0P__1874  (.L_HI(net1874));
 sg13g2_tiehi \soc_I.tx_uart_i.tx_data_reg[1]$_SDFFE_PN0P__1875  (.L_HI(net1875));
 sg13g2_tiehi \soc_I.tx_uart_i.tx_data_reg[2]$_SDFFE_PN0P__1876  (.L_HI(net1876));
 sg13g2_tiehi \soc_I.tx_uart_i.tx_data_reg[3]$_SDFFE_PN0P__1877  (.L_HI(net1877));
 sg13g2_tiehi \soc_I.tx_uart_i.tx_data_reg[4]$_SDFFE_PN0P__1878  (.L_HI(net1878));
 sg13g2_tiehi \soc_I.tx_uart_i.tx_data_reg[5]$_SDFFE_PN0P__1879  (.L_HI(net1879));
 sg13g2_tiehi \soc_I.tx_uart_i.tx_data_reg[6]$_SDFFE_PN0P__1880  (.L_HI(net1880));
 sg13g2_tiehi \soc_I.tx_uart_i.tx_data_reg[7]$_SDFFE_PN0P__1881  (.L_HI(net1881));
 sg13g2_tiehi \soc_I.tx_uart_i.tx_out$_SDFFE_PN1N__1882  (.L_HI(net1882));
 sg13g2_tiehi \soc_I.tx_uart_i.txfer_done$_SDFFE_PN0P__1883  (.L_HI(net1883));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[0]$_SDFFCE_PP1P__1884  (.L_HI(net1884));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[10]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[11]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[12]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[13]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[14]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[15]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[1]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[2]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[3]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[4]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[5]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[6]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[7]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[8]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \soc_I.tx_uart_i.wait_states[9]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \soc_I.uart_lsr_rdy$_SDFF_PN0__1900  (.L_HI(net1900));
 sg13g2_tiehi \soc_I.uart_rx_ready$_SDFF_PN0__1901  (.L_HI(net1901));
 sg13g2_tiehi \soc_I.uart_tx_ready$_SDFF_PN0__1902  (.L_HI(net1902));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_5_0__f_clk (.X(clknet_5_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_5_1__f_clk (.X(clknet_5_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_5_2__f_clk (.X(clknet_5_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_5_3__f_clk (.X(clknet_5_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_5_4__f_clk (.X(clknet_5_4__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_5_5__f_clk (.X(clknet_5_5__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_5_6__f_clk (.X(clknet_5_6__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_5_7__f_clk (.X(clknet_5_7__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_5_8__f_clk (.X(clknet_5_8__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_5_9__f_clk (.X(clknet_5_9__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_5_10__f_clk (.X(clknet_5_10__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_5_11__f_clk (.X(clknet_5_11__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_5_12__f_clk (.X(clknet_5_12__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_5_13__f_clk (.X(clknet_5_13__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_5_14__f_clk (.X(clknet_5_14__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_5_15__f_clk (.X(clknet_5_15__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_5_16__f_clk (.X(clknet_5_16__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_5_17__f_clk (.X(clknet_5_17__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_5_18__f_clk (.X(clknet_5_18__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_5_19__f_clk (.X(clknet_5_19__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_5_20__f_clk (.X(clknet_5_20__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_5_21__f_clk (.X(clknet_5_21__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_5_22__f_clk (.X(clknet_5_22__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_5_23__f_clk (.X(clknet_5_23__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_5_24__f_clk (.X(clknet_5_24__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_5_25__f_clk (.X(clknet_5_25__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_5_26__f_clk (.X(clknet_5_26__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_5_27__f_clk (.X(clknet_5_27__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_5_28__f_clk (.X(clknet_5_28__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_5_29__f_clk (.X(clknet_5_29__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_5_30__f_clk (.X(clknet_5_30__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_5_31__f_clk (.X(clknet_5_31__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_buf_16 clkload1 (.A(clknet_5_2__leaf_clk));
 sg13g2_buf_16 clkload2 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_162_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_30_clk));
 sg13g2_buf_16 clkload12 (.A(clknet_leaf_31_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_45_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_139_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_140_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_leaf_119_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_82_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_76_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_68_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00220_));
 sg13g2_antennanp ANTENNA_2 (.A(_00220_));
 sg13g2_antennanp ANTENNA_3 (.A(_00222_));
 sg13g2_antennanp ANTENNA_4 (.A(_00224_));
 sg13g2_antennanp ANTENNA_5 (.A(_00262_));
 sg13g2_antennanp ANTENNA_6 (.A(_00263_));
 sg13g2_antennanp ANTENNA_7 (.A(_00264_));
 sg13g2_antennanp ANTENNA_8 (.A(_00922_));
 sg13g2_antennanp ANTENNA_9 (.A(_00922_));
 sg13g2_antennanp ANTENNA_10 (.A(_01573_));
 sg13g2_antennanp ANTENNA_11 (.A(_01573_));
 sg13g2_antennanp ANTENNA_12 (.A(_01573_));
 sg13g2_antennanp ANTENNA_13 (.A(_01573_));
 sg13g2_antennanp ANTENNA_14 (.A(_01573_));
 sg13g2_antennanp ANTENNA_15 (.A(_01573_));
 sg13g2_antennanp ANTENNA_16 (.A(_01903_));
 sg13g2_antennanp ANTENNA_17 (.A(_01903_));
 sg13g2_antennanp ANTENNA_18 (.A(_01903_));
 sg13g2_antennanp ANTENNA_19 (.A(_01903_));
 sg13g2_antennanp ANTENNA_20 (.A(_01903_));
 sg13g2_antennanp ANTENNA_21 (.A(_01903_));
 sg13g2_antennanp ANTENNA_22 (.A(_02081_));
 sg13g2_antennanp ANTENNA_23 (.A(_02081_));
 sg13g2_antennanp ANTENNA_24 (.A(_02081_));
 sg13g2_antennanp ANTENNA_25 (.A(_02081_));
 sg13g2_antennanp ANTENNA_26 (.A(_02081_));
 sg13g2_antennanp ANTENNA_27 (.A(_02081_));
 sg13g2_antennanp ANTENNA_28 (.A(_02081_));
 sg13g2_antennanp ANTENNA_29 (.A(_02081_));
 sg13g2_antennanp ANTENNA_30 (.A(_02081_));
 sg13g2_antennanp ANTENNA_31 (.A(_02081_));
 sg13g2_antennanp ANTENNA_32 (.A(_02081_));
 sg13g2_antennanp ANTENNA_33 (.A(_02081_));
 sg13g2_antennanp ANTENNA_34 (.A(_02081_));
 sg13g2_antennanp ANTENNA_35 (.A(_02081_));
 sg13g2_antennanp ANTENNA_36 (.A(_02277_));
 sg13g2_antennanp ANTENNA_37 (.A(_02277_));
 sg13g2_antennanp ANTENNA_38 (.A(_02277_));
 sg13g2_antennanp ANTENNA_39 (.A(_02277_));
 sg13g2_antennanp ANTENNA_40 (.A(_02277_));
 sg13g2_antennanp ANTENNA_41 (.A(_02537_));
 sg13g2_antennanp ANTENNA_42 (.A(_02558_));
 sg13g2_antennanp ANTENNA_43 (.A(_03712_));
 sg13g2_antennanp ANTENNA_44 (.A(_03714_));
 sg13g2_antennanp ANTENNA_45 (.A(_03714_));
 sg13g2_antennanp ANTENNA_46 (.A(_03714_));
 sg13g2_antennanp ANTENNA_47 (.A(_03714_));
 sg13g2_antennanp ANTENNA_48 (.A(_03720_));
 sg13g2_antennanp ANTENNA_49 (.A(_03760_));
 sg13g2_antennanp ANTENNA_50 (.A(_03975_));
 sg13g2_antennanp ANTENNA_51 (.A(_04266_));
 sg13g2_antennanp ANTENNA_52 (.A(_04266_));
 sg13g2_antennanp ANTENNA_53 (.A(_04266_));
 sg13g2_antennanp ANTENNA_54 (.A(_04693_));
 sg13g2_antennanp ANTENNA_55 (.A(_04693_));
 sg13g2_antennanp ANTENNA_56 (.A(_04693_));
 sg13g2_antennanp ANTENNA_57 (.A(_04693_));
 sg13g2_antennanp ANTENNA_58 (.A(_04727_));
 sg13g2_antennanp ANTENNA_59 (.A(_04727_));
 sg13g2_antennanp ANTENNA_60 (.A(_04727_));
 sg13g2_antennanp ANTENNA_61 (.A(_04727_));
 sg13g2_antennanp ANTENNA_62 (.A(_04763_));
 sg13g2_antennanp ANTENNA_63 (.A(_04763_));
 sg13g2_antennanp ANTENNA_64 (.A(_04763_));
 sg13g2_antennanp ANTENNA_65 (.A(_04763_));
 sg13g2_antennanp ANTENNA_66 (.A(_04798_));
 sg13g2_antennanp ANTENNA_67 (.A(_04798_));
 sg13g2_antennanp ANTENNA_68 (.A(_04798_));
 sg13g2_antennanp ANTENNA_69 (.A(_04798_));
 sg13g2_antennanp ANTENNA_70 (.A(_04832_));
 sg13g2_antennanp ANTENNA_71 (.A(_04832_));
 sg13g2_antennanp ANTENNA_72 (.A(_04832_));
 sg13g2_antennanp ANTENNA_73 (.A(_04832_));
 sg13g2_antennanp ANTENNA_74 (.A(_04866_));
 sg13g2_antennanp ANTENNA_75 (.A(_04866_));
 sg13g2_antennanp ANTENNA_76 (.A(_04866_));
 sg13g2_antennanp ANTENNA_77 (.A(_04866_));
 sg13g2_antennanp ANTENNA_78 (.A(_04900_));
 sg13g2_antennanp ANTENNA_79 (.A(_04900_));
 sg13g2_antennanp ANTENNA_80 (.A(_04900_));
 sg13g2_antennanp ANTENNA_81 (.A(_04900_));
 sg13g2_antennanp ANTENNA_82 (.A(_05003_));
 sg13g2_antennanp ANTENNA_83 (.A(_05003_));
 sg13g2_antennanp ANTENNA_84 (.A(_05003_));
 sg13g2_antennanp ANTENNA_85 (.A(_05037_));
 sg13g2_antennanp ANTENNA_86 (.A(_05037_));
 sg13g2_antennanp ANTENNA_87 (.A(_05037_));
 sg13g2_antennanp ANTENNA_88 (.A(_05037_));
 sg13g2_antennanp ANTENNA_89 (.A(_05139_));
 sg13g2_antennanp ANTENNA_90 (.A(_05139_));
 sg13g2_antennanp ANTENNA_91 (.A(_05139_));
 sg13g2_antennanp ANTENNA_92 (.A(_05139_));
 sg13g2_antennanp ANTENNA_93 (.A(_05173_));
 sg13g2_antennanp ANTENNA_94 (.A(_05173_));
 sg13g2_antennanp ANTENNA_95 (.A(_05173_));
 sg13g2_antennanp ANTENNA_96 (.A(_06134_));
 sg13g2_antennanp ANTENNA_97 (.A(_06145_));
 sg13g2_antennanp ANTENNA_98 (.A(_06246_));
 sg13g2_antennanp ANTENNA_99 (.A(_06251_));
 sg13g2_antennanp ANTENNA_100 (.A(_07613_));
 sg13g2_antennanp ANTENNA_101 (.A(_07613_));
 sg13g2_antennanp ANTENNA_102 (.A(_07613_));
 sg13g2_antennanp ANTENNA_103 (.A(_07613_));
 sg13g2_antennanp ANTENNA_104 (.A(clk));
 sg13g2_antennanp ANTENNA_105 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_106 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_107 (.A(sclk));
 sg13g2_antennanp ANTENNA_108 (.A(sclk));
 sg13g2_antennanp ANTENNA_109 (.A(sclk));
 sg13g2_antennanp ANTENNA_110 (.A(sclk));
 sg13g2_antennanp ANTENNA_111 (.A(sclk));
 sg13g2_antennanp ANTENNA_112 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_113 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_114 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_115 (.A(\soc_I.kianv_I.datapath_unit_I.A1[0] ));
 sg13g2_antennanp ANTENNA_116 (.A(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_antennanp ANTENNA_117 (.A(\soc_I.kianv_I.datapath_unit_I.A1[14] ));
 sg13g2_antennanp ANTENNA_118 (.A(\soc_I.kianv_I.datapath_unit_I.A1[15] ));
 sg13g2_antennanp ANTENNA_119 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_120 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_121 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_122 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_123 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_124 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_125 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_126 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_127 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_128 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_129 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_130 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_131 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_132 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_133 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_134 (.A(net2));
 sg13g2_antennanp ANTENNA_135 (.A(net3));
 sg13g2_antennanp ANTENNA_136 (.A(net4));
 sg13g2_antennanp ANTENNA_137 (.A(net4));
 sg13g2_antennanp ANTENNA_138 (.A(net6));
 sg13g2_antennanp ANTENNA_139 (.A(net7));
 sg13g2_antennanp ANTENNA_140 (.A(net398));
 sg13g2_antennanp ANTENNA_141 (.A(net398));
 sg13g2_antennanp ANTENNA_142 (.A(net398));
 sg13g2_antennanp ANTENNA_143 (.A(net398));
 sg13g2_antennanp ANTENNA_144 (.A(net398));
 sg13g2_antennanp ANTENNA_145 (.A(net398));
 sg13g2_antennanp ANTENNA_146 (.A(net398));
 sg13g2_antennanp ANTENNA_147 (.A(net398));
 sg13g2_antennanp ANTENNA_148 (.A(net398));
 sg13g2_antennanp ANTENNA_149 (.A(net438));
 sg13g2_antennanp ANTENNA_150 (.A(net438));
 sg13g2_antennanp ANTENNA_151 (.A(net438));
 sg13g2_antennanp ANTENNA_152 (.A(net438));
 sg13g2_antennanp ANTENNA_153 (.A(net438));
 sg13g2_antennanp ANTENNA_154 (.A(net438));
 sg13g2_antennanp ANTENNA_155 (.A(net438));
 sg13g2_antennanp ANTENNA_156 (.A(net438));
 sg13g2_antennanp ANTENNA_157 (.A(net438));
 sg13g2_antennanp ANTENNA_158 (.A(net619));
 sg13g2_antennanp ANTENNA_159 (.A(net619));
 sg13g2_antennanp ANTENNA_160 (.A(net619));
 sg13g2_antennanp ANTENNA_161 (.A(net619));
 sg13g2_antennanp ANTENNA_162 (.A(net619));
 sg13g2_antennanp ANTENNA_163 (.A(net619));
 sg13g2_antennanp ANTENNA_164 (.A(net619));
 sg13g2_antennanp ANTENNA_165 (.A(net619));
 sg13g2_antennanp ANTENNA_166 (.A(net619));
 sg13g2_antennanp ANTENNA_167 (.A(net619));
 sg13g2_antennanp ANTENNA_168 (.A(net619));
 sg13g2_antennanp ANTENNA_169 (.A(net619));
 sg13g2_antennanp ANTENNA_170 (.A(net619));
 sg13g2_antennanp ANTENNA_171 (.A(net619));
 sg13g2_antennanp ANTENNA_172 (.A(net619));
 sg13g2_antennanp ANTENNA_173 (.A(net619));
 sg13g2_antennanp ANTENNA_174 (.A(net620));
 sg13g2_antennanp ANTENNA_175 (.A(net620));
 sg13g2_antennanp ANTENNA_176 (.A(net620));
 sg13g2_antennanp ANTENNA_177 (.A(net620));
 sg13g2_antennanp ANTENNA_178 (.A(net620));
 sg13g2_antennanp ANTENNA_179 (.A(net620));
 sg13g2_antennanp ANTENNA_180 (.A(net620));
 sg13g2_antennanp ANTENNA_181 (.A(net620));
 sg13g2_antennanp ANTENNA_182 (.A(net620));
 sg13g2_antennanp ANTENNA_183 (.A(net620));
 sg13g2_antennanp ANTENNA_184 (.A(net620));
 sg13g2_antennanp ANTENNA_185 (.A(net620));
 sg13g2_antennanp ANTENNA_186 (.A(net620));
 sg13g2_antennanp ANTENNA_187 (.A(net620));
 sg13g2_antennanp ANTENNA_188 (.A(net620));
 sg13g2_antennanp ANTENNA_189 (.A(net620));
 sg13g2_antennanp ANTENNA_190 (.A(net621));
 sg13g2_antennanp ANTENNA_191 (.A(net621));
 sg13g2_antennanp ANTENNA_192 (.A(net621));
 sg13g2_antennanp ANTENNA_193 (.A(net621));
 sg13g2_antennanp ANTENNA_194 (.A(net621));
 sg13g2_antennanp ANTENNA_195 (.A(net621));
 sg13g2_antennanp ANTENNA_196 (.A(net621));
 sg13g2_antennanp ANTENNA_197 (.A(net621));
 sg13g2_antennanp ANTENNA_198 (.A(net621));
 sg13g2_antennanp ANTENNA_199 (.A(net621));
 sg13g2_antennanp ANTENNA_200 (.A(net621));
 sg13g2_antennanp ANTENNA_201 (.A(net621));
 sg13g2_antennanp ANTENNA_202 (.A(_00220_));
 sg13g2_antennanp ANTENNA_203 (.A(_00220_));
 sg13g2_antennanp ANTENNA_204 (.A(_00222_));
 sg13g2_antennanp ANTENNA_205 (.A(_00224_));
 sg13g2_antennanp ANTENNA_206 (.A(_00262_));
 sg13g2_antennanp ANTENNA_207 (.A(_00263_));
 sg13g2_antennanp ANTENNA_208 (.A(_00263_));
 sg13g2_antennanp ANTENNA_209 (.A(_00264_));
 sg13g2_antennanp ANTENNA_210 (.A(_00264_));
 sg13g2_antennanp ANTENNA_211 (.A(_00922_));
 sg13g2_antennanp ANTENNA_212 (.A(_00922_));
 sg13g2_antennanp ANTENNA_213 (.A(_01573_));
 sg13g2_antennanp ANTENNA_214 (.A(_01573_));
 sg13g2_antennanp ANTENNA_215 (.A(_01573_));
 sg13g2_antennanp ANTENNA_216 (.A(_01573_));
 sg13g2_antennanp ANTENNA_217 (.A(_01573_));
 sg13g2_antennanp ANTENNA_218 (.A(_01573_));
 sg13g2_antennanp ANTENNA_219 (.A(_01840_));
 sg13g2_antennanp ANTENNA_220 (.A(_01840_));
 sg13g2_antennanp ANTENNA_221 (.A(_01840_));
 sg13g2_antennanp ANTENNA_222 (.A(_01840_));
 sg13g2_antennanp ANTENNA_223 (.A(_01840_));
 sg13g2_antennanp ANTENNA_224 (.A(_01840_));
 sg13g2_antennanp ANTENNA_225 (.A(_01903_));
 sg13g2_antennanp ANTENNA_226 (.A(_01903_));
 sg13g2_antennanp ANTENNA_227 (.A(_01903_));
 sg13g2_antennanp ANTENNA_228 (.A(_01903_));
 sg13g2_antennanp ANTENNA_229 (.A(_01903_));
 sg13g2_antennanp ANTENNA_230 (.A(_01903_));
 sg13g2_antennanp ANTENNA_231 (.A(_02081_));
 sg13g2_antennanp ANTENNA_232 (.A(_02081_));
 sg13g2_antennanp ANTENNA_233 (.A(_02081_));
 sg13g2_antennanp ANTENNA_234 (.A(_02081_));
 sg13g2_antennanp ANTENNA_235 (.A(_02081_));
 sg13g2_antennanp ANTENNA_236 (.A(_02081_));
 sg13g2_antennanp ANTENNA_237 (.A(_02081_));
 sg13g2_antennanp ANTENNA_238 (.A(_02081_));
 sg13g2_antennanp ANTENNA_239 (.A(_02081_));
 sg13g2_antennanp ANTENNA_240 (.A(_02081_));
 sg13g2_antennanp ANTENNA_241 (.A(_02081_));
 sg13g2_antennanp ANTENNA_242 (.A(_02081_));
 sg13g2_antennanp ANTENNA_243 (.A(_02081_));
 sg13g2_antennanp ANTENNA_244 (.A(_02537_));
 sg13g2_antennanp ANTENNA_245 (.A(_02558_));
 sg13g2_antennanp ANTENNA_246 (.A(_03712_));
 sg13g2_antennanp ANTENNA_247 (.A(_03714_));
 sg13g2_antennanp ANTENNA_248 (.A(_03714_));
 sg13g2_antennanp ANTENNA_249 (.A(_03714_));
 sg13g2_antennanp ANTENNA_250 (.A(_03714_));
 sg13g2_antennanp ANTENNA_251 (.A(_03720_));
 sg13g2_antennanp ANTENNA_252 (.A(_03760_));
 sg13g2_antennanp ANTENNA_253 (.A(_03975_));
 sg13g2_antennanp ANTENNA_254 (.A(_04266_));
 sg13g2_antennanp ANTENNA_255 (.A(_04266_));
 sg13g2_antennanp ANTENNA_256 (.A(_04266_));
 sg13g2_antennanp ANTENNA_257 (.A(_04693_));
 sg13g2_antennanp ANTENNA_258 (.A(_04693_));
 sg13g2_antennanp ANTENNA_259 (.A(_04693_));
 sg13g2_antennanp ANTENNA_260 (.A(_04693_));
 sg13g2_antennanp ANTENNA_261 (.A(_04727_));
 sg13g2_antennanp ANTENNA_262 (.A(_04727_));
 sg13g2_antennanp ANTENNA_263 (.A(_04727_));
 sg13g2_antennanp ANTENNA_264 (.A(_04727_));
 sg13g2_antennanp ANTENNA_265 (.A(_04763_));
 sg13g2_antennanp ANTENNA_266 (.A(_04763_));
 sg13g2_antennanp ANTENNA_267 (.A(_04763_));
 sg13g2_antennanp ANTENNA_268 (.A(_04763_));
 sg13g2_antennanp ANTENNA_269 (.A(_04798_));
 sg13g2_antennanp ANTENNA_270 (.A(_04798_));
 sg13g2_antennanp ANTENNA_271 (.A(_04798_));
 sg13g2_antennanp ANTENNA_272 (.A(_04798_));
 sg13g2_antennanp ANTENNA_273 (.A(_04832_));
 sg13g2_antennanp ANTENNA_274 (.A(_04832_));
 sg13g2_antennanp ANTENNA_275 (.A(_04832_));
 sg13g2_antennanp ANTENNA_276 (.A(_04832_));
 sg13g2_antennanp ANTENNA_277 (.A(_04900_));
 sg13g2_antennanp ANTENNA_278 (.A(_04900_));
 sg13g2_antennanp ANTENNA_279 (.A(_04900_));
 sg13g2_antennanp ANTENNA_280 (.A(_04900_));
 sg13g2_antennanp ANTENNA_281 (.A(_05910_));
 sg13g2_antennanp ANTENNA_282 (.A(_05910_));
 sg13g2_antennanp ANTENNA_283 (.A(_06134_));
 sg13g2_antennanp ANTENNA_284 (.A(_06246_));
 sg13g2_antennanp ANTENNA_285 (.A(_06251_));
 sg13g2_antennanp ANTENNA_286 (.A(_06253_));
 sg13g2_antennanp ANTENNA_287 (.A(_06253_));
 sg13g2_antennanp ANTENNA_288 (.A(_06253_));
 sg13g2_antennanp ANTENNA_289 (.A(_06253_));
 sg13g2_antennanp ANTENNA_290 (.A(_07613_));
 sg13g2_antennanp ANTENNA_291 (.A(_07613_));
 sg13g2_antennanp ANTENNA_292 (.A(_07613_));
 sg13g2_antennanp ANTENNA_293 (.A(_07613_));
 sg13g2_antennanp ANTENNA_294 (.A(clk));
 sg13g2_antennanp ANTENNA_295 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_296 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_297 (.A(sclk));
 sg13g2_antennanp ANTENNA_298 (.A(sclk));
 sg13g2_antennanp ANTENNA_299 (.A(sclk));
 sg13g2_antennanp ANTENNA_300 (.A(sclk));
 sg13g2_antennanp ANTENNA_301 (.A(sclk));
 sg13g2_antennanp ANTENNA_302 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_303 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_304 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_305 (.A(\soc_I.kianv_I.datapath_unit_I.A1[0] ));
 sg13g2_antennanp ANTENNA_306 (.A(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_antennanp ANTENNA_307 (.A(\soc_I.kianv_I.datapath_unit_I.A1[12] ));
 sg13g2_antennanp ANTENNA_308 (.A(\soc_I.kianv_I.datapath_unit_I.A1[15] ));
 sg13g2_antennanp ANTENNA_309 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_310 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_311 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_312 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_313 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_314 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_315 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_316 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_317 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_318 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_319 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_320 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_321 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_322 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_323 (.A(net2));
 sg13g2_antennanp ANTENNA_324 (.A(net4));
 sg13g2_antennanp ANTENNA_325 (.A(net6));
 sg13g2_antennanp ANTENNA_326 (.A(net6));
 sg13g2_antennanp ANTENNA_327 (.A(net398));
 sg13g2_antennanp ANTENNA_328 (.A(net398));
 sg13g2_antennanp ANTENNA_329 (.A(net398));
 sg13g2_antennanp ANTENNA_330 (.A(net398));
 sg13g2_antennanp ANTENNA_331 (.A(net398));
 sg13g2_antennanp ANTENNA_332 (.A(net398));
 sg13g2_antennanp ANTENNA_333 (.A(net398));
 sg13g2_antennanp ANTENNA_334 (.A(net398));
 sg13g2_antennanp ANTENNA_335 (.A(net398));
 sg13g2_antennanp ANTENNA_336 (.A(net438));
 sg13g2_antennanp ANTENNA_337 (.A(net438));
 sg13g2_antennanp ANTENNA_338 (.A(net438));
 sg13g2_antennanp ANTENNA_339 (.A(net438));
 sg13g2_antennanp ANTENNA_340 (.A(net438));
 sg13g2_antennanp ANTENNA_341 (.A(net438));
 sg13g2_antennanp ANTENNA_342 (.A(net438));
 sg13g2_antennanp ANTENNA_343 (.A(net438));
 sg13g2_antennanp ANTENNA_344 (.A(net438));
 sg13g2_antennanp ANTENNA_345 (.A(net619));
 sg13g2_antennanp ANTENNA_346 (.A(net619));
 sg13g2_antennanp ANTENNA_347 (.A(net619));
 sg13g2_antennanp ANTENNA_348 (.A(net619));
 sg13g2_antennanp ANTENNA_349 (.A(net619));
 sg13g2_antennanp ANTENNA_350 (.A(net619));
 sg13g2_antennanp ANTENNA_351 (.A(net619));
 sg13g2_antennanp ANTENNA_352 (.A(net619));
 sg13g2_antennanp ANTENNA_353 (.A(net619));
 sg13g2_antennanp ANTENNA_354 (.A(net619));
 sg13g2_antennanp ANTENNA_355 (.A(net619));
 sg13g2_antennanp ANTENNA_356 (.A(net619));
 sg13g2_antennanp ANTENNA_357 (.A(net619));
 sg13g2_antennanp ANTENNA_358 (.A(net619));
 sg13g2_antennanp ANTENNA_359 (.A(net620));
 sg13g2_antennanp ANTENNA_360 (.A(net620));
 sg13g2_antennanp ANTENNA_361 (.A(net620));
 sg13g2_antennanp ANTENNA_362 (.A(net620));
 sg13g2_antennanp ANTENNA_363 (.A(net620));
 sg13g2_antennanp ANTENNA_364 (.A(net620));
 sg13g2_antennanp ANTENNA_365 (.A(net620));
 sg13g2_antennanp ANTENNA_366 (.A(net620));
 sg13g2_antennanp ANTENNA_367 (.A(net620));
 sg13g2_antennanp ANTENNA_368 (.A(net621));
 sg13g2_antennanp ANTENNA_369 (.A(net621));
 sg13g2_antennanp ANTENNA_370 (.A(net621));
 sg13g2_antennanp ANTENNA_371 (.A(net621));
 sg13g2_antennanp ANTENNA_372 (.A(net621));
 sg13g2_antennanp ANTENNA_373 (.A(net621));
 sg13g2_antennanp ANTENNA_374 (.A(net621));
 sg13g2_antennanp ANTENNA_375 (.A(net621));
 sg13g2_antennanp ANTENNA_376 (.A(net621));
 sg13g2_antennanp ANTENNA_377 (.A(net621));
 sg13g2_antennanp ANTENNA_378 (.A(net621));
 sg13g2_antennanp ANTENNA_379 (.A(net621));
 sg13g2_antennanp ANTENNA_380 (.A(net621));
 sg13g2_antennanp ANTENNA_381 (.A(_00220_));
 sg13g2_antennanp ANTENNA_382 (.A(_00220_));
 sg13g2_antennanp ANTENNA_383 (.A(_00222_));
 sg13g2_antennanp ANTENNA_384 (.A(_00224_));
 sg13g2_antennanp ANTENNA_385 (.A(_00262_));
 sg13g2_antennanp ANTENNA_386 (.A(_00263_));
 sg13g2_antennanp ANTENNA_387 (.A(_00263_));
 sg13g2_antennanp ANTENNA_388 (.A(_00922_));
 sg13g2_antennanp ANTENNA_389 (.A(_00922_));
 sg13g2_antennanp ANTENNA_390 (.A(_01573_));
 sg13g2_antennanp ANTENNA_391 (.A(_01573_));
 sg13g2_antennanp ANTENNA_392 (.A(_01573_));
 sg13g2_antennanp ANTENNA_393 (.A(_01573_));
 sg13g2_antennanp ANTENNA_394 (.A(_01573_));
 sg13g2_antennanp ANTENNA_395 (.A(_01573_));
 sg13g2_antennanp ANTENNA_396 (.A(_01840_));
 sg13g2_antennanp ANTENNA_397 (.A(_01840_));
 sg13g2_antennanp ANTENNA_398 (.A(_01840_));
 sg13g2_antennanp ANTENNA_399 (.A(_01840_));
 sg13g2_antennanp ANTENNA_400 (.A(_01840_));
 sg13g2_antennanp ANTENNA_401 (.A(_01903_));
 sg13g2_antennanp ANTENNA_402 (.A(_01903_));
 sg13g2_antennanp ANTENNA_403 (.A(_01903_));
 sg13g2_antennanp ANTENNA_404 (.A(_01903_));
 sg13g2_antennanp ANTENNA_405 (.A(_01903_));
 sg13g2_antennanp ANTENNA_406 (.A(_01903_));
 sg13g2_antennanp ANTENNA_407 (.A(_02081_));
 sg13g2_antennanp ANTENNA_408 (.A(_02081_));
 sg13g2_antennanp ANTENNA_409 (.A(_02081_));
 sg13g2_antennanp ANTENNA_410 (.A(_02081_));
 sg13g2_antennanp ANTENNA_411 (.A(_02081_));
 sg13g2_antennanp ANTENNA_412 (.A(_02081_));
 sg13g2_antennanp ANTENNA_413 (.A(_02081_));
 sg13g2_antennanp ANTENNA_414 (.A(_02081_));
 sg13g2_antennanp ANTENNA_415 (.A(_02081_));
 sg13g2_antennanp ANTENNA_416 (.A(_02081_));
 sg13g2_antennanp ANTENNA_417 (.A(_02081_));
 sg13g2_antennanp ANTENNA_418 (.A(_02081_));
 sg13g2_antennanp ANTENNA_419 (.A(_02081_));
 sg13g2_antennanp ANTENNA_420 (.A(_02537_));
 sg13g2_antennanp ANTENNA_421 (.A(_02558_));
 sg13g2_antennanp ANTENNA_422 (.A(_03712_));
 sg13g2_antennanp ANTENNA_423 (.A(_03714_));
 sg13g2_antennanp ANTENNA_424 (.A(_03714_));
 sg13g2_antennanp ANTENNA_425 (.A(_03714_));
 sg13g2_antennanp ANTENNA_426 (.A(_03714_));
 sg13g2_antennanp ANTENNA_427 (.A(_03720_));
 sg13g2_antennanp ANTENNA_428 (.A(_03760_));
 sg13g2_antennanp ANTENNA_429 (.A(_03975_));
 sg13g2_antennanp ANTENNA_430 (.A(_04273_));
 sg13g2_antennanp ANTENNA_431 (.A(_04273_));
 sg13g2_antennanp ANTENNA_432 (.A(_04273_));
 sg13g2_antennanp ANTENNA_433 (.A(_04273_));
 sg13g2_antennanp ANTENNA_434 (.A(_04693_));
 sg13g2_antennanp ANTENNA_435 (.A(_04693_));
 sg13g2_antennanp ANTENNA_436 (.A(_04693_));
 sg13g2_antennanp ANTENNA_437 (.A(_04693_));
 sg13g2_antennanp ANTENNA_438 (.A(_04727_));
 sg13g2_antennanp ANTENNA_439 (.A(_04727_));
 sg13g2_antennanp ANTENNA_440 (.A(_04727_));
 sg13g2_antennanp ANTENNA_441 (.A(_04727_));
 sg13g2_antennanp ANTENNA_442 (.A(_04763_));
 sg13g2_antennanp ANTENNA_443 (.A(_04763_));
 sg13g2_antennanp ANTENNA_444 (.A(_04763_));
 sg13g2_antennanp ANTENNA_445 (.A(_04763_));
 sg13g2_antennanp ANTENNA_446 (.A(_04798_));
 sg13g2_antennanp ANTENNA_447 (.A(_04798_));
 sg13g2_antennanp ANTENNA_448 (.A(_04798_));
 sg13g2_antennanp ANTENNA_449 (.A(_04798_));
 sg13g2_antennanp ANTENNA_450 (.A(_04832_));
 sg13g2_antennanp ANTENNA_451 (.A(_04832_));
 sg13g2_antennanp ANTENNA_452 (.A(_04832_));
 sg13g2_antennanp ANTENNA_453 (.A(_04832_));
 sg13g2_antennanp ANTENNA_454 (.A(_04900_));
 sg13g2_antennanp ANTENNA_455 (.A(_04900_));
 sg13g2_antennanp ANTENNA_456 (.A(_04900_));
 sg13g2_antennanp ANTENNA_457 (.A(_04900_));
 sg13g2_antennanp ANTENNA_458 (.A(_05910_));
 sg13g2_antennanp ANTENNA_459 (.A(_05910_));
 sg13g2_antennanp ANTENNA_460 (.A(_06251_));
 sg13g2_antennanp ANTENNA_461 (.A(_07613_));
 sg13g2_antennanp ANTENNA_462 (.A(_07613_));
 sg13g2_antennanp ANTENNA_463 (.A(_07613_));
 sg13g2_antennanp ANTENNA_464 (.A(_07613_));
 sg13g2_antennanp ANTENNA_465 (.A(clk));
 sg13g2_antennanp ANTENNA_466 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_467 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_468 (.A(sclk));
 sg13g2_antennanp ANTENNA_469 (.A(sclk));
 sg13g2_antennanp ANTENNA_470 (.A(sclk));
 sg13g2_antennanp ANTENNA_471 (.A(sclk));
 sg13g2_antennanp ANTENNA_472 (.A(sclk));
 sg13g2_antennanp ANTENNA_473 (.A(sclk));
 sg13g2_antennanp ANTENNA_474 (.A(sclk));
 sg13g2_antennanp ANTENNA_475 (.A(sclk));
 sg13g2_antennanp ANTENNA_476 (.A(sclk));
 sg13g2_antennanp ANTENNA_477 (.A(sclk));
 sg13g2_antennanp ANTENNA_478 (.A(sclk));
 sg13g2_antennanp ANTENNA_479 (.A(sclk));
 sg13g2_antennanp ANTENNA_480 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_481 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_482 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_483 (.A(\soc_I.kianv_I.datapath_unit_I.A1[0] ));
 sg13g2_antennanp ANTENNA_484 (.A(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_antennanp ANTENNA_485 (.A(\soc_I.kianv_I.datapath_unit_I.A1[12] ));
 sg13g2_antennanp ANTENNA_486 (.A(\soc_I.kianv_I.datapath_unit_I.A1[15] ));
 sg13g2_antennanp ANTENNA_487 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_488 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_489 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_490 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_491 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_492 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_493 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_494 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_495 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_496 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_497 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_498 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_499 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_500 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_501 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_502 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_503 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_504 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_505 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_506 (.A(net398));
 sg13g2_antennanp ANTENNA_507 (.A(net398));
 sg13g2_antennanp ANTENNA_508 (.A(net398));
 sg13g2_antennanp ANTENNA_509 (.A(net398));
 sg13g2_antennanp ANTENNA_510 (.A(net398));
 sg13g2_antennanp ANTENNA_511 (.A(net398));
 sg13g2_antennanp ANTENNA_512 (.A(net398));
 sg13g2_antennanp ANTENNA_513 (.A(net398));
 sg13g2_antennanp ANTENNA_514 (.A(net398));
 sg13g2_antennanp ANTENNA_515 (.A(net438));
 sg13g2_antennanp ANTENNA_516 (.A(net438));
 sg13g2_antennanp ANTENNA_517 (.A(net438));
 sg13g2_antennanp ANTENNA_518 (.A(net438));
 sg13g2_antennanp ANTENNA_519 (.A(net438));
 sg13g2_antennanp ANTENNA_520 (.A(net438));
 sg13g2_antennanp ANTENNA_521 (.A(net438));
 sg13g2_antennanp ANTENNA_522 (.A(net438));
 sg13g2_antennanp ANTENNA_523 (.A(net438));
 sg13g2_antennanp ANTENNA_524 (.A(net619));
 sg13g2_antennanp ANTENNA_525 (.A(net619));
 sg13g2_antennanp ANTENNA_526 (.A(net619));
 sg13g2_antennanp ANTENNA_527 (.A(net619));
 sg13g2_antennanp ANTENNA_528 (.A(net619));
 sg13g2_antennanp ANTENNA_529 (.A(net619));
 sg13g2_antennanp ANTENNA_530 (.A(net619));
 sg13g2_antennanp ANTENNA_531 (.A(net619));
 sg13g2_antennanp ANTENNA_532 (.A(net619));
 sg13g2_antennanp ANTENNA_533 (.A(net619));
 sg13g2_antennanp ANTENNA_534 (.A(net619));
 sg13g2_antennanp ANTENNA_535 (.A(net619));
 sg13g2_antennanp ANTENNA_536 (.A(net619));
 sg13g2_antennanp ANTENNA_537 (.A(net619));
 sg13g2_antennanp ANTENNA_538 (.A(net619));
 sg13g2_antennanp ANTENNA_539 (.A(net619));
 sg13g2_antennanp ANTENNA_540 (.A(net620));
 sg13g2_antennanp ANTENNA_541 (.A(net620));
 sg13g2_antennanp ANTENNA_542 (.A(net620));
 sg13g2_antennanp ANTENNA_543 (.A(net620));
 sg13g2_antennanp ANTENNA_544 (.A(net620));
 sg13g2_antennanp ANTENNA_545 (.A(net620));
 sg13g2_antennanp ANTENNA_546 (.A(net620));
 sg13g2_antennanp ANTENNA_547 (.A(net620));
 sg13g2_antennanp ANTENNA_548 (.A(net620));
 sg13g2_antennanp ANTENNA_549 (.A(_00220_));
 sg13g2_antennanp ANTENNA_550 (.A(_00222_));
 sg13g2_antennanp ANTENNA_551 (.A(_00224_));
 sg13g2_antennanp ANTENNA_552 (.A(_00262_));
 sg13g2_antennanp ANTENNA_553 (.A(_00263_));
 sg13g2_antennanp ANTENNA_554 (.A(_00263_));
 sg13g2_antennanp ANTENNA_555 (.A(_00922_));
 sg13g2_antennanp ANTENNA_556 (.A(_00922_));
 sg13g2_antennanp ANTENNA_557 (.A(_01573_));
 sg13g2_antennanp ANTENNA_558 (.A(_01573_));
 sg13g2_antennanp ANTENNA_559 (.A(_01573_));
 sg13g2_antennanp ANTENNA_560 (.A(_01573_));
 sg13g2_antennanp ANTENNA_561 (.A(_01573_));
 sg13g2_antennanp ANTENNA_562 (.A(_01573_));
 sg13g2_antennanp ANTENNA_563 (.A(_01840_));
 sg13g2_antennanp ANTENNA_564 (.A(_01840_));
 sg13g2_antennanp ANTENNA_565 (.A(_01840_));
 sg13g2_antennanp ANTENNA_566 (.A(_01840_));
 sg13g2_antennanp ANTENNA_567 (.A(_01840_));
 sg13g2_antennanp ANTENNA_568 (.A(_01840_));
 sg13g2_antennanp ANTENNA_569 (.A(_01840_));
 sg13g2_antennanp ANTENNA_570 (.A(_01840_));
 sg13g2_antennanp ANTENNA_571 (.A(_01840_));
 sg13g2_antennanp ANTENNA_572 (.A(_01840_));
 sg13g2_antennanp ANTENNA_573 (.A(_01903_));
 sg13g2_antennanp ANTENNA_574 (.A(_01903_));
 sg13g2_antennanp ANTENNA_575 (.A(_01903_));
 sg13g2_antennanp ANTENNA_576 (.A(_01903_));
 sg13g2_antennanp ANTENNA_577 (.A(_01903_));
 sg13g2_antennanp ANTENNA_578 (.A(_01903_));
 sg13g2_antennanp ANTENNA_579 (.A(_02081_));
 sg13g2_antennanp ANTENNA_580 (.A(_02081_));
 sg13g2_antennanp ANTENNA_581 (.A(_02081_));
 sg13g2_antennanp ANTENNA_582 (.A(_02081_));
 sg13g2_antennanp ANTENNA_583 (.A(_02081_));
 sg13g2_antennanp ANTENNA_584 (.A(_02081_));
 sg13g2_antennanp ANTENNA_585 (.A(_02081_));
 sg13g2_antennanp ANTENNA_586 (.A(_02081_));
 sg13g2_antennanp ANTENNA_587 (.A(_02081_));
 sg13g2_antennanp ANTENNA_588 (.A(_02081_));
 sg13g2_antennanp ANTENNA_589 (.A(_02081_));
 sg13g2_antennanp ANTENNA_590 (.A(_02081_));
 sg13g2_antennanp ANTENNA_591 (.A(_02081_));
 sg13g2_antennanp ANTENNA_592 (.A(_02081_));
 sg13g2_antennanp ANTENNA_593 (.A(_02081_));
 sg13g2_antennanp ANTENNA_594 (.A(_02081_));
 sg13g2_antennanp ANTENNA_595 (.A(_02537_));
 sg13g2_antennanp ANTENNA_596 (.A(_02558_));
 sg13g2_antennanp ANTENNA_597 (.A(_03712_));
 sg13g2_antennanp ANTENNA_598 (.A(_03714_));
 sg13g2_antennanp ANTENNA_599 (.A(_03714_));
 sg13g2_antennanp ANTENNA_600 (.A(_03714_));
 sg13g2_antennanp ANTENNA_601 (.A(_03714_));
 sg13g2_antennanp ANTENNA_602 (.A(_03720_));
 sg13g2_antennanp ANTENNA_603 (.A(_03760_));
 sg13g2_antennanp ANTENNA_604 (.A(_03975_));
 sg13g2_antennanp ANTENNA_605 (.A(_04273_));
 sg13g2_antennanp ANTENNA_606 (.A(_04273_));
 sg13g2_antennanp ANTENNA_607 (.A(_04273_));
 sg13g2_antennanp ANTENNA_608 (.A(_04273_));
 sg13g2_antennanp ANTENNA_609 (.A(_04273_));
 sg13g2_antennanp ANTENNA_610 (.A(_04273_));
 sg13g2_antennanp ANTENNA_611 (.A(_04693_));
 sg13g2_antennanp ANTENNA_612 (.A(_04693_));
 sg13g2_antennanp ANTENNA_613 (.A(_04693_));
 sg13g2_antennanp ANTENNA_614 (.A(_04693_));
 sg13g2_antennanp ANTENNA_615 (.A(_04727_));
 sg13g2_antennanp ANTENNA_616 (.A(_04727_));
 sg13g2_antennanp ANTENNA_617 (.A(_04727_));
 sg13g2_antennanp ANTENNA_618 (.A(_04727_));
 sg13g2_antennanp ANTENNA_619 (.A(_04763_));
 sg13g2_antennanp ANTENNA_620 (.A(_04763_));
 sg13g2_antennanp ANTENNA_621 (.A(_04763_));
 sg13g2_antennanp ANTENNA_622 (.A(_04763_));
 sg13g2_antennanp ANTENNA_623 (.A(_04798_));
 sg13g2_antennanp ANTENNA_624 (.A(_04798_));
 sg13g2_antennanp ANTENNA_625 (.A(_04798_));
 sg13g2_antennanp ANTENNA_626 (.A(_04798_));
 sg13g2_antennanp ANTENNA_627 (.A(_04832_));
 sg13g2_antennanp ANTENNA_628 (.A(_04832_));
 sg13g2_antennanp ANTENNA_629 (.A(_04832_));
 sg13g2_antennanp ANTENNA_630 (.A(_04832_));
 sg13g2_antennanp ANTENNA_631 (.A(_04900_));
 sg13g2_antennanp ANTENNA_632 (.A(_04900_));
 sg13g2_antennanp ANTENNA_633 (.A(_04900_));
 sg13g2_antennanp ANTENNA_634 (.A(_04900_));
 sg13g2_antennanp ANTENNA_635 (.A(_05910_));
 sg13g2_antennanp ANTENNA_636 (.A(_05910_));
 sg13g2_antennanp ANTENNA_637 (.A(_06251_));
 sg13g2_antennanp ANTENNA_638 (.A(_07613_));
 sg13g2_antennanp ANTENNA_639 (.A(_07613_));
 sg13g2_antennanp ANTENNA_640 (.A(_07613_));
 sg13g2_antennanp ANTENNA_641 (.A(clk));
 sg13g2_antennanp ANTENNA_642 (.A(clk));
 sg13g2_antennanp ANTENNA_643 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_644 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_645 (.A(sclk));
 sg13g2_antennanp ANTENNA_646 (.A(sclk));
 sg13g2_antennanp ANTENNA_647 (.A(sclk));
 sg13g2_antennanp ANTENNA_648 (.A(sclk));
 sg13g2_antennanp ANTENNA_649 (.A(sclk));
 sg13g2_antennanp ANTENNA_650 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_651 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_652 (.A(sio2_o));
 sg13g2_antennanp ANTENNA_653 (.A(\soc_I.kianv_I.datapath_unit_I.A1[0] ));
 sg13g2_antennanp ANTENNA_654 (.A(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_antennanp ANTENNA_655 (.A(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_antennanp ANTENNA_656 (.A(\soc_I.kianv_I.datapath_unit_I.A1[12] ));
 sg13g2_antennanp ANTENNA_657 (.A(\soc_I.kianv_I.datapath_unit_I.A1[15] ));
 sg13g2_antennanp ANTENNA_658 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_659 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_660 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_661 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_662 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_663 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_664 (.A(\soc_I.spi0_I.cen ));
 sg13g2_antennanp ANTENNA_665 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_666 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_667 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_668 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_669 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_670 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_671 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_672 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_673 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_674 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_675 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_676 (.A(net438));
 sg13g2_antennanp ANTENNA_677 (.A(net438));
 sg13g2_antennanp ANTENNA_678 (.A(net438));
 sg13g2_antennanp ANTENNA_679 (.A(net438));
 sg13g2_antennanp ANTENNA_680 (.A(net438));
 sg13g2_antennanp ANTENNA_681 (.A(net438));
 sg13g2_antennanp ANTENNA_682 (.A(net438));
 sg13g2_antennanp ANTENNA_683 (.A(net438));
 sg13g2_antennanp ANTENNA_684 (.A(net438));
 sg13g2_antennanp ANTENNA_685 (.A(net619));
 sg13g2_antennanp ANTENNA_686 (.A(net619));
 sg13g2_antennanp ANTENNA_687 (.A(net619));
 sg13g2_antennanp ANTENNA_688 (.A(net619));
 sg13g2_antennanp ANTENNA_689 (.A(net619));
 sg13g2_antennanp ANTENNA_690 (.A(net619));
 sg13g2_antennanp ANTENNA_691 (.A(net619));
 sg13g2_antennanp ANTENNA_692 (.A(net619));
 sg13g2_antennanp ANTENNA_693 (.A(net619));
 sg13g2_antennanp ANTENNA_694 (.A(net619));
 sg13g2_antennanp ANTENNA_695 (.A(net619));
 sg13g2_antennanp ANTENNA_696 (.A(net619));
 sg13g2_antennanp ANTENNA_697 (.A(net619));
 sg13g2_antennanp ANTENNA_698 (.A(net619));
 sg13g2_antennanp ANTENNA_699 (.A(net619));
 sg13g2_antennanp ANTENNA_700 (.A(net619));
 sg13g2_antennanp ANTENNA_701 (.A(_00220_));
 sg13g2_antennanp ANTENNA_702 (.A(_00222_));
 sg13g2_antennanp ANTENNA_703 (.A(_00224_));
 sg13g2_antennanp ANTENNA_704 (.A(_00262_));
 sg13g2_antennanp ANTENNA_705 (.A(_00263_));
 sg13g2_antennanp ANTENNA_706 (.A(_00263_));
 sg13g2_antennanp ANTENNA_707 (.A(_00922_));
 sg13g2_antennanp ANTENNA_708 (.A(_00922_));
 sg13g2_antennanp ANTENNA_709 (.A(_01573_));
 sg13g2_antennanp ANTENNA_710 (.A(_01573_));
 sg13g2_antennanp ANTENNA_711 (.A(_01573_));
 sg13g2_antennanp ANTENNA_712 (.A(_01573_));
 sg13g2_antennanp ANTENNA_713 (.A(_01573_));
 sg13g2_antennanp ANTENNA_714 (.A(_01573_));
 sg13g2_antennanp ANTENNA_715 (.A(_01840_));
 sg13g2_antennanp ANTENNA_716 (.A(_01840_));
 sg13g2_antennanp ANTENNA_717 (.A(_01840_));
 sg13g2_antennanp ANTENNA_718 (.A(_01840_));
 sg13g2_antennanp ANTENNA_719 (.A(_01840_));
 sg13g2_antennanp ANTENNA_720 (.A(_01840_));
 sg13g2_antennanp ANTENNA_721 (.A(_01903_));
 sg13g2_antennanp ANTENNA_722 (.A(_01903_));
 sg13g2_antennanp ANTENNA_723 (.A(_01903_));
 sg13g2_antennanp ANTENNA_724 (.A(_01903_));
 sg13g2_antennanp ANTENNA_725 (.A(_01903_));
 sg13g2_antennanp ANTENNA_726 (.A(_01903_));
 sg13g2_antennanp ANTENNA_727 (.A(_02081_));
 sg13g2_antennanp ANTENNA_728 (.A(_02081_));
 sg13g2_antennanp ANTENNA_729 (.A(_02081_));
 sg13g2_antennanp ANTENNA_730 (.A(_02081_));
 sg13g2_antennanp ANTENNA_731 (.A(_02081_));
 sg13g2_antennanp ANTENNA_732 (.A(_02081_));
 sg13g2_antennanp ANTENNA_733 (.A(_02081_));
 sg13g2_antennanp ANTENNA_734 (.A(_02081_));
 sg13g2_antennanp ANTENNA_735 (.A(_02081_));
 sg13g2_antennanp ANTENNA_736 (.A(_02081_));
 sg13g2_antennanp ANTENNA_737 (.A(_02081_));
 sg13g2_antennanp ANTENNA_738 (.A(_02081_));
 sg13g2_antennanp ANTENNA_739 (.A(_02081_));
 sg13g2_antennanp ANTENNA_740 (.A(_02081_));
 sg13g2_antennanp ANTENNA_741 (.A(_02081_));
 sg13g2_antennanp ANTENNA_742 (.A(_02081_));
 sg13g2_antennanp ANTENNA_743 (.A(_02081_));
 sg13g2_antennanp ANTENNA_744 (.A(_02537_));
 sg13g2_antennanp ANTENNA_745 (.A(_02558_));
 sg13g2_antennanp ANTENNA_746 (.A(_03712_));
 sg13g2_antennanp ANTENNA_747 (.A(_03714_));
 sg13g2_antennanp ANTENNA_748 (.A(_03714_));
 sg13g2_antennanp ANTENNA_749 (.A(_03714_));
 sg13g2_antennanp ANTENNA_750 (.A(_03714_));
 sg13g2_antennanp ANTENNA_751 (.A(_03720_));
 sg13g2_antennanp ANTENNA_752 (.A(_03760_));
 sg13g2_antennanp ANTENNA_753 (.A(_03975_));
 sg13g2_antennanp ANTENNA_754 (.A(_04273_));
 sg13g2_antennanp ANTENNA_755 (.A(_04273_));
 sg13g2_antennanp ANTENNA_756 (.A(_04273_));
 sg13g2_antennanp ANTENNA_757 (.A(_04273_));
 sg13g2_antennanp ANTENNA_758 (.A(_04273_));
 sg13g2_antennanp ANTENNA_759 (.A(_04273_));
 sg13g2_antennanp ANTENNA_760 (.A(_04693_));
 sg13g2_antennanp ANTENNA_761 (.A(_04693_));
 sg13g2_antennanp ANTENNA_762 (.A(_04693_));
 sg13g2_antennanp ANTENNA_763 (.A(_04693_));
 sg13g2_antennanp ANTENNA_764 (.A(_04727_));
 sg13g2_antennanp ANTENNA_765 (.A(_04727_));
 sg13g2_antennanp ANTENNA_766 (.A(_04727_));
 sg13g2_antennanp ANTENNA_767 (.A(_04727_));
 sg13g2_antennanp ANTENNA_768 (.A(_04763_));
 sg13g2_antennanp ANTENNA_769 (.A(_04763_));
 sg13g2_antennanp ANTENNA_770 (.A(_04763_));
 sg13g2_antennanp ANTENNA_771 (.A(_04763_));
 sg13g2_antennanp ANTENNA_772 (.A(_04798_));
 sg13g2_antennanp ANTENNA_773 (.A(_04798_));
 sg13g2_antennanp ANTENNA_774 (.A(_04798_));
 sg13g2_antennanp ANTENNA_775 (.A(_04798_));
 sg13g2_antennanp ANTENNA_776 (.A(_04832_));
 sg13g2_antennanp ANTENNA_777 (.A(_04832_));
 sg13g2_antennanp ANTENNA_778 (.A(_04832_));
 sg13g2_antennanp ANTENNA_779 (.A(_04832_));
 sg13g2_antennanp ANTENNA_780 (.A(_04900_));
 sg13g2_antennanp ANTENNA_781 (.A(_04900_));
 sg13g2_antennanp ANTENNA_782 (.A(_04900_));
 sg13g2_antennanp ANTENNA_783 (.A(_04900_));
 sg13g2_antennanp ANTENNA_784 (.A(_05910_));
 sg13g2_antennanp ANTENNA_785 (.A(_05910_));
 sg13g2_antennanp ANTENNA_786 (.A(_06251_));
 sg13g2_antennanp ANTENNA_787 (.A(_07613_));
 sg13g2_antennanp ANTENNA_788 (.A(_07613_));
 sg13g2_antennanp ANTENNA_789 (.A(_07613_));
 sg13g2_antennanp ANTENNA_790 (.A(clk));
 sg13g2_antennanp ANTENNA_791 (.A(clk));
 sg13g2_antennanp ANTENNA_792 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_793 (.A(pwm_o));
 sg13g2_antennanp ANTENNA_794 (.A(sclk));
 sg13g2_antennanp ANTENNA_795 (.A(sclk));
 sg13g2_antennanp ANTENNA_796 (.A(sclk));
 sg13g2_antennanp ANTENNA_797 (.A(sclk));
 sg13g2_antennanp ANTENNA_798 (.A(sclk));
 sg13g2_antennanp ANTENNA_799 (.A(\soc_I.kianv_I.datapath_unit_I.A1[0] ));
 sg13g2_antennanp ANTENNA_800 (.A(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_antennanp ANTENNA_801 (.A(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_antennanp ANTENNA_802 (.A(\soc_I.kianv_I.datapath_unit_I.A1[12] ));
 sg13g2_antennanp ANTENNA_803 (.A(\soc_I.kianv_I.datapath_unit_I.A1[15] ));
 sg13g2_antennanp ANTENNA_804 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_805 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_806 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_807 (.A(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_antennanp ANTENNA_808 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_809 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_810 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_811 (.A(\soc_I.spi0_I.sclk ));
 sg13g2_antennanp ANTENNA_812 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_813 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_814 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_815 (.A(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_antennanp ANTENNA_816 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_817 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_818 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_819 (.A(\soc_I.tx_uart_i.tx_out ));
 sg13g2_antennanp ANTENNA_820 (.A(net619));
 sg13g2_antennanp ANTENNA_821 (.A(net619));
 sg13g2_antennanp ANTENNA_822 (.A(net619));
 sg13g2_antennanp ANTENNA_823 (.A(net619));
 sg13g2_antennanp ANTENNA_824 (.A(net619));
 sg13g2_antennanp ANTENNA_825 (.A(net619));
 sg13g2_antennanp ANTENNA_826 (.A(net619));
 sg13g2_antennanp ANTENNA_827 (.A(net619));
 sg13g2_antennanp ANTENNA_828 (.A(net619));
 sg13g2_antennanp ANTENNA_829 (.A(net619));
 sg13g2_antennanp ANTENNA_830 (.A(net619));
 sg13g2_antennanp ANTENNA_831 (.A(net619));
 sg13g2_antennanp ANTENNA_832 (.A(net619));
 sg13g2_antennanp ANTENNA_833 (.A(net619));
 sg13g2_antennanp ANTENNA_834 (.A(net619));
 sg13g2_antennanp ANTENNA_835 (.A(net619));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_4 FILLER_0_63 ();
 sg13g2_fill_2 FILLER_0_97 ();
 sg13g2_decap_8 FILLER_0_129 ();
 sg13g2_decap_8 FILLER_0_136 ();
 sg13g2_decap_8 FILLER_0_143 ();
 sg13g2_decap_4 FILLER_0_150 ();
 sg13g2_fill_1 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_190 ();
 sg13g2_decap_8 FILLER_0_197 ();
 sg13g2_decap_8 FILLER_0_204 ();
 sg13g2_fill_1 FILLER_0_211 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_fill_2 FILLER_0_228 ();
 sg13g2_fill_1 FILLER_0_230 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_fill_1 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_4 FILLER_0_268 ();
 sg13g2_fill_2 FILLER_0_272 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_fill_2 FILLER_0_297 ();
 sg13g2_fill_1 FILLER_0_299 ();
 sg13g2_fill_2 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_4 FILLER_0_322 ();
 sg13g2_fill_1 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_340 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_4 FILLER_0_354 ();
 sg13g2_fill_2 FILLER_0_362 ();
 sg13g2_fill_1 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_decap_8 FILLER_0_422 ();
 sg13g2_decap_4 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_fill_2 FILLER_0_462 ();
 sg13g2_fill_1 FILLER_0_464 ();
 sg13g2_decap_4 FILLER_0_495 ();
 sg13g2_decap_8 FILLER_0_503 ();
 sg13g2_decap_8 FILLER_0_510 ();
 sg13g2_decap_8 FILLER_0_517 ();
 sg13g2_fill_2 FILLER_0_524 ();
 sg13g2_fill_1 FILLER_0_526 ();
 sg13g2_decap_8 FILLER_0_561 ();
 sg13g2_decap_8 FILLER_0_568 ();
 sg13g2_decap_8 FILLER_0_575 ();
 sg13g2_fill_1 FILLER_0_582 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_4 FILLER_0_616 ();
 sg13g2_fill_1 FILLER_0_620 ();
 sg13g2_fill_2 FILLER_0_647 ();
 sg13g2_fill_2 FILLER_0_679 ();
 sg13g2_fill_1 FILLER_0_692 ();
 sg13g2_fill_1 FILLER_0_697 ();
 sg13g2_fill_1 FILLER_0_702 ();
 sg13g2_fill_1 FILLER_0_708 ();
 sg13g2_fill_1 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_761 ();
 sg13g2_decap_8 FILLER_0_768 ();
 sg13g2_decap_8 FILLER_0_775 ();
 sg13g2_decap_8 FILLER_0_782 ();
 sg13g2_fill_2 FILLER_0_789 ();
 sg13g2_decap_8 FILLER_0_795 ();
 sg13g2_fill_1 FILLER_0_802 ();
 sg13g2_fill_2 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_4 FILLER_0_826 ();
 sg13g2_decap_4 FILLER_0_860 ();
 sg13g2_decap_4 FILLER_0_873 ();
 sg13g2_decap_8 FILLER_0_886 ();
 sg13g2_fill_1 FILLER_0_893 ();
 sg13g2_fill_2 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_909 ();
 sg13g2_decap_8 FILLER_0_916 ();
 sg13g2_decap_8 FILLER_0_923 ();
 sg13g2_fill_1 FILLER_0_930 ();
 sg13g2_decap_8 FILLER_0_965 ();
 sg13g2_decap_8 FILLER_0_972 ();
 sg13g2_decap_8 FILLER_0_979 ();
 sg13g2_fill_2 FILLER_0_986 ();
 sg13g2_fill_1 FILLER_0_988 ();
 sg13g2_fill_1 FILLER_0_993 ();
 sg13g2_decap_4 FILLER_0_999 ();
 sg13g2_fill_1 FILLER_0_1012 ();
 sg13g2_decap_8 FILLER_0_1017 ();
 sg13g2_decap_8 FILLER_0_1024 ();
 sg13g2_decap_8 FILLER_0_1031 ();
 sg13g2_fill_2 FILLER_0_1038 ();
 sg13g2_decap_8 FILLER_0_1045 ();
 sg13g2_decap_8 FILLER_0_1082 ();
 sg13g2_fill_1 FILLER_0_1089 ();
 sg13g2_decap_8 FILLER_0_1099 ();
 sg13g2_fill_2 FILLER_0_1106 ();
 sg13g2_fill_1 FILLER_0_1108 ();
 sg13g2_fill_2 FILLER_0_1118 ();
 sg13g2_fill_1 FILLER_0_1120 ();
 sg13g2_decap_8 FILLER_0_1125 ();
 sg13g2_decap_8 FILLER_0_1132 ();
 sg13g2_decap_8 FILLER_0_1139 ();
 sg13g2_decap_8 FILLER_0_1146 ();
 sg13g2_decap_8 FILLER_0_1153 ();
 sg13g2_decap_8 FILLER_0_1160 ();
 sg13g2_decap_8 FILLER_0_1167 ();
 sg13g2_decap_8 FILLER_0_1174 ();
 sg13g2_decap_8 FILLER_0_1181 ();
 sg13g2_decap_8 FILLER_0_1188 ();
 sg13g2_decap_8 FILLER_0_1195 ();
 sg13g2_decap_8 FILLER_0_1202 ();
 sg13g2_decap_8 FILLER_0_1209 ();
 sg13g2_decap_8 FILLER_0_1216 ();
 sg13g2_decap_8 FILLER_0_1223 ();
 sg13g2_decap_8 FILLER_0_1230 ();
 sg13g2_decap_8 FILLER_0_1237 ();
 sg13g2_decap_8 FILLER_0_1244 ();
 sg13g2_decap_8 FILLER_0_1251 ();
 sg13g2_decap_8 FILLER_0_1258 ();
 sg13g2_decap_8 FILLER_0_1265 ();
 sg13g2_decap_8 FILLER_0_1272 ();
 sg13g2_decap_8 FILLER_0_1279 ();
 sg13g2_decap_8 FILLER_0_1286 ();
 sg13g2_decap_8 FILLER_0_1293 ();
 sg13g2_decap_8 FILLER_0_1300 ();
 sg13g2_decap_8 FILLER_0_1307 ();
 sg13g2_decap_8 FILLER_0_1314 ();
 sg13g2_decap_8 FILLER_0_1321 ();
 sg13g2_decap_8 FILLER_0_1328 ();
 sg13g2_decap_8 FILLER_0_1335 ();
 sg13g2_decap_8 FILLER_0_1342 ();
 sg13g2_decap_8 FILLER_0_1349 ();
 sg13g2_decap_8 FILLER_0_1356 ();
 sg13g2_decap_8 FILLER_0_1363 ();
 sg13g2_decap_8 FILLER_0_1370 ();
 sg13g2_decap_8 FILLER_0_1377 ();
 sg13g2_decap_8 FILLER_0_1384 ();
 sg13g2_decap_8 FILLER_0_1391 ();
 sg13g2_decap_8 FILLER_0_1398 ();
 sg13g2_decap_8 FILLER_0_1405 ();
 sg13g2_decap_8 FILLER_0_1412 ();
 sg13g2_decap_8 FILLER_0_1419 ();
 sg13g2_decap_8 FILLER_0_1426 ();
 sg13g2_decap_8 FILLER_0_1433 ();
 sg13g2_decap_8 FILLER_0_1440 ();
 sg13g2_decap_8 FILLER_0_1447 ();
 sg13g2_decap_8 FILLER_0_1454 ();
 sg13g2_decap_8 FILLER_0_1461 ();
 sg13g2_decap_8 FILLER_0_1468 ();
 sg13g2_decap_8 FILLER_0_1475 ();
 sg13g2_decap_8 FILLER_0_1482 ();
 sg13g2_decap_8 FILLER_0_1489 ();
 sg13g2_decap_8 FILLER_0_1496 ();
 sg13g2_decap_8 FILLER_0_1503 ();
 sg13g2_decap_8 FILLER_0_1510 ();
 sg13g2_decap_8 FILLER_0_1517 ();
 sg13g2_decap_8 FILLER_0_1524 ();
 sg13g2_decap_8 FILLER_0_1531 ();
 sg13g2_decap_8 FILLER_0_1538 ();
 sg13g2_decap_8 FILLER_0_1545 ();
 sg13g2_decap_8 FILLER_0_1552 ();
 sg13g2_decap_8 FILLER_0_1559 ();
 sg13g2_decap_8 FILLER_0_1566 ();
 sg13g2_decap_8 FILLER_0_1573 ();
 sg13g2_decap_8 FILLER_0_1580 ();
 sg13g2_decap_8 FILLER_0_1587 ();
 sg13g2_decap_8 FILLER_0_1594 ();
 sg13g2_decap_8 FILLER_0_1601 ();
 sg13g2_decap_8 FILLER_0_1608 ();
 sg13g2_decap_8 FILLER_0_1615 ();
 sg13g2_decap_8 FILLER_0_1622 ();
 sg13g2_decap_8 FILLER_0_1629 ();
 sg13g2_decap_8 FILLER_0_1636 ();
 sg13g2_decap_8 FILLER_0_1643 ();
 sg13g2_decap_8 FILLER_0_1650 ();
 sg13g2_decap_8 FILLER_0_1657 ();
 sg13g2_decap_8 FILLER_0_1664 ();
 sg13g2_decap_8 FILLER_0_1671 ();
 sg13g2_decap_8 FILLER_0_1678 ();
 sg13g2_decap_8 FILLER_0_1685 ();
 sg13g2_decap_8 FILLER_0_1692 ();
 sg13g2_decap_8 FILLER_0_1699 ();
 sg13g2_decap_8 FILLER_0_1706 ();
 sg13g2_decap_8 FILLER_0_1713 ();
 sg13g2_decap_8 FILLER_0_1720 ();
 sg13g2_decap_8 FILLER_0_1727 ();
 sg13g2_decap_8 FILLER_0_1734 ();
 sg13g2_decap_8 FILLER_0_1741 ();
 sg13g2_decap_8 FILLER_0_1748 ();
 sg13g2_decap_8 FILLER_0_1755 ();
 sg13g2_decap_8 FILLER_0_1762 ();
 sg13g2_decap_4 FILLER_0_1769 ();
 sg13g2_fill_1 FILLER_0_1773 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_75 ();
 sg13g2_fill_1 FILLER_1_81 ();
 sg13g2_fill_2 FILLER_1_86 ();
 sg13g2_decap_8 FILLER_1_118 ();
 sg13g2_decap_8 FILLER_1_125 ();
 sg13g2_fill_1 FILLER_1_132 ();
 sg13g2_fill_2 FILLER_1_137 ();
 sg13g2_decap_4 FILLER_1_144 ();
 sg13g2_fill_1 FILLER_1_148 ();
 sg13g2_decap_8 FILLER_1_262 ();
 sg13g2_fill_2 FILLER_1_269 ();
 sg13g2_fill_1 FILLER_1_271 ();
 sg13g2_decap_4 FILLER_1_376 ();
 sg13g2_fill_2 FILLER_1_380 ();
 sg13g2_fill_2 FILLER_1_392 ();
 sg13g2_fill_1 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_409 ();
 sg13g2_decap_8 FILLER_1_416 ();
 sg13g2_fill_2 FILLER_1_423 ();
 sg13g2_decap_8 FILLER_1_456 ();
 sg13g2_decap_4 FILLER_1_463 ();
 sg13g2_fill_1 FILLER_1_481 ();
 sg13g2_fill_2 FILLER_1_486 ();
 sg13g2_decap_4 FILLER_1_519 ();
 sg13g2_fill_1 FILLER_1_528 ();
 sg13g2_decap_4 FILLER_1_533 ();
 sg13g2_fill_1 FILLER_1_537 ();
 sg13g2_fill_1 FILLER_1_543 ();
 sg13g2_fill_1 FILLER_1_557 ();
 sg13g2_decap_8 FILLER_1_566 ();
 sg13g2_decap_8 FILLER_1_573 ();
 sg13g2_fill_1 FILLER_1_580 ();
 sg13g2_fill_1 FILLER_1_590 ();
 sg13g2_decap_4 FILLER_1_595 ();
 sg13g2_fill_2 FILLER_1_599 ();
 sg13g2_decap_8 FILLER_1_605 ();
 sg13g2_decap_4 FILLER_1_612 ();
 sg13g2_decap_4 FILLER_1_626 ();
 sg13g2_decap_8 FILLER_1_634 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_4 FILLER_1_662 ();
 sg13g2_fill_1 FILLER_1_692 ();
 sg13g2_fill_1 FILLER_1_696 ();
 sg13g2_fill_2 FILLER_1_725 ();
 sg13g2_fill_1 FILLER_1_739 ();
 sg13g2_fill_1 FILLER_1_743 ();
 sg13g2_fill_2 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_925 ();
 sg13g2_fill_1 FILLER_1_932 ();
 sg13g2_fill_2 FILLER_1_942 ();
 sg13g2_fill_1 FILLER_1_944 ();
 sg13g2_fill_2 FILLER_1_1067 ();
 sg13g2_fill_1 FILLER_1_1069 ();
 sg13g2_decap_8 FILLER_1_1074 ();
 sg13g2_decap_4 FILLER_1_1081 ();
 sg13g2_decap_8 FILLER_1_1137 ();
 sg13g2_decap_8 FILLER_1_1144 ();
 sg13g2_decap_8 FILLER_1_1151 ();
 sg13g2_decap_8 FILLER_1_1158 ();
 sg13g2_decap_8 FILLER_1_1165 ();
 sg13g2_decap_8 FILLER_1_1172 ();
 sg13g2_decap_8 FILLER_1_1179 ();
 sg13g2_decap_8 FILLER_1_1186 ();
 sg13g2_decap_8 FILLER_1_1193 ();
 sg13g2_decap_8 FILLER_1_1200 ();
 sg13g2_decap_8 FILLER_1_1207 ();
 sg13g2_decap_8 FILLER_1_1214 ();
 sg13g2_decap_8 FILLER_1_1221 ();
 sg13g2_decap_8 FILLER_1_1228 ();
 sg13g2_decap_8 FILLER_1_1235 ();
 sg13g2_decap_8 FILLER_1_1242 ();
 sg13g2_decap_8 FILLER_1_1249 ();
 sg13g2_decap_8 FILLER_1_1256 ();
 sg13g2_decap_8 FILLER_1_1263 ();
 sg13g2_decap_8 FILLER_1_1270 ();
 sg13g2_decap_8 FILLER_1_1277 ();
 sg13g2_decap_8 FILLER_1_1284 ();
 sg13g2_decap_8 FILLER_1_1291 ();
 sg13g2_decap_8 FILLER_1_1298 ();
 sg13g2_decap_8 FILLER_1_1305 ();
 sg13g2_decap_8 FILLER_1_1312 ();
 sg13g2_decap_8 FILLER_1_1319 ();
 sg13g2_decap_8 FILLER_1_1326 ();
 sg13g2_decap_8 FILLER_1_1333 ();
 sg13g2_decap_8 FILLER_1_1340 ();
 sg13g2_decap_8 FILLER_1_1347 ();
 sg13g2_decap_8 FILLER_1_1354 ();
 sg13g2_decap_8 FILLER_1_1361 ();
 sg13g2_decap_8 FILLER_1_1368 ();
 sg13g2_decap_8 FILLER_1_1375 ();
 sg13g2_decap_8 FILLER_1_1382 ();
 sg13g2_decap_8 FILLER_1_1389 ();
 sg13g2_decap_8 FILLER_1_1396 ();
 sg13g2_decap_8 FILLER_1_1403 ();
 sg13g2_decap_8 FILLER_1_1410 ();
 sg13g2_decap_8 FILLER_1_1417 ();
 sg13g2_decap_8 FILLER_1_1424 ();
 sg13g2_decap_8 FILLER_1_1431 ();
 sg13g2_decap_8 FILLER_1_1438 ();
 sg13g2_decap_8 FILLER_1_1445 ();
 sg13g2_decap_8 FILLER_1_1452 ();
 sg13g2_decap_8 FILLER_1_1459 ();
 sg13g2_decap_8 FILLER_1_1466 ();
 sg13g2_decap_8 FILLER_1_1473 ();
 sg13g2_decap_8 FILLER_1_1480 ();
 sg13g2_decap_8 FILLER_1_1487 ();
 sg13g2_decap_8 FILLER_1_1494 ();
 sg13g2_decap_8 FILLER_1_1501 ();
 sg13g2_decap_8 FILLER_1_1508 ();
 sg13g2_decap_8 FILLER_1_1515 ();
 sg13g2_decap_8 FILLER_1_1522 ();
 sg13g2_decap_8 FILLER_1_1529 ();
 sg13g2_decap_8 FILLER_1_1536 ();
 sg13g2_decap_8 FILLER_1_1543 ();
 sg13g2_decap_8 FILLER_1_1550 ();
 sg13g2_decap_8 FILLER_1_1557 ();
 sg13g2_decap_8 FILLER_1_1564 ();
 sg13g2_decap_8 FILLER_1_1571 ();
 sg13g2_decap_8 FILLER_1_1578 ();
 sg13g2_decap_8 FILLER_1_1585 ();
 sg13g2_decap_8 FILLER_1_1592 ();
 sg13g2_decap_8 FILLER_1_1599 ();
 sg13g2_decap_8 FILLER_1_1606 ();
 sg13g2_decap_8 FILLER_1_1613 ();
 sg13g2_decap_8 FILLER_1_1620 ();
 sg13g2_decap_8 FILLER_1_1627 ();
 sg13g2_decap_8 FILLER_1_1634 ();
 sg13g2_decap_8 FILLER_1_1641 ();
 sg13g2_decap_8 FILLER_1_1648 ();
 sg13g2_decap_8 FILLER_1_1655 ();
 sg13g2_decap_8 FILLER_1_1662 ();
 sg13g2_decap_8 FILLER_1_1669 ();
 sg13g2_decap_8 FILLER_1_1676 ();
 sg13g2_decap_8 FILLER_1_1683 ();
 sg13g2_decap_8 FILLER_1_1690 ();
 sg13g2_decap_8 FILLER_1_1697 ();
 sg13g2_decap_8 FILLER_1_1704 ();
 sg13g2_decap_8 FILLER_1_1711 ();
 sg13g2_decap_8 FILLER_1_1718 ();
 sg13g2_decap_8 FILLER_1_1725 ();
 sg13g2_decap_8 FILLER_1_1732 ();
 sg13g2_decap_8 FILLER_1_1739 ();
 sg13g2_decap_8 FILLER_1_1746 ();
 sg13g2_decap_8 FILLER_1_1753 ();
 sg13g2_decap_8 FILLER_1_1760 ();
 sg13g2_decap_8 FILLER_1_1767 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_fill_1 FILLER_2_35 ();
 sg13g2_decap_4 FILLER_2_41 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_83 ();
 sg13g2_fill_2 FILLER_2_90 ();
 sg13g2_fill_1 FILLER_2_92 ();
 sg13g2_decap_8 FILLER_2_114 ();
 sg13g2_decap_4 FILLER_2_121 ();
 sg13g2_fill_1 FILLER_2_125 ();
 sg13g2_fill_2 FILLER_2_156 ();
 sg13g2_fill_1 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_184 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_decap_4 FILLER_2_198 ();
 sg13g2_fill_2 FILLER_2_202 ();
 sg13g2_decap_4 FILLER_2_213 ();
 sg13g2_decap_4 FILLER_2_242 ();
 sg13g2_fill_2 FILLER_2_255 ();
 sg13g2_fill_1 FILLER_2_257 ();
 sg13g2_decap_8 FILLER_2_262 ();
 sg13g2_decap_8 FILLER_2_269 ();
 sg13g2_decap_4 FILLER_2_276 ();
 sg13g2_fill_2 FILLER_2_280 ();
 sg13g2_fill_2 FILLER_2_303 ();
 sg13g2_fill_1 FILLER_2_305 ();
 sg13g2_fill_2 FILLER_2_327 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_4 FILLER_2_354 ();
 sg13g2_fill_2 FILLER_2_368 ();
 sg13g2_decap_4 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_425 ();
 sg13g2_fill_2 FILLER_2_432 ();
 sg13g2_fill_1 FILLER_2_443 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_fill_2 FILLER_2_455 ();
 sg13g2_fill_2 FILLER_2_483 ();
 sg13g2_fill_2 FILLER_2_506 ();
 sg13g2_fill_1 FILLER_2_508 ();
 sg13g2_fill_2 FILLER_2_513 ();
 sg13g2_fill_1 FILLER_2_515 ();
 sg13g2_fill_2 FILLER_2_542 ();
 sg13g2_fill_1 FILLER_2_544 ();
 sg13g2_decap_4 FILLER_2_576 ();
 sg13g2_fill_2 FILLER_2_585 ();
 sg13g2_fill_1 FILLER_2_618 ();
 sg13g2_decap_8 FILLER_2_649 ();
 sg13g2_decap_8 FILLER_2_656 ();
 sg13g2_decap_4 FILLER_2_663 ();
 sg13g2_fill_1 FILLER_2_688 ();
 sg13g2_fill_1 FILLER_2_739 ();
 sg13g2_decap_4 FILLER_2_750 ();
 sg13g2_decap_8 FILLER_2_764 ();
 sg13g2_fill_2 FILLER_2_771 ();
 sg13g2_decap_4 FILLER_2_800 ();
 sg13g2_decap_8 FILLER_2_825 ();
 sg13g2_decap_8 FILLER_2_832 ();
 sg13g2_fill_2 FILLER_2_839 ();
 sg13g2_decap_4 FILLER_2_851 ();
 sg13g2_decap_4 FILLER_2_880 ();
 sg13g2_fill_2 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_895 ();
 sg13g2_decap_4 FILLER_2_902 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_fill_1 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_948 ();
 sg13g2_decap_8 FILLER_2_955 ();
 sg13g2_decap_8 FILLER_2_962 ();
 sg13g2_decap_8 FILLER_2_969 ();
 sg13g2_fill_2 FILLER_2_976 ();
 sg13g2_fill_1 FILLER_2_978 ();
 sg13g2_fill_2 FILLER_2_997 ();
 sg13g2_fill_1 FILLER_2_999 ();
 sg13g2_decap_8 FILLER_2_1004 ();
 sg13g2_decap_8 FILLER_2_1011 ();
 sg13g2_fill_2 FILLER_2_1023 ();
 sg13g2_fill_1 FILLER_2_1025 ();
 sg13g2_decap_4 FILLER_2_1030 ();
 sg13g2_fill_1 FILLER_2_1034 ();
 sg13g2_decap_4 FILLER_2_1039 ();
 sg13g2_fill_1 FILLER_2_1043 ();
 sg13g2_fill_2 FILLER_2_1048 ();
 sg13g2_fill_1 FILLER_2_1050 ();
 sg13g2_decap_8 FILLER_2_1082 ();
 sg13g2_decap_4 FILLER_2_1089 ();
 sg13g2_decap_8 FILLER_2_1097 ();
 sg13g2_decap_8 FILLER_2_1125 ();
 sg13g2_decap_8 FILLER_2_1158 ();
 sg13g2_decap_8 FILLER_2_1165 ();
 sg13g2_decap_8 FILLER_2_1172 ();
 sg13g2_decap_8 FILLER_2_1179 ();
 sg13g2_decap_8 FILLER_2_1186 ();
 sg13g2_decap_8 FILLER_2_1193 ();
 sg13g2_decap_8 FILLER_2_1200 ();
 sg13g2_decap_8 FILLER_2_1207 ();
 sg13g2_decap_8 FILLER_2_1214 ();
 sg13g2_decap_8 FILLER_2_1221 ();
 sg13g2_decap_8 FILLER_2_1228 ();
 sg13g2_decap_8 FILLER_2_1235 ();
 sg13g2_decap_8 FILLER_2_1242 ();
 sg13g2_decap_8 FILLER_2_1249 ();
 sg13g2_decap_8 FILLER_2_1256 ();
 sg13g2_decap_8 FILLER_2_1263 ();
 sg13g2_decap_8 FILLER_2_1270 ();
 sg13g2_decap_8 FILLER_2_1277 ();
 sg13g2_decap_8 FILLER_2_1284 ();
 sg13g2_decap_8 FILLER_2_1291 ();
 sg13g2_decap_8 FILLER_2_1298 ();
 sg13g2_decap_8 FILLER_2_1305 ();
 sg13g2_decap_8 FILLER_2_1312 ();
 sg13g2_decap_8 FILLER_2_1319 ();
 sg13g2_decap_8 FILLER_2_1326 ();
 sg13g2_decap_8 FILLER_2_1333 ();
 sg13g2_decap_8 FILLER_2_1340 ();
 sg13g2_decap_8 FILLER_2_1347 ();
 sg13g2_decap_8 FILLER_2_1354 ();
 sg13g2_decap_8 FILLER_2_1361 ();
 sg13g2_decap_8 FILLER_2_1368 ();
 sg13g2_decap_8 FILLER_2_1375 ();
 sg13g2_decap_8 FILLER_2_1382 ();
 sg13g2_decap_8 FILLER_2_1389 ();
 sg13g2_decap_8 FILLER_2_1396 ();
 sg13g2_decap_8 FILLER_2_1403 ();
 sg13g2_decap_8 FILLER_2_1410 ();
 sg13g2_decap_8 FILLER_2_1417 ();
 sg13g2_decap_8 FILLER_2_1424 ();
 sg13g2_decap_8 FILLER_2_1431 ();
 sg13g2_decap_8 FILLER_2_1438 ();
 sg13g2_decap_8 FILLER_2_1445 ();
 sg13g2_decap_8 FILLER_2_1452 ();
 sg13g2_decap_8 FILLER_2_1459 ();
 sg13g2_decap_8 FILLER_2_1466 ();
 sg13g2_decap_8 FILLER_2_1473 ();
 sg13g2_decap_8 FILLER_2_1480 ();
 sg13g2_decap_8 FILLER_2_1487 ();
 sg13g2_decap_8 FILLER_2_1494 ();
 sg13g2_decap_8 FILLER_2_1501 ();
 sg13g2_decap_8 FILLER_2_1508 ();
 sg13g2_decap_8 FILLER_2_1515 ();
 sg13g2_decap_8 FILLER_2_1522 ();
 sg13g2_decap_8 FILLER_2_1529 ();
 sg13g2_decap_8 FILLER_2_1536 ();
 sg13g2_decap_8 FILLER_2_1543 ();
 sg13g2_decap_8 FILLER_2_1550 ();
 sg13g2_decap_8 FILLER_2_1557 ();
 sg13g2_decap_8 FILLER_2_1564 ();
 sg13g2_decap_8 FILLER_2_1571 ();
 sg13g2_decap_8 FILLER_2_1578 ();
 sg13g2_decap_8 FILLER_2_1585 ();
 sg13g2_decap_8 FILLER_2_1592 ();
 sg13g2_decap_8 FILLER_2_1599 ();
 sg13g2_decap_8 FILLER_2_1606 ();
 sg13g2_decap_8 FILLER_2_1613 ();
 sg13g2_decap_8 FILLER_2_1620 ();
 sg13g2_decap_8 FILLER_2_1627 ();
 sg13g2_decap_8 FILLER_2_1634 ();
 sg13g2_decap_8 FILLER_2_1641 ();
 sg13g2_decap_8 FILLER_2_1648 ();
 sg13g2_decap_8 FILLER_2_1655 ();
 sg13g2_decap_8 FILLER_2_1662 ();
 sg13g2_decap_8 FILLER_2_1669 ();
 sg13g2_decap_8 FILLER_2_1676 ();
 sg13g2_decap_8 FILLER_2_1683 ();
 sg13g2_decap_8 FILLER_2_1690 ();
 sg13g2_decap_8 FILLER_2_1697 ();
 sg13g2_decap_8 FILLER_2_1704 ();
 sg13g2_decap_8 FILLER_2_1711 ();
 sg13g2_decap_8 FILLER_2_1718 ();
 sg13g2_decap_8 FILLER_2_1725 ();
 sg13g2_decap_8 FILLER_2_1732 ();
 sg13g2_decap_8 FILLER_2_1739 ();
 sg13g2_decap_8 FILLER_2_1746 ();
 sg13g2_decap_8 FILLER_2_1753 ();
 sg13g2_decap_8 FILLER_2_1760 ();
 sg13g2_decap_8 FILLER_2_1767 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_fill_2 FILLER_3_21 ();
 sg13g2_fill_1 FILLER_3_23 ();
 sg13g2_fill_2 FILLER_3_50 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_fill_2 FILLER_3_63 ();
 sg13g2_fill_1 FILLER_3_79 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_fill_2 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_104 ();
 sg13g2_decap_8 FILLER_3_111 ();
 sg13g2_decap_4 FILLER_3_118 ();
 sg13g2_fill_1 FILLER_3_122 ();
 sg13g2_decap_8 FILLER_3_127 ();
 sg13g2_decap_8 FILLER_3_134 ();
 sg13g2_decap_4 FILLER_3_141 ();
 sg13g2_fill_2 FILLER_3_145 ();
 sg13g2_decap_4 FILLER_3_152 ();
 sg13g2_decap_8 FILLER_3_177 ();
 sg13g2_fill_2 FILLER_3_184 ();
 sg13g2_decap_4 FILLER_3_216 ();
 sg13g2_fill_1 FILLER_3_220 ();
 sg13g2_decap_4 FILLER_3_242 ();
 sg13g2_fill_2 FILLER_3_246 ();
 sg13g2_fill_1 FILLER_3_278 ();
 sg13g2_fill_2 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_328 ();
 sg13g2_decap_4 FILLER_3_335 ();
 sg13g2_decap_4 FILLER_3_365 ();
 sg13g2_fill_1 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_fill_1 FILLER_3_398 ();
 sg13g2_decap_8 FILLER_3_412 ();
 sg13g2_decap_8 FILLER_3_419 ();
 sg13g2_fill_1 FILLER_3_426 ();
 sg13g2_decap_8 FILLER_3_453 ();
 sg13g2_fill_2 FILLER_3_460 ();
 sg13g2_decap_8 FILLER_3_466 ();
 sg13g2_decap_8 FILLER_3_473 ();
 sg13g2_decap_4 FILLER_3_480 ();
 sg13g2_fill_2 FILLER_3_484 ();
 sg13g2_decap_8 FILLER_3_507 ();
 sg13g2_decap_8 FILLER_3_514 ();
 sg13g2_fill_2 FILLER_3_521 ();
 sg13g2_decap_4 FILLER_3_528 ();
 sg13g2_fill_1 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_537 ();
 sg13g2_fill_2 FILLER_3_544 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_fill_2 FILLER_3_574 ();
 sg13g2_decap_4 FILLER_3_606 ();
 sg13g2_fill_1 FILLER_3_610 ();
 sg13g2_decap_8 FILLER_3_615 ();
 sg13g2_fill_2 FILLER_3_622 ();
 sg13g2_decap_4 FILLER_3_634 ();
 sg13g2_fill_1 FILLER_3_638 ();
 sg13g2_fill_2 FILLER_3_689 ();
 sg13g2_fill_1 FILLER_3_730 ();
 sg13g2_fill_1 FILLER_3_778 ();
 sg13g2_fill_1 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_827 ();
 sg13g2_fill_1 FILLER_3_834 ();
 sg13g2_fill_2 FILLER_3_882 ();
 sg13g2_fill_1 FILLER_3_884 ();
 sg13g2_decap_8 FILLER_3_916 ();
 sg13g2_decap_8 FILLER_3_928 ();
 sg13g2_decap_8 FILLER_3_935 ();
 sg13g2_fill_2 FILLER_3_946 ();
 sg13g2_fill_1 FILLER_3_969 ();
 sg13g2_fill_2 FILLER_3_1017 ();
 sg13g2_decap_8 FILLER_3_1045 ();
 sg13g2_fill_2 FILLER_3_1077 ();
 sg13g2_fill_1 FILLER_3_1079 ();
 sg13g2_decap_8 FILLER_3_1140 ();
 sg13g2_decap_8 FILLER_3_1147 ();
 sg13g2_decap_8 FILLER_3_1154 ();
 sg13g2_decap_8 FILLER_3_1161 ();
 sg13g2_decap_8 FILLER_3_1168 ();
 sg13g2_decap_8 FILLER_3_1175 ();
 sg13g2_decap_8 FILLER_3_1182 ();
 sg13g2_decap_8 FILLER_3_1189 ();
 sg13g2_decap_8 FILLER_3_1196 ();
 sg13g2_decap_8 FILLER_3_1203 ();
 sg13g2_decap_8 FILLER_3_1210 ();
 sg13g2_decap_8 FILLER_3_1217 ();
 sg13g2_decap_8 FILLER_3_1224 ();
 sg13g2_decap_8 FILLER_3_1231 ();
 sg13g2_decap_8 FILLER_3_1238 ();
 sg13g2_decap_8 FILLER_3_1245 ();
 sg13g2_decap_8 FILLER_3_1252 ();
 sg13g2_decap_8 FILLER_3_1259 ();
 sg13g2_decap_8 FILLER_3_1266 ();
 sg13g2_decap_8 FILLER_3_1273 ();
 sg13g2_decap_8 FILLER_3_1280 ();
 sg13g2_decap_8 FILLER_3_1287 ();
 sg13g2_decap_8 FILLER_3_1294 ();
 sg13g2_decap_8 FILLER_3_1301 ();
 sg13g2_decap_8 FILLER_3_1308 ();
 sg13g2_decap_8 FILLER_3_1315 ();
 sg13g2_decap_8 FILLER_3_1322 ();
 sg13g2_decap_8 FILLER_3_1329 ();
 sg13g2_decap_8 FILLER_3_1336 ();
 sg13g2_decap_8 FILLER_3_1343 ();
 sg13g2_decap_8 FILLER_3_1350 ();
 sg13g2_decap_8 FILLER_3_1357 ();
 sg13g2_decap_8 FILLER_3_1364 ();
 sg13g2_decap_8 FILLER_3_1371 ();
 sg13g2_decap_8 FILLER_3_1378 ();
 sg13g2_decap_8 FILLER_3_1385 ();
 sg13g2_decap_8 FILLER_3_1392 ();
 sg13g2_decap_8 FILLER_3_1399 ();
 sg13g2_decap_8 FILLER_3_1406 ();
 sg13g2_decap_8 FILLER_3_1413 ();
 sg13g2_decap_8 FILLER_3_1420 ();
 sg13g2_decap_8 FILLER_3_1427 ();
 sg13g2_decap_8 FILLER_3_1434 ();
 sg13g2_decap_8 FILLER_3_1441 ();
 sg13g2_decap_8 FILLER_3_1448 ();
 sg13g2_decap_8 FILLER_3_1455 ();
 sg13g2_decap_8 FILLER_3_1462 ();
 sg13g2_decap_8 FILLER_3_1469 ();
 sg13g2_decap_8 FILLER_3_1476 ();
 sg13g2_decap_8 FILLER_3_1483 ();
 sg13g2_decap_8 FILLER_3_1490 ();
 sg13g2_decap_8 FILLER_3_1497 ();
 sg13g2_decap_8 FILLER_3_1504 ();
 sg13g2_decap_8 FILLER_3_1511 ();
 sg13g2_decap_8 FILLER_3_1518 ();
 sg13g2_decap_8 FILLER_3_1525 ();
 sg13g2_decap_8 FILLER_3_1532 ();
 sg13g2_decap_8 FILLER_3_1539 ();
 sg13g2_decap_8 FILLER_3_1546 ();
 sg13g2_decap_8 FILLER_3_1553 ();
 sg13g2_decap_8 FILLER_3_1560 ();
 sg13g2_decap_8 FILLER_3_1567 ();
 sg13g2_decap_8 FILLER_3_1574 ();
 sg13g2_decap_8 FILLER_3_1581 ();
 sg13g2_decap_8 FILLER_3_1588 ();
 sg13g2_decap_8 FILLER_3_1595 ();
 sg13g2_decap_8 FILLER_3_1602 ();
 sg13g2_decap_8 FILLER_3_1609 ();
 sg13g2_decap_8 FILLER_3_1616 ();
 sg13g2_decap_8 FILLER_3_1623 ();
 sg13g2_decap_8 FILLER_3_1630 ();
 sg13g2_decap_8 FILLER_3_1637 ();
 sg13g2_decap_8 FILLER_3_1644 ();
 sg13g2_decap_8 FILLER_3_1651 ();
 sg13g2_decap_8 FILLER_3_1658 ();
 sg13g2_decap_8 FILLER_3_1665 ();
 sg13g2_decap_8 FILLER_3_1672 ();
 sg13g2_decap_8 FILLER_3_1679 ();
 sg13g2_decap_8 FILLER_3_1686 ();
 sg13g2_decap_8 FILLER_3_1693 ();
 sg13g2_decap_8 FILLER_3_1700 ();
 sg13g2_decap_8 FILLER_3_1707 ();
 sg13g2_decap_8 FILLER_3_1714 ();
 sg13g2_decap_8 FILLER_3_1721 ();
 sg13g2_decap_8 FILLER_3_1728 ();
 sg13g2_decap_8 FILLER_3_1735 ();
 sg13g2_decap_8 FILLER_3_1742 ();
 sg13g2_decap_8 FILLER_3_1749 ();
 sg13g2_decap_8 FILLER_3_1756 ();
 sg13g2_decap_8 FILLER_3_1763 ();
 sg13g2_decap_4 FILLER_3_1770 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_4 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_36 ();
 sg13g2_fill_2 FILLER_4_43 ();
 sg13g2_fill_1 FILLER_4_45 ();
 sg13g2_fill_2 FILLER_4_72 ();
 sg13g2_decap_8 FILLER_4_100 ();
 sg13g2_decap_8 FILLER_4_107 ();
 sg13g2_fill_2 FILLER_4_114 ();
 sg13g2_decap_8 FILLER_4_142 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_decap_4 FILLER_4_214 ();
 sg13g2_fill_1 FILLER_4_249 ();
 sg13g2_decap_8 FILLER_4_276 ();
 sg13g2_fill_2 FILLER_4_283 ();
 sg13g2_fill_2 FILLER_4_290 ();
 sg13g2_fill_1 FILLER_4_292 ();
 sg13g2_decap_8 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_304 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_4 FILLER_4_318 ();
 sg13g2_fill_2 FILLER_4_331 ();
 sg13g2_fill_1 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_fill_2 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_4 FILLER_4_358 ();
 sg13g2_fill_2 FILLER_4_371 ();
 sg13g2_fill_1 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_fill_2 FILLER_4_385 ();
 sg13g2_fill_1 FILLER_4_387 ();
 sg13g2_fill_1 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_402 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_decap_4 FILLER_4_434 ();
 sg13g2_fill_1 FILLER_4_438 ();
 sg13g2_decap_4 FILLER_4_460 ();
 sg13g2_fill_1 FILLER_4_464 ();
 sg13g2_decap_4 FILLER_4_478 ();
 sg13g2_fill_1 FILLER_4_482 ();
 sg13g2_decap_8 FILLER_4_496 ();
 sg13g2_decap_8 FILLER_4_503 ();
 sg13g2_decap_4 FILLER_4_510 ();
 sg13g2_fill_2 FILLER_4_514 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_4 FILLER_4_581 ();
 sg13g2_fill_1 FILLER_4_585 ();
 sg13g2_decap_4 FILLER_4_595 ();
 sg13g2_fill_1 FILLER_4_599 ();
 sg13g2_decap_8 FILLER_4_621 ();
 sg13g2_fill_2 FILLER_4_641 ();
 sg13g2_fill_1 FILLER_4_643 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_4 FILLER_4_676 ();
 sg13g2_fill_2 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_761 ();
 sg13g2_decap_8 FILLER_4_768 ();
 sg13g2_decap_4 FILLER_4_775 ();
 sg13g2_fill_2 FILLER_4_779 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_4 FILLER_4_826 ();
 sg13g2_fill_1 FILLER_4_830 ();
 sg13g2_decap_8 FILLER_4_835 ();
 sg13g2_fill_1 FILLER_4_842 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_decap_8 FILLER_4_875 ();
 sg13g2_decap_4 FILLER_4_882 ();
 sg13g2_fill_1 FILLER_4_886 ();
 sg13g2_decap_8 FILLER_4_891 ();
 sg13g2_fill_1 FILLER_4_898 ();
 sg13g2_decap_8 FILLER_4_920 ();
 sg13g2_fill_1 FILLER_4_927 ();
 sg13g2_decap_4 FILLER_4_933 ();
 sg13g2_fill_2 FILLER_4_937 ();
 sg13g2_decap_4 FILLER_4_943 ();
 sg13g2_fill_1 FILLER_4_947 ();
 sg13g2_decap_8 FILLER_4_969 ();
 sg13g2_fill_1 FILLER_4_976 ();
 sg13g2_decap_8 FILLER_4_981 ();
 sg13g2_fill_2 FILLER_4_988 ();
 sg13g2_decap_4 FILLER_4_994 ();
 sg13g2_fill_1 FILLER_4_998 ();
 sg13g2_fill_1 FILLER_4_1020 ();
 sg13g2_decap_8 FILLER_4_1025 ();
 sg13g2_decap_4 FILLER_4_1032 ();
 sg13g2_fill_1 FILLER_4_1036 ();
 sg13g2_fill_2 FILLER_4_1046 ();
 sg13g2_fill_1 FILLER_4_1048 ();
 sg13g2_fill_2 FILLER_4_1053 ();
 sg13g2_decap_4 FILLER_4_1076 ();
 sg13g2_fill_2 FILLER_4_1085 ();
 sg13g2_decap_8 FILLER_4_1095 ();
 sg13g2_decap_8 FILLER_4_1102 ();
 sg13g2_fill_2 FILLER_4_1109 ();
 sg13g2_decap_4 FILLER_4_1120 ();
 sg13g2_fill_1 FILLER_4_1124 ();
 sg13g2_decap_4 FILLER_4_1151 ();
 sg13g2_fill_1 FILLER_4_1155 ();
 sg13g2_decap_8 FILLER_4_1160 ();
 sg13g2_decap_8 FILLER_4_1167 ();
 sg13g2_decap_8 FILLER_4_1174 ();
 sg13g2_decap_8 FILLER_4_1181 ();
 sg13g2_decap_8 FILLER_4_1188 ();
 sg13g2_decap_8 FILLER_4_1195 ();
 sg13g2_decap_8 FILLER_4_1202 ();
 sg13g2_decap_8 FILLER_4_1209 ();
 sg13g2_decap_8 FILLER_4_1216 ();
 sg13g2_decap_8 FILLER_4_1223 ();
 sg13g2_decap_8 FILLER_4_1230 ();
 sg13g2_decap_8 FILLER_4_1237 ();
 sg13g2_decap_8 FILLER_4_1244 ();
 sg13g2_decap_8 FILLER_4_1251 ();
 sg13g2_decap_8 FILLER_4_1258 ();
 sg13g2_decap_8 FILLER_4_1265 ();
 sg13g2_decap_8 FILLER_4_1272 ();
 sg13g2_decap_8 FILLER_4_1279 ();
 sg13g2_decap_8 FILLER_4_1286 ();
 sg13g2_decap_8 FILLER_4_1293 ();
 sg13g2_decap_8 FILLER_4_1300 ();
 sg13g2_decap_8 FILLER_4_1307 ();
 sg13g2_decap_8 FILLER_4_1314 ();
 sg13g2_decap_8 FILLER_4_1321 ();
 sg13g2_decap_8 FILLER_4_1328 ();
 sg13g2_decap_8 FILLER_4_1335 ();
 sg13g2_decap_8 FILLER_4_1342 ();
 sg13g2_decap_8 FILLER_4_1349 ();
 sg13g2_decap_8 FILLER_4_1356 ();
 sg13g2_decap_8 FILLER_4_1363 ();
 sg13g2_decap_8 FILLER_4_1370 ();
 sg13g2_decap_8 FILLER_4_1377 ();
 sg13g2_decap_8 FILLER_4_1384 ();
 sg13g2_decap_8 FILLER_4_1391 ();
 sg13g2_decap_8 FILLER_4_1398 ();
 sg13g2_decap_8 FILLER_4_1405 ();
 sg13g2_decap_8 FILLER_4_1412 ();
 sg13g2_decap_8 FILLER_4_1419 ();
 sg13g2_decap_8 FILLER_4_1426 ();
 sg13g2_decap_8 FILLER_4_1433 ();
 sg13g2_decap_8 FILLER_4_1440 ();
 sg13g2_decap_8 FILLER_4_1447 ();
 sg13g2_decap_8 FILLER_4_1454 ();
 sg13g2_decap_8 FILLER_4_1461 ();
 sg13g2_decap_8 FILLER_4_1468 ();
 sg13g2_decap_8 FILLER_4_1475 ();
 sg13g2_decap_8 FILLER_4_1482 ();
 sg13g2_decap_8 FILLER_4_1489 ();
 sg13g2_decap_8 FILLER_4_1496 ();
 sg13g2_decap_8 FILLER_4_1503 ();
 sg13g2_decap_8 FILLER_4_1510 ();
 sg13g2_decap_8 FILLER_4_1517 ();
 sg13g2_decap_8 FILLER_4_1524 ();
 sg13g2_decap_8 FILLER_4_1531 ();
 sg13g2_decap_8 FILLER_4_1538 ();
 sg13g2_decap_8 FILLER_4_1545 ();
 sg13g2_decap_8 FILLER_4_1552 ();
 sg13g2_decap_8 FILLER_4_1559 ();
 sg13g2_decap_8 FILLER_4_1566 ();
 sg13g2_decap_8 FILLER_4_1573 ();
 sg13g2_decap_8 FILLER_4_1580 ();
 sg13g2_decap_8 FILLER_4_1587 ();
 sg13g2_decap_8 FILLER_4_1594 ();
 sg13g2_decap_8 FILLER_4_1601 ();
 sg13g2_decap_8 FILLER_4_1608 ();
 sg13g2_decap_8 FILLER_4_1615 ();
 sg13g2_decap_8 FILLER_4_1622 ();
 sg13g2_decap_8 FILLER_4_1629 ();
 sg13g2_decap_8 FILLER_4_1636 ();
 sg13g2_decap_8 FILLER_4_1643 ();
 sg13g2_decap_8 FILLER_4_1650 ();
 sg13g2_decap_8 FILLER_4_1657 ();
 sg13g2_decap_8 FILLER_4_1664 ();
 sg13g2_decap_8 FILLER_4_1671 ();
 sg13g2_decap_8 FILLER_4_1678 ();
 sg13g2_decap_8 FILLER_4_1685 ();
 sg13g2_decap_8 FILLER_4_1692 ();
 sg13g2_decap_8 FILLER_4_1699 ();
 sg13g2_decap_8 FILLER_4_1706 ();
 sg13g2_decap_8 FILLER_4_1713 ();
 sg13g2_decap_8 FILLER_4_1720 ();
 sg13g2_decap_8 FILLER_4_1727 ();
 sg13g2_decap_8 FILLER_4_1734 ();
 sg13g2_decap_8 FILLER_4_1741 ();
 sg13g2_decap_8 FILLER_4_1748 ();
 sg13g2_decap_8 FILLER_4_1755 ();
 sg13g2_decap_8 FILLER_4_1762 ();
 sg13g2_decap_4 FILLER_4_1769 ();
 sg13g2_fill_1 FILLER_4_1773 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_fill_1 FILLER_5_40 ();
 sg13g2_decap_8 FILLER_5_45 ();
 sg13g2_decap_8 FILLER_5_52 ();
 sg13g2_decap_4 FILLER_5_59 ();
 sg13g2_decap_8 FILLER_5_72 ();
 sg13g2_decap_8 FILLER_5_79 ();
 sg13g2_decap_4 FILLER_5_86 ();
 sg13g2_fill_1 FILLER_5_90 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_fill_1 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_129 ();
 sg13g2_fill_1 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_138 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_4 FILLER_5_151 ();
 sg13g2_fill_1 FILLER_5_155 ();
 sg13g2_decap_8 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_202 ();
 sg13g2_fill_1 FILLER_5_235 ();
 sg13g2_fill_1 FILLER_5_244 ();
 sg13g2_fill_1 FILLER_5_272 ();
 sg13g2_decap_4 FILLER_5_278 ();
 sg13g2_fill_1 FILLER_5_282 ();
 sg13g2_fill_2 FILLER_5_287 ();
 sg13g2_fill_2 FILLER_5_323 ();
 sg13g2_decap_4 FILLER_5_351 ();
 sg13g2_fill_1 FILLER_5_359 ();
 sg13g2_fill_2 FILLER_5_386 ();
 sg13g2_fill_2 FILLER_5_414 ();
 sg13g2_fill_2 FILLER_5_420 ();
 sg13g2_decap_4 FILLER_5_431 ();
 sg13g2_fill_2 FILLER_5_435 ();
 sg13g2_decap_4 FILLER_5_462 ();
 sg13g2_fill_1 FILLER_5_500 ();
 sg13g2_decap_8 FILLER_5_505 ();
 sg13g2_decap_8 FILLER_5_516 ();
 sg13g2_fill_1 FILLER_5_523 ();
 sg13g2_decap_8 FILLER_5_528 ();
 sg13g2_decap_4 FILLER_5_535 ();
 sg13g2_decap_4 FILLER_5_543 ();
 sg13g2_decap_8 FILLER_5_551 ();
 sg13g2_decap_4 FILLER_5_558 ();
 sg13g2_fill_1 FILLER_5_562 ();
 sg13g2_fill_1 FILLER_5_568 ();
 sg13g2_fill_1 FILLER_5_599 ();
 sg13g2_decap_4 FILLER_5_621 ();
 sg13g2_fill_1 FILLER_5_716 ();
 sg13g2_fill_1 FILLER_5_733 ();
 sg13g2_decap_8 FILLER_5_755 ();
 sg13g2_decap_8 FILLER_5_762 ();
 sg13g2_decap_8 FILLER_5_769 ();
 sg13g2_decap_8 FILLER_5_776 ();
 sg13g2_fill_1 FILLER_5_783 ();
 sg13g2_fill_1 FILLER_5_824 ();
 sg13g2_decap_8 FILLER_5_856 ();
 sg13g2_decap_8 FILLER_5_867 ();
 sg13g2_decap_8 FILLER_5_874 ();
 sg13g2_fill_1 FILLER_5_881 ();
 sg13g2_fill_1 FILLER_5_892 ();
 sg13g2_fill_1 FILLER_5_897 ();
 sg13g2_fill_1 FILLER_5_903 ();
 sg13g2_fill_2 FILLER_5_925 ();
 sg13g2_fill_1 FILLER_5_927 ();
 sg13g2_decap_8 FILLER_5_958 ();
 sg13g2_decap_8 FILLER_5_965 ();
 sg13g2_decap_4 FILLER_5_972 ();
 sg13g2_fill_2 FILLER_5_976 ();
 sg13g2_fill_1 FILLER_5_982 ();
 sg13g2_fill_1 FILLER_5_988 ();
 sg13g2_fill_2 FILLER_5_993 ();
 sg13g2_decap_8 FILLER_5_1021 ();
 sg13g2_fill_2 FILLER_5_1028 ();
 sg13g2_fill_1 FILLER_5_1030 ();
 sg13g2_decap_8 FILLER_5_1070 ();
 sg13g2_decap_8 FILLER_5_1077 ();
 sg13g2_decap_4 FILLER_5_1084 ();
 sg13g2_fill_2 FILLER_5_1088 ();
 sg13g2_fill_2 FILLER_5_1099 ();
 sg13g2_fill_1 FILLER_5_1101 ();
 sg13g2_decap_8 FILLER_5_1106 ();
 sg13g2_decap_4 FILLER_5_1113 ();
 sg13g2_decap_4 FILLER_5_1143 ();
 sg13g2_fill_2 FILLER_5_1147 ();
 sg13g2_decap_8 FILLER_5_1179 ();
 sg13g2_decap_8 FILLER_5_1186 ();
 sg13g2_decap_8 FILLER_5_1193 ();
 sg13g2_decap_8 FILLER_5_1200 ();
 sg13g2_decap_8 FILLER_5_1207 ();
 sg13g2_decap_8 FILLER_5_1214 ();
 sg13g2_decap_8 FILLER_5_1221 ();
 sg13g2_decap_8 FILLER_5_1228 ();
 sg13g2_decap_8 FILLER_5_1235 ();
 sg13g2_decap_8 FILLER_5_1242 ();
 sg13g2_decap_8 FILLER_5_1249 ();
 sg13g2_decap_8 FILLER_5_1256 ();
 sg13g2_decap_8 FILLER_5_1263 ();
 sg13g2_decap_8 FILLER_5_1270 ();
 sg13g2_decap_8 FILLER_5_1277 ();
 sg13g2_decap_8 FILLER_5_1284 ();
 sg13g2_decap_8 FILLER_5_1291 ();
 sg13g2_decap_8 FILLER_5_1298 ();
 sg13g2_decap_8 FILLER_5_1305 ();
 sg13g2_decap_8 FILLER_5_1312 ();
 sg13g2_decap_8 FILLER_5_1319 ();
 sg13g2_decap_8 FILLER_5_1326 ();
 sg13g2_decap_8 FILLER_5_1333 ();
 sg13g2_decap_8 FILLER_5_1340 ();
 sg13g2_decap_8 FILLER_5_1347 ();
 sg13g2_decap_8 FILLER_5_1354 ();
 sg13g2_decap_8 FILLER_5_1361 ();
 sg13g2_decap_8 FILLER_5_1368 ();
 sg13g2_decap_8 FILLER_5_1375 ();
 sg13g2_decap_8 FILLER_5_1382 ();
 sg13g2_decap_8 FILLER_5_1389 ();
 sg13g2_decap_8 FILLER_5_1396 ();
 sg13g2_decap_8 FILLER_5_1403 ();
 sg13g2_decap_8 FILLER_5_1410 ();
 sg13g2_decap_8 FILLER_5_1417 ();
 sg13g2_decap_8 FILLER_5_1424 ();
 sg13g2_decap_8 FILLER_5_1431 ();
 sg13g2_decap_8 FILLER_5_1438 ();
 sg13g2_decap_8 FILLER_5_1445 ();
 sg13g2_decap_8 FILLER_5_1452 ();
 sg13g2_decap_8 FILLER_5_1459 ();
 sg13g2_decap_8 FILLER_5_1466 ();
 sg13g2_decap_8 FILLER_5_1473 ();
 sg13g2_decap_8 FILLER_5_1480 ();
 sg13g2_decap_8 FILLER_5_1487 ();
 sg13g2_decap_4 FILLER_5_1494 ();
 sg13g2_decap_8 FILLER_5_1502 ();
 sg13g2_decap_8 FILLER_5_1509 ();
 sg13g2_decap_8 FILLER_5_1516 ();
 sg13g2_decap_8 FILLER_5_1523 ();
 sg13g2_decap_8 FILLER_5_1530 ();
 sg13g2_decap_8 FILLER_5_1537 ();
 sg13g2_decap_8 FILLER_5_1544 ();
 sg13g2_decap_8 FILLER_5_1551 ();
 sg13g2_decap_8 FILLER_5_1558 ();
 sg13g2_decap_8 FILLER_5_1565 ();
 sg13g2_decap_8 FILLER_5_1572 ();
 sg13g2_decap_8 FILLER_5_1579 ();
 sg13g2_decap_8 FILLER_5_1586 ();
 sg13g2_decap_4 FILLER_5_1593 ();
 sg13g2_decap_4 FILLER_5_1634 ();
 sg13g2_fill_2 FILLER_5_1638 ();
 sg13g2_decap_8 FILLER_5_1644 ();
 sg13g2_decap_8 FILLER_5_1651 ();
 sg13g2_decap_8 FILLER_5_1658 ();
 sg13g2_fill_2 FILLER_5_1665 ();
 sg13g2_decap_8 FILLER_5_1693 ();
 sg13g2_decap_8 FILLER_5_1700 ();
 sg13g2_decap_8 FILLER_5_1707 ();
 sg13g2_decap_8 FILLER_5_1714 ();
 sg13g2_decap_8 FILLER_5_1721 ();
 sg13g2_decap_8 FILLER_5_1728 ();
 sg13g2_decap_8 FILLER_5_1735 ();
 sg13g2_decap_8 FILLER_5_1742 ();
 sg13g2_decap_8 FILLER_5_1749 ();
 sg13g2_decap_8 FILLER_5_1756 ();
 sg13g2_decap_8 FILLER_5_1763 ();
 sg13g2_decap_4 FILLER_5_1770 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_18 ();
 sg13g2_fill_1 FILLER_6_45 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_decap_8 FILLER_6_79 ();
 sg13g2_decap_4 FILLER_6_86 ();
 sg13g2_fill_1 FILLER_6_90 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_4 FILLER_6_119 ();
 sg13g2_fill_1 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_155 ();
 sg13g2_fill_2 FILLER_6_162 ();
 sg13g2_fill_1 FILLER_6_164 ();
 sg13g2_decap_8 FILLER_6_169 ();
 sg13g2_decap_8 FILLER_6_176 ();
 sg13g2_fill_1 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_219 ();
 sg13g2_fill_2 FILLER_6_237 ();
 sg13g2_fill_2 FILLER_6_309 ();
 sg13g2_fill_1 FILLER_6_315 ();
 sg13g2_decap_4 FILLER_6_337 ();
 sg13g2_fill_1 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_fill_1 FILLER_6_360 ();
 sg13g2_fill_1 FILLER_6_370 ();
 sg13g2_fill_2 FILLER_6_376 ();
 sg13g2_fill_1 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_409 ();
 sg13g2_decap_8 FILLER_6_416 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_fill_2 FILLER_6_430 ();
 sg13g2_fill_1 FILLER_6_432 ();
 sg13g2_fill_2 FILLER_6_438 ();
 sg13g2_fill_1 FILLER_6_440 ();
 sg13g2_decap_8 FILLER_6_454 ();
 sg13g2_fill_2 FILLER_6_461 ();
 sg13g2_fill_1 FILLER_6_463 ();
 sg13g2_decap_4 FILLER_6_473 ();
 sg13g2_fill_2 FILLER_6_477 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_4 FILLER_6_490 ();
 sg13g2_fill_2 FILLER_6_525 ();
 sg13g2_decap_4 FILLER_6_531 ();
 sg13g2_decap_8 FILLER_6_570 ();
 sg13g2_decap_4 FILLER_6_577 ();
 sg13g2_fill_2 FILLER_6_585 ();
 sg13g2_fill_1 FILLER_6_587 ();
 sg13g2_fill_2 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_615 ();
 sg13g2_decap_8 FILLER_6_622 ();
 sg13g2_fill_2 FILLER_6_629 ();
 sg13g2_fill_1 FILLER_6_631 ();
 sg13g2_fill_1 FILLER_6_642 ();
 sg13g2_decap_8 FILLER_6_647 ();
 sg13g2_decap_8 FILLER_6_654 ();
 sg13g2_decap_8 FILLER_6_661 ();
 sg13g2_fill_2 FILLER_6_694 ();
 sg13g2_fill_1 FILLER_6_700 ();
 sg13g2_fill_1 FILLER_6_705 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_4 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_755 ();
 sg13g2_decap_8 FILLER_6_762 ();
 sg13g2_fill_1 FILLER_6_769 ();
 sg13g2_fill_1 FILLER_6_780 ();
 sg13g2_decap_8 FILLER_6_811 ();
 sg13g2_decap_4 FILLER_6_839 ();
 sg13g2_fill_2 FILLER_6_882 ();
 sg13g2_fill_1 FILLER_6_884 ();
 sg13g2_decap_4 FILLER_6_933 ();
 sg13g2_decap_4 FILLER_6_942 ();
 sg13g2_decap_8 FILLER_6_950 ();
 sg13g2_decap_4 FILLER_6_957 ();
 sg13g2_fill_1 FILLER_6_961 ();
 sg13g2_decap_4 FILLER_6_997 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_fill_1 FILLER_6_1012 ();
 sg13g2_decap_4 FILLER_6_1018 ();
 sg13g2_fill_1 FILLER_6_1022 ();
 sg13g2_decap_8 FILLER_6_1049 ();
 sg13g2_decap_4 FILLER_6_1056 ();
 sg13g2_decap_8 FILLER_6_1065 ();
 sg13g2_decap_8 FILLER_6_1076 ();
 sg13g2_decap_8 FILLER_6_1083 ();
 sg13g2_fill_1 FILLER_6_1090 ();
 sg13g2_decap_8 FILLER_6_1138 ();
 sg13g2_decap_8 FILLER_6_1145 ();
 sg13g2_fill_2 FILLER_6_1152 ();
 sg13g2_decap_8 FILLER_6_1190 ();
 sg13g2_decap_4 FILLER_6_1197 ();
 sg13g2_fill_2 FILLER_6_1201 ();
 sg13g2_fill_2 FILLER_6_1213 ();
 sg13g2_fill_1 FILLER_6_1215 ();
 sg13g2_decap_8 FILLER_6_1220 ();
 sg13g2_decap_8 FILLER_6_1227 ();
 sg13g2_decap_8 FILLER_6_1234 ();
 sg13g2_decap_8 FILLER_6_1241 ();
 sg13g2_decap_8 FILLER_6_1248 ();
 sg13g2_decap_8 FILLER_6_1255 ();
 sg13g2_decap_8 FILLER_6_1262 ();
 sg13g2_decap_8 FILLER_6_1269 ();
 sg13g2_decap_8 FILLER_6_1276 ();
 sg13g2_decap_8 FILLER_6_1283 ();
 sg13g2_decap_8 FILLER_6_1290 ();
 sg13g2_decap_8 FILLER_6_1297 ();
 sg13g2_decap_8 FILLER_6_1304 ();
 sg13g2_decap_8 FILLER_6_1311 ();
 sg13g2_decap_8 FILLER_6_1318 ();
 sg13g2_decap_8 FILLER_6_1325 ();
 sg13g2_decap_8 FILLER_6_1332 ();
 sg13g2_decap_8 FILLER_6_1339 ();
 sg13g2_decap_8 FILLER_6_1346 ();
 sg13g2_decap_8 FILLER_6_1353 ();
 sg13g2_decap_8 FILLER_6_1360 ();
 sg13g2_decap_8 FILLER_6_1367 ();
 sg13g2_decap_8 FILLER_6_1374 ();
 sg13g2_decap_8 FILLER_6_1381 ();
 sg13g2_decap_8 FILLER_6_1388 ();
 sg13g2_decap_8 FILLER_6_1395 ();
 sg13g2_decap_8 FILLER_6_1402 ();
 sg13g2_decap_8 FILLER_6_1409 ();
 sg13g2_decap_8 FILLER_6_1416 ();
 sg13g2_decap_8 FILLER_6_1423 ();
 sg13g2_decap_8 FILLER_6_1430 ();
 sg13g2_decap_8 FILLER_6_1437 ();
 sg13g2_decap_8 FILLER_6_1444 ();
 sg13g2_decap_8 FILLER_6_1451 ();
 sg13g2_decap_8 FILLER_6_1458 ();
 sg13g2_decap_8 FILLER_6_1465 ();
 sg13g2_decap_8 FILLER_6_1472 ();
 sg13g2_decap_8 FILLER_6_1479 ();
 sg13g2_decap_4 FILLER_6_1486 ();
 sg13g2_fill_2 FILLER_6_1490 ();
 sg13g2_decap_4 FILLER_6_1528 ();
 sg13g2_decap_8 FILLER_6_1536 ();
 sg13g2_decap_8 FILLER_6_1543 ();
 sg13g2_decap_4 FILLER_6_1550 ();
 sg13g2_fill_2 FILLER_6_1554 ();
 sg13g2_decap_4 FILLER_6_1560 ();
 sg13g2_decap_4 FILLER_6_1574 ();
 sg13g2_fill_1 FILLER_6_1604 ();
 sg13g2_fill_1 FILLER_6_1631 ();
 sg13g2_fill_1 FILLER_6_1658 ();
 sg13g2_fill_1 FILLER_6_1669 ();
 sg13g2_fill_1 FILLER_6_1674 ();
 sg13g2_decap_8 FILLER_6_1679 ();
 sg13g2_fill_1 FILLER_6_1686 ();
 sg13g2_decap_4 FILLER_6_1708 ();
 sg13g2_decap_8 FILLER_6_1716 ();
 sg13g2_decap_8 FILLER_6_1723 ();
 sg13g2_decap_8 FILLER_6_1730 ();
 sg13g2_decap_8 FILLER_6_1737 ();
 sg13g2_decap_8 FILLER_6_1744 ();
 sg13g2_decap_8 FILLER_6_1751 ();
 sg13g2_decap_8 FILLER_6_1758 ();
 sg13g2_decap_8 FILLER_6_1765 ();
 sg13g2_fill_2 FILLER_6_1772 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_16 ();
 sg13g2_decap_4 FILLER_7_21 ();
 sg13g2_fill_2 FILLER_7_25 ();
 sg13g2_decap_4 FILLER_7_31 ();
 sg13g2_decap_8 FILLER_7_61 ();
 sg13g2_fill_1 FILLER_7_68 ();
 sg13g2_fill_1 FILLER_7_104 ();
 sg13g2_decap_8 FILLER_7_136 ();
 sg13g2_decap_4 FILLER_7_143 ();
 sg13g2_fill_2 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_209 ();
 sg13g2_fill_2 FILLER_7_240 ();
 sg13g2_fill_2 FILLER_7_263 ();
 sg13g2_fill_2 FILLER_7_269 ();
 sg13g2_fill_1 FILLER_7_271 ();
 sg13g2_fill_2 FILLER_7_277 ();
 sg13g2_fill_1 FILLER_7_279 ();
 sg13g2_decap_4 FILLER_7_285 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_4 FILLER_7_305 ();
 sg13g2_fill_1 FILLER_7_309 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_4 FILLER_7_343 ();
 sg13g2_fill_2 FILLER_7_347 ();
 sg13g2_fill_2 FILLER_7_375 ();
 sg13g2_fill_1 FILLER_7_377 ();
 sg13g2_fill_1 FILLER_7_399 ();
 sg13g2_fill_1 FILLER_7_430 ();
 sg13g2_fill_1 FILLER_7_435 ();
 sg13g2_fill_2 FILLER_7_462 ();
 sg13g2_fill_2 FILLER_7_503 ();
 sg13g2_decap_8 FILLER_7_552 ();
 sg13g2_decap_4 FILLER_7_559 ();
 sg13g2_fill_1 FILLER_7_563 ();
 sg13g2_decap_8 FILLER_7_576 ();
 sg13g2_decap_4 FILLER_7_583 ();
 sg13g2_fill_2 FILLER_7_587 ();
 sg13g2_fill_2 FILLER_7_624 ();
 sg13g2_fill_1 FILLER_7_693 ();
 sg13g2_decap_4 FILLER_7_712 ();
 sg13g2_fill_1 FILLER_7_729 ();
 sg13g2_decap_4 FILLER_7_739 ();
 sg13g2_fill_1 FILLER_7_748 ();
 sg13g2_decap_4 FILLER_7_753 ();
 sg13g2_fill_2 FILLER_7_767 ();
 sg13g2_fill_1 FILLER_7_769 ();
 sg13g2_fill_2 FILLER_7_779 ();
 sg13g2_fill_1 FILLER_7_781 ();
 sg13g2_decap_4 FILLER_7_843 ();
 sg13g2_fill_1 FILLER_7_847 ();
 sg13g2_fill_1 FILLER_7_853 ();
 sg13g2_fill_1 FILLER_7_858 ();
 sg13g2_decap_8 FILLER_7_863 ();
 sg13g2_fill_2 FILLER_7_870 ();
 sg13g2_fill_1 FILLER_7_872 ();
 sg13g2_decap_8 FILLER_7_877 ();
 sg13g2_fill_1 FILLER_7_884 ();
 sg13g2_decap_4 FILLER_7_898 ();
 sg13g2_fill_1 FILLER_7_902 ();
 sg13g2_decap_4 FILLER_7_907 ();
 sg13g2_fill_2 FILLER_7_911 ();
 sg13g2_fill_2 FILLER_7_939 ();
 sg13g2_decap_8 FILLER_7_967 ();
 sg13g2_decap_8 FILLER_7_974 ();
 sg13g2_fill_1 FILLER_7_981 ();
 sg13g2_decap_8 FILLER_7_1007 ();
 sg13g2_fill_2 FILLER_7_1014 ();
 sg13g2_fill_1 FILLER_7_1021 ();
 sg13g2_fill_2 FILLER_7_1026 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_decap_8 FILLER_7_1033 ();
 sg13g2_decap_4 FILLER_7_1040 ();
 sg13g2_fill_1 FILLER_7_1044 ();
 sg13g2_fill_1 FILLER_7_1054 ();
 sg13g2_fill_2 FILLER_7_1059 ();
 sg13g2_fill_1 FILLER_7_1065 ();
 sg13g2_fill_2 FILLER_7_1092 ();
 sg13g2_decap_8 FILLER_7_1129 ();
 sg13g2_decap_4 FILLER_7_1136 ();
 sg13g2_decap_8 FILLER_7_1150 ();
 sg13g2_decap_8 FILLER_7_1157 ();
 sg13g2_decap_8 FILLER_7_1164 ();
 sg13g2_decap_8 FILLER_7_1171 ();
 sg13g2_decap_4 FILLER_7_1178 ();
 sg13g2_decap_8 FILLER_7_1203 ();
 sg13g2_decap_8 FILLER_7_1262 ();
 sg13g2_decap_8 FILLER_7_1269 ();
 sg13g2_decap_8 FILLER_7_1276 ();
 sg13g2_decap_8 FILLER_7_1283 ();
 sg13g2_decap_8 FILLER_7_1290 ();
 sg13g2_decap_8 FILLER_7_1297 ();
 sg13g2_decap_8 FILLER_7_1304 ();
 sg13g2_decap_8 FILLER_7_1311 ();
 sg13g2_decap_8 FILLER_7_1318 ();
 sg13g2_fill_2 FILLER_7_1325 ();
 sg13g2_fill_1 FILLER_7_1327 ();
 sg13g2_decap_8 FILLER_7_1338 ();
 sg13g2_decap_8 FILLER_7_1345 ();
 sg13g2_decap_8 FILLER_7_1352 ();
 sg13g2_decap_8 FILLER_7_1359 ();
 sg13g2_fill_2 FILLER_7_1366 ();
 sg13g2_fill_1 FILLER_7_1368 ();
 sg13g2_decap_8 FILLER_7_1399 ();
 sg13g2_decap_8 FILLER_7_1406 ();
 sg13g2_decap_8 FILLER_7_1417 ();
 sg13g2_decap_8 FILLER_7_1424 ();
 sg13g2_decap_8 FILLER_7_1431 ();
 sg13g2_decap_8 FILLER_7_1438 ();
 sg13g2_decap_8 FILLER_7_1445 ();
 sg13g2_decap_8 FILLER_7_1452 ();
 sg13g2_decap_8 FILLER_7_1459 ();
 sg13g2_decap_8 FILLER_7_1466 ();
 sg13g2_decap_8 FILLER_7_1473 ();
 sg13g2_decap_8 FILLER_7_1480 ();
 sg13g2_decap_8 FILLER_7_1487 ();
 sg13g2_decap_8 FILLER_7_1494 ();
 sg13g2_fill_2 FILLER_7_1521 ();
 sg13g2_fill_2 FILLER_7_1575 ();
 sg13g2_decap_8 FILLER_7_1610 ();
 sg13g2_decap_4 FILLER_7_1617 ();
 sg13g2_fill_1 FILLER_7_1621 ();
 sg13g2_decap_8 FILLER_7_1643 ();
 sg13g2_fill_2 FILLER_7_1650 ();
 sg13g2_fill_1 FILLER_7_1652 ();
 sg13g2_decap_4 FILLER_7_1689 ();
 sg13g2_fill_2 FILLER_7_1693 ();
 sg13g2_decap_4 FILLER_7_1731 ();
 sg13g2_fill_2 FILLER_7_1735 ();
 sg13g2_decap_8 FILLER_7_1741 ();
 sg13g2_decap_8 FILLER_7_1748 ();
 sg13g2_decap_8 FILLER_7_1755 ();
 sg13g2_decap_8 FILLER_7_1762 ();
 sg13g2_decap_4 FILLER_7_1769 ();
 sg13g2_fill_1 FILLER_7_1773 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_37 ();
 sg13g2_fill_1 FILLER_8_83 ();
 sg13g2_fill_1 FILLER_8_88 ();
 sg13g2_fill_2 FILLER_8_110 ();
 sg13g2_fill_2 FILLER_8_116 ();
 sg13g2_fill_2 FILLER_8_122 ();
 sg13g2_decap_8 FILLER_8_145 ();
 sg13g2_decap_8 FILLER_8_152 ();
 sg13g2_fill_2 FILLER_8_159 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_fill_2 FILLER_8_179 ();
 sg13g2_fill_1 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_fill_2 FILLER_8_238 ();
 sg13g2_fill_1 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_272 ();
 sg13g2_fill_2 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_307 ();
 sg13g2_fill_1 FILLER_8_309 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_fill_2 FILLER_8_321 ();
 sg13g2_fill_1 FILLER_8_323 ();
 sg13g2_fill_2 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_4 FILLER_8_367 ();
 sg13g2_fill_1 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_8_421 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_8_461 ();
 sg13g2_decap_8 FILLER_8_468 ();
 sg13g2_decap_4 FILLER_8_475 ();
 sg13g2_fill_2 FILLER_8_489 ();
 sg13g2_decap_4 FILLER_8_505 ();
 sg13g2_fill_1 FILLER_8_509 ();
 sg13g2_decap_8 FILLER_8_514 ();
 sg13g2_fill_1 FILLER_8_521 ();
 sg13g2_fill_2 FILLER_8_573 ();
 sg13g2_fill_1 FILLER_8_575 ();
 sg13g2_decap_8 FILLER_8_580 ();
 sg13g2_fill_1 FILLER_8_587 ();
 sg13g2_fill_1 FILLER_8_596 ();
 sg13g2_fill_1 FILLER_8_601 ();
 sg13g2_decap_4 FILLER_8_612 ();
 sg13g2_fill_1 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_631 ();
 sg13g2_decap_8 FILLER_8_638 ();
 sg13g2_decap_8 FILLER_8_645 ();
 sg13g2_decap_8 FILLER_8_652 ();
 sg13g2_decap_4 FILLER_8_659 ();
 sg13g2_decap_4 FILLER_8_677 ();
 sg13g2_fill_2 FILLER_8_686 ();
 sg13g2_fill_1 FILLER_8_688 ();
 sg13g2_fill_1 FILLER_8_698 ();
 sg13g2_fill_1 FILLER_8_725 ();
 sg13g2_decap_8 FILLER_8_752 ();
 sg13g2_decap_8 FILLER_8_795 ();
 sg13g2_decap_4 FILLER_8_802 ();
 sg13g2_fill_2 FILLER_8_810 ();
 sg13g2_fill_1 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_821 ();
 sg13g2_fill_1 FILLER_8_828 ();
 sg13g2_decap_8 FILLER_8_834 ();
 sg13g2_decap_4 FILLER_8_841 ();
 sg13g2_fill_2 FILLER_8_876 ();
 sg13g2_fill_1 FILLER_8_878 ();
 sg13g2_decap_8 FILLER_8_909 ();
 sg13g2_decap_4 FILLER_8_916 ();
 sg13g2_decap_4 FILLER_8_924 ();
 sg13g2_fill_1 FILLER_8_928 ();
 sg13g2_fill_1 FILLER_8_933 ();
 sg13g2_decap_8 FILLER_8_938 ();
 sg13g2_fill_2 FILLER_8_945 ();
 sg13g2_fill_1 FILLER_8_947 ();
 sg13g2_decap_4 FILLER_8_952 ();
 sg13g2_fill_1 FILLER_8_987 ();
 sg13g2_fill_2 FILLER_8_1009 ();
 sg13g2_fill_1 FILLER_8_1015 ();
 sg13g2_fill_2 FILLER_8_1042 ();
 sg13g2_decap_8 FILLER_8_1070 ();
 sg13g2_fill_2 FILLER_8_1077 ();
 sg13g2_fill_1 FILLER_8_1079 ();
 sg13g2_decap_4 FILLER_8_1106 ();
 sg13g2_decap_8 FILLER_8_1139 ();
 sg13g2_fill_1 FILLER_8_1146 ();
 sg13g2_decap_8 FILLER_8_1173 ();
 sg13g2_fill_2 FILLER_8_1180 ();
 sg13g2_decap_8 FILLER_8_1203 ();
 sg13g2_fill_1 FILLER_8_1210 ();
 sg13g2_decap_4 FILLER_8_1215 ();
 sg13g2_fill_1 FILLER_8_1219 ();
 sg13g2_decap_8 FILLER_8_1230 ();
 sg13g2_decap_8 FILLER_8_1237 ();
 sg13g2_fill_1 FILLER_8_1244 ();
 sg13g2_decap_8 FILLER_8_1249 ();
 sg13g2_decap_8 FILLER_8_1256 ();
 sg13g2_fill_2 FILLER_8_1263 ();
 sg13g2_decap_8 FILLER_8_1278 ();
 sg13g2_decap_8 FILLER_8_1285 ();
 sg13g2_decap_8 FILLER_8_1292 ();
 sg13g2_decap_8 FILLER_8_1299 ();
 sg13g2_fill_2 FILLER_8_1336 ();
 sg13g2_fill_1 FILLER_8_1338 ();
 sg13g2_decap_8 FILLER_8_1365 ();
 sg13g2_decap_4 FILLER_8_1372 ();
 sg13g2_fill_1 FILLER_8_1376 ();
 sg13g2_decap_8 FILLER_8_1387 ();
 sg13g2_fill_2 FILLER_8_1394 ();
 sg13g2_fill_2 FILLER_8_1442 ();
 sg13g2_fill_1 FILLER_8_1444 ();
 sg13g2_decap_8 FILLER_8_1449 ();
 sg13g2_decap_4 FILLER_8_1456 ();
 sg13g2_fill_2 FILLER_8_1460 ();
 sg13g2_fill_2 FILLER_8_1472 ();
 sg13g2_decap_8 FILLER_8_1478 ();
 sg13g2_decap_4 FILLER_8_1485 ();
 sg13g2_fill_2 FILLER_8_1489 ();
 sg13g2_decap_8 FILLER_8_1538 ();
 sg13g2_decap_4 FILLER_8_1545 ();
 sg13g2_fill_2 FILLER_8_1549 ();
 sg13g2_decap_8 FILLER_8_1561 ();
 sg13g2_fill_2 FILLER_8_1568 ();
 sg13g2_fill_1 FILLER_8_1570 ();
 sg13g2_decap_4 FILLER_8_1596 ();
 sg13g2_fill_1 FILLER_8_1600 ();
 sg13g2_decap_4 FILLER_8_1627 ();
 sg13g2_fill_2 FILLER_8_1631 ();
 sg13g2_decap_8 FILLER_8_1659 ();
 sg13g2_decap_8 FILLER_8_1666 ();
 sg13g2_fill_1 FILLER_8_1673 ();
 sg13g2_decap_4 FILLER_8_1678 ();
 sg13g2_fill_1 FILLER_8_1682 ();
 sg13g2_decap_8 FILLER_8_1696 ();
 sg13g2_decap_8 FILLER_8_1703 ();
 sg13g2_decap_8 FILLER_8_1710 ();
 sg13g2_fill_2 FILLER_8_1717 ();
 sg13g2_fill_1 FILLER_8_1719 ();
 sg13g2_decap_8 FILLER_8_1756 ();
 sg13g2_decap_8 FILLER_8_1763 ();
 sg13g2_decap_4 FILLER_8_1770 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_fill_1 FILLER_9_33 ();
 sg13g2_fill_2 FILLER_9_43 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_79 ();
 sg13g2_fill_2 FILLER_9_86 ();
 sg13g2_fill_1 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_110 ();
 sg13g2_decap_8 FILLER_9_117 ();
 sg13g2_decap_4 FILLER_9_124 ();
 sg13g2_fill_2 FILLER_9_184 ();
 sg13g2_fill_1 FILLER_9_186 ();
 sg13g2_decap_4 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_229 ();
 sg13g2_fill_2 FILLER_9_234 ();
 sg13g2_decap_4 FILLER_9_240 ();
 sg13g2_fill_2 FILLER_9_244 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_fill_2 FILLER_9_287 ();
 sg13g2_fill_2 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_fill_2 FILLER_9_364 ();
 sg13g2_decap_4 FILLER_9_428 ();
 sg13g2_fill_1 FILLER_9_432 ();
 sg13g2_fill_1 FILLER_9_446 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_4 FILLER_9_466 ();
 sg13g2_fill_1 FILLER_9_470 ();
 sg13g2_fill_1 FILLER_9_497 ();
 sg13g2_fill_2 FILLER_9_524 ();
 sg13g2_fill_1 FILLER_9_526 ();
 sg13g2_fill_1 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_537 ();
 sg13g2_decap_8 FILLER_9_544 ();
 sg13g2_decap_8 FILLER_9_551 ();
 sg13g2_fill_2 FILLER_9_563 ();
 sg13g2_fill_1 FILLER_9_565 ();
 sg13g2_fill_1 FILLER_9_579 ();
 sg13g2_decap_8 FILLER_9_606 ();
 sg13g2_fill_2 FILLER_9_617 ();
 sg13g2_fill_1 FILLER_9_619 ();
 sg13g2_decap_4 FILLER_9_624 ();
 sg13g2_fill_1 FILLER_9_628 ();
 sg13g2_fill_1 FILLER_9_650 ();
 sg13g2_fill_2 FILLER_9_656 ();
 sg13g2_fill_1 FILLER_9_684 ();
 sg13g2_fill_2 FILLER_9_689 ();
 sg13g2_decap_8 FILLER_9_695 ();
 sg13g2_fill_2 FILLER_9_702 ();
 sg13g2_decap_4 FILLER_9_712 ();
 sg13g2_fill_2 FILLER_9_716 ();
 sg13g2_decap_8 FILLER_9_739 ();
 sg13g2_decap_8 FILLER_9_746 ();
 sg13g2_fill_1 FILLER_9_753 ();
 sg13g2_decap_8 FILLER_9_758 ();
 sg13g2_decap_4 FILLER_9_765 ();
 sg13g2_decap_4 FILLER_9_786 ();
 sg13g2_fill_2 FILLER_9_790 ();
 sg13g2_fill_2 FILLER_9_802 ();
 sg13g2_fill_1 FILLER_9_804 ();
 sg13g2_decap_8 FILLER_9_831 ();
 sg13g2_decap_8 FILLER_9_842 ();
 sg13g2_decap_8 FILLER_9_849 ();
 sg13g2_fill_2 FILLER_9_865 ();
 sg13g2_fill_1 FILLER_9_867 ();
 sg13g2_fill_1 FILLER_9_872 ();
 sg13g2_decap_4 FILLER_9_877 ();
 sg13g2_fill_2 FILLER_9_881 ();
 sg13g2_fill_2 FILLER_9_919 ();
 sg13g2_fill_1 FILLER_9_921 ();
 sg13g2_fill_2 FILLER_9_958 ();
 sg13g2_fill_1 FILLER_9_964 ();
 sg13g2_fill_2 FILLER_9_969 ();
 sg13g2_fill_1 FILLER_9_971 ();
 sg13g2_fill_2 FILLER_9_976 ();
 sg13g2_fill_1 FILLER_9_978 ();
 sg13g2_decap_4 FILLER_9_988 ();
 sg13g2_decap_8 FILLER_9_1005 ();
 sg13g2_decap_8 FILLER_9_1012 ();
 sg13g2_decap_8 FILLER_9_1019 ();
 sg13g2_decap_8 FILLER_9_1026 ();
 sg13g2_decap_8 FILLER_9_1037 ();
 sg13g2_decap_8 FILLER_9_1044 ();
 sg13g2_fill_1 FILLER_9_1051 ();
 sg13g2_fill_2 FILLER_9_1083 ();
 sg13g2_fill_1 FILLER_9_1085 ();
 sg13g2_decap_8 FILLER_9_1099 ();
 sg13g2_decap_4 FILLER_9_1106 ();
 sg13g2_decap_4 FILLER_9_1119 ();
 sg13g2_fill_1 FILLER_9_1123 ();
 sg13g2_decap_4 FILLER_9_1150 ();
 sg13g2_decap_8 FILLER_9_1168 ();
 sg13g2_decap_8 FILLER_9_1175 ();
 sg13g2_fill_2 FILLER_9_1203 ();
 sg13g2_fill_2 FILLER_9_1215 ();
 sg13g2_fill_1 FILLER_9_1227 ();
 sg13g2_decap_8 FILLER_9_1254 ();
 sg13g2_decap_4 FILLER_9_1261 ();
 sg13g2_decap_8 FILLER_9_1278 ();
 sg13g2_decap_8 FILLER_9_1285 ();
 sg13g2_decap_8 FILLER_9_1292 ();
 sg13g2_decap_8 FILLER_9_1299 ();
 sg13g2_decap_8 FILLER_9_1306 ();
 sg13g2_decap_8 FILLER_9_1313 ();
 sg13g2_decap_8 FILLER_9_1320 ();
 sg13g2_fill_1 FILLER_9_1327 ();
 sg13g2_fill_2 FILLER_9_1336 ();
 sg13g2_fill_2 FILLER_9_1348 ();
 sg13g2_fill_1 FILLER_9_1350 ();
 sg13g2_decap_4 FILLER_9_1355 ();
 sg13g2_fill_2 FILLER_9_1359 ();
 sg13g2_decap_4 FILLER_9_1397 ();
 sg13g2_fill_1 FILLER_9_1401 ();
 sg13g2_fill_2 FILLER_9_1412 ();
 sg13g2_fill_1 FILLER_9_1414 ();
 sg13g2_decap_4 FILLER_9_1419 ();
 sg13g2_fill_2 FILLER_9_1436 ();
 sg13g2_fill_2 FILLER_9_1464 ();
 sg13g2_fill_1 FILLER_9_1466 ();
 sg13g2_decap_8 FILLER_9_1493 ();
 sg13g2_decap_8 FILLER_9_1504 ();
 sg13g2_decap_4 FILLER_9_1511 ();
 sg13g2_fill_1 FILLER_9_1551 ();
 sg13g2_decap_8 FILLER_9_1578 ();
 sg13g2_decap_4 FILLER_9_1585 ();
 sg13g2_fill_1 FILLER_9_1589 ();
 sg13g2_decap_8 FILLER_9_1594 ();
 sg13g2_decap_8 FILLER_9_1601 ();
 sg13g2_decap_8 FILLER_9_1612 ();
 sg13g2_decap_8 FILLER_9_1619 ();
 sg13g2_decap_4 FILLER_9_1636 ();
 sg13g2_decap_8 FILLER_9_1644 ();
 sg13g2_decap_4 FILLER_9_1651 ();
 sg13g2_fill_2 FILLER_9_1655 ();
 sg13g2_decap_4 FILLER_9_1693 ();
 sg13g2_fill_2 FILLER_9_1697 ();
 sg13g2_decap_4 FILLER_9_1709 ();
 sg13g2_fill_2 FILLER_9_1713 ();
 sg13g2_decap_4 FILLER_9_1719 ();
 sg13g2_decap_8 FILLER_9_1759 ();
 sg13g2_decap_8 FILLER_9_1766 ();
 sg13g2_fill_1 FILLER_9_1773 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_27 ();
 sg13g2_fill_2 FILLER_10_33 ();
 sg13g2_fill_2 FILLER_10_61 ();
 sg13g2_decap_4 FILLER_10_67 ();
 sg13g2_fill_2 FILLER_10_71 ();
 sg13g2_decap_8 FILLER_10_78 ();
 sg13g2_fill_2 FILLER_10_85 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_4 FILLER_10_105 ();
 sg13g2_fill_1 FILLER_10_109 ();
 sg13g2_fill_2 FILLER_10_145 ();
 sg13g2_decap_4 FILLER_10_169 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_281 ();
 sg13g2_decap_4 FILLER_10_292 ();
 sg13g2_decap_4 FILLER_10_300 ();
 sg13g2_fill_2 FILLER_10_304 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_fill_2 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_fill_2 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_411 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_decap_8 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_10_436 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_4 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_488 ();
 sg13g2_decap_4 FILLER_10_495 ();
 sg13g2_fill_1 FILLER_10_499 ();
 sg13g2_decap_4 FILLER_10_505 ();
 sg13g2_fill_1 FILLER_10_509 ();
 sg13g2_decap_4 FILLER_10_514 ();
 sg13g2_fill_2 FILLER_10_522 ();
 sg13g2_fill_1 FILLER_10_524 ();
 sg13g2_decap_8 FILLER_10_586 ();
 sg13g2_fill_2 FILLER_10_597 ();
 sg13g2_fill_1 FILLER_10_599 ();
 sg13g2_decap_8 FILLER_10_657 ();
 sg13g2_fill_1 FILLER_10_721 ();
 sg13g2_fill_1 FILLER_10_748 ();
 sg13g2_fill_2 FILLER_10_757 ();
 sg13g2_fill_1 FILLER_10_759 ();
 sg13g2_decap_4 FILLER_10_764 ();
 sg13g2_decap_8 FILLER_10_794 ();
 sg13g2_decap_8 FILLER_10_801 ();
 sg13g2_fill_2 FILLER_10_808 ();
 sg13g2_fill_1 FILLER_10_810 ();
 sg13g2_fill_1 FILLER_10_847 ();
 sg13g2_fill_2 FILLER_10_874 ();
 sg13g2_fill_1 FILLER_10_881 ();
 sg13g2_fill_2 FILLER_10_887 ();
 sg13g2_decap_8 FILLER_10_897 ();
 sg13g2_decap_8 FILLER_10_904 ();
 sg13g2_decap_4 FILLER_10_911 ();
 sg13g2_fill_1 FILLER_10_915 ();
 sg13g2_decap_8 FILLER_10_942 ();
 sg13g2_decap_4 FILLER_10_949 ();
 sg13g2_fill_2 FILLER_10_953 ();
 sg13g2_decap_8 FILLER_10_1011 ();
 sg13g2_fill_2 FILLER_10_1022 ();
 sg13g2_fill_1 FILLER_10_1024 ();
 sg13g2_decap_8 FILLER_10_1029 ();
 sg13g2_fill_2 FILLER_10_1036 ();
 sg13g2_fill_1 FILLER_10_1038 ();
 sg13g2_fill_1 FILLER_10_1077 ();
 sg13g2_fill_2 FILLER_10_1083 ();
 sg13g2_fill_1 FILLER_10_1085 ();
 sg13g2_decap_4 FILLER_10_1090 ();
 sg13g2_decap_4 FILLER_10_1098 ();
 sg13g2_fill_1 FILLER_10_1102 ();
 sg13g2_fill_2 FILLER_10_1108 ();
 sg13g2_fill_1 FILLER_10_1110 ();
 sg13g2_decap_4 FILLER_10_1119 ();
 sg13g2_fill_1 FILLER_10_1128 ();
 sg13g2_decap_4 FILLER_10_1133 ();
 sg13g2_decap_8 FILLER_10_1141 ();
 sg13g2_decap_8 FILLER_10_1148 ();
 sg13g2_fill_2 FILLER_10_1155 ();
 sg13g2_fill_2 FILLER_10_1212 ();
 sg13g2_fill_1 FILLER_10_1214 ();
 sg13g2_decap_8 FILLER_10_1245 ();
 sg13g2_decap_8 FILLER_10_1252 ();
 sg13g2_decap_8 FILLER_10_1259 ();
 sg13g2_decap_8 FILLER_10_1266 ();
 sg13g2_decap_8 FILLER_10_1273 ();
 sg13g2_decap_8 FILLER_10_1280 ();
 sg13g2_decap_8 FILLER_10_1287 ();
 sg13g2_fill_2 FILLER_10_1294 ();
 sg13g2_decap_8 FILLER_10_1332 ();
 sg13g2_decap_4 FILLER_10_1361 ();
 sg13g2_decap_4 FILLER_10_1373 ();
 sg13g2_fill_2 FILLER_10_1377 ();
 sg13g2_decap_4 FILLER_10_1383 ();
 sg13g2_decap_8 FILLER_10_1434 ();
 sg13g2_fill_2 FILLER_10_1441 ();
 sg13g2_decap_8 FILLER_10_1447 ();
 sg13g2_decap_4 FILLER_10_1454 ();
 sg13g2_fill_2 FILLER_10_1458 ();
 sg13g2_fill_2 FILLER_10_1481 ();
 sg13g2_decap_8 FILLER_10_1487 ();
 sg13g2_decap_4 FILLER_10_1494 ();
 sg13g2_fill_1 FILLER_10_1498 ();
 sg13g2_fill_2 FILLER_10_1509 ();
 sg13g2_fill_1 FILLER_10_1511 ();
 sg13g2_fill_2 FILLER_10_1516 ();
 sg13g2_decap_8 FILLER_10_1528 ();
 sg13g2_decap_8 FILLER_10_1539 ();
 sg13g2_decap_8 FILLER_10_1546 ();
 sg13g2_decap_4 FILLER_10_1567 ();
 sg13g2_fill_2 FILLER_10_1571 ();
 sg13g2_decap_8 FILLER_10_1609 ();
 sg13g2_fill_2 FILLER_10_1616 ();
 sg13g2_fill_2 FILLER_10_1628 ();
 sg13g2_decap_8 FILLER_10_1634 ();
 sg13g2_decap_8 FILLER_10_1641 ();
 sg13g2_fill_1 FILLER_10_1658 ();
 sg13g2_fill_1 FILLER_10_1685 ();
 sg13g2_decap_4 FILLER_10_1733 ();
 sg13g2_fill_1 FILLER_10_1737 ();
 sg13g2_decap_8 FILLER_10_1742 ();
 sg13g2_decap_8 FILLER_10_1749 ();
 sg13g2_decap_8 FILLER_10_1756 ();
 sg13g2_decap_8 FILLER_10_1763 ();
 sg13g2_decap_4 FILLER_10_1770 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_fill_2 FILLER_11_25 ();
 sg13g2_fill_1 FILLER_11_27 ();
 sg13g2_decap_4 FILLER_11_37 ();
 sg13g2_fill_2 FILLER_11_41 ();
 sg13g2_fill_2 FILLER_11_47 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_decap_4 FILLER_11_60 ();
 sg13g2_fill_2 FILLER_11_64 ();
 sg13g2_fill_2 FILLER_11_92 ();
 sg13g2_decap_8 FILLER_11_115 ();
 sg13g2_decap_4 FILLER_11_122 ();
 sg13g2_fill_1 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_131 ();
 sg13g2_fill_1 FILLER_11_138 ();
 sg13g2_fill_2 FILLER_11_212 ();
 sg13g2_fill_1 FILLER_11_244 ();
 sg13g2_fill_2 FILLER_11_273 ();
 sg13g2_fill_1 FILLER_11_275 ();
 sg13g2_fill_1 FILLER_11_341 ();
 sg13g2_fill_1 FILLER_11_404 ();
 sg13g2_decap_8 FILLER_11_436 ();
 sg13g2_decap_4 FILLER_11_443 ();
 sg13g2_fill_1 FILLER_11_447 ();
 sg13g2_fill_1 FILLER_11_456 ();
 sg13g2_decap_4 FILLER_11_462 ();
 sg13g2_fill_1 FILLER_11_471 ();
 sg13g2_fill_2 FILLER_11_507 ();
 sg13g2_fill_1 FILLER_11_509 ();
 sg13g2_fill_2 FILLER_11_519 ();
 sg13g2_fill_1 FILLER_11_521 ();
 sg13g2_fill_2 FILLER_11_527 ();
 sg13g2_fill_1 FILLER_11_529 ();
 sg13g2_decap_4 FILLER_11_534 ();
 sg13g2_fill_2 FILLER_11_538 ();
 sg13g2_decap_8 FILLER_11_545 ();
 sg13g2_decap_4 FILLER_11_552 ();
 sg13g2_fill_2 FILLER_11_556 ();
 sg13g2_fill_1 FILLER_11_563 ();
 sg13g2_decap_8 FILLER_11_603 ();
 sg13g2_fill_1 FILLER_11_610 ();
 sg13g2_fill_2 FILLER_11_621 ();
 sg13g2_fill_1 FILLER_11_628 ();
 sg13g2_fill_2 FILLER_11_633 ();
 sg13g2_fill_1 FILLER_11_635 ();
 sg13g2_decap_4 FILLER_11_640 ();
 sg13g2_fill_1 FILLER_11_703 ();
 sg13g2_decap_8 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_decap_8 FILLER_11_739 ();
 sg13g2_fill_2 FILLER_11_746 ();
 sg13g2_fill_1 FILLER_11_748 ();
 sg13g2_fill_2 FILLER_11_785 ();
 sg13g2_fill_1 FILLER_11_787 ();
 sg13g2_decap_4 FILLER_11_836 ();
 sg13g2_fill_2 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_4 FILLER_11_854 ();
 sg13g2_fill_2 FILLER_11_879 ();
 sg13g2_fill_1 FILLER_11_881 ();
 sg13g2_decap_4 FILLER_11_908 ();
 sg13g2_fill_1 FILLER_11_912 ();
 sg13g2_fill_2 FILLER_11_922 ();
 sg13g2_decap_4 FILLER_11_928 ();
 sg13g2_decap_8 FILLER_11_953 ();
 sg13g2_decap_4 FILLER_11_960 ();
 sg13g2_fill_1 FILLER_11_964 ();
 sg13g2_decap_8 FILLER_11_973 ();
 sg13g2_decap_8 FILLER_11_980 ();
 sg13g2_decap_8 FILLER_11_987 ();
 sg13g2_decap_8 FILLER_11_994 ();
 sg13g2_decap_4 FILLER_11_1001 ();
 sg13g2_fill_2 FILLER_11_1005 ();
 sg13g2_decap_8 FILLER_11_1038 ();
 sg13g2_fill_1 FILLER_11_1045 ();
 sg13g2_fill_1 FILLER_11_1050 ();
 sg13g2_decap_8 FILLER_11_1060 ();
 sg13g2_fill_2 FILLER_11_1067 ();
 sg13g2_decap_4 FILLER_11_1073 ();
 sg13g2_fill_2 FILLER_11_1077 ();
 sg13g2_decap_4 FILLER_11_1157 ();
 sg13g2_fill_1 FILLER_11_1161 ();
 sg13g2_decap_8 FILLER_11_1166 ();
 sg13g2_decap_8 FILLER_11_1173 ();
 sg13g2_fill_1 FILLER_11_1180 ();
 sg13g2_fill_1 FILLER_11_1194 ();
 sg13g2_decap_8 FILLER_11_1228 ();
 sg13g2_decap_8 FILLER_11_1235 ();
 sg13g2_decap_8 FILLER_11_1242 ();
 sg13g2_decap_8 FILLER_11_1249 ();
 sg13g2_decap_8 FILLER_11_1256 ();
 sg13g2_decap_8 FILLER_11_1263 ();
 sg13g2_decap_8 FILLER_11_1270 ();
 sg13g2_decap_8 FILLER_11_1277 ();
 sg13g2_decap_8 FILLER_11_1284 ();
 sg13g2_decap_8 FILLER_11_1291 ();
 sg13g2_decap_4 FILLER_11_1298 ();
 sg13g2_decap_8 FILLER_11_1306 ();
 sg13g2_decap_8 FILLER_11_1313 ();
 sg13g2_fill_2 FILLER_11_1320 ();
 sg13g2_fill_1 FILLER_11_1322 ();
 sg13g2_fill_2 FILLER_11_1344 ();
 sg13g2_decap_8 FILLER_11_1372 ();
 sg13g2_fill_2 FILLER_11_1379 ();
 sg13g2_fill_1 FILLER_11_1381 ();
 sg13g2_decap_8 FILLER_11_1387 ();
 sg13g2_fill_1 FILLER_11_1394 ();
 sg13g2_fill_2 FILLER_11_1405 ();
 sg13g2_fill_1 FILLER_11_1407 ();
 sg13g2_decap_4 FILLER_11_1421 ();
 sg13g2_fill_1 FILLER_11_1425 ();
 sg13g2_decap_4 FILLER_11_1462 ();
 sg13g2_fill_2 FILLER_11_1554 ();
 sg13g2_fill_1 FILLER_11_1556 ();
 sg13g2_decap_4 FILLER_11_1583 ();
 sg13g2_fill_2 FILLER_11_1587 ();
 sg13g2_fill_2 FILLER_11_1620 ();
 sg13g2_fill_1 FILLER_11_1622 ();
 sg13g2_fill_1 FILLER_11_1649 ();
 sg13g2_fill_1 FILLER_11_1660 ();
 sg13g2_fill_1 FILLER_11_1666 ();
 sg13g2_decap_8 FILLER_11_1675 ();
 sg13g2_decap_8 FILLER_11_1682 ();
 sg13g2_fill_1 FILLER_11_1689 ();
 sg13g2_decap_8 FILLER_11_1694 ();
 sg13g2_decap_8 FILLER_11_1701 ();
 sg13g2_fill_2 FILLER_11_1708 ();
 sg13g2_decap_8 FILLER_11_1720 ();
 sg13g2_decap_8 FILLER_11_1727 ();
 sg13g2_decap_8 FILLER_11_1734 ();
 sg13g2_decap_8 FILLER_11_1741 ();
 sg13g2_decap_8 FILLER_11_1748 ();
 sg13g2_decap_8 FILLER_11_1755 ();
 sg13g2_decap_8 FILLER_11_1762 ();
 sg13g2_decap_4 FILLER_11_1769 ();
 sg13g2_fill_1 FILLER_11_1773 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_4 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_fill_1 FILLER_12_123 ();
 sg13g2_fill_2 FILLER_12_129 ();
 sg13g2_decap_8 FILLER_12_135 ();
 sg13g2_decap_4 FILLER_12_142 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_176 ();
 sg13g2_decap_4 FILLER_12_183 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_240 ();
 sg13g2_decap_4 FILLER_12_268 ();
 sg13g2_fill_2 FILLER_12_272 ();
 sg13g2_fill_2 FILLER_12_312 ();
 sg13g2_fill_1 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_fill_1 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_fill_2 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_4 FILLER_12_393 ();
 sg13g2_fill_2 FILLER_12_432 ();
 sg13g2_fill_1 FILLER_12_434 ();
 sg13g2_fill_1 FILLER_12_466 ();
 sg13g2_decap_4 FILLER_12_493 ();
 sg13g2_fill_1 FILLER_12_523 ();
 sg13g2_fill_2 FILLER_12_550 ();
 sg13g2_fill_2 FILLER_12_578 ();
 sg13g2_fill_1 FILLER_12_580 ();
 sg13g2_decap_8 FILLER_12_585 ();
 sg13g2_fill_2 FILLER_12_592 ();
 sg13g2_fill_1 FILLER_12_624 ();
 sg13g2_decap_4 FILLER_12_651 ();
 sg13g2_fill_2 FILLER_12_655 ();
 sg13g2_fill_2 FILLER_12_696 ();
 sg13g2_decap_4 FILLER_12_729 ();
 sg13g2_fill_1 FILLER_12_733 ();
 sg13g2_fill_2 FILLER_12_738 ();
 sg13g2_fill_1 FILLER_12_740 ();
 sg13g2_fill_1 FILLER_12_767 ();
 sg13g2_fill_2 FILLER_12_772 ();
 sg13g2_fill_1 FILLER_12_774 ();
 sg13g2_decap_8 FILLER_12_796 ();
 sg13g2_fill_2 FILLER_12_803 ();
 sg13g2_fill_1 FILLER_12_830 ();
 sg13g2_decap_4 FILLER_12_878 ();
 sg13g2_fill_1 FILLER_12_882 ();
 sg13g2_fill_1 FILLER_12_892 ();
 sg13g2_decap_8 FILLER_12_914 ();
 sg13g2_decap_4 FILLER_12_921 ();
 sg13g2_fill_1 FILLER_12_925 ();
 sg13g2_decap_8 FILLER_12_947 ();
 sg13g2_decap_4 FILLER_12_954 ();
 sg13g2_decap_8 FILLER_12_984 ();
 sg13g2_decap_8 FILLER_12_991 ();
 sg13g2_decap_8 FILLER_12_998 ();
 sg13g2_decap_4 FILLER_12_1010 ();
 sg13g2_fill_2 FILLER_12_1014 ();
 sg13g2_fill_2 FILLER_12_1020 ();
 sg13g2_fill_1 FILLER_12_1022 ();
 sg13g2_decap_8 FILLER_12_1044 ();
 sg13g2_fill_2 FILLER_12_1051 ();
 sg13g2_decap_8 FILLER_12_1074 ();
 sg13g2_decap_8 FILLER_12_1081 ();
 sg13g2_fill_2 FILLER_12_1088 ();
 sg13g2_fill_2 FILLER_12_1111 ();
 sg13g2_fill_1 FILLER_12_1113 ();
 sg13g2_fill_2 FILLER_12_1119 ();
 sg13g2_fill_1 FILLER_12_1121 ();
 sg13g2_fill_1 FILLER_12_1143 ();
 sg13g2_decap_8 FILLER_12_1148 ();
 sg13g2_fill_2 FILLER_12_1155 ();
 sg13g2_fill_2 FILLER_12_1167 ();
 sg13g2_fill_1 FILLER_12_1169 ();
 sg13g2_fill_2 FILLER_12_1196 ();
 sg13g2_fill_1 FILLER_12_1198 ();
 sg13g2_fill_1 FILLER_12_1225 ();
 sg13g2_decap_8 FILLER_12_1252 ();
 sg13g2_decap_8 FILLER_12_1259 ();
 sg13g2_fill_2 FILLER_12_1266 ();
 sg13g2_fill_1 FILLER_12_1268 ();
 sg13g2_decap_8 FILLER_12_1295 ();
 sg13g2_fill_2 FILLER_12_1312 ();
 sg13g2_fill_1 FILLER_12_1314 ();
 sg13g2_decap_8 FILLER_12_1344 ();
 sg13g2_fill_2 FILLER_12_1351 ();
 sg13g2_decap_4 FILLER_12_1357 ();
 sg13g2_fill_1 FILLER_12_1361 ();
 sg13g2_fill_2 FILLER_12_1398 ();
 sg13g2_fill_1 FILLER_12_1400 ();
 sg13g2_fill_1 FILLER_12_1427 ();
 sg13g2_decap_8 FILLER_12_1471 ();
 sg13g2_decap_8 FILLER_12_1478 ();
 sg13g2_decap_8 FILLER_12_1485 ();
 sg13g2_fill_1 FILLER_12_1492 ();
 sg13g2_decap_8 FILLER_12_1503 ();
 sg13g2_fill_1 FILLER_12_1510 ();
 sg13g2_decap_4 FILLER_12_1532 ();
 sg13g2_decap_8 FILLER_12_1540 ();
 sg13g2_decap_4 FILLER_12_1547 ();
 sg13g2_fill_2 FILLER_12_1561 ();
 sg13g2_fill_1 FILLER_12_1563 ();
 sg13g2_decap_4 FILLER_12_1568 ();
 sg13g2_fill_1 FILLER_12_1572 ();
 sg13g2_decap_8 FILLER_12_1583 ();
 sg13g2_decap_4 FILLER_12_1590 ();
 sg13g2_fill_1 FILLER_12_1594 ();
 sg13g2_decap_4 FILLER_12_1599 ();
 sg13g2_decap_8 FILLER_12_1613 ();
 sg13g2_decap_4 FILLER_12_1654 ();
 sg13g2_fill_2 FILLER_12_1658 ();
 sg13g2_fill_1 FILLER_12_1686 ();
 sg13g2_fill_2 FILLER_12_1695 ();
 sg13g2_fill_2 FILLER_12_1707 ();
 sg13g2_decap_8 FILLER_12_1739 ();
 sg13g2_decap_8 FILLER_12_1746 ();
 sg13g2_decap_8 FILLER_12_1753 ();
 sg13g2_decap_8 FILLER_12_1760 ();
 sg13g2_decap_8 FILLER_12_1767 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_15 ();
 sg13g2_fill_2 FILLER_13_47 ();
 sg13g2_fill_2 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_73 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_fill_2 FILLER_13_150 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_4 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_fill_2 FILLER_13_210 ();
 sg13g2_fill_2 FILLER_13_227 ();
 sg13g2_fill_2 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_fill_1 FILLER_13_305 ();
 sg13g2_fill_1 FILLER_13_315 ();
 sg13g2_fill_2 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_fill_2 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_fill_2 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_418 ();
 sg13g2_decap_4 FILLER_13_425 ();
 sg13g2_fill_2 FILLER_13_429 ();
 sg13g2_decap_4 FILLER_13_436 ();
 sg13g2_fill_1 FILLER_13_440 ();
 sg13g2_decap_8 FILLER_13_445 ();
 sg13g2_fill_1 FILLER_13_477 ();
 sg13g2_decap_4 FILLER_13_507 ();
 sg13g2_fill_1 FILLER_13_511 ();
 sg13g2_decap_4 FILLER_13_520 ();
 sg13g2_decap_8 FILLER_13_549 ();
 sg13g2_decap_4 FILLER_13_556 ();
 sg13g2_fill_1 FILLER_13_564 ();
 sg13g2_decap_8 FILLER_13_586 ();
 sg13g2_fill_1 FILLER_13_593 ();
 sg13g2_decap_4 FILLER_13_598 ();
 sg13g2_fill_1 FILLER_13_602 ();
 sg13g2_fill_2 FILLER_13_612 ();
 sg13g2_fill_1 FILLER_13_614 ();
 sg13g2_fill_1 FILLER_13_619 ();
 sg13g2_fill_2 FILLER_13_641 ();
 sg13g2_fill_2 FILLER_13_648 ();
 sg13g2_fill_1 FILLER_13_650 ();
 sg13g2_fill_1 FILLER_13_664 ();
 sg13g2_fill_1 FILLER_13_670 ();
 sg13g2_fill_1 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_741 ();
 sg13g2_decap_4 FILLER_13_752 ();
 sg13g2_fill_1 FILLER_13_760 ();
 sg13g2_decap_4 FILLER_13_771 ();
 sg13g2_decap_8 FILLER_13_796 ();
 sg13g2_decap_8 FILLER_13_803 ();
 sg13g2_fill_1 FILLER_13_810 ();
 sg13g2_decap_8 FILLER_13_832 ();
 sg13g2_decap_8 FILLER_13_843 ();
 sg13g2_fill_1 FILLER_13_850 ();
 sg13g2_decap_4 FILLER_13_855 ();
 sg13g2_decap_8 FILLER_13_867 ();
 sg13g2_decap_4 FILLER_13_874 ();
 sg13g2_fill_2 FILLER_13_883 ();
 sg13g2_fill_1 FILLER_13_885 ();
 sg13g2_fill_2 FILLER_13_894 ();
 sg13g2_decap_4 FILLER_13_917 ();
 sg13g2_fill_1 FILLER_13_921 ();
 sg13g2_decap_8 FILLER_13_926 ();
 sg13g2_decap_8 FILLER_13_933 ();
 sg13g2_decap_8 FILLER_13_940 ();
 sg13g2_decap_4 FILLER_13_947 ();
 sg13g2_fill_2 FILLER_13_960 ();
 sg13g2_decap_4 FILLER_13_996 ();
 sg13g2_fill_2 FILLER_13_1047 ();
 sg13g2_fill_1 FILLER_13_1049 ();
 sg13g2_fill_2 FILLER_13_1054 ();
 sg13g2_fill_1 FILLER_13_1056 ();
 sg13g2_fill_2 FILLER_13_1083 ();
 sg13g2_fill_1 FILLER_13_1089 ();
 sg13g2_fill_2 FILLER_13_1162 ();
 sg13g2_fill_2 FILLER_13_1174 ();
 sg13g2_fill_1 FILLER_13_1176 ();
 sg13g2_decap_8 FILLER_13_1181 ();
 sg13g2_decap_4 FILLER_13_1188 ();
 sg13g2_decap_4 FILLER_13_1217 ();
 sg13g2_fill_1 FILLER_13_1221 ();
 sg13g2_decap_8 FILLER_13_1252 ();
 sg13g2_decap_8 FILLER_13_1259 ();
 sg13g2_decap_8 FILLER_13_1266 ();
 sg13g2_fill_2 FILLER_13_1273 ();
 sg13g2_decap_8 FILLER_13_1279 ();
 sg13g2_decap_8 FILLER_13_1286 ();
 sg13g2_fill_1 FILLER_13_1323 ();
 sg13g2_fill_2 FILLER_13_1334 ();
 sg13g2_fill_1 FILLER_13_1346 ();
 sg13g2_decap_4 FILLER_13_1373 ();
 sg13g2_fill_1 FILLER_13_1377 ();
 sg13g2_decap_4 FILLER_13_1382 ();
 sg13g2_fill_1 FILLER_13_1386 ();
 sg13g2_decap_8 FILLER_13_1416 ();
 sg13g2_decap_8 FILLER_13_1423 ();
 sg13g2_decap_8 FILLER_13_1430 ();
 sg13g2_fill_1 FILLER_13_1437 ();
 sg13g2_decap_8 FILLER_13_1448 ();
 sg13g2_decap_8 FILLER_13_1455 ();
 sg13g2_decap_8 FILLER_13_1462 ();
 sg13g2_decap_8 FILLER_13_1521 ();
 sg13g2_fill_2 FILLER_13_1528 ();
 sg13g2_decap_8 FILLER_13_1534 ();
 sg13g2_decap_4 FILLER_13_1541 ();
 sg13g2_fill_1 FILLER_13_1545 ();
 sg13g2_decap_8 FILLER_13_1572 ();
 sg13g2_fill_2 FILLER_13_1579 ();
 sg13g2_decap_4 FILLER_13_1607 ();
 sg13g2_fill_1 FILLER_13_1611 ();
 sg13g2_fill_1 FILLER_13_1624 ();
 sg13g2_decap_8 FILLER_13_1661 ();
 sg13g2_decap_4 FILLER_13_1668 ();
 sg13g2_fill_1 FILLER_13_1672 ();
 sg13g2_fill_2 FILLER_13_1677 ();
 sg13g2_fill_1 FILLER_13_1679 ();
 sg13g2_fill_1 FILLER_13_1684 ();
 sg13g2_decap_8 FILLER_13_1706 ();
 sg13g2_decap_4 FILLER_13_1713 ();
 sg13g2_fill_2 FILLER_13_1717 ();
 sg13g2_decap_8 FILLER_13_1749 ();
 sg13g2_decap_8 FILLER_13_1756 ();
 sg13g2_decap_8 FILLER_13_1763 ();
 sg13g2_decap_4 FILLER_13_1770 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_29 ();
 sg13g2_decap_8 FILLER_14_36 ();
 sg13g2_fill_1 FILLER_14_43 ();
 sg13g2_fill_1 FILLER_14_48 ();
 sg13g2_fill_1 FILLER_14_75 ();
 sg13g2_fill_1 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_86 ();
 sg13g2_fill_2 FILLER_14_93 ();
 sg13g2_decap_8 FILLER_14_120 ();
 sg13g2_decap_8 FILLER_14_131 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_fill_1 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_fill_2 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_fill_2 FILLER_14_203 ();
 sg13g2_fill_1 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_211 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_decap_8 FILLER_14_225 ();
 sg13g2_fill_2 FILLER_14_232 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_240 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_fill_1 FILLER_14_253 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_fill_1 FILLER_14_269 ();
 sg13g2_fill_2 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_decap_4 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_302 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_332 ();
 sg13g2_fill_1 FILLER_14_337 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_fill_2 FILLER_14_360 ();
 sg13g2_fill_2 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_369 ();
 sg13g2_fill_2 FILLER_14_374 ();
 sg13g2_fill_1 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_fill_2 FILLER_14_403 ();
 sg13g2_fill_1 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_fill_2 FILLER_14_430 ();
 sg13g2_fill_2 FILLER_14_437 ();
 sg13g2_decap_8 FILLER_14_443 ();
 sg13g2_decap_4 FILLER_14_450 ();
 sg13g2_fill_1 FILLER_14_454 ();
 sg13g2_decap_4 FILLER_14_476 ();
 sg13g2_fill_2 FILLER_14_480 ();
 sg13g2_decap_4 FILLER_14_524 ();
 sg13g2_decap_8 FILLER_14_549 ();
 sg13g2_decap_4 FILLER_14_556 ();
 sg13g2_decap_4 FILLER_14_565 ();
 sg13g2_decap_4 FILLER_14_590 ();
 sg13g2_fill_1 FILLER_14_594 ();
 sg13g2_fill_2 FILLER_14_621 ();
 sg13g2_fill_1 FILLER_14_623 ();
 sg13g2_decap_4 FILLER_14_645 ();
 sg13g2_fill_1 FILLER_14_649 ();
 sg13g2_fill_1 FILLER_14_679 ();
 sg13g2_fill_2 FILLER_14_701 ();
 sg13g2_decap_8 FILLER_14_740 ();
 sg13g2_fill_2 FILLER_14_747 ();
 sg13g2_decap_8 FILLER_14_757 ();
 sg13g2_decap_4 FILLER_14_764 ();
 sg13g2_fill_2 FILLER_14_768 ();
 sg13g2_fill_1 FILLER_14_784 ();
 sg13g2_fill_2 FILLER_14_837 ();
 sg13g2_fill_1 FILLER_14_839 ();
 sg13g2_decap_8 FILLER_14_871 ();
 sg13g2_fill_1 FILLER_14_878 ();
 sg13g2_decap_4 FILLER_14_905 ();
 sg13g2_fill_2 FILLER_14_909 ();
 sg13g2_fill_2 FILLER_14_942 ();
 sg13g2_fill_1 FILLER_14_944 ();
 sg13g2_fill_1 FILLER_14_976 ();
 sg13g2_decap_8 FILLER_14_998 ();
 sg13g2_fill_2 FILLER_14_1005 ();
 sg13g2_decap_8 FILLER_14_1011 ();
 sg13g2_decap_8 FILLER_14_1018 ();
 sg13g2_decap_8 FILLER_14_1025 ();
 sg13g2_decap_8 FILLER_14_1032 ();
 sg13g2_decap_4 FILLER_14_1039 ();
 sg13g2_fill_2 FILLER_14_1048 ();
 sg13g2_fill_1 FILLER_14_1050 ();
 sg13g2_decap_8 FILLER_14_1055 ();
 sg13g2_decap_4 FILLER_14_1062 ();
 sg13g2_decap_8 FILLER_14_1096 ();
 sg13g2_decap_8 FILLER_14_1103 ();
 sg13g2_decap_4 FILLER_14_1115 ();
 sg13g2_fill_2 FILLER_14_1119 ();
 sg13g2_decap_8 FILLER_14_1147 ();
 sg13g2_decap_8 FILLER_14_1154 ();
 sg13g2_fill_1 FILLER_14_1191 ();
 sg13g2_fill_2 FILLER_14_1218 ();
 sg13g2_fill_1 FILLER_14_1220 ();
 sg13g2_fill_1 FILLER_14_1231 ();
 sg13g2_decap_8 FILLER_14_1240 ();
 sg13g2_decap_8 FILLER_14_1247 ();
 sg13g2_decap_8 FILLER_14_1254 ();
 sg13g2_fill_2 FILLER_14_1261 ();
 sg13g2_decap_8 FILLER_14_1276 ();
 sg13g2_decap_8 FILLER_14_1283 ();
 sg13g2_decap_8 FILLER_14_1290 ();
 sg13g2_decap_8 FILLER_14_1297 ();
 sg13g2_decap_8 FILLER_14_1304 ();
 sg13g2_decap_8 FILLER_14_1311 ();
 sg13g2_decap_8 FILLER_14_1318 ();
 sg13g2_fill_1 FILLER_14_1325 ();
 sg13g2_fill_2 FILLER_14_1352 ();
 sg13g2_fill_1 FILLER_14_1354 ();
 sg13g2_fill_2 FILLER_14_1363 ();
 sg13g2_decap_4 FILLER_14_1391 ();
 sg13g2_fill_2 FILLER_14_1395 ();
 sg13g2_decap_8 FILLER_14_1402 ();
 sg13g2_decap_4 FILLER_14_1409 ();
 sg13g2_fill_2 FILLER_14_1413 ();
 sg13g2_decap_8 FILLER_14_1419 ();
 sg13g2_fill_2 FILLER_14_1426 ();
 sg13g2_fill_1 FILLER_14_1428 ();
 sg13g2_fill_2 FILLER_14_1439 ();
 sg13g2_fill_2 FILLER_14_1450 ();
 sg13g2_fill_1 FILLER_14_1452 ();
 sg13g2_decap_4 FILLER_14_1474 ();
 sg13g2_decap_8 FILLER_14_1482 ();
 sg13g2_decap_8 FILLER_14_1489 ();
 sg13g2_fill_1 FILLER_14_1496 ();
 sg13g2_decap_8 FILLER_14_1505 ();
 sg13g2_fill_2 FILLER_14_1512 ();
 sg13g2_decap_8 FILLER_14_1554 ();
 sg13g2_decap_4 FILLER_14_1561 ();
 sg13g2_fill_2 FILLER_14_1565 ();
 sg13g2_decap_8 FILLER_14_1592 ();
 sg13g2_fill_1 FILLER_14_1599 ();
 sg13g2_decap_4 FILLER_14_1636 ();
 sg13g2_fill_2 FILLER_14_1640 ();
 sg13g2_decap_8 FILLER_14_1646 ();
 sg13g2_decap_4 FILLER_14_1653 ();
 sg13g2_decap_4 FILLER_14_1769 ();
 sg13g2_fill_1 FILLER_14_1773 ();
 sg13g2_fill_2 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_55 ();
 sg13g2_decap_8 FILLER_15_62 ();
 sg13g2_decap_4 FILLER_15_69 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_decap_4 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_87 ();
 sg13g2_decap_8 FILLER_15_92 ();
 sg13g2_decap_8 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_106 ();
 sg13g2_fill_2 FILLER_15_113 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_fill_2 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_decap_8 FILLER_15_157 ();
 sg13g2_decap_8 FILLER_15_164 ();
 sg13g2_fill_1 FILLER_15_171 ();
 sg13g2_fill_1 FILLER_15_259 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_307 ();
 sg13g2_decap_4 FILLER_15_318 ();
 sg13g2_fill_1 FILLER_15_322 ();
 sg13g2_decap_4 FILLER_15_344 ();
 sg13g2_fill_2 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_458 ();
 sg13g2_decap_8 FILLER_15_465 ();
 sg13g2_decap_8 FILLER_15_472 ();
 sg13g2_decap_4 FILLER_15_479 ();
 sg13g2_decap_4 FILLER_15_496 ();
 sg13g2_decap_8 FILLER_15_531 ();
 sg13g2_fill_1 FILLER_15_538 ();
 sg13g2_decap_4 FILLER_15_581 ();
 sg13g2_fill_1 FILLER_15_585 ();
 sg13g2_decap_8 FILLER_15_591 ();
 sg13g2_decap_4 FILLER_15_598 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_fill_1 FILLER_15_613 ();
 sg13g2_decap_4 FILLER_15_619 ();
 sg13g2_fill_1 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_628 ();
 sg13g2_decap_8 FILLER_15_635 ();
 sg13g2_decap_8 FILLER_15_642 ();
 sg13g2_decap_8 FILLER_15_649 ();
 sg13g2_fill_2 FILLER_15_660 ();
 sg13g2_fill_2 FILLER_15_674 ();
 sg13g2_fill_2 FILLER_15_706 ();
 sg13g2_fill_1 FILLER_15_731 ();
 sg13g2_decap_8 FILLER_15_736 ();
 sg13g2_decap_4 FILLER_15_743 ();
 sg13g2_fill_1 FILLER_15_747 ();
 sg13g2_fill_1 FILLER_15_764 ();
 sg13g2_decap_8 FILLER_15_769 ();
 sg13g2_fill_2 FILLER_15_780 ();
 sg13g2_decap_4 FILLER_15_786 ();
 sg13g2_fill_2 FILLER_15_790 ();
 sg13g2_decap_8 FILLER_15_796 ();
 sg13g2_decap_4 FILLER_15_803 ();
 sg13g2_fill_1 FILLER_15_807 ();
 sg13g2_fill_1 FILLER_15_823 ();
 sg13g2_decap_8 FILLER_15_828 ();
 sg13g2_decap_8 FILLER_15_835 ();
 sg13g2_decap_8 FILLER_15_842 ();
 sg13g2_fill_2 FILLER_15_849 ();
 sg13g2_decap_4 FILLER_15_855 ();
 sg13g2_fill_1 FILLER_15_859 ();
 sg13g2_fill_1 FILLER_15_865 ();
 sg13g2_decap_8 FILLER_15_870 ();
 sg13g2_decap_4 FILLER_15_877 ();
 sg13g2_fill_1 FILLER_15_881 ();
 sg13g2_decap_4 FILLER_15_887 ();
 sg13g2_fill_2 FILLER_15_891 ();
 sg13g2_decap_4 FILLER_15_897 ();
 sg13g2_decap_8 FILLER_15_905 ();
 sg13g2_decap_4 FILLER_15_917 ();
 sg13g2_decap_4 FILLER_15_925 ();
 sg13g2_decap_8 FILLER_15_933 ();
 sg13g2_decap_8 FILLER_15_940 ();
 sg13g2_decap_8 FILLER_15_947 ();
 sg13g2_decap_4 FILLER_15_954 ();
 sg13g2_fill_2 FILLER_15_988 ();
 sg13g2_fill_1 FILLER_15_990 ();
 sg13g2_decap_8 FILLER_15_1021 ();
 sg13g2_decap_8 FILLER_15_1028 ();
 sg13g2_decap_4 FILLER_15_1035 ();
 sg13g2_fill_1 FILLER_15_1039 ();
 sg13g2_decap_8 FILLER_15_1066 ();
 sg13g2_decap_8 FILLER_15_1073 ();
 sg13g2_decap_8 FILLER_15_1080 ();
 sg13g2_fill_2 FILLER_15_1087 ();
 sg13g2_fill_1 FILLER_15_1089 ();
 sg13g2_fill_2 FILLER_15_1095 ();
 sg13g2_decap_4 FILLER_15_1101 ();
 sg13g2_fill_2 FILLER_15_1110 ();
 sg13g2_fill_1 FILLER_15_1112 ();
 sg13g2_fill_1 FILLER_15_1126 ();
 sg13g2_decap_4 FILLER_15_1131 ();
 sg13g2_decap_8 FILLER_15_1148 ();
 sg13g2_decap_8 FILLER_15_1155 ();
 sg13g2_decap_8 FILLER_15_1162 ();
 sg13g2_decap_8 FILLER_15_1169 ();
 sg13g2_decap_8 FILLER_15_1176 ();
 sg13g2_decap_8 FILLER_15_1183 ();
 sg13g2_decap_8 FILLER_15_1190 ();
 sg13g2_decap_8 FILLER_15_1197 ();
 sg13g2_decap_8 FILLER_15_1204 ();
 sg13g2_decap_8 FILLER_15_1211 ();
 sg13g2_fill_1 FILLER_15_1228 ();
 sg13g2_decap_8 FILLER_15_1255 ();
 sg13g2_fill_2 FILLER_15_1262 ();
 sg13g2_fill_2 FILLER_15_1294 ();
 sg13g2_decap_8 FILLER_15_1306 ();
 sg13g2_fill_2 FILLER_15_1313 ();
 sg13g2_fill_1 FILLER_15_1320 ();
 sg13g2_decap_8 FILLER_15_1339 ();
 sg13g2_decap_4 FILLER_15_1346 ();
 sg13g2_fill_1 FILLER_15_1358 ();
 sg13g2_decap_4 FILLER_15_1376 ();
 sg13g2_fill_2 FILLER_15_1390 ();
 sg13g2_fill_2 FILLER_15_1396 ();
 sg13g2_fill_1 FILLER_15_1460 ();
 sg13g2_decap_8 FILLER_15_1475 ();
 sg13g2_decap_4 FILLER_15_1482 ();
 sg13g2_decap_8 FILLER_15_1531 ();
 sg13g2_decap_8 FILLER_15_1538 ();
 sg13g2_decap_8 FILLER_15_1545 ();
 sg13g2_fill_2 FILLER_15_1552 ();
 sg13g2_decap_8 FILLER_15_1590 ();
 sg13g2_fill_1 FILLER_15_1597 ();
 sg13g2_decap_4 FILLER_15_1602 ();
 sg13g2_decap_4 FILLER_15_1616 ();
 sg13g2_fill_2 FILLER_15_1620 ();
 sg13g2_fill_2 FILLER_15_1632 ();
 sg13g2_decap_8 FILLER_15_1638 ();
 sg13g2_decap_4 FILLER_15_1645 ();
 sg13g2_fill_1 FILLER_15_1649 ();
 sg13g2_fill_2 FILLER_15_1707 ();
 sg13g2_decap_8 FILLER_15_1728 ();
 sg13g2_fill_2 FILLER_15_1735 ();
 sg13g2_fill_1 FILLER_15_1737 ();
 sg13g2_decap_4 FILLER_15_1768 ();
 sg13g2_fill_2 FILLER_15_1772 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_32 ();
 sg13g2_fill_1 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_fill_1 FILLER_16_207 ();
 sg13g2_fill_2 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_227 ();
 sg13g2_fill_2 FILLER_16_253 ();
 sg13g2_fill_1 FILLER_16_255 ();
 sg13g2_decap_4 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_fill_2 FILLER_16_288 ();
 sg13g2_fill_1 FILLER_16_290 ();
 sg13g2_fill_2 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_351 ();
 sg13g2_fill_2 FILLER_16_360 ();
 sg13g2_fill_2 FILLER_16_393 ();
 sg13g2_fill_1 FILLER_16_395 ();
 sg13g2_decap_4 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_404 ();
 sg13g2_decap_8 FILLER_16_410 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_fill_2 FILLER_16_424 ();
 sg13g2_decap_8 FILLER_16_431 ();
 sg13g2_decap_8 FILLER_16_438 ();
 sg13g2_decap_8 FILLER_16_445 ();
 sg13g2_decap_8 FILLER_16_452 ();
 sg13g2_fill_1 FILLER_16_459 ();
 sg13g2_decap_4 FILLER_16_465 ();
 sg13g2_fill_2 FILLER_16_473 ();
 sg13g2_fill_1 FILLER_16_475 ();
 sg13g2_fill_1 FILLER_16_485 ();
 sg13g2_fill_2 FILLER_16_490 ();
 sg13g2_fill_2 FILLER_16_510 ();
 sg13g2_decap_4 FILLER_16_517 ();
 sg13g2_fill_1 FILLER_16_521 ();
 sg13g2_decap_8 FILLER_16_530 ();
 sg13g2_fill_2 FILLER_16_537 ();
 sg13g2_fill_1 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_544 ();
 sg13g2_decap_8 FILLER_16_551 ();
 sg13g2_fill_2 FILLER_16_558 ();
 sg13g2_fill_1 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_566 ();
 sg13g2_decap_8 FILLER_16_573 ();
 sg13g2_decap_4 FILLER_16_580 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_4 FILLER_16_602 ();
 sg13g2_fill_2 FILLER_16_606 ();
 sg13g2_fill_1 FILLER_16_638 ();
 sg13g2_fill_1 FILLER_16_675 ();
 sg13g2_fill_1 FILLER_16_702 ();
 sg13g2_decap_8 FILLER_16_762 ();
 sg13g2_decap_4 FILLER_16_769 ();
 sg13g2_fill_1 FILLER_16_809 ();
 sg13g2_fill_2 FILLER_16_815 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_fill_1 FILLER_16_850 ();
 sg13g2_decap_4 FILLER_16_877 ();
 sg13g2_fill_1 FILLER_16_881 ();
 sg13g2_fill_1 FILLER_16_908 ();
 sg13g2_fill_1 FILLER_16_940 ();
 sg13g2_fill_2 FILLER_16_950 ();
 sg13g2_fill_2 FILLER_16_957 ();
 sg13g2_fill_2 FILLER_16_964 ();
 sg13g2_fill_1 FILLER_16_966 ();
 sg13g2_fill_1 FILLER_16_971 ();
 sg13g2_decap_8 FILLER_16_976 ();
 sg13g2_decap_8 FILLER_16_983 ();
 sg13g2_decap_8 FILLER_16_990 ();
 sg13g2_decap_4 FILLER_16_1007 ();
 sg13g2_fill_1 FILLER_16_1024 ();
 sg13g2_decap_8 FILLER_16_1029 ();
 sg13g2_decap_4 FILLER_16_1036 ();
 sg13g2_fill_1 FILLER_16_1040 ();
 sg13g2_decap_8 FILLER_16_1072 ();
 sg13g2_fill_1 FILLER_16_1105 ();
 sg13g2_decap_8 FILLER_16_1132 ();
 sg13g2_decap_8 FILLER_16_1139 ();
 sg13g2_decap_8 FILLER_16_1146 ();
 sg13g2_decap_8 FILLER_16_1153 ();
 sg13g2_decap_8 FILLER_16_1196 ();
 sg13g2_decap_8 FILLER_16_1203 ();
 sg13g2_decap_8 FILLER_16_1210 ();
 sg13g2_fill_2 FILLER_16_1217 ();
 sg13g2_decap_8 FILLER_16_1255 ();
 sg13g2_decap_8 FILLER_16_1262 ();
 sg13g2_fill_1 FILLER_16_1269 ();
 sg13g2_decap_8 FILLER_16_1274 ();
 sg13g2_fill_2 FILLER_16_1281 ();
 sg13g2_decap_8 FILLER_16_1319 ();
 sg13g2_decap_8 FILLER_16_1326 ();
 sg13g2_decap_8 FILLER_16_1333 ();
 sg13g2_decap_4 FILLER_16_1340 ();
 sg13g2_fill_1 FILLER_16_1344 ();
 sg13g2_decap_4 FILLER_16_1353 ();
 sg13g2_fill_1 FILLER_16_1357 ();
 sg13g2_decap_8 FILLER_16_1394 ();
 sg13g2_decap_8 FILLER_16_1401 ();
 sg13g2_decap_8 FILLER_16_1408 ();
 sg13g2_decap_8 FILLER_16_1415 ();
 sg13g2_decap_8 FILLER_16_1422 ();
 sg13g2_fill_2 FILLER_16_1429 ();
 sg13g2_fill_1 FILLER_16_1431 ();
 sg13g2_decap_4 FILLER_16_1442 ();
 sg13g2_fill_1 FILLER_16_1446 ();
 sg13g2_fill_2 FILLER_16_1487 ();
 sg13g2_fill_1 FILLER_16_1489 ();
 sg13g2_fill_1 FILLER_16_1521 ();
 sg13g2_decap_8 FILLER_16_1548 ();
 sg13g2_decap_8 FILLER_16_1555 ();
 sg13g2_fill_2 FILLER_16_1562 ();
 sg13g2_fill_2 FILLER_16_1572 ();
 sg13g2_fill_1 FILLER_16_1574 ();
 sg13g2_decap_8 FILLER_16_1618 ();
 sg13g2_fill_2 FILLER_16_1625 ();
 sg13g2_decap_8 FILLER_16_1653 ();
 sg13g2_decap_4 FILLER_16_1660 ();
 sg13g2_decap_8 FILLER_16_1672 ();
 sg13g2_decap_4 FILLER_16_1679 ();
 sg13g2_fill_1 FILLER_16_1683 ();
 sg13g2_decap_4 FILLER_16_1697 ();
 sg13g2_fill_1 FILLER_16_1701 ();
 sg13g2_fill_2 FILLER_16_1710 ();
 sg13g2_fill_1 FILLER_16_1712 ();
 sg13g2_decap_8 FILLER_16_1766 ();
 sg13g2_fill_1 FILLER_16_1773 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_12 ();
 sg13g2_decap_8 FILLER_17_19 ();
 sg13g2_fill_1 FILLER_17_26 ();
 sg13g2_fill_2 FILLER_17_31 ();
 sg13g2_fill_1 FILLER_17_33 ();
 sg13g2_decap_4 FILLER_17_65 ();
 sg13g2_fill_1 FILLER_17_69 ();
 sg13g2_decap_8 FILLER_17_74 ();
 sg13g2_decap_8 FILLER_17_81 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_90 ();
 sg13g2_decap_4 FILLER_17_112 ();
 sg13g2_decap_4 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_decap_8 FILLER_17_129 ();
 sg13g2_decap_4 FILLER_17_136 ();
 sg13g2_decap_8 FILLER_17_144 ();
 sg13g2_decap_8 FILLER_17_151 ();
 sg13g2_fill_2 FILLER_17_158 ();
 sg13g2_fill_1 FILLER_17_160 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_decap_4 FILLER_17_224 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_4 FILLER_17_287 ();
 sg13g2_fill_1 FILLER_17_291 ();
 sg13g2_fill_2 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_fill_2 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_4 FILLER_17_362 ();
 sg13g2_fill_2 FILLER_17_366 ();
 sg13g2_fill_1 FILLER_17_373 ();
 sg13g2_fill_1 FILLER_17_378 ();
 sg13g2_fill_1 FILLER_17_383 ();
 sg13g2_fill_1 FILLER_17_397 ();
 sg13g2_fill_1 FILLER_17_424 ();
 sg13g2_fill_1 FILLER_17_451 ();
 sg13g2_fill_1 FILLER_17_478 ();
 sg13g2_decap_8 FILLER_17_505 ();
 sg13g2_fill_2 FILLER_17_538 ();
 sg13g2_fill_2 FILLER_17_571 ();
 sg13g2_fill_1 FILLER_17_573 ();
 sg13g2_decap_8 FILLER_17_608 ();
 sg13g2_fill_1 FILLER_17_672 ();
 sg13g2_fill_1 FILLER_17_713 ();
 sg13g2_fill_2 FILLER_17_732 ();
 sg13g2_fill_1 FILLER_17_734 ();
 sg13g2_decap_8 FILLER_17_740 ();
 sg13g2_fill_1 FILLER_17_747 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_4 FILLER_17_770 ();
 sg13g2_fill_2 FILLER_17_774 ();
 sg13g2_decap_4 FILLER_17_780 ();
 sg13g2_fill_1 FILLER_17_784 ();
 sg13g2_fill_2 FILLER_17_794 ();
 sg13g2_fill_1 FILLER_17_796 ();
 sg13g2_fill_2 FILLER_17_801 ();
 sg13g2_fill_1 FILLER_17_803 ();
 sg13g2_decap_4 FILLER_17_825 ();
 sg13g2_decap_8 FILLER_17_850 ();
 sg13g2_fill_2 FILLER_17_857 ();
 sg13g2_decap_4 FILLER_17_863 ();
 sg13g2_fill_1 FILLER_17_867 ();
 sg13g2_fill_2 FILLER_17_872 ();
 sg13g2_fill_1 FILLER_17_874 ();
 sg13g2_decap_4 FILLER_17_911 ();
 sg13g2_fill_2 FILLER_17_915 ();
 sg13g2_decap_8 FILLER_17_921 ();
 sg13g2_fill_1 FILLER_17_928 ();
 sg13g2_decap_8 FILLER_17_967 ();
 sg13g2_decap_4 FILLER_17_1009 ();
 sg13g2_fill_1 FILLER_17_1013 ();
 sg13g2_decap_4 FILLER_17_1040 ();
 sg13g2_decap_4 FILLER_17_1065 ();
 sg13g2_decap_8 FILLER_17_1074 ();
 sg13g2_fill_2 FILLER_17_1085 ();
 sg13g2_fill_2 FILLER_17_1137 ();
 sg13g2_fill_1 FILLER_17_1139 ();
 sg13g2_decap_8 FILLER_17_1161 ();
 sg13g2_decap_8 FILLER_17_1168 ();
 sg13g2_decap_4 FILLER_17_1175 ();
 sg13g2_fill_1 FILLER_17_1179 ();
 sg13g2_decap_8 FILLER_17_1184 ();
 sg13g2_fill_1 FILLER_17_1191 ();
 sg13g2_fill_1 FILLER_17_1213 ();
 sg13g2_fill_1 FILLER_17_1224 ();
 sg13g2_decap_4 FILLER_17_1255 ();
 sg13g2_fill_1 FILLER_17_1259 ();
 sg13g2_fill_1 FILLER_17_1264 ();
 sg13g2_fill_2 FILLER_17_1291 ();
 sg13g2_fill_1 FILLER_17_1303 ();
 sg13g2_fill_2 FILLER_17_1325 ();
 sg13g2_decap_8 FILLER_17_1348 ();
 sg13g2_fill_1 FILLER_17_1355 ();
 sg13g2_decap_4 FILLER_17_1370 ();
 sg13g2_fill_1 FILLER_17_1374 ();
 sg13g2_decap_8 FILLER_17_1379 ();
 sg13g2_decap_8 FILLER_17_1386 ();
 sg13g2_decap_4 FILLER_17_1393 ();
 sg13g2_decap_8 FILLER_17_1459 ();
 sg13g2_decap_8 FILLER_17_1466 ();
 sg13g2_decap_8 FILLER_17_1473 ();
 sg13g2_decap_8 FILLER_17_1480 ();
 sg13g2_decap_8 FILLER_17_1487 ();
 sg13g2_decap_4 FILLER_17_1494 ();
 sg13g2_fill_2 FILLER_17_1498 ();
 sg13g2_decap_8 FILLER_17_1510 ();
 sg13g2_fill_1 FILLER_17_1517 ();
 sg13g2_decap_8 FILLER_17_1543 ();
 sg13g2_fill_1 FILLER_17_1550 ();
 sg13g2_fill_1 FILLER_17_1556 ();
 sg13g2_decap_8 FILLER_17_1587 ();
 sg13g2_fill_2 FILLER_17_1609 ();
 sg13g2_decap_4 FILLER_17_1615 ();
 sg13g2_decap_8 FILLER_17_1640 ();
 sg13g2_decap_4 FILLER_17_1647 ();
 sg13g2_fill_2 FILLER_17_1687 ();
 sg13g2_fill_1 FILLER_17_1689 ();
 sg13g2_fill_1 FILLER_17_1721 ();
 sg13g2_fill_2 FILLER_17_1732 ();
 sg13g2_decap_4 FILLER_17_1738 ();
 sg13g2_decap_4 FILLER_17_1768 ();
 sg13g2_fill_2 FILLER_17_1772 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_47 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_84 ();
 sg13g2_fill_1 FILLER_18_86 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_4 FILLER_18_189 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_229 ();
 sg13g2_fill_2 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_fill_2 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_4 FILLER_18_392 ();
 sg13g2_decap_4 FILLER_18_417 ();
 sg13g2_fill_1 FILLER_18_421 ();
 sg13g2_fill_1 FILLER_18_426 ();
 sg13g2_decap_8 FILLER_18_432 ();
 sg13g2_fill_1 FILLER_18_439 ();
 sg13g2_decap_8 FILLER_18_444 ();
 sg13g2_decap_4 FILLER_18_451 ();
 sg13g2_fill_2 FILLER_18_455 ();
 sg13g2_decap_4 FILLER_18_466 ();
 sg13g2_fill_2 FILLER_18_474 ();
 sg13g2_decap_8 FILLER_18_522 ();
 sg13g2_decap_8 FILLER_18_529 ();
 sg13g2_decap_8 FILLER_18_536 ();
 sg13g2_decap_8 FILLER_18_582 ();
 sg13g2_decap_8 FILLER_18_589 ();
 sg13g2_decap_4 FILLER_18_596 ();
 sg13g2_fill_2 FILLER_18_600 ();
 sg13g2_decap_8 FILLER_18_606 ();
 sg13g2_fill_1 FILLER_18_613 ();
 sg13g2_decap_4 FILLER_18_619 ();
 sg13g2_fill_2 FILLER_18_649 ();
 sg13g2_fill_1 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_656 ();
 sg13g2_fill_2 FILLER_18_663 ();
 sg13g2_decap_8 FILLER_18_674 ();
 sg13g2_fill_2 FILLER_18_681 ();
 sg13g2_fill_1 FILLER_18_683 ();
 sg13g2_fill_1 FILLER_18_699 ();
 sg13g2_decap_4 FILLER_18_747 ();
 sg13g2_fill_1 FILLER_18_751 ();
 sg13g2_decap_4 FILLER_18_797 ();
 sg13g2_fill_2 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_824 ();
 sg13g2_decap_8 FILLER_18_831 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_fill_1 FILLER_18_859 ();
 sg13g2_decap_4 FILLER_18_864 ();
 sg13g2_fill_2 FILLER_18_873 ();
 sg13g2_decap_8 FILLER_18_879 ();
 sg13g2_decap_8 FILLER_18_886 ();
 sg13g2_fill_1 FILLER_18_893 ();
 sg13g2_decap_4 FILLER_18_898 ();
 sg13g2_decap_4 FILLER_18_906 ();
 sg13g2_fill_2 FILLER_18_910 ();
 sg13g2_fill_1 FILLER_18_955 ();
 sg13g2_fill_2 FILLER_18_977 ();
 sg13g2_fill_1 FILLER_18_979 ();
 sg13g2_fill_1 FILLER_18_984 ();
 sg13g2_decap_4 FILLER_18_989 ();
 sg13g2_fill_2 FILLER_18_993 ();
 sg13g2_fill_1 FILLER_18_1000 ();
 sg13g2_decap_4 FILLER_18_1005 ();
 sg13g2_fill_1 FILLER_18_1009 ();
 sg13g2_fill_1 FILLER_18_1031 ();
 sg13g2_decap_8 FILLER_18_1053 ();
 sg13g2_fill_2 FILLER_18_1060 ();
 sg13g2_fill_2 FILLER_18_1088 ();
 sg13g2_fill_1 FILLER_18_1090 ();
 sg13g2_decap_4 FILLER_18_1133 ();
 sg13g2_fill_2 FILLER_18_1137 ();
 sg13g2_decap_8 FILLER_18_1160 ();
 sg13g2_decap_4 FILLER_18_1167 ();
 sg13g2_fill_1 FILLER_18_1171 ();
 sg13g2_decap_8 FILLER_18_1176 ();
 sg13g2_decap_8 FILLER_18_1183 ();
 sg13g2_fill_1 FILLER_18_1190 ();
 sg13g2_decap_8 FILLER_18_1219 ();
 sg13g2_decap_4 FILLER_18_1226 ();
 sg13g2_fill_1 FILLER_18_1230 ();
 sg13g2_decap_8 FILLER_18_1235 ();
 sg13g2_decap_8 FILLER_18_1246 ();
 sg13g2_decap_8 FILLER_18_1253 ();
 sg13g2_decap_8 FILLER_18_1260 ();
 sg13g2_decap_8 FILLER_18_1267 ();
 sg13g2_decap_4 FILLER_18_1274 ();
 sg13g2_fill_1 FILLER_18_1278 ();
 sg13g2_decap_8 FILLER_18_1331 ();
 sg13g2_decap_8 FILLER_18_1338 ();
 sg13g2_decap_4 FILLER_18_1345 ();
 sg13g2_fill_2 FILLER_18_1357 ();
 sg13g2_decap_8 FILLER_18_1406 ();
 sg13g2_fill_1 FILLER_18_1413 ();
 sg13g2_decap_8 FILLER_18_1418 ();
 sg13g2_decap_8 FILLER_18_1425 ();
 sg13g2_decap_8 FILLER_18_1432 ();
 sg13g2_fill_2 FILLER_18_1439 ();
 sg13g2_fill_1 FILLER_18_1441 ();
 sg13g2_fill_2 FILLER_18_1446 ();
 sg13g2_fill_1 FILLER_18_1448 ();
 sg13g2_fill_2 FILLER_18_1485 ();
 sg13g2_fill_1 FILLER_18_1487 ();
 sg13g2_decap_8 FILLER_18_1535 ();
 sg13g2_decap_8 FILLER_18_1542 ();
 sg13g2_fill_2 FILLER_18_1549 ();
 sg13g2_decap_8 FILLER_18_1571 ();
 sg13g2_decap_8 FILLER_18_1578 ();
 sg13g2_decap_8 FILLER_18_1585 ();
 sg13g2_decap_8 FILLER_18_1592 ();
 sg13g2_fill_1 FILLER_18_1599 ();
 sg13g2_decap_8 FILLER_18_1626 ();
 sg13g2_decap_4 FILLER_18_1654 ();
 sg13g2_fill_2 FILLER_18_1658 ();
 sg13g2_decap_4 FILLER_18_1670 ();
 sg13g2_fill_1 FILLER_18_1674 ();
 sg13g2_decap_8 FILLER_18_1679 ();
 sg13g2_fill_2 FILLER_18_1686 ();
 sg13g2_fill_1 FILLER_18_1688 ();
 sg13g2_decap_4 FILLER_18_1745 ();
 sg13g2_decap_8 FILLER_18_1753 ();
 sg13g2_decap_8 FILLER_18_1760 ();
 sg13g2_decap_8 FILLER_18_1767 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_33 ();
 sg13g2_decap_8 FILLER_19_44 ();
 sg13g2_decap_4 FILLER_19_51 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_decap_4 FILLER_19_66 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_fill_2 FILLER_19_173 ();
 sg13g2_fill_1 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_4 FILLER_19_194 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_decap_4 FILLER_19_237 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_271 ();
 sg13g2_decap_4 FILLER_19_302 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_decap_4 FILLER_19_311 ();
 sg13g2_fill_2 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_4 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_fill_2 FILLER_19_374 ();
 sg13g2_fill_1 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_fill_2 FILLER_19_409 ();
 sg13g2_fill_2 FILLER_19_436 ();
 sg13g2_fill_2 FILLER_19_450 ();
 sg13g2_fill_1 FILLER_19_452 ();
 sg13g2_decap_4 FILLER_19_457 ();
 sg13g2_decap_4 FILLER_19_470 ();
 sg13g2_fill_2 FILLER_19_474 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_fill_1 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_577 ();
 sg13g2_decap_4 FILLER_19_584 ();
 sg13g2_fill_2 FILLER_19_588 ();
 sg13g2_fill_2 FILLER_19_631 ();
 sg13g2_decap_4 FILLER_19_658 ();
 sg13g2_fill_2 FILLER_19_662 ();
 sg13g2_fill_2 FILLER_19_677 ();
 sg13g2_fill_1 FILLER_19_706 ();
 sg13g2_decap_8 FILLER_19_722 ();
 sg13g2_fill_2 FILLER_19_729 ();
 sg13g2_fill_2 FILLER_19_735 ();
 sg13g2_fill_2 FILLER_19_741 ();
 sg13g2_decap_4 FILLER_19_747 ();
 sg13g2_fill_2 FILLER_19_755 ();
 sg13g2_fill_2 FILLER_19_761 ();
 sg13g2_decap_8 FILLER_19_776 ();
 sg13g2_fill_1 FILLER_19_783 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_decap_4 FILLER_19_817 ();
 sg13g2_fill_1 FILLER_19_821 ();
 sg13g2_decap_4 FILLER_19_843 ();
 sg13g2_fill_2 FILLER_19_847 ();
 sg13g2_fill_2 FILLER_19_906 ();
 sg13g2_decap_8 FILLER_19_976 ();
 sg13g2_fill_2 FILLER_19_1009 ();
 sg13g2_decap_8 FILLER_19_1032 ();
 sg13g2_decap_8 FILLER_19_1039 ();
 sg13g2_fill_2 FILLER_19_1051 ();
 sg13g2_decap_4 FILLER_19_1062 ();
 sg13g2_fill_2 FILLER_19_1079 ();
 sg13g2_decap_8 FILLER_19_1097 ();
 sg13g2_fill_1 FILLER_19_1104 ();
 sg13g2_fill_2 FILLER_19_1118 ();
 sg13g2_fill_1 FILLER_19_1120 ();
 sg13g2_decap_8 FILLER_19_1142 ();
 sg13g2_decap_8 FILLER_19_1149 ();
 sg13g2_decap_8 FILLER_19_1156 ();
 sg13g2_fill_2 FILLER_19_1163 ();
 sg13g2_fill_2 FILLER_19_1212 ();
 sg13g2_fill_1 FILLER_19_1214 ();
 sg13g2_decap_8 FILLER_19_1251 ();
 sg13g2_decap_8 FILLER_19_1258 ();
 sg13g2_decap_8 FILLER_19_1265 ();
 sg13g2_decap_8 FILLER_19_1272 ();
 sg13g2_decap_8 FILLER_19_1279 ();
 sg13g2_decap_8 FILLER_19_1286 ();
 sg13g2_decap_8 FILLER_19_1301 ();
 sg13g2_fill_2 FILLER_19_1308 ();
 sg13g2_fill_2 FILLER_19_1322 ();
 sg13g2_fill_2 FILLER_19_1355 ();
 sg13g2_decap_8 FILLER_19_1361 ();
 sg13g2_decap_8 FILLER_19_1394 ();
 sg13g2_decap_8 FILLER_19_1422 ();
 sg13g2_decap_4 FILLER_19_1429 ();
 sg13g2_fill_2 FILLER_19_1460 ();
 sg13g2_decap_8 FILLER_19_1487 ();
 sg13g2_decap_4 FILLER_19_1494 ();
 sg13g2_fill_1 FILLER_19_1498 ();
 sg13g2_decap_8 FILLER_19_1503 ();
 sg13g2_decap_8 FILLER_19_1510 ();
 sg13g2_decap_8 FILLER_19_1517 ();
 sg13g2_decap_8 FILLER_19_1524 ();
 sg13g2_fill_2 FILLER_19_1531 ();
 sg13g2_decap_8 FILLER_19_1594 ();
 sg13g2_decap_8 FILLER_19_1605 ();
 sg13g2_fill_1 FILLER_19_1612 ();
 sg13g2_decap_4 FILLER_19_1639 ();
 sg13g2_fill_1 FILLER_19_1643 ();
 sg13g2_fill_1 FILLER_19_1667 ();
 sg13g2_decap_8 FILLER_19_1715 ();
 sg13g2_decap_8 FILLER_19_1722 ();
 sg13g2_decap_8 FILLER_19_1729 ();
 sg13g2_decap_8 FILLER_19_1736 ();
 sg13g2_decap_8 FILLER_19_1743 ();
 sg13g2_decap_8 FILLER_19_1750 ();
 sg13g2_decap_8 FILLER_19_1757 ();
 sg13g2_decap_8 FILLER_19_1764 ();
 sg13g2_fill_2 FILLER_19_1771 ();
 sg13g2_fill_1 FILLER_19_1773 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_fill_2 FILLER_20_69 ();
 sg13g2_fill_1 FILLER_20_71 ();
 sg13g2_decap_4 FILLER_20_76 ();
 sg13g2_fill_1 FILLER_20_80 ();
 sg13g2_decap_4 FILLER_20_102 ();
 sg13g2_fill_1 FILLER_20_106 ();
 sg13g2_decap_4 FILLER_20_128 ();
 sg13g2_decap_4 FILLER_20_137 ();
 sg13g2_fill_1 FILLER_20_141 ();
 sg13g2_fill_2 FILLER_20_146 ();
 sg13g2_fill_1 FILLER_20_148 ();
 sg13g2_decap_8 FILLER_20_153 ();
 sg13g2_decap_4 FILLER_20_160 ();
 sg13g2_fill_1 FILLER_20_164 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_4 FILLER_20_193 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_207 ();
 sg13g2_fill_1 FILLER_20_209 ();
 sg13g2_fill_2 FILLER_20_222 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_decap_4 FILLER_20_251 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_fill_2 FILLER_20_299 ();
 sg13g2_fill_1 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_306 ();
 sg13g2_decap_4 FILLER_20_313 ();
 sg13g2_fill_2 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_4 FILLER_20_347 ();
 sg13g2_fill_2 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_fill_1 FILLER_20_419 ();
 sg13g2_fill_2 FILLER_20_472 ();
 sg13g2_fill_1 FILLER_20_474 ();
 sg13g2_decap_4 FILLER_20_540 ();
 sg13g2_fill_2 FILLER_20_544 ();
 sg13g2_decap_8 FILLER_20_551 ();
 sg13g2_fill_2 FILLER_20_562 ();
 sg13g2_fill_1 FILLER_20_564 ();
 sg13g2_decap_8 FILLER_20_586 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_fill_2 FILLER_20_609 ();
 sg13g2_fill_1 FILLER_20_611 ();
 sg13g2_fill_2 FILLER_20_616 ();
 sg13g2_fill_1 FILLER_20_618 ();
 sg13g2_fill_2 FILLER_20_705 ();
 sg13g2_decap_4 FILLER_20_711 ();
 sg13g2_fill_1 FILLER_20_754 ();
 sg13g2_fill_1 FILLER_20_759 ();
 sg13g2_decap_4 FILLER_20_764 ();
 sg13g2_fill_1 FILLER_20_768 ();
 sg13g2_fill_1 FILLER_20_773 ();
 sg13g2_fill_2 FILLER_20_807 ();
 sg13g2_decap_8 FILLER_20_817 ();
 sg13g2_decap_8 FILLER_20_824 ();
 sg13g2_fill_2 FILLER_20_831 ();
 sg13g2_fill_2 FILLER_20_859 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_20_865 ();
 sg13g2_decap_8 FILLER_20_872 ();
 sg13g2_decap_4 FILLER_20_884 ();
 sg13g2_fill_1 FILLER_20_888 ();
 sg13g2_decap_4 FILLER_20_918 ();
 sg13g2_fill_2 FILLER_20_922 ();
 sg13g2_decap_8 FILLER_20_932 ();
 sg13g2_decap_8 FILLER_20_939 ();
 sg13g2_decap_8 FILLER_20_946 ();
 sg13g2_decap_8 FILLER_20_953 ();
 sg13g2_decap_8 FILLER_20_960 ();
 sg13g2_decap_8 FILLER_20_967 ();
 sg13g2_decap_8 FILLER_20_974 ();
 sg13g2_decap_8 FILLER_20_981 ();
 sg13g2_fill_2 FILLER_20_988 ();
 sg13g2_fill_1 FILLER_20_990 ();
 sg13g2_decap_8 FILLER_20_995 ();
 sg13g2_decap_8 FILLER_20_1002 ();
 sg13g2_decap_8 FILLER_20_1009 ();
 sg13g2_decap_8 FILLER_20_1016 ();
 sg13g2_fill_1 FILLER_20_1023 ();
 sg13g2_decap_4 FILLER_20_1049 ();
 sg13g2_fill_1 FILLER_20_1053 ();
 sg13g2_fill_2 FILLER_20_1080 ();
 sg13g2_fill_1 FILLER_20_1082 ();
 sg13g2_fill_1 FILLER_20_1087 ();
 sg13g2_decap_8 FILLER_20_1092 ();
 sg13g2_decap_4 FILLER_20_1099 ();
 sg13g2_fill_1 FILLER_20_1103 ();
 sg13g2_decap_8 FILLER_20_1129 ();
 sg13g2_decap_8 FILLER_20_1136 ();
 sg13g2_fill_1 FILLER_20_1143 ();
 sg13g2_fill_2 FILLER_20_1154 ();
 sg13g2_fill_1 FILLER_20_1156 ();
 sg13g2_decap_8 FILLER_20_1167 ();
 sg13g2_fill_1 FILLER_20_1174 ();
 sg13g2_decap_4 FILLER_20_1202 ();
 sg13g2_decap_8 FILLER_20_1242 ();
 sg13g2_decap_8 FILLER_20_1249 ();
 sg13g2_decap_8 FILLER_20_1256 ();
 sg13g2_decap_8 FILLER_20_1263 ();
 sg13g2_decap_8 FILLER_20_1270 ();
 sg13g2_fill_1 FILLER_20_1277 ();
 sg13g2_fill_2 FILLER_20_1304 ();
 sg13g2_decap_4 FILLER_20_1310 ();
 sg13g2_fill_1 FILLER_20_1314 ();
 sg13g2_fill_1 FILLER_20_1320 ();
 sg13g2_fill_1 FILLER_20_1325 ();
 sg13g2_fill_1 FILLER_20_1330 ();
 sg13g2_fill_2 FILLER_20_1350 ();
 sg13g2_fill_2 FILLER_20_1357 ();
 sg13g2_fill_1 FILLER_20_1359 ();
 sg13g2_decap_8 FILLER_20_1365 ();
 sg13g2_decap_4 FILLER_20_1372 ();
 sg13g2_fill_1 FILLER_20_1376 ();
 sg13g2_decap_8 FILLER_20_1415 ();
 sg13g2_decap_8 FILLER_20_1422 ();
 sg13g2_fill_1 FILLER_20_1429 ();
 sg13g2_decap_8 FILLER_20_1513 ();
 sg13g2_decap_8 FILLER_20_1524 ();
 sg13g2_decap_4 FILLER_20_1531 ();
 sg13g2_fill_2 FILLER_20_1535 ();
 sg13g2_fill_1 FILLER_20_1624 ();
 sg13g2_decap_8 FILLER_20_1635 ();
 sg13g2_decap_8 FILLER_20_1642 ();
 sg13g2_fill_2 FILLER_20_1649 ();
 sg13g2_decap_4 FILLER_20_1681 ();
 sg13g2_fill_1 FILLER_20_1685 ();
 sg13g2_fill_2 FILLER_20_1690 ();
 sg13g2_fill_1 FILLER_20_1692 ();
 sg13g2_decap_8 FILLER_20_1754 ();
 sg13g2_decap_8 FILLER_20_1761 ();
 sg13g2_decap_4 FILLER_20_1768 ();
 sg13g2_fill_2 FILLER_20_1772 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_8 ();
 sg13g2_decap_8 FILLER_21_19 ();
 sg13g2_decap_8 FILLER_21_26 ();
 sg13g2_fill_1 FILLER_21_33 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_44 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_fill_2 FILLER_21_78 ();
 sg13g2_fill_1 FILLER_21_148 ();
 sg13g2_decap_8 FILLER_21_170 ();
 sg13g2_fill_1 FILLER_21_177 ();
 sg13g2_decap_4 FILLER_21_207 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_fill_1 FILLER_21_235 ();
 sg13g2_decap_4 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_4 FILLER_21_266 ();
 sg13g2_fill_1 FILLER_21_275 ();
 sg13g2_fill_2 FILLER_21_280 ();
 sg13g2_fill_2 FILLER_21_286 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_4 FILLER_21_326 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_fill_2 FILLER_21_353 ();
 sg13g2_decap_4 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_21_409 ();
 sg13g2_decap_4 FILLER_21_416 ();
 sg13g2_fill_1 FILLER_21_420 ();
 sg13g2_fill_2 FILLER_21_435 ();
 sg13g2_fill_1 FILLER_21_437 ();
 sg13g2_decap_8 FILLER_21_459 ();
 sg13g2_decap_4 FILLER_21_466 ();
 sg13g2_fill_2 FILLER_21_470 ();
 sg13g2_fill_2 FILLER_21_502 ();
 sg13g2_fill_1 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_514 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_4 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_566 ();
 sg13g2_decap_8 FILLER_21_573 ();
 sg13g2_decap_4 FILLER_21_580 ();
 sg13g2_fill_1 FILLER_21_584 ();
 sg13g2_decap_4 FILLER_21_615 ();
 sg13g2_decap_8 FILLER_21_660 ();
 sg13g2_decap_4 FILLER_21_667 ();
 sg13g2_decap_4 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_704 ();
 sg13g2_decap_8 FILLER_21_711 ();
 sg13g2_decap_8 FILLER_21_718 ();
 sg13g2_fill_2 FILLER_21_725 ();
 sg13g2_fill_2 FILLER_21_753 ();
 sg13g2_decap_4 FILLER_21_760 ();
 sg13g2_decap_8 FILLER_21_774 ();
 sg13g2_decap_8 FILLER_21_781 ();
 sg13g2_fill_2 FILLER_21_788 ();
 sg13g2_decap_8 FILLER_21_794 ();
 sg13g2_fill_1 FILLER_21_801 ();
 sg13g2_decap_4 FILLER_21_828 ();
 sg13g2_decap_4 FILLER_21_837 ();
 sg13g2_fill_1 FILLER_21_841 ();
 sg13g2_decap_4 FILLER_21_846 ();
 sg13g2_fill_1 FILLER_21_850 ();
 sg13g2_fill_1 FILLER_21_855 ();
 sg13g2_decap_8 FILLER_21_882 ();
 sg13g2_decap_8 FILLER_21_889 ();
 sg13g2_fill_1 FILLER_21_938 ();
 sg13g2_fill_2 FILLER_21_944 ();
 sg13g2_fill_2 FILLER_21_950 ();
 sg13g2_fill_1 FILLER_21_952 ();
 sg13g2_fill_2 FILLER_21_961 ();
 sg13g2_fill_1 FILLER_21_963 ();
 sg13g2_fill_2 FILLER_21_968 ();
 sg13g2_fill_1 FILLER_21_970 ();
 sg13g2_fill_2 FILLER_21_1013 ();
 sg13g2_fill_1 FILLER_21_1015 ();
 sg13g2_fill_2 FILLER_21_1021 ();
 sg13g2_fill_1 FILLER_21_1023 ();
 sg13g2_decap_8 FILLER_21_1028 ();
 sg13g2_decap_8 FILLER_21_1035 ();
 sg13g2_fill_1 FILLER_21_1042 ();
 sg13g2_fill_1 FILLER_21_1064 ();
 sg13g2_decap_8 FILLER_21_1069 ();
 sg13g2_fill_1 FILLER_21_1076 ();
 sg13g2_decap_4 FILLER_21_1108 ();
 sg13g2_decap_4 FILLER_21_1151 ();
 sg13g2_fill_2 FILLER_21_1215 ();
 sg13g2_decap_4 FILLER_21_1234 ();
 sg13g2_decap_4 FILLER_21_1281 ();
 sg13g2_decap_8 FILLER_21_1289 ();
 sg13g2_decap_8 FILLER_21_1296 ();
 sg13g2_fill_2 FILLER_21_1303 ();
 sg13g2_decap_4 FILLER_21_1314 ();
 sg13g2_fill_1 FILLER_21_1318 ();
 sg13g2_fill_1 FILLER_21_1324 ();
 sg13g2_fill_1 FILLER_21_1329 ();
 sg13g2_fill_1 FILLER_21_1338 ();
 sg13g2_fill_2 FILLER_21_1345 ();
 sg13g2_fill_2 FILLER_21_1352 ();
 sg13g2_fill_2 FILLER_21_1359 ();
 sg13g2_fill_2 FILLER_21_1369 ();
 sg13g2_fill_1 FILLER_21_1397 ();
 sg13g2_decap_8 FILLER_21_1434 ();
 sg13g2_decap_4 FILLER_21_1441 ();
 sg13g2_decap_8 FILLER_21_1455 ();
 sg13g2_decap_8 FILLER_21_1462 ();
 sg13g2_decap_8 FILLER_21_1469 ();
 sg13g2_decap_8 FILLER_21_1476 ();
 sg13g2_fill_2 FILLER_21_1483 ();
 sg13g2_decap_8 FILLER_21_1488 ();
 sg13g2_fill_2 FILLER_21_1495 ();
 sg13g2_fill_1 FILLER_21_1497 ();
 sg13g2_fill_1 FILLER_21_1502 ();
 sg13g2_decap_8 FILLER_21_1539 ();
 sg13g2_decap_8 FILLER_21_1546 ();
 sg13g2_decap_8 FILLER_21_1553 ();
 sg13g2_decap_8 FILLER_21_1560 ();
 sg13g2_decap_8 FILLER_21_1567 ();
 sg13g2_decap_8 FILLER_21_1574 ();
 sg13g2_decap_8 FILLER_21_1581 ();
 sg13g2_fill_2 FILLER_21_1588 ();
 sg13g2_decap_8 FILLER_21_1626 ();
 sg13g2_decap_8 FILLER_21_1633 ();
 sg13g2_decap_8 FILLER_21_1640 ();
 sg13g2_decap_4 FILLER_21_1647 ();
 sg13g2_fill_2 FILLER_21_1651 ();
 sg13g2_decap_8 FILLER_21_1663 ();
 sg13g2_decap_4 FILLER_21_1670 ();
 sg13g2_fill_2 FILLER_21_1674 ();
 sg13g2_decap_8 FILLER_21_1697 ();
 sg13g2_fill_1 FILLER_21_1704 ();
 sg13g2_fill_1 FILLER_21_1715 ();
 sg13g2_decap_8 FILLER_21_1742 ();
 sg13g2_decap_8 FILLER_21_1749 ();
 sg13g2_decap_8 FILLER_21_1756 ();
 sg13g2_decap_8 FILLER_21_1763 ();
 sg13g2_decap_4 FILLER_21_1770 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_fill_1 FILLER_22_37 ();
 sg13g2_fill_2 FILLER_22_64 ();
 sg13g2_decap_8 FILLER_22_87 ();
 sg13g2_decap_8 FILLER_22_94 ();
 sg13g2_fill_2 FILLER_22_101 ();
 sg13g2_decap_4 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_132 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_4 FILLER_22_144 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_2 FILLER_22_170 ();
 sg13g2_decap_4 FILLER_22_197 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_fill_1 FILLER_22_211 ();
 sg13g2_decap_4 FILLER_22_233 ();
 sg13g2_fill_2 FILLER_22_237 ();
 sg13g2_decap_4 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_fill_2 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_368 ();
 sg13g2_decap_4 FILLER_22_399 ();
 sg13g2_fill_1 FILLER_22_403 ();
 sg13g2_fill_1 FILLER_22_455 ();
 sg13g2_fill_2 FILLER_22_477 ();
 sg13g2_fill_1 FILLER_22_479 ();
 sg13g2_decap_4 FILLER_22_483 ();
 sg13g2_fill_1 FILLER_22_500 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_fill_1 FILLER_22_592 ();
 sg13g2_decap_8 FILLER_22_597 ();
 sg13g2_fill_2 FILLER_22_604 ();
 sg13g2_decap_4 FILLER_22_646 ();
 sg13g2_fill_2 FILLER_22_650 ();
 sg13g2_decap_4 FILLER_22_673 ();
 sg13g2_fill_1 FILLER_22_677 ();
 sg13g2_fill_2 FILLER_22_762 ();
 sg13g2_decap_8 FILLER_22_794 ();
 sg13g2_decap_8 FILLER_22_822 ();
 sg13g2_decap_8 FILLER_22_829 ();
 sg13g2_fill_2 FILLER_22_836 ();
 sg13g2_fill_2 FILLER_22_843 ();
 sg13g2_fill_1 FILLER_22_845 ();
 sg13g2_fill_1 FILLER_22_862 ();
 sg13g2_fill_2 FILLER_22_889 ();
 sg13g2_fill_1 FILLER_22_891 ();
 sg13g2_fill_1 FILLER_22_897 ();
 sg13g2_decap_8 FILLER_22_902 ();
 sg13g2_decap_8 FILLER_22_909 ();
 sg13g2_decap_8 FILLER_22_916 ();
 sg13g2_decap_8 FILLER_22_923 ();
 sg13g2_decap_8 FILLER_22_930 ();
 sg13g2_fill_2 FILLER_22_937 ();
 sg13g2_fill_1 FILLER_22_939 ();
 sg13g2_decap_4 FILLER_22_966 ();
 sg13g2_fill_1 FILLER_22_970 ();
 sg13g2_decap_8 FILLER_22_992 ();
 sg13g2_decap_8 FILLER_22_999 ();
 sg13g2_decap_8 FILLER_22_1006 ();
 sg13g2_fill_1 FILLER_22_1064 ();
 sg13g2_decap_8 FILLER_22_1086 ();
 sg13g2_fill_2 FILLER_22_1093 ();
 sg13g2_decap_4 FILLER_22_1104 ();
 sg13g2_fill_1 FILLER_22_1108 ();
 sg13g2_decap_8 FILLER_22_1144 ();
 sg13g2_decap_8 FILLER_22_1151 ();
 sg13g2_fill_2 FILLER_22_1158 ();
 sg13g2_decap_8 FILLER_22_1164 ();
 sg13g2_decap_4 FILLER_22_1171 ();
 sg13g2_fill_1 FILLER_22_1205 ();
 sg13g2_fill_2 FILLER_22_1211 ();
 sg13g2_decap_8 FILLER_22_1223 ();
 sg13g2_fill_2 FILLER_22_1230 ();
 sg13g2_fill_1 FILLER_22_1232 ();
 sg13g2_decap_4 FILLER_22_1259 ();
 sg13g2_decap_8 FILLER_22_1267 ();
 sg13g2_decap_8 FILLER_22_1274 ();
 sg13g2_decap_4 FILLER_22_1281 ();
 sg13g2_decap_8 FILLER_22_1289 ();
 sg13g2_decap_8 FILLER_22_1296 ();
 sg13g2_decap_4 FILLER_22_1303 ();
 sg13g2_fill_1 FILLER_22_1307 ();
 sg13g2_fill_1 FILLER_22_1320 ();
 sg13g2_fill_1 FILLER_22_1326 ();
 sg13g2_fill_2 FILLER_22_1336 ();
 sg13g2_fill_2 FILLER_22_1354 ();
 sg13g2_fill_1 FILLER_22_1356 ();
 sg13g2_decap_8 FILLER_22_1362 ();
 sg13g2_decap_8 FILLER_22_1369 ();
 sg13g2_fill_1 FILLER_22_1376 ();
 sg13g2_fill_1 FILLER_22_1381 ();
 sg13g2_decap_8 FILLER_22_1400 ();
 sg13g2_decap_4 FILLER_22_1407 ();
 sg13g2_fill_1 FILLER_22_1415 ();
 sg13g2_decap_4 FILLER_22_1420 ();
 sg13g2_fill_2 FILLER_22_1424 ();
 sg13g2_fill_1 FILLER_22_1452 ();
 sg13g2_decap_8 FILLER_22_1478 ();
 sg13g2_decap_8 FILLER_22_1485 ();
 sg13g2_decap_8 FILLER_22_1518 ();
 sg13g2_decap_8 FILLER_22_1525 ();
 sg13g2_decap_8 FILLER_22_1532 ();
 sg13g2_decap_8 FILLER_22_1539 ();
 sg13g2_decap_4 FILLER_22_1603 ();
 sg13g2_decap_8 FILLER_22_1611 ();
 sg13g2_fill_2 FILLER_22_1618 ();
 sg13g2_decap_8 FILLER_22_1686 ();
 sg13g2_decap_8 FILLER_22_1693 ();
 sg13g2_decap_8 FILLER_22_1700 ();
 sg13g2_decap_8 FILLER_22_1707 ();
 sg13g2_decap_4 FILLER_22_1714 ();
 sg13g2_fill_2 FILLER_22_1718 ();
 sg13g2_decap_8 FILLER_22_1728 ();
 sg13g2_decap_8 FILLER_22_1735 ();
 sg13g2_decap_8 FILLER_22_1742 ();
 sg13g2_decap_8 FILLER_22_1749 ();
 sg13g2_decap_8 FILLER_22_1756 ();
 sg13g2_decap_8 FILLER_22_1763 ();
 sg13g2_decap_4 FILLER_22_1770 ();
 sg13g2_fill_2 FILLER_23_31 ();
 sg13g2_fill_2 FILLER_23_37 ();
 sg13g2_fill_1 FILLER_23_39 ();
 sg13g2_fill_2 FILLER_23_44 ();
 sg13g2_fill_1 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_85 ();
 sg13g2_decap_4 FILLER_23_92 ();
 sg13g2_decap_4 FILLER_23_117 ();
 sg13g2_fill_1 FILLER_23_121 ();
 sg13g2_decap_8 FILLER_23_127 ();
 sg13g2_decap_4 FILLER_23_134 ();
 sg13g2_decap_8 FILLER_23_142 ();
 sg13g2_decap_8 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_156 ();
 sg13g2_decap_4 FILLER_23_163 ();
 sg13g2_fill_2 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_173 ();
 sg13g2_decap_8 FILLER_23_180 ();
 sg13g2_decap_8 FILLER_23_187 ();
 sg13g2_decap_4 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_198 ();
 sg13g2_decap_8 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_240 ();
 sg13g2_decap_8 FILLER_23_247 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_265 ();
 sg13g2_decap_4 FILLER_23_280 ();
 sg13g2_decap_4 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_318 ();
 sg13g2_decap_4 FILLER_23_340 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_fill_1 FILLER_23_391 ();
 sg13g2_fill_2 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_23_422 ();
 sg13g2_fill_2 FILLER_23_429 ();
 sg13g2_fill_2 FILLER_23_488 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_fill_2 FILLER_23_518 ();
 sg13g2_fill_2 FILLER_23_541 ();
 sg13g2_fill_2 FILLER_23_564 ();
 sg13g2_fill_1 FILLER_23_566 ();
 sg13g2_fill_2 FILLER_23_598 ();
 sg13g2_fill_1 FILLER_23_600 ();
 sg13g2_fill_2 FILLER_23_622 ();
 sg13g2_decap_4 FILLER_23_642 ();
 sg13g2_decap_8 FILLER_23_670 ();
 sg13g2_decap_8 FILLER_23_677 ();
 sg13g2_fill_2 FILLER_23_684 ();
 sg13g2_fill_2 FILLER_23_689 ();
 sg13g2_fill_1 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_755 ();
 sg13g2_fill_2 FILLER_23_762 ();
 sg13g2_fill_1 FILLER_23_764 ();
 sg13g2_fill_2 FILLER_23_775 ();
 sg13g2_fill_1 FILLER_23_777 ();
 sg13g2_decap_4 FILLER_23_782 ();
 sg13g2_fill_2 FILLER_23_786 ();
 sg13g2_fill_2 FILLER_23_809 ();
 sg13g2_fill_1 FILLER_23_811 ();
 sg13g2_fill_2 FILLER_23_865 ();
 sg13g2_fill_2 FILLER_23_891 ();
 sg13g2_decap_8 FILLER_23_919 ();
 sg13g2_fill_2 FILLER_23_926 ();
 sg13g2_fill_1 FILLER_23_928 ();
 sg13g2_decap_8 FILLER_23_955 ();
 sg13g2_decap_8 FILLER_23_962 ();
 sg13g2_fill_2 FILLER_23_973 ();
 sg13g2_decap_8 FILLER_23_979 ();
 sg13g2_decap_8 FILLER_23_986 ();
 sg13g2_fill_2 FILLER_23_993 ();
 sg13g2_fill_1 FILLER_23_995 ();
 sg13g2_decap_8 FILLER_23_1017 ();
 sg13g2_decap_8 FILLER_23_1024 ();
 sg13g2_decap_4 FILLER_23_1031 ();
 sg13g2_decap_8 FILLER_23_1052 ();
 sg13g2_decap_8 FILLER_23_1059 ();
 sg13g2_fill_2 FILLER_23_1066 ();
 sg13g2_fill_1 FILLER_23_1068 ();
 sg13g2_decap_4 FILLER_23_1132 ();
 sg13g2_fill_2 FILLER_23_1136 ();
 sg13g2_fill_1 FILLER_23_1177 ();
 sg13g2_fill_2 FILLER_23_1187 ();
 sg13g2_fill_1 FILLER_23_1277 ();
 sg13g2_fill_1 FILLER_23_1316 ();
 sg13g2_decap_4 FILLER_23_1321 ();
 sg13g2_decap_4 FILLER_23_1337 ();
 sg13g2_fill_1 FILLER_23_1341 ();
 sg13g2_fill_2 FILLER_23_1346 ();
 sg13g2_fill_1 FILLER_23_1348 ();
 sg13g2_decap_8 FILLER_23_1375 ();
 sg13g2_decap_8 FILLER_23_1382 ();
 sg13g2_decap_4 FILLER_23_1389 ();
 sg13g2_fill_1 FILLER_23_1393 ();
 sg13g2_decap_4 FILLER_23_1430 ();
 sg13g2_decap_8 FILLER_23_1438 ();
 sg13g2_decap_8 FILLER_23_1445 ();
 sg13g2_decap_4 FILLER_23_1452 ();
 sg13g2_fill_1 FILLER_23_1456 ();
 sg13g2_decap_8 FILLER_23_1493 ();
 sg13g2_decap_4 FILLER_23_1514 ();
 sg13g2_fill_2 FILLER_23_1518 ();
 sg13g2_fill_2 FILLER_23_1560 ();
 sg13g2_fill_1 FILLER_23_1562 ();
 sg13g2_decap_8 FILLER_23_1567 ();
 sg13g2_decap_8 FILLER_23_1574 ();
 sg13g2_decap_8 FILLER_23_1581 ();
 sg13g2_fill_1 FILLER_23_1588 ();
 sg13g2_decap_4 FILLER_23_1625 ();
 sg13g2_fill_1 FILLER_23_1629 ();
 sg13g2_decap_8 FILLER_23_1643 ();
 sg13g2_decap_8 FILLER_23_1650 ();
 sg13g2_decap_8 FILLER_23_1657 ();
 sg13g2_decap_4 FILLER_23_1664 ();
 sg13g2_decap_8 FILLER_23_1672 ();
 sg13g2_decap_8 FILLER_23_1679 ();
 sg13g2_decap_8 FILLER_23_1686 ();
 sg13g2_decap_8 FILLER_23_1693 ();
 sg13g2_fill_2 FILLER_23_1700 ();
 sg13g2_fill_1 FILLER_23_1702 ();
 sg13g2_fill_1 FILLER_23_1713 ();
 sg13g2_decap_8 FILLER_23_1740 ();
 sg13g2_decap_8 FILLER_23_1747 ();
 sg13g2_decap_8 FILLER_23_1754 ();
 sg13g2_decap_8 FILLER_23_1761 ();
 sg13g2_decap_4 FILLER_23_1768 ();
 sg13g2_fill_2 FILLER_23_1772 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_fill_2 FILLER_24_25 ();
 sg13g2_decap_4 FILLER_24_32 ();
 sg13g2_fill_1 FILLER_24_36 ();
 sg13g2_decap_8 FILLER_24_41 ();
 sg13g2_fill_2 FILLER_24_48 ();
 sg13g2_fill_1 FILLER_24_50 ();
 sg13g2_decap_8 FILLER_24_64 ();
 sg13g2_decap_8 FILLER_24_71 ();
 sg13g2_decap_8 FILLER_24_78 ();
 sg13g2_decap_8 FILLER_24_85 ();
 sg13g2_decap_8 FILLER_24_92 ();
 sg13g2_decap_8 FILLER_24_99 ();
 sg13g2_decap_8 FILLER_24_106 ();
 sg13g2_decap_8 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_157 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_decap_8 FILLER_24_255 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_decap_4 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_324 ();
 sg13g2_decap_4 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_351 ();
 sg13g2_fill_1 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_381 ();
 sg13g2_fill_2 FILLER_24_404 ();
 sg13g2_decap_4 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_4 FILLER_24_434 ();
 sg13g2_fill_1 FILLER_24_438 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_decap_8 FILLER_24_459 ();
 sg13g2_decap_8 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_473 ();
 sg13g2_fill_2 FILLER_24_480 ();
 sg13g2_fill_1 FILLER_24_482 ();
 sg13g2_decap_4 FILLER_24_509 ();
 sg13g2_fill_2 FILLER_24_513 ();
 sg13g2_fill_2 FILLER_24_519 ();
 sg13g2_fill_2 FILLER_24_542 ();
 sg13g2_decap_4 FILLER_24_565 ();
 sg13g2_fill_1 FILLER_24_573 ();
 sg13g2_decap_8 FILLER_24_578 ();
 sg13g2_decap_8 FILLER_24_585 ();
 sg13g2_fill_2 FILLER_24_622 ();
 sg13g2_decap_8 FILLER_24_648 ();
 sg13g2_fill_1 FILLER_24_655 ();
 sg13g2_fill_1 FILLER_24_695 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_fill_1 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_760 ();
 sg13g2_fill_1 FILLER_24_767 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_fill_1 FILLER_24_812 ();
 sg13g2_fill_2 FILLER_24_834 ();
 sg13g2_fill_1 FILLER_24_836 ();
 sg13g2_fill_2 FILLER_24_846 ();
 sg13g2_fill_1 FILLER_24_873 ();
 sg13g2_decap_4 FILLER_24_895 ();
 sg13g2_fill_1 FILLER_24_899 ();
 sg13g2_fill_2 FILLER_24_904 ();
 sg13g2_fill_2 FILLER_24_927 ();
 sg13g2_fill_1 FILLER_24_929 ();
 sg13g2_fill_2 FILLER_24_935 ();
 sg13g2_decap_4 FILLER_24_941 ();
 sg13g2_fill_1 FILLER_24_945 ();
 sg13g2_decap_4 FILLER_24_950 ();
 sg13g2_fill_1 FILLER_24_954 ();
 sg13g2_fill_2 FILLER_24_986 ();
 sg13g2_fill_1 FILLER_24_988 ();
 sg13g2_fill_1 FILLER_24_1020 ();
 sg13g2_decap_8 FILLER_24_1052 ();
 sg13g2_decap_8 FILLER_24_1059 ();
 sg13g2_decap_8 FILLER_24_1066 ();
 sg13g2_decap_4 FILLER_24_1073 ();
 sg13g2_fill_1 FILLER_24_1077 ();
 sg13g2_decap_8 FILLER_24_1083 ();
 sg13g2_fill_2 FILLER_24_1090 ();
 sg13g2_fill_1 FILLER_24_1096 ();
 sg13g2_decap_8 FILLER_24_1101 ();
 sg13g2_decap_8 FILLER_24_1108 ();
 sg13g2_decap_8 FILLER_24_1115 ();
 sg13g2_decap_8 FILLER_24_1122 ();
 sg13g2_decap_4 FILLER_24_1129 ();
 sg13g2_decap_8 FILLER_24_1143 ();
 sg13g2_decap_8 FILLER_24_1150 ();
 sg13g2_decap_8 FILLER_24_1157 ();
 sg13g2_decap_4 FILLER_24_1168 ();
 sg13g2_fill_2 FILLER_24_1172 ();
 sg13g2_decap_8 FILLER_24_1219 ();
 sg13g2_fill_2 FILLER_24_1226 ();
 sg13g2_decap_8 FILLER_24_1232 ();
 sg13g2_decap_8 FILLER_24_1239 ();
 sg13g2_decap_8 FILLER_24_1246 ();
 sg13g2_decap_8 FILLER_24_1253 ();
 sg13g2_decap_8 FILLER_24_1264 ();
 sg13g2_fill_1 FILLER_24_1271 ();
 sg13g2_fill_1 FILLER_24_1310 ();
 sg13g2_fill_2 FILLER_24_1350 ();
 sg13g2_decap_4 FILLER_24_1362 ();
 sg13g2_fill_1 FILLER_24_1366 ();
 sg13g2_fill_1 FILLER_24_1393 ();
 sg13g2_decap_8 FILLER_24_1430 ();
 sg13g2_fill_1 FILLER_24_1437 ();
 sg13g2_decap_4 FILLER_24_1442 ();
 sg13g2_decap_4 FILLER_24_1456 ();
 sg13g2_decap_8 FILLER_24_1487 ();
 sg13g2_fill_2 FILLER_24_1494 ();
 sg13g2_fill_1 FILLER_24_1510 ();
 sg13g2_decap_4 FILLER_24_1532 ();
 sg13g2_decap_8 FILLER_24_1540 ();
 sg13g2_decap_8 FILLER_24_1547 ();
 sg13g2_decap_8 FILLER_24_1554 ();
 sg13g2_decap_8 FILLER_24_1561 ();
 sg13g2_decap_4 FILLER_24_1568 ();
 sg13g2_fill_1 FILLER_24_1572 ();
 sg13g2_fill_2 FILLER_24_1583 ();
 sg13g2_fill_2 FILLER_24_1595 ();
 sg13g2_fill_1 FILLER_24_1597 ();
 sg13g2_fill_2 FILLER_24_1602 ();
 sg13g2_fill_1 FILLER_24_1604 ();
 sg13g2_decap_4 FILLER_24_1609 ();
 sg13g2_fill_2 FILLER_24_1613 ();
 sg13g2_fill_2 FILLER_24_1636 ();
 sg13g2_fill_1 FILLER_24_1638 ();
 sg13g2_decap_4 FILLER_24_1643 ();
 sg13g2_fill_2 FILLER_24_1647 ();
 sg13g2_decap_8 FILLER_24_1659 ();
 sg13g2_decap_8 FILLER_24_1666 ();
 sg13g2_fill_1 FILLER_24_1673 ();
 sg13g2_decap_8 FILLER_24_1721 ();
 sg13g2_decap_8 FILLER_24_1728 ();
 sg13g2_decap_8 FILLER_24_1735 ();
 sg13g2_decap_8 FILLER_24_1742 ();
 sg13g2_decap_8 FILLER_24_1749 ();
 sg13g2_decap_8 FILLER_24_1756 ();
 sg13g2_decap_8 FILLER_24_1763 ();
 sg13g2_decap_4 FILLER_24_1770 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_27 ();
 sg13g2_fill_1 FILLER_25_32 ();
 sg13g2_fill_2 FILLER_25_59 ();
 sg13g2_decap_8 FILLER_25_82 ();
 sg13g2_decap_4 FILLER_25_89 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_decap_4 FILLER_25_115 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_decap_8 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_177 ();
 sg13g2_decap_4 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_decap_4 FILLER_25_215 ();
 sg13g2_fill_2 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_230 ();
 sg13g2_decap_8 FILLER_25_237 ();
 sg13g2_decap_8 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_283 ();
 sg13g2_decap_8 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_fill_1 FILLER_25_307 ();
 sg13g2_fill_1 FILLER_25_313 ();
 sg13g2_fill_2 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_4 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_fill_1 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_426 ();
 sg13g2_decap_4 FILLER_25_433 ();
 sg13g2_fill_1 FILLER_25_437 ();
 sg13g2_decap_8 FILLER_25_464 ();
 sg13g2_decap_8 FILLER_25_471 ();
 sg13g2_decap_8 FILLER_25_478 ();
 sg13g2_fill_2 FILLER_25_485 ();
 sg13g2_fill_1 FILLER_25_487 ();
 sg13g2_decap_8 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_decap_4 FILLER_25_543 ();
 sg13g2_fill_1 FILLER_25_547 ();
 sg13g2_fill_2 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_fill_1 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_572 ();
 sg13g2_decap_4 FILLER_25_579 ();
 sg13g2_decap_8 FILLER_25_643 ();
 sg13g2_decap_4 FILLER_25_650 ();
 sg13g2_fill_2 FILLER_25_654 ();
 sg13g2_decap_8 FILLER_25_661 ();
 sg13g2_decap_4 FILLER_25_668 ();
 sg13g2_fill_2 FILLER_25_672 ();
 sg13g2_fill_1 FILLER_25_687 ();
 sg13g2_decap_8 FILLER_25_696 ();
 sg13g2_fill_2 FILLER_25_703 ();
 sg13g2_decap_8 FILLER_25_715 ();
 sg13g2_fill_2 FILLER_25_722 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_fill_2 FILLER_25_750 ();
 sg13g2_fill_2 FILLER_25_760 ();
 sg13g2_fill_1 FILLER_25_762 ();
 sg13g2_fill_2 FILLER_25_767 ();
 sg13g2_decap_8 FILLER_25_773 ();
 sg13g2_decap_8 FILLER_25_780 ();
 sg13g2_fill_1 FILLER_25_787 ();
 sg13g2_decap_8 FILLER_25_824 ();
 sg13g2_fill_1 FILLER_25_835 ();
 sg13g2_fill_1 FILLER_25_865 ();
 sg13g2_decap_4 FILLER_25_874 ();
 sg13g2_fill_2 FILLER_25_878 ();
 sg13g2_decap_8 FILLER_25_913 ();
 sg13g2_decap_4 FILLER_25_920 ();
 sg13g2_fill_2 FILLER_25_924 ();
 sg13g2_decap_8 FILLER_25_952 ();
 sg13g2_decap_4 FILLER_25_959 ();
 sg13g2_fill_2 FILLER_25_963 ();
 sg13g2_decap_8 FILLER_25_970 ();
 sg13g2_decap_8 FILLER_25_981 ();
 sg13g2_decap_4 FILLER_25_988 ();
 sg13g2_fill_2 FILLER_25_997 ();
 sg13g2_fill_1 FILLER_25_999 ();
 sg13g2_fill_2 FILLER_25_1004 ();
 sg13g2_fill_2 FILLER_25_1010 ();
 sg13g2_fill_2 FILLER_25_1016 ();
 sg13g2_fill_2 FILLER_25_1039 ();
 sg13g2_fill_1 FILLER_25_1041 ();
 sg13g2_fill_1 FILLER_25_1046 ();
 sg13g2_fill_2 FILLER_25_1073 ();
 sg13g2_fill_1 FILLER_25_1075 ();
 sg13g2_fill_2 FILLER_25_1127 ();
 sg13g2_fill_1 FILLER_25_1129 ();
 sg13g2_decap_8 FILLER_25_1169 ();
 sg13g2_decap_4 FILLER_25_1176 ();
 sg13g2_fill_2 FILLER_25_1180 ();
 sg13g2_decap_8 FILLER_25_1218 ();
 sg13g2_fill_2 FILLER_25_1225 ();
 sg13g2_fill_1 FILLER_25_1227 ();
 sg13g2_decap_8 FILLER_25_1232 ();
 sg13g2_fill_2 FILLER_25_1239 ();
 sg13g2_fill_1 FILLER_25_1241 ();
 sg13g2_decap_4 FILLER_25_1268 ();
 sg13g2_fill_1 FILLER_25_1280 ();
 sg13g2_decap_4 FILLER_25_1285 ();
 sg13g2_fill_2 FILLER_25_1293 ();
 sg13g2_fill_2 FILLER_25_1299 ();
 sg13g2_fill_1 FILLER_25_1301 ();
 sg13g2_decap_4 FILLER_25_1310 ();
 sg13g2_decap_8 FILLER_25_1319 ();
 sg13g2_fill_2 FILLER_25_1330 ();
 sg13g2_fill_1 FILLER_25_1332 ();
 sg13g2_decap_8 FILLER_25_1337 ();
 sg13g2_fill_1 FILLER_25_1348 ();
 sg13g2_decap_8 FILLER_25_1387 ();
 sg13g2_decap_4 FILLER_25_1404 ();
 sg13g2_decap_8 FILLER_25_1412 ();
 sg13g2_decap_8 FILLER_25_1419 ();
 sg13g2_decap_4 FILLER_25_1426 ();
 sg13g2_fill_1 FILLER_25_1430 ();
 sg13g2_decap_4 FILLER_25_1457 ();
 sg13g2_fill_2 FILLER_25_1461 ();
 sg13g2_decap_8 FILLER_25_1515 ();
 sg13g2_fill_2 FILLER_25_1522 ();
 sg13g2_fill_1 FILLER_25_1524 ();
 sg13g2_fill_2 FILLER_25_1535 ();
 sg13g2_fill_2 FILLER_25_1563 ();
 sg13g2_fill_1 FILLER_25_1565 ();
 sg13g2_fill_1 FILLER_25_1592 ();
 sg13g2_fill_2 FILLER_25_1619 ();
 sg13g2_fill_1 FILLER_25_1621 ();
 sg13g2_decap_4 FILLER_25_1708 ();
 sg13g2_fill_1 FILLER_25_1712 ();
 sg13g2_decap_8 FILLER_25_1739 ();
 sg13g2_decap_8 FILLER_25_1746 ();
 sg13g2_decap_8 FILLER_25_1753 ();
 sg13g2_decap_8 FILLER_25_1760 ();
 sg13g2_decap_8 FILLER_25_1767 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_7 ();
 sg13g2_decap_4 FILLER_26_12 ();
 sg13g2_fill_2 FILLER_26_16 ();
 sg13g2_fill_1 FILLER_26_23 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_decap_4 FILLER_26_39 ();
 sg13g2_fill_2 FILLER_26_43 ();
 sg13g2_fill_2 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_fill_2 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_58 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_fill_2 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_194 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_fill_2 FILLER_26_307 ();
 sg13g2_fill_2 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_fill_2 FILLER_26_403 ();
 sg13g2_fill_1 FILLER_26_405 ();
 sg13g2_fill_2 FILLER_26_419 ();
 sg13g2_decap_4 FILLER_26_430 ();
 sg13g2_fill_1 FILLER_26_434 ();
 sg13g2_fill_2 FILLER_26_440 ();
 sg13g2_fill_1 FILLER_26_442 ();
 sg13g2_fill_2 FILLER_26_464 ();
 sg13g2_decap_8 FILLER_26_496 ();
 sg13g2_fill_1 FILLER_26_503 ();
 sg13g2_decap_8 FILLER_26_523 ();
 sg13g2_fill_2 FILLER_26_556 ();
 sg13g2_fill_2 FILLER_26_563 ();
 sg13g2_decap_8 FILLER_26_573 ();
 sg13g2_decap_4 FILLER_26_580 ();
 sg13g2_fill_1 FILLER_26_589 ();
 sg13g2_fill_2 FILLER_26_603 ();
 sg13g2_fill_1 FILLER_26_605 ();
 sg13g2_fill_2 FILLER_26_611 ();
 sg13g2_fill_1 FILLER_26_613 ();
 sg13g2_fill_2 FILLER_26_639 ();
 sg13g2_fill_1 FILLER_26_641 ();
 sg13g2_fill_2 FILLER_26_647 ();
 sg13g2_fill_1 FILLER_26_649 ();
 sg13g2_fill_2 FILLER_26_654 ();
 sg13g2_fill_1 FILLER_26_664 ();
 sg13g2_fill_2 FILLER_26_704 ();
 sg13g2_fill_1 FILLER_26_706 ();
 sg13g2_fill_1 FILLER_26_744 ();
 sg13g2_fill_2 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_764 ();
 sg13g2_decap_8 FILLER_26_771 ();
 sg13g2_fill_2 FILLER_26_778 ();
 sg13g2_fill_1 FILLER_26_780 ();
 sg13g2_decap_8 FILLER_26_785 ();
 sg13g2_decap_8 FILLER_26_792 ();
 sg13g2_fill_1 FILLER_26_799 ();
 sg13g2_fill_2 FILLER_26_805 ();
 sg13g2_fill_1 FILLER_26_807 ();
 sg13g2_fill_2 FILLER_26_843 ();
 sg13g2_fill_2 FILLER_26_866 ();
 sg13g2_decap_8 FILLER_26_915 ();
 sg13g2_fill_2 FILLER_26_922 ();
 sg13g2_fill_2 FILLER_26_929 ();
 sg13g2_fill_1 FILLER_26_931 ();
 sg13g2_fill_1 FILLER_26_965 ();
 sg13g2_fill_1 FILLER_26_992 ();
 sg13g2_fill_1 FILLER_26_1040 ();
 sg13g2_fill_2 FILLER_26_1050 ();
 sg13g2_fill_1 FILLER_26_1052 ();
 sg13g2_fill_2 FILLER_26_1057 ();
 sg13g2_fill_2 FILLER_26_1080 ();
 sg13g2_decap_8 FILLER_26_1094 ();
 sg13g2_decap_8 FILLER_26_1101 ();
 sg13g2_fill_2 FILLER_26_1108 ();
 sg13g2_decap_8 FILLER_26_1131 ();
 sg13g2_decap_8 FILLER_26_1138 ();
 sg13g2_decap_4 FILLER_26_1145 ();
 sg13g2_fill_1 FILLER_26_1149 ();
 sg13g2_decap_4 FILLER_26_1154 ();
 sg13g2_fill_2 FILLER_26_1158 ();
 sg13g2_decap_8 FILLER_26_1164 ();
 sg13g2_decap_4 FILLER_26_1171 ();
 sg13g2_fill_1 FILLER_26_1175 ();
 sg13g2_fill_2 FILLER_26_1209 ();
 sg13g2_decap_4 FILLER_26_1245 ();
 sg13g2_decap_8 FILLER_26_1257 ();
 sg13g2_decap_8 FILLER_26_1264 ();
 sg13g2_fill_1 FILLER_26_1271 ();
 sg13g2_decap_8 FILLER_26_1278 ();
 sg13g2_decap_4 FILLER_26_1285 ();
 sg13g2_decap_8 FILLER_26_1315 ();
 sg13g2_decap_4 FILLER_26_1322 ();
 sg13g2_fill_1 FILLER_26_1326 ();
 sg13g2_decap_8 FILLER_26_1331 ();
 sg13g2_decap_8 FILLER_26_1364 ();
 sg13g2_decap_8 FILLER_26_1371 ();
 sg13g2_decap_4 FILLER_26_1378 ();
 sg13g2_decap_8 FILLER_26_1386 ();
 sg13g2_decap_4 FILLER_26_1393 ();
 sg13g2_fill_1 FILLER_26_1397 ();
 sg13g2_fill_2 FILLER_26_1428 ();
 sg13g2_fill_1 FILLER_26_1430 ();
 sg13g2_decap_8 FILLER_26_1435 ();
 sg13g2_decap_8 FILLER_26_1442 ();
 sg13g2_decap_8 FILLER_26_1449 ();
 sg13g2_decap_8 FILLER_26_1456 ();
 sg13g2_decap_4 FILLER_26_1463 ();
 sg13g2_fill_1 FILLER_26_1467 ();
 sg13g2_decap_4 FILLER_26_1472 ();
 sg13g2_fill_2 FILLER_26_1476 ();
 sg13g2_decap_8 FILLER_26_1488 ();
 sg13g2_decap_8 FILLER_26_1495 ();
 sg13g2_decap_4 FILLER_26_1502 ();
 sg13g2_decap_8 FILLER_26_1511 ();
 sg13g2_decap_4 FILLER_26_1522 ();
 sg13g2_fill_1 FILLER_26_1526 ();
 sg13g2_decap_8 FILLER_26_1532 ();
 sg13g2_fill_2 FILLER_26_1539 ();
 sg13g2_decap_8 FILLER_26_1558 ();
 sg13g2_decap_8 FILLER_26_1565 ();
 sg13g2_decap_8 FILLER_26_1576 ();
 sg13g2_decap_8 FILLER_26_1583 ();
 sg13g2_fill_2 FILLER_26_1590 ();
 sg13g2_decap_8 FILLER_26_1628 ();
 sg13g2_decap_8 FILLER_26_1635 ();
 sg13g2_decap_8 FILLER_26_1642 ();
 sg13g2_decap_4 FILLER_26_1649 ();
 sg13g2_fill_2 FILLER_26_1663 ();
 sg13g2_fill_1 FILLER_26_1665 ();
 sg13g2_decap_8 FILLER_26_1670 ();
 sg13g2_fill_2 FILLER_26_1677 ();
 sg13g2_fill_1 FILLER_26_1679 ();
 sg13g2_decap_8 FILLER_26_1693 ();
 sg13g2_fill_2 FILLER_26_1700 ();
 sg13g2_fill_1 FILLER_26_1702 ();
 sg13g2_decap_8 FILLER_26_1713 ();
 sg13g2_decap_8 FILLER_26_1724 ();
 sg13g2_decap_8 FILLER_26_1731 ();
 sg13g2_decap_8 FILLER_26_1738 ();
 sg13g2_decap_8 FILLER_26_1745 ();
 sg13g2_decap_8 FILLER_26_1752 ();
 sg13g2_decap_8 FILLER_26_1759 ();
 sg13g2_decap_8 FILLER_26_1766 ();
 sg13g2_fill_1 FILLER_26_1773 ();
 sg13g2_decap_8 FILLER_27_26 ();
 sg13g2_decap_4 FILLER_27_33 ();
 sg13g2_fill_2 FILLER_27_37 ();
 sg13g2_fill_2 FILLER_27_78 ();
 sg13g2_decap_8 FILLER_27_101 ();
 sg13g2_decap_8 FILLER_27_108 ();
 sg13g2_decap_8 FILLER_27_115 ();
 sg13g2_fill_2 FILLER_27_122 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_150 ();
 sg13g2_decap_8 FILLER_27_156 ();
 sg13g2_decap_4 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_fill_2 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_320 ();
 sg13g2_decap_8 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_334 ();
 sg13g2_decap_8 FILLER_27_341 ();
 sg13g2_decap_4 FILLER_27_348 ();
 sg13g2_fill_1 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_fill_1 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_fill_1 FILLER_27_383 ();
 sg13g2_fill_2 FILLER_27_405 ();
 sg13g2_fill_1 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_27_443 ();
 sg13g2_fill_1 FILLER_27_447 ();
 sg13g2_decap_8 FILLER_27_461 ();
 sg13g2_fill_2 FILLER_27_468 ();
 sg13g2_fill_1 FILLER_27_470 ();
 sg13g2_decap_8 FILLER_27_475 ();
 sg13g2_fill_2 FILLER_27_482 ();
 sg13g2_fill_1 FILLER_27_484 ();
 sg13g2_decap_8 FILLER_27_506 ();
 sg13g2_decap_8 FILLER_27_513 ();
 sg13g2_decap_8 FILLER_27_520 ();
 sg13g2_decap_8 FILLER_27_527 ();
 sg13g2_decap_4 FILLER_27_534 ();
 sg13g2_decap_8 FILLER_27_542 ();
 sg13g2_fill_1 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_575 ();
 sg13g2_decap_4 FILLER_27_582 ();
 sg13g2_fill_1 FILLER_27_586 ();
 sg13g2_fill_2 FILLER_27_679 ();
 sg13g2_decap_4 FILLER_27_702 ();
 sg13g2_fill_1 FILLER_27_706 ();
 sg13g2_fill_2 FILLER_27_711 ();
 sg13g2_decap_4 FILLER_27_738 ();
 sg13g2_fill_1 FILLER_27_742 ();
 sg13g2_decap_4 FILLER_27_748 ();
 sg13g2_fill_2 FILLER_27_752 ();
 sg13g2_fill_2 FILLER_27_762 ();
 sg13g2_fill_2 FILLER_27_804 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_867 ();
 sg13g2_decap_8 FILLER_27_882 ();
 sg13g2_decap_4 FILLER_27_889 ();
 sg13g2_fill_1 FILLER_27_893 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_912 ();
 sg13g2_decap_8 FILLER_27_919 ();
 sg13g2_decap_4 FILLER_27_926 ();
 sg13g2_decap_8 FILLER_27_964 ();
 sg13g2_decap_4 FILLER_27_971 ();
 sg13g2_fill_1 FILLER_27_975 ();
 sg13g2_fill_2 FILLER_27_980 ();
 sg13g2_decap_8 FILLER_27_1003 ();
 sg13g2_decap_8 FILLER_27_1018 ();
 sg13g2_decap_8 FILLER_27_1025 ();
 sg13g2_decap_8 FILLER_27_1032 ();
 sg13g2_decap_8 FILLER_27_1039 ();
 sg13g2_decap_8 FILLER_27_1046 ();
 sg13g2_fill_1 FILLER_27_1053 ();
 sg13g2_decap_8 FILLER_27_1075 ();
 sg13g2_fill_1 FILLER_27_1082 ();
 sg13g2_decap_8 FILLER_27_1118 ();
 sg13g2_decap_4 FILLER_27_1125 ();
 sg13g2_fill_2 FILLER_27_1137 ();
 sg13g2_fill_2 FILLER_27_1175 ();
 sg13g2_fill_1 FILLER_27_1177 ();
 sg13g2_fill_1 FILLER_27_1199 ();
 sg13g2_fill_2 FILLER_27_1230 ();
 sg13g2_fill_1 FILLER_27_1232 ();
 sg13g2_decap_8 FILLER_27_1293 ();
 sg13g2_decap_4 FILLER_27_1334 ();
 sg13g2_decap_4 FILLER_27_1342 ();
 sg13g2_decap_8 FILLER_27_1350 ();
 sg13g2_decap_8 FILLER_27_1357 ();
 sg13g2_fill_1 FILLER_27_1364 ();
 sg13g2_decap_8 FILLER_27_1414 ();
 sg13g2_fill_2 FILLER_27_1421 ();
 sg13g2_fill_2 FILLER_27_1458 ();
 sg13g2_fill_1 FILLER_27_1460 ();
 sg13g2_fill_1 FILLER_27_1487 ();
 sg13g2_fill_1 FILLER_27_1498 ();
 sg13g2_fill_1 FILLER_27_1509 ();
 sg13g2_fill_1 FILLER_27_1536 ();
 sg13g2_fill_2 FILLER_27_1573 ();
 sg13g2_decap_8 FILLER_27_1601 ();
 sg13g2_fill_2 FILLER_27_1608 ();
 sg13g2_decap_4 FILLER_27_1614 ();
 sg13g2_fill_2 FILLER_27_1618 ();
 sg13g2_fill_2 FILLER_27_1656 ();
 sg13g2_fill_1 FILLER_27_1658 ();
 sg13g2_decap_4 FILLER_27_1685 ();
 sg13g2_fill_2 FILLER_27_1689 ();
 sg13g2_decap_8 FILLER_27_1717 ();
 sg13g2_decap_8 FILLER_27_1724 ();
 sg13g2_decap_8 FILLER_27_1731 ();
 sg13g2_decap_8 FILLER_27_1738 ();
 sg13g2_decap_8 FILLER_27_1745 ();
 sg13g2_decap_8 FILLER_27_1752 ();
 sg13g2_decap_8 FILLER_27_1759 ();
 sg13g2_decap_8 FILLER_27_1766 ();
 sg13g2_fill_1 FILLER_27_1773 ();
 sg13g2_fill_1 FILLER_28_26 ();
 sg13g2_fill_1 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_37 ();
 sg13g2_fill_2 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_46 ();
 sg13g2_decap_4 FILLER_28_51 ();
 sg13g2_fill_2 FILLER_28_55 ();
 sg13g2_fill_2 FILLER_28_75 ();
 sg13g2_decap_8 FILLER_28_90 ();
 sg13g2_decap_4 FILLER_28_97 ();
 sg13g2_fill_2 FILLER_28_101 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_117 ();
 sg13g2_decap_8 FILLER_28_124 ();
 sg13g2_fill_2 FILLER_28_136 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_fill_2 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_173 ();
 sg13g2_fill_2 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_decap_4 FILLER_28_228 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_fill_2 FILLER_28_266 ();
 sg13g2_fill_1 FILLER_28_268 ();
 sg13g2_decap_4 FILLER_28_295 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_decap_4 FILLER_28_325 ();
 sg13g2_decap_8 FILLER_28_333 ();
 sg13g2_decap_4 FILLER_28_340 ();
 sg13g2_fill_2 FILLER_28_344 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_382 ();
 sg13g2_fill_1 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_decap_4 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_431 ();
 sg13g2_fill_2 FILLER_28_437 ();
 sg13g2_fill_1 FILLER_28_443 ();
 sg13g2_fill_1 FILLER_28_465 ();
 sg13g2_fill_1 FILLER_28_471 ();
 sg13g2_fill_2 FILLER_28_476 ();
 sg13g2_fill_2 FILLER_28_482 ();
 sg13g2_fill_2 FILLER_28_505 ();
 sg13g2_fill_2 FILLER_28_515 ();
 sg13g2_decap_8 FILLER_28_530 ();
 sg13g2_fill_2 FILLER_28_541 ();
 sg13g2_fill_1 FILLER_28_548 ();
 sg13g2_decap_8 FILLER_28_574 ();
 sg13g2_decap_4 FILLER_28_581 ();
 sg13g2_fill_2 FILLER_28_585 ();
 sg13g2_fill_2 FILLER_28_592 ();
 sg13g2_decap_8 FILLER_28_598 ();
 sg13g2_decap_4 FILLER_28_605 ();
 sg13g2_decap_8 FILLER_28_613 ();
 sg13g2_decap_8 FILLER_28_620 ();
 sg13g2_fill_2 FILLER_28_627 ();
 sg13g2_fill_1 FILLER_28_629 ();
 sg13g2_fill_1 FILLER_28_643 ();
 sg13g2_decap_8 FILLER_28_660 ();
 sg13g2_fill_1 FILLER_28_696 ();
 sg13g2_decap_4 FILLER_28_706 ();
 sg13g2_fill_2 FILLER_28_710 ();
 sg13g2_decap_8 FILLER_28_716 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_773 ();
 sg13g2_fill_2 FILLER_28_780 ();
 sg13g2_fill_1 FILLER_28_782 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_fill_1 FILLER_28_826 ();
 sg13g2_fill_2 FILLER_28_831 ();
 sg13g2_fill_1 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_fill_1 FILLER_28_854 ();
 sg13g2_decap_4 FILLER_28_860 ();
 sg13g2_fill_2 FILLER_28_864 ();
 sg13g2_fill_1 FILLER_28_878 ();
 sg13g2_decap_8 FILLER_28_884 ();
 sg13g2_fill_1 FILLER_28_891 ();
 sg13g2_fill_1 FILLER_28_923 ();
 sg13g2_decap_8 FILLER_28_960 ();
 sg13g2_decap_4 FILLER_28_967 ();
 sg13g2_fill_1 FILLER_28_971 ();
 sg13g2_decap_4 FILLER_28_976 ();
 sg13g2_decap_8 FILLER_28_1001 ();
 sg13g2_fill_1 FILLER_28_1008 ();
 sg13g2_decap_8 FILLER_28_1040 ();
 sg13g2_decap_4 FILLER_28_1047 ();
 sg13g2_decap_8 FILLER_28_1060 ();
 sg13g2_decap_8 FILLER_28_1067 ();
 sg13g2_decap_4 FILLER_28_1074 ();
 sg13g2_decap_8 FILLER_28_1083 ();
 sg13g2_decap_4 FILLER_28_1090 ();
 sg13g2_fill_1 FILLER_28_1094 ();
 sg13g2_decap_8 FILLER_28_1103 ();
 sg13g2_fill_1 FILLER_28_1110 ();
 sg13g2_fill_1 FILLER_28_1120 ();
 sg13g2_decap_8 FILLER_28_1151 ();
 sg13g2_fill_1 FILLER_28_1158 ();
 sg13g2_decap_8 FILLER_28_1163 ();
 sg13g2_decap_8 FILLER_28_1170 ();
 sg13g2_fill_2 FILLER_28_1177 ();
 sg13g2_decap_4 FILLER_28_1200 ();
 sg13g2_fill_2 FILLER_28_1204 ();
 sg13g2_fill_1 FILLER_28_1216 ();
 sg13g2_decap_8 FILLER_28_1243 ();
 sg13g2_decap_8 FILLER_28_1250 ();
 sg13g2_fill_1 FILLER_28_1257 ();
 sg13g2_decap_4 FILLER_28_1275 ();
 sg13g2_decap_4 FILLER_28_1309 ();
 sg13g2_fill_1 FILLER_28_1313 ();
 sg13g2_fill_2 FILLER_28_1323 ();
 sg13g2_fill_2 FILLER_28_1337 ();
 sg13g2_decap_8 FILLER_28_1369 ();
 sg13g2_decap_8 FILLER_28_1376 ();
 sg13g2_decap_4 FILLER_28_1383 ();
 sg13g2_fill_2 FILLER_28_1387 ();
 sg13g2_decap_4 FILLER_28_1393 ();
 sg13g2_fill_1 FILLER_28_1397 ();
 sg13g2_decap_4 FILLER_28_1402 ();
 sg13g2_fill_2 FILLER_28_1447 ();
 sg13g2_decap_8 FILLER_28_1459 ();
 sg13g2_decap_4 FILLER_28_1466 ();
 sg13g2_fill_1 FILLER_28_1470 ();
 sg13g2_decap_8 FILLER_28_1475 ();
 sg13g2_decap_8 FILLER_28_1482 ();
 sg13g2_fill_1 FILLER_28_1489 ();
 sg13g2_fill_1 FILLER_28_1502 ();
 sg13g2_fill_1 FILLER_28_1516 ();
 sg13g2_decap_8 FILLER_28_1527 ();
 sg13g2_fill_2 FILLER_28_1544 ();
 sg13g2_fill_2 FILLER_28_1550 ();
 sg13g2_fill_1 FILLER_28_1562 ();
 sg13g2_fill_2 FILLER_28_1583 ();
 sg13g2_decap_4 FILLER_28_1589 ();
 sg13g2_fill_2 FILLER_28_1593 ();
 sg13g2_decap_8 FILLER_28_1600 ();
 sg13g2_decap_4 FILLER_28_1607 ();
 sg13g2_fill_2 FILLER_28_1611 ();
 sg13g2_decap_8 FILLER_28_1617 ();
 sg13g2_fill_1 FILLER_28_1624 ();
 sg13g2_decap_8 FILLER_28_1630 ();
 sg13g2_decap_8 FILLER_28_1641 ();
 sg13g2_decap_8 FILLER_28_1648 ();
 sg13g2_decap_8 FILLER_28_1655 ();
 sg13g2_decap_4 FILLER_28_1662 ();
 sg13g2_decap_8 FILLER_28_1670 ();
 sg13g2_decap_8 FILLER_28_1677 ();
 sg13g2_decap_8 FILLER_28_1684 ();
 sg13g2_decap_4 FILLER_28_1691 ();
 sg13g2_fill_2 FILLER_28_1695 ();
 sg13g2_decap_8 FILLER_28_1701 ();
 sg13g2_decap_8 FILLER_28_1708 ();
 sg13g2_decap_8 FILLER_28_1715 ();
 sg13g2_decap_8 FILLER_28_1722 ();
 sg13g2_decap_8 FILLER_28_1729 ();
 sg13g2_decap_8 FILLER_28_1736 ();
 sg13g2_decap_8 FILLER_28_1743 ();
 sg13g2_decap_8 FILLER_28_1750 ();
 sg13g2_decap_8 FILLER_28_1757 ();
 sg13g2_decap_8 FILLER_28_1764 ();
 sg13g2_fill_2 FILLER_28_1771 ();
 sg13g2_fill_1 FILLER_28_1773 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_15 ();
 sg13g2_fill_1 FILLER_29_17 ();
 sg13g2_fill_1 FILLER_29_101 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_213 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_392 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_29_456 ();
 sg13g2_fill_2 FILLER_29_463 ();
 sg13g2_fill_1 FILLER_29_465 ();
 sg13g2_decap_8 FILLER_29_492 ();
 sg13g2_decap_8 FILLER_29_516 ();
 sg13g2_fill_2 FILLER_29_523 ();
 sg13g2_fill_1 FILLER_29_525 ();
 sg13g2_fill_2 FILLER_29_557 ();
 sg13g2_fill_1 FILLER_29_559 ();
 sg13g2_decap_8 FILLER_29_564 ();
 sg13g2_decap_8 FILLER_29_571 ();
 sg13g2_fill_1 FILLER_29_609 ();
 sg13g2_fill_1 FILLER_29_615 ();
 sg13g2_fill_1 FILLER_29_620 ();
 sg13g2_fill_2 FILLER_29_625 ();
 sg13g2_fill_1 FILLER_29_637 ();
 sg13g2_fill_1 FILLER_29_690 ();
 sg13g2_fill_2 FILLER_29_730 ();
 sg13g2_fill_2 FILLER_29_736 ();
 sg13g2_fill_2 FILLER_29_747 ();
 sg13g2_decap_8 FILLER_29_758 ();
 sg13g2_fill_2 FILLER_29_801 ();
 sg13g2_fill_1 FILLER_29_803 ();
 sg13g2_decap_8 FILLER_29_808 ();
 sg13g2_decap_8 FILLER_29_815 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_fill_1 FILLER_29_847 ();
 sg13g2_decap_4 FILLER_29_857 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_4 FILLER_29_893 ();
 sg13g2_fill_2 FILLER_29_901 ();
 sg13g2_fill_1 FILLER_29_903 ();
 sg13g2_decap_8 FILLER_29_912 ();
 sg13g2_decap_8 FILLER_29_919 ();
 sg13g2_fill_2 FILLER_29_926 ();
 sg13g2_fill_1 FILLER_29_928 ();
 sg13g2_decap_4 FILLER_29_934 ();
 sg13g2_decap_4 FILLER_29_950 ();
 sg13g2_decap_8 FILLER_29_984 ();
 sg13g2_decap_8 FILLER_29_991 ();
 sg13g2_decap_8 FILLER_29_998 ();
 sg13g2_fill_2 FILLER_29_1005 ();
 sg13g2_decap_4 FILLER_29_1033 ();
 sg13g2_fill_1 FILLER_29_1037 ();
 sg13g2_decap_4 FILLER_29_1068 ();
 sg13g2_decap_4 FILLER_29_1102 ();
 sg13g2_fill_1 FILLER_29_1106 ();
 sg13g2_decap_8 FILLER_29_1133 ();
 sg13g2_fill_2 FILLER_29_1140 ();
 sg13g2_fill_1 FILLER_29_1178 ();
 sg13g2_fill_1 FILLER_29_1200 ();
 sg13g2_fill_1 FILLER_29_1211 ();
 sg13g2_fill_1 FILLER_29_1238 ();
 sg13g2_fill_2 FILLER_29_1243 ();
 sg13g2_fill_1 FILLER_29_1245 ();
 sg13g2_fill_2 FILLER_29_1277 ();
 sg13g2_fill_1 FILLER_29_1279 ();
 sg13g2_decap_8 FILLER_29_1295 ();
 sg13g2_decap_8 FILLER_29_1302 ();
 sg13g2_decap_8 FILLER_29_1309 ();
 sg13g2_decap_4 FILLER_29_1316 ();
 sg13g2_fill_2 FILLER_29_1336 ();
 sg13g2_decap_8 FILLER_29_1349 ();
 sg13g2_fill_1 FILLER_29_1356 ();
 sg13g2_fill_1 FILLER_29_1367 ();
 sg13g2_fill_1 FILLER_29_1371 ();
 sg13g2_fill_1 FILLER_29_1376 ();
 sg13g2_fill_1 FILLER_29_1382 ();
 sg13g2_fill_1 FILLER_29_1391 ();
 sg13g2_fill_1 FILLER_29_1418 ();
 sg13g2_fill_1 FILLER_29_1441 ();
 sg13g2_decap_8 FILLER_29_1446 ();
 sg13g2_decap_8 FILLER_29_1453 ();
 sg13g2_fill_1 FILLER_29_1460 ();
 sg13g2_decap_8 FILLER_29_1465 ();
 sg13g2_fill_2 FILLER_29_1472 ();
 sg13g2_fill_2 FILLER_29_1490 ();
 sg13g2_decap_4 FILLER_29_1496 ();
 sg13g2_fill_1 FILLER_29_1500 ();
 sg13g2_fill_1 FILLER_29_1505 ();
 sg13g2_decap_8 FILLER_29_1513 ();
 sg13g2_fill_1 FILLER_29_1520 ();
 sg13g2_decap_4 FILLER_29_1526 ();
 sg13g2_fill_2 FILLER_29_1530 ();
 sg13g2_decap_8 FILLER_29_1536 ();
 sg13g2_decap_8 FILLER_29_1543 ();
 sg13g2_decap_8 FILLER_29_1550 ();
 sg13g2_decap_8 FILLER_29_1557 ();
 sg13g2_decap_4 FILLER_29_1564 ();
 sg13g2_fill_1 FILLER_29_1568 ();
 sg13g2_decap_4 FILLER_29_1578 ();
 sg13g2_decap_8 FILLER_29_1586 ();
 sg13g2_decap_4 FILLER_29_1593 ();
 sg13g2_fill_2 FILLER_29_1597 ();
 sg13g2_decap_8 FILLER_29_1638 ();
 sg13g2_fill_2 FILLER_29_1645 ();
 sg13g2_fill_1 FILLER_29_1647 ();
 sg13g2_decap_8 FILLER_29_1656 ();
 sg13g2_decap_8 FILLER_29_1663 ();
 sg13g2_decap_8 FILLER_29_1670 ();
 sg13g2_decap_8 FILLER_29_1677 ();
 sg13g2_decap_8 FILLER_29_1684 ();
 sg13g2_decap_8 FILLER_29_1691 ();
 sg13g2_decap_8 FILLER_29_1698 ();
 sg13g2_decap_8 FILLER_29_1705 ();
 sg13g2_decap_8 FILLER_29_1712 ();
 sg13g2_decap_8 FILLER_29_1719 ();
 sg13g2_decap_8 FILLER_29_1726 ();
 sg13g2_decap_8 FILLER_29_1733 ();
 sg13g2_decap_8 FILLER_29_1740 ();
 sg13g2_decap_8 FILLER_29_1747 ();
 sg13g2_decap_8 FILLER_29_1754 ();
 sg13g2_decap_8 FILLER_29_1761 ();
 sg13g2_decap_4 FILLER_29_1768 ();
 sg13g2_fill_2 FILLER_29_1772 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_decap_4 FILLER_30_51 ();
 sg13g2_fill_2 FILLER_30_59 ();
 sg13g2_decap_8 FILLER_30_65 ();
 sg13g2_decap_8 FILLER_30_72 ();
 sg13g2_decap_4 FILLER_30_88 ();
 sg13g2_decap_8 FILLER_30_113 ();
 sg13g2_decap_4 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_124 ();
 sg13g2_decap_4 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_decap_8 FILLER_30_183 ();
 sg13g2_decap_4 FILLER_30_190 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_decap_8 FILLER_30_204 ();
 sg13g2_decap_4 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_246 ();
 sg13g2_decap_8 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_decap_4 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_fill_1 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_fill_1 FILLER_30_401 ();
 sg13g2_decap_4 FILLER_30_406 ();
 sg13g2_fill_2 FILLER_30_410 ();
 sg13g2_decap_8 FILLER_30_416 ();
 sg13g2_decap_8 FILLER_30_423 ();
 sg13g2_decap_4 FILLER_30_430 ();
 sg13g2_fill_2 FILLER_30_434 ();
 sg13g2_fill_2 FILLER_30_440 ();
 sg13g2_fill_1 FILLER_30_442 ();
 sg13g2_decap_8 FILLER_30_456 ();
 sg13g2_decap_8 FILLER_30_463 ();
 sg13g2_decap_4 FILLER_30_470 ();
 sg13g2_fill_2 FILLER_30_500 ();
 sg13g2_fill_1 FILLER_30_502 ();
 sg13g2_decap_8 FILLER_30_537 ();
 sg13g2_decap_8 FILLER_30_544 ();
 sg13g2_fill_2 FILLER_30_551 ();
 sg13g2_fill_1 FILLER_30_553 ();
 sg13g2_fill_2 FILLER_30_580 ();
 sg13g2_decap_4 FILLER_30_603 ();
 sg13g2_decap_4 FILLER_30_633 ();
 sg13g2_fill_2 FILLER_30_662 ();
 sg13g2_fill_2 FILLER_30_669 ();
 sg13g2_fill_1 FILLER_30_671 ();
 sg13g2_decap_8 FILLER_30_676 ();
 sg13g2_fill_1 FILLER_30_683 ();
 sg13g2_fill_2 FILLER_30_706 ();
 sg13g2_fill_1 FILLER_30_765 ();
 sg13g2_decap_4 FILLER_30_779 ();
 sg13g2_decap_8 FILLER_30_792 ();
 sg13g2_decap_4 FILLER_30_799 ();
 sg13g2_decap_8 FILLER_30_865 ();
 sg13g2_decap_8 FILLER_30_876 ();
 sg13g2_decap_8 FILLER_30_883 ();
 sg13g2_fill_2 FILLER_30_890 ();
 sg13g2_decap_8 FILLER_30_923 ();
 sg13g2_fill_1 FILLER_30_930 ();
 sg13g2_decap_8 FILLER_30_957 ();
 sg13g2_decap_8 FILLER_30_964 ();
 sg13g2_decap_4 FILLER_30_971 ();
 sg13g2_fill_2 FILLER_30_975 ();
 sg13g2_fill_2 FILLER_30_982 ();
 sg13g2_fill_1 FILLER_30_984 ();
 sg13g2_decap_4 FILLER_30_1015 ();
 sg13g2_fill_2 FILLER_30_1045 ();
 sg13g2_decap_8 FILLER_30_1060 ();
 sg13g2_decap_8 FILLER_30_1067 ();
 sg13g2_decap_4 FILLER_30_1074 ();
 sg13g2_fill_2 FILLER_30_1083 ();
 sg13g2_fill_1 FILLER_30_1085 ();
 sg13g2_fill_2 FILLER_30_1132 ();
 sg13g2_decap_8 FILLER_30_1160 ();
 sg13g2_decap_8 FILLER_30_1167 ();
 sg13g2_fill_1 FILLER_30_1174 ();
 sg13g2_decap_8 FILLER_30_1179 ();
 sg13g2_decap_4 FILLER_30_1186 ();
 sg13g2_fill_2 FILLER_30_1190 ();
 sg13g2_decap_8 FILLER_30_1228 ();
 sg13g2_decap_8 FILLER_30_1235 ();
 sg13g2_decap_8 FILLER_30_1242 ();
 sg13g2_decap_4 FILLER_30_1249 ();
 sg13g2_fill_2 FILLER_30_1253 ();
 sg13g2_decap_8 FILLER_30_1259 ();
 sg13g2_decap_4 FILLER_30_1266 ();
 sg13g2_decap_4 FILLER_30_1274 ();
 sg13g2_fill_2 FILLER_30_1278 ();
 sg13g2_fill_2 FILLER_30_1294 ();
 sg13g2_decap_4 FILLER_30_1300 ();
 sg13g2_fill_1 FILLER_30_1304 ();
 sg13g2_fill_2 FILLER_30_1308 ();
 sg13g2_fill_1 FILLER_30_1310 ();
 sg13g2_decap_4 FILLER_30_1319 ();
 sg13g2_decap_8 FILLER_30_1328 ();
 sg13g2_decap_8 FILLER_30_1335 ();
 sg13g2_decap_8 FILLER_30_1342 ();
 sg13g2_decap_8 FILLER_30_1349 ();
 sg13g2_decap_4 FILLER_30_1373 ();
 sg13g2_fill_2 FILLER_30_1394 ();
 sg13g2_fill_1 FILLER_30_1396 ();
 sg13g2_decap_8 FILLER_30_1427 ();
 sg13g2_fill_1 FILLER_30_1434 ();
 sg13g2_fill_1 FILLER_30_1466 ();
 sg13g2_fill_1 FILLER_30_1472 ();
 sg13g2_fill_1 FILLER_30_1477 ();
 sg13g2_fill_2 FILLER_30_1483 ();
 sg13g2_decap_8 FILLER_30_1511 ();
 sg13g2_fill_2 FILLER_30_1518 ();
 sg13g2_fill_1 FILLER_30_1525 ();
 sg13g2_decap_8 FILLER_30_1552 ();
 sg13g2_decap_4 FILLER_30_1559 ();
 sg13g2_fill_1 FILLER_30_1563 ();
 sg13g2_decap_4 FILLER_30_1567 ();
 sg13g2_decap_8 FILLER_30_1602 ();
 sg13g2_decap_4 FILLER_30_1609 ();
 sg13g2_decap_8 FILLER_30_1617 ();
 sg13g2_fill_1 FILLER_30_1624 ();
 sg13g2_decap_8 FILLER_30_1629 ();
 sg13g2_fill_2 FILLER_30_1636 ();
 sg13g2_decap_8 FILLER_30_1664 ();
 sg13g2_decap_8 FILLER_30_1675 ();
 sg13g2_decap_8 FILLER_30_1682 ();
 sg13g2_decap_8 FILLER_30_1689 ();
 sg13g2_decap_8 FILLER_30_1696 ();
 sg13g2_decap_8 FILLER_30_1703 ();
 sg13g2_decap_8 FILLER_30_1710 ();
 sg13g2_decap_8 FILLER_30_1717 ();
 sg13g2_decap_8 FILLER_30_1724 ();
 sg13g2_decap_8 FILLER_30_1731 ();
 sg13g2_decap_8 FILLER_30_1738 ();
 sg13g2_decap_8 FILLER_30_1745 ();
 sg13g2_decap_8 FILLER_30_1752 ();
 sg13g2_decap_8 FILLER_30_1759 ();
 sg13g2_decap_8 FILLER_30_1766 ();
 sg13g2_fill_1 FILLER_30_1773 ();
 sg13g2_decap_4 FILLER_31_31 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_decap_4 FILLER_31_114 ();
 sg13g2_fill_2 FILLER_31_144 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_decap_4 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_decap_4 FILLER_31_335 ();
 sg13g2_fill_2 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_421 ();
 sg13g2_decap_8 FILLER_31_428 ();
 sg13g2_decap_4 FILLER_31_435 ();
 sg13g2_fill_2 FILLER_31_439 ();
 sg13g2_decap_8 FILLER_31_467 ();
 sg13g2_fill_2 FILLER_31_474 ();
 sg13g2_fill_1 FILLER_31_476 ();
 sg13g2_fill_2 FILLER_31_486 ();
 sg13g2_decap_4 FILLER_31_495 ();
 sg13g2_fill_2 FILLER_31_499 ();
 sg13g2_decap_4 FILLER_31_511 ();
 sg13g2_fill_1 FILLER_31_519 ();
 sg13g2_fill_2 FILLER_31_545 ();
 sg13g2_decap_8 FILLER_31_551 ();
 sg13g2_decap_8 FILLER_31_558 ();
 sg13g2_decap_8 FILLER_31_565 ();
 sg13g2_fill_2 FILLER_31_572 ();
 sg13g2_fill_1 FILLER_31_574 ();
 sg13g2_fill_2 FILLER_31_601 ();
 sg13g2_fill_1 FILLER_31_603 ();
 sg13g2_fill_2 FILLER_31_609 ();
 sg13g2_fill_1 FILLER_31_611 ();
 sg13g2_fill_2 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_622 ();
 sg13g2_decap_8 FILLER_31_629 ();
 sg13g2_fill_2 FILLER_31_636 ();
 sg13g2_decap_4 FILLER_31_659 ();
 sg13g2_fill_1 FILLER_31_663 ();
 sg13g2_decap_8 FILLER_31_668 ();
 sg13g2_decap_8 FILLER_31_675 ();
 sg13g2_fill_2 FILLER_31_682 ();
 sg13g2_fill_2 FILLER_31_693 ();
 sg13g2_fill_2 FILLER_31_717 ();
 sg13g2_fill_1 FILLER_31_726 ();
 sg13g2_decap_4 FILLER_31_739 ();
 sg13g2_fill_2 FILLER_31_743 ();
 sg13g2_fill_2 FILLER_31_759 ();
 sg13g2_fill_1 FILLER_31_766 ();
 sg13g2_fill_2 FILLER_31_797 ();
 sg13g2_fill_1 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_821 ();
 sg13g2_decap_8 FILLER_31_828 ();
 sg13g2_decap_8 FILLER_31_835 ();
 sg13g2_decap_4 FILLER_31_842 ();
 sg13g2_fill_1 FILLER_31_864 ();
 sg13g2_fill_2 FILLER_31_891 ();
 sg13g2_fill_1 FILLER_31_893 ();
 sg13g2_fill_2 FILLER_31_925 ();
 sg13g2_fill_1 FILLER_31_927 ();
 sg13g2_decap_4 FILLER_31_964 ();
 sg13g2_fill_2 FILLER_31_968 ();
 sg13g2_decap_8 FILLER_31_974 ();
 sg13g2_fill_2 FILLER_31_981 ();
 sg13g2_decap_8 FILLER_31_988 ();
 sg13g2_fill_2 FILLER_31_995 ();
 sg13g2_fill_1 FILLER_31_997 ();
 sg13g2_decap_8 FILLER_31_1002 ();
 sg13g2_decap_8 FILLER_31_1009 ();
 sg13g2_decap_8 FILLER_31_1016 ();
 sg13g2_fill_1 FILLER_31_1023 ();
 sg13g2_decap_8 FILLER_31_1032 ();
 sg13g2_decap_8 FILLER_31_1039 ();
 sg13g2_fill_2 FILLER_31_1046 ();
 sg13g2_fill_1 FILLER_31_1048 ();
 sg13g2_decap_4 FILLER_31_1075 ();
 sg13g2_decap_8 FILLER_31_1144 ();
 sg13g2_decap_8 FILLER_31_1151 ();
 sg13g2_fill_2 FILLER_31_1207 ();
 sg13g2_decap_8 FILLER_31_1213 ();
 sg13g2_decap_8 FILLER_31_1220 ();
 sg13g2_decap_4 FILLER_31_1227 ();
 sg13g2_fill_2 FILLER_31_1231 ();
 sg13g2_fill_1 FILLER_31_1332 ();
 sg13g2_fill_1 FILLER_31_1354 ();
 sg13g2_fill_2 FILLER_31_1359 ();
 sg13g2_fill_1 FILLER_31_1376 ();
 sg13g2_decap_8 FILLER_31_1381 ();
 sg13g2_fill_2 FILLER_31_1388 ();
 sg13g2_fill_1 FILLER_31_1390 ();
 sg13g2_decap_8 FILLER_31_1395 ();
 sg13g2_decap_4 FILLER_31_1402 ();
 sg13g2_fill_1 FILLER_31_1406 ();
 sg13g2_fill_2 FILLER_31_1420 ();
 sg13g2_decap_8 FILLER_31_1426 ();
 sg13g2_decap_8 FILLER_31_1433 ();
 sg13g2_decap_4 FILLER_31_1440 ();
 sg13g2_fill_2 FILLER_31_1444 ();
 sg13g2_decap_8 FILLER_31_1450 ();
 sg13g2_decap_8 FILLER_31_1457 ();
 sg13g2_decap_4 FILLER_31_1464 ();
 sg13g2_fill_2 FILLER_31_1479 ();
 sg13g2_fill_1 FILLER_31_1481 ();
 sg13g2_fill_2 FILLER_31_1515 ();
 sg13g2_fill_1 FILLER_31_1517 ();
 sg13g2_decap_8 FILLER_31_1528 ();
 sg13g2_decap_4 FILLER_31_1535 ();
 sg13g2_decap_8 FILLER_31_1574 ();
 sg13g2_decap_8 FILLER_31_1581 ();
 sg13g2_fill_2 FILLER_31_1661 ();
 sg13g2_fill_1 FILLER_31_1663 ();
 sg13g2_decap_8 FILLER_31_1716 ();
 sg13g2_decap_8 FILLER_31_1723 ();
 sg13g2_decap_8 FILLER_31_1730 ();
 sg13g2_decap_8 FILLER_31_1737 ();
 sg13g2_decap_8 FILLER_31_1744 ();
 sg13g2_decap_8 FILLER_31_1751 ();
 sg13g2_decap_8 FILLER_31_1758 ();
 sg13g2_decap_8 FILLER_31_1765 ();
 sg13g2_fill_2 FILLER_31_1772 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_18 ();
 sg13g2_fill_1 FILLER_32_25 ();
 sg13g2_decap_4 FILLER_32_39 ();
 sg13g2_fill_1 FILLER_32_43 ();
 sg13g2_decap_8 FILLER_32_48 ();
 sg13g2_decap_8 FILLER_32_55 ();
 sg13g2_decap_8 FILLER_32_62 ();
 sg13g2_decap_4 FILLER_32_69 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_decap_8 FILLER_32_78 ();
 sg13g2_decap_8 FILLER_32_85 ();
 sg13g2_decap_8 FILLER_32_92 ();
 sg13g2_decap_8 FILLER_32_99 ();
 sg13g2_decap_8 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_113 ();
 sg13g2_decap_4 FILLER_32_120 ();
 sg13g2_fill_1 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_138 ();
 sg13g2_fill_1 FILLER_32_140 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_decap_8 FILLER_32_188 ();
 sg13g2_decap_4 FILLER_32_195 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_decap_4 FILLER_32_214 ();
 sg13g2_fill_2 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_fill_1 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_decap_8 FILLER_32_275 ();
 sg13g2_decap_4 FILLER_32_282 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_343 ();
 sg13g2_fill_1 FILLER_32_345 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_4 FILLER_32_357 ();
 sg13g2_fill_1 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_4 FILLER_32_395 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_436 ();
 sg13g2_fill_1 FILLER_32_438 ();
 sg13g2_decap_4 FILLER_32_470 ();
 sg13g2_fill_1 FILLER_32_482 ();
 sg13g2_fill_2 FILLER_32_488 ();
 sg13g2_fill_2 FILLER_32_522 ();
 sg13g2_fill_1 FILLER_32_545 ();
 sg13g2_decap_8 FILLER_32_585 ();
 sg13g2_decap_4 FILLER_32_592 ();
 sg13g2_fill_2 FILLER_32_596 ();
 sg13g2_decap_8 FILLER_32_633 ();
 sg13g2_decap_8 FILLER_32_640 ();
 sg13g2_fill_1 FILLER_32_709 ();
 sg13g2_fill_2 FILLER_32_727 ();
 sg13g2_decap_8 FILLER_32_733 ();
 sg13g2_decap_8 FILLER_32_740 ();
 sg13g2_decap_8 FILLER_32_747 ();
 sg13g2_fill_1 FILLER_32_754 ();
 sg13g2_fill_2 FILLER_32_759 ();
 sg13g2_fill_1 FILLER_32_761 ();
 sg13g2_decap_8 FILLER_32_766 ();
 sg13g2_decap_4 FILLER_32_773 ();
 sg13g2_fill_1 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_782 ();
 sg13g2_decap_8 FILLER_32_789 ();
 sg13g2_decap_4 FILLER_32_822 ();
 sg13g2_decap_4 FILLER_32_852 ();
 sg13g2_decap_4 FILLER_32_882 ();
 sg13g2_fill_1 FILLER_32_886 ();
 sg13g2_fill_1 FILLER_32_897 ();
 sg13g2_decap_4 FILLER_32_902 ();
 sg13g2_decap_8 FILLER_32_910 ();
 sg13g2_decap_8 FILLER_32_917 ();
 sg13g2_decap_8 FILLER_32_924 ();
 sg13g2_fill_1 FILLER_32_931 ();
 sg13g2_decap_4 FILLER_32_936 ();
 sg13g2_decap_4 FILLER_32_944 ();
 sg13g2_fill_2 FILLER_32_956 ();
 sg13g2_fill_1 FILLER_32_958 ();
 sg13g2_fill_1 FILLER_32_989 ();
 sg13g2_decap_8 FILLER_32_994 ();
 sg13g2_decap_8 FILLER_32_1001 ();
 sg13g2_decap_8 FILLER_32_1008 ();
 sg13g2_decap_8 FILLER_32_1046 ();
 sg13g2_fill_1 FILLER_32_1053 ();
 sg13g2_fill_1 FILLER_32_1063 ();
 sg13g2_decap_8 FILLER_32_1073 ();
 sg13g2_decap_4 FILLER_32_1080 ();
 sg13g2_fill_1 FILLER_32_1084 ();
 sg13g2_fill_2 FILLER_32_1107 ();
 sg13g2_fill_1 FILLER_32_1109 ();
 sg13g2_fill_2 FILLER_32_1114 ();
 sg13g2_decap_8 FILLER_32_1120 ();
 sg13g2_decap_8 FILLER_32_1127 ();
 sg13g2_decap_8 FILLER_32_1134 ();
 sg13g2_decap_8 FILLER_32_1141 ();
 sg13g2_decap_8 FILLER_32_1148 ();
 sg13g2_fill_2 FILLER_32_1155 ();
 sg13g2_fill_1 FILLER_32_1157 ();
 sg13g2_fill_1 FILLER_32_1168 ();
 sg13g2_fill_2 FILLER_32_1195 ();
 sg13g2_fill_1 FILLER_32_1197 ();
 sg13g2_fill_2 FILLER_32_1228 ();
 sg13g2_fill_1 FILLER_32_1234 ();
 sg13g2_fill_1 FILLER_32_1243 ();
 sg13g2_decap_8 FILLER_32_1248 ();
 sg13g2_decap_8 FILLER_32_1255 ();
 sg13g2_fill_2 FILLER_32_1262 ();
 sg13g2_decap_4 FILLER_32_1268 ();
 sg13g2_decap_8 FILLER_32_1276 ();
 sg13g2_fill_1 FILLER_32_1283 ();
 sg13g2_decap_8 FILLER_32_1288 ();
 sg13g2_decap_8 FILLER_32_1295 ();
 sg13g2_decap_8 FILLER_32_1302 ();
 sg13g2_decap_4 FILLER_32_1309 ();
 sg13g2_fill_2 FILLER_32_1313 ();
 sg13g2_decap_8 FILLER_32_1320 ();
 sg13g2_decap_4 FILLER_32_1327 ();
 sg13g2_decap_4 FILLER_32_1339 ();
 sg13g2_fill_1 FILLER_32_1343 ();
 sg13g2_decap_8 FILLER_32_1355 ();
 sg13g2_decap_8 FILLER_32_1362 ();
 sg13g2_fill_1 FILLER_32_1369 ();
 sg13g2_fill_2 FILLER_32_1396 ();
 sg13g2_fill_2 FILLER_32_1436 ();
 sg13g2_fill_1 FILLER_32_1438 ();
 sg13g2_fill_2 FILLER_32_1465 ();
 sg13g2_fill_1 FILLER_32_1467 ();
 sg13g2_fill_2 FILLER_32_1472 ();
 sg13g2_fill_1 FILLER_32_1474 ();
 sg13g2_decap_8 FILLER_32_1483 ();
 sg13g2_fill_1 FILLER_32_1490 ();
 sg13g2_decap_4 FILLER_32_1528 ();
 sg13g2_fill_1 FILLER_32_1532 ();
 sg13g2_fill_1 FILLER_32_1538 ();
 sg13g2_fill_2 FILLER_32_1544 ();
 sg13g2_decap_4 FILLER_32_1550 ();
 sg13g2_fill_1 FILLER_32_1554 ();
 sg13g2_decap_8 FILLER_32_1581 ();
 sg13g2_decap_8 FILLER_32_1588 ();
 sg13g2_decap_4 FILLER_32_1595 ();
 sg13g2_fill_1 FILLER_32_1599 ();
 sg13g2_decap_4 FILLER_32_1604 ();
 sg13g2_fill_2 FILLER_32_1608 ();
 sg13g2_fill_2 FILLER_32_1616 ();
 sg13g2_decap_8 FILLER_32_1622 ();
 sg13g2_decap_4 FILLER_32_1629 ();
 sg13g2_decap_8 FILLER_32_1671 ();
 sg13g2_decap_4 FILLER_32_1678 ();
 sg13g2_fill_2 FILLER_32_1682 ();
 sg13g2_fill_1 FILLER_32_1702 ();
 sg13g2_decap_8 FILLER_32_1733 ();
 sg13g2_decap_8 FILLER_32_1740 ();
 sg13g2_decap_8 FILLER_32_1747 ();
 sg13g2_decap_8 FILLER_32_1754 ();
 sg13g2_decap_8 FILLER_32_1761 ();
 sg13g2_decap_4 FILLER_32_1768 ();
 sg13g2_fill_2 FILLER_32_1772 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_11 ();
 sg13g2_fill_1 FILLER_33_13 ();
 sg13g2_fill_1 FILLER_33_18 ();
 sg13g2_fill_2 FILLER_33_45 ();
 sg13g2_fill_1 FILLER_33_47 ();
 sg13g2_fill_2 FILLER_33_57 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_4 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_74 ();
 sg13g2_fill_2 FILLER_33_96 ();
 sg13g2_fill_2 FILLER_33_103 ();
 sg13g2_fill_1 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_110 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_161 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_184 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_decap_8 FILLER_33_222 ();
 sg13g2_decap_8 FILLER_33_229 ();
 sg13g2_decap_4 FILLER_33_236 ();
 sg13g2_fill_1 FILLER_33_240 ();
 sg13g2_decap_4 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_decap_4 FILLER_33_276 ();
 sg13g2_decap_8 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_292 ();
 sg13g2_fill_2 FILLER_33_297 ();
 sg13g2_decap_4 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_decap_4 FILLER_33_348 ();
 sg13g2_decap_8 FILLER_33_356 ();
 sg13g2_fill_2 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_393 ();
 sg13g2_fill_2 FILLER_33_408 ();
 sg13g2_fill_1 FILLER_33_410 ();
 sg13g2_fill_1 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_425 ();
 sg13g2_fill_2 FILLER_33_432 ();
 sg13g2_fill_1 FILLER_33_434 ();
 sg13g2_fill_2 FILLER_33_445 ();
 sg13g2_fill_2 FILLER_33_460 ();
 sg13g2_fill_1 FILLER_33_462 ();
 sg13g2_decap_4 FILLER_33_508 ();
 sg13g2_decap_4 FILLER_33_521 ();
 sg13g2_decap_8 FILLER_33_529 ();
 sg13g2_decap_8 FILLER_33_536 ();
 sg13g2_fill_2 FILLER_33_543 ();
 sg13g2_fill_2 FILLER_33_550 ();
 sg13g2_fill_1 FILLER_33_552 ();
 sg13g2_fill_1 FILLER_33_562 ();
 sg13g2_fill_2 FILLER_33_568 ();
 sg13g2_fill_1 FILLER_33_570 ();
 sg13g2_decap_4 FILLER_33_597 ();
 sg13g2_fill_2 FILLER_33_601 ();
 sg13g2_fill_2 FILLER_33_607 ();
 sg13g2_fill_1 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_621 ();
 sg13g2_fill_2 FILLER_33_628 ();
 sg13g2_fill_1 FILLER_33_630 ();
 sg13g2_fill_2 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_657 ();
 sg13g2_decap_8 FILLER_33_664 ();
 sg13g2_fill_1 FILLER_33_689 ();
 sg13g2_fill_1 FILLER_33_699 ();
 sg13g2_fill_1 FILLER_33_703 ();
 sg13g2_fill_2 FILLER_33_713 ();
 sg13g2_decap_4 FILLER_33_745 ();
 sg13g2_fill_2 FILLER_33_749 ();
 sg13g2_fill_1 FILLER_33_755 ();
 sg13g2_fill_2 FILLER_33_760 ();
 sg13g2_fill_1 FILLER_33_772 ();
 sg13g2_fill_2 FILLER_33_799 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_fill_2 FILLER_33_829 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_4 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_856 ();
 sg13g2_fill_1 FILLER_33_863 ();
 sg13g2_decap_8 FILLER_33_868 ();
 sg13g2_decap_4 FILLER_33_875 ();
 sg13g2_fill_2 FILLER_33_879 ();
 sg13g2_fill_2 FILLER_33_886 ();
 sg13g2_fill_1 FILLER_33_888 ();
 sg13g2_decap_4 FILLER_33_893 ();
 sg13g2_fill_2 FILLER_33_897 ();
 sg13g2_fill_1 FILLER_33_925 ();
 sg13g2_fill_1 FILLER_33_931 ();
 sg13g2_fill_2 FILLER_33_936 ();
 sg13g2_fill_1 FILLER_33_953 ();
 sg13g2_decap_8 FILLER_33_971 ();
 sg13g2_decap_8 FILLER_33_1014 ();
 sg13g2_fill_2 FILLER_33_1021 ();
 sg13g2_fill_1 FILLER_33_1023 ();
 sg13g2_fill_1 FILLER_33_1033 ();
 sg13g2_fill_2 FILLER_33_1043 ();
 sg13g2_fill_2 FILLER_33_1049 ();
 sg13g2_fill_2 FILLER_33_1056 ();
 sg13g2_fill_1 FILLER_33_1058 ();
 sg13g2_fill_1 FILLER_33_1085 ();
 sg13g2_decap_8 FILLER_33_1120 ();
 sg13g2_fill_2 FILLER_33_1127 ();
 sg13g2_fill_2 FILLER_33_1134 ();
 sg13g2_fill_1 FILLER_33_1136 ();
 sg13g2_fill_2 FILLER_33_1142 ();
 sg13g2_fill_1 FILLER_33_1144 ();
 sg13g2_fill_2 FILLER_33_1149 ();
 sg13g2_fill_1 FILLER_33_1151 ();
 sg13g2_decap_8 FILLER_33_1156 ();
 sg13g2_decap_8 FILLER_33_1163 ();
 sg13g2_decap_4 FILLER_33_1170 ();
 sg13g2_fill_1 FILLER_33_1174 ();
 sg13g2_decap_8 FILLER_33_1179 ();
 sg13g2_decap_4 FILLER_33_1186 ();
 sg13g2_decap_8 FILLER_33_1194 ();
 sg13g2_decap_8 FILLER_33_1201 ();
 sg13g2_decap_8 FILLER_33_1208 ();
 sg13g2_decap_8 FILLER_33_1215 ();
 sg13g2_decap_8 FILLER_33_1222 ();
 sg13g2_fill_1 FILLER_33_1245 ();
 sg13g2_decap_8 FILLER_33_1257 ();
 sg13g2_decap_8 FILLER_33_1264 ();
 sg13g2_fill_1 FILLER_33_1271 ();
 sg13g2_fill_2 FILLER_33_1280 ();
 sg13g2_fill_2 FILLER_33_1286 ();
 sg13g2_fill_2 FILLER_33_1314 ();
 sg13g2_fill_1 FILLER_33_1316 ();
 sg13g2_fill_1 FILLER_33_1372 ();
 sg13g2_fill_2 FILLER_33_1385 ();
 sg13g2_fill_1 FILLER_33_1387 ();
 sg13g2_decap_8 FILLER_33_1392 ();
 sg13g2_decap_8 FILLER_33_1399 ();
 sg13g2_decap_8 FILLER_33_1406 ();
 sg13g2_fill_2 FILLER_33_1413 ();
 sg13g2_fill_2 FILLER_33_1421 ();
 sg13g2_decap_8 FILLER_33_1440 ();
 sg13g2_fill_2 FILLER_33_1447 ();
 sg13g2_fill_1 FILLER_33_1449 ();
 sg13g2_decap_8 FILLER_33_1484 ();
 sg13g2_decap_8 FILLER_33_1491 ();
 sg13g2_decap_8 FILLER_33_1512 ();
 sg13g2_fill_2 FILLER_33_1519 ();
 sg13g2_fill_1 FILLER_33_1521 ();
 sg13g2_fill_1 FILLER_33_1555 ();
 sg13g2_decap_8 FILLER_33_1579 ();
 sg13g2_decap_8 FILLER_33_1586 ();
 sg13g2_decap_8 FILLER_33_1593 ();
 sg13g2_decap_8 FILLER_33_1600 ();
 sg13g2_decap_4 FILLER_33_1607 ();
 sg13g2_fill_2 FILLER_33_1622 ();
 sg13g2_decap_4 FILLER_33_1628 ();
 sg13g2_fill_1 FILLER_33_1659 ();
 sg13g2_decap_4 FILLER_33_1677 ();
 sg13g2_decap_8 FILLER_33_1703 ();
 sg13g2_decap_4 FILLER_33_1710 ();
 sg13g2_decap_8 FILLER_33_1718 ();
 sg13g2_decap_4 FILLER_33_1725 ();
 sg13g2_decap_8 FILLER_33_1733 ();
 sg13g2_decap_8 FILLER_33_1740 ();
 sg13g2_decap_8 FILLER_33_1747 ();
 sg13g2_decap_8 FILLER_33_1754 ();
 sg13g2_decap_8 FILLER_33_1761 ();
 sg13g2_decap_4 FILLER_33_1768 ();
 sg13g2_fill_2 FILLER_33_1772 ();
 sg13g2_decap_4 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_135 ();
 sg13g2_decap_8 FILLER_34_142 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_fill_2 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_fill_2 FILLER_34_309 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_4 FILLER_34_322 ();
 sg13g2_fill_2 FILLER_34_326 ();
 sg13g2_decap_4 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_decap_4 FILLER_34_370 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_453 ();
 sg13g2_decap_8 FILLER_34_460 ();
 sg13g2_fill_2 FILLER_34_467 ();
 sg13g2_fill_1 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_474 ();
 sg13g2_decap_4 FILLER_34_481 ();
 sg13g2_decap_4 FILLER_34_506 ();
 sg13g2_fill_1 FILLER_34_510 ();
 sg13g2_decap_8 FILLER_34_537 ();
 sg13g2_decap_4 FILLER_34_544 ();
 sg13g2_decap_8 FILLER_34_552 ();
 sg13g2_decap_4 FILLER_34_559 ();
 sg13g2_decap_4 FILLER_34_568 ();
 sg13g2_fill_2 FILLER_34_572 ();
 sg13g2_fill_2 FILLER_34_578 ();
 sg13g2_decap_8 FILLER_34_584 ();
 sg13g2_fill_2 FILLER_34_591 ();
 sg13g2_fill_1 FILLER_34_717 ();
 sg13g2_decap_8 FILLER_34_723 ();
 sg13g2_fill_1 FILLER_34_735 ();
 sg13g2_decap_4 FILLER_34_743 ();
 sg13g2_fill_1 FILLER_34_747 ();
 sg13g2_decap_8 FILLER_34_768 ();
 sg13g2_decap_4 FILLER_34_775 ();
 sg13g2_fill_1 FILLER_34_779 ();
 sg13g2_decap_8 FILLER_34_820 ();
 sg13g2_fill_2 FILLER_34_827 ();
 sg13g2_fill_1 FILLER_34_829 ();
 sg13g2_decap_4 FILLER_34_835 ();
 sg13g2_decap_4 FILLER_34_844 ();
 sg13g2_fill_2 FILLER_34_848 ();
 sg13g2_fill_2 FILLER_34_880 ();
 sg13g2_decap_8 FILLER_34_912 ();
 sg13g2_fill_2 FILLER_34_919 ();
 sg13g2_fill_2 FILLER_34_950 ();
 sg13g2_decap_8 FILLER_34_978 ();
 sg13g2_decap_8 FILLER_34_989 ();
 sg13g2_decap_8 FILLER_34_996 ();
 sg13g2_fill_1 FILLER_34_1003 ();
 sg13g2_fill_2 FILLER_34_1073 ();
 sg13g2_decap_4 FILLER_34_1125 ();
 sg13g2_fill_2 FILLER_34_1135 ();
 sg13g2_fill_1 FILLER_34_1137 ();
 sg13g2_fill_1 FILLER_34_1164 ();
 sg13g2_fill_1 FILLER_34_1191 ();
 sg13g2_fill_1 FILLER_34_1196 ();
 sg13g2_fill_1 FILLER_34_1205 ();
 sg13g2_decap_4 FILLER_34_1232 ();
 sg13g2_fill_2 FILLER_34_1236 ();
 sg13g2_fill_2 FILLER_34_1268 ();
 sg13g2_fill_1 FILLER_34_1304 ();
 sg13g2_fill_2 FILLER_34_1309 ();
 sg13g2_fill_1 FILLER_34_1311 ();
 sg13g2_fill_2 FILLER_34_1324 ();
 sg13g2_fill_2 FILLER_34_1330 ();
 sg13g2_fill_2 FILLER_34_1335 ();
 sg13g2_fill_2 FILLER_34_1373 ();
 sg13g2_fill_2 FILLER_34_1379 ();
 sg13g2_fill_1 FILLER_34_1421 ();
 sg13g2_decap_4 FILLER_34_1448 ();
 sg13g2_fill_2 FILLER_34_1452 ();
 sg13g2_decap_8 FILLER_34_1462 ();
 sg13g2_decap_8 FILLER_34_1469 ();
 sg13g2_fill_2 FILLER_34_1476 ();
 sg13g2_fill_2 FILLER_34_1482 ();
 sg13g2_fill_1 FILLER_34_1484 ();
 sg13g2_decap_8 FILLER_34_1489 ();
 sg13g2_decap_8 FILLER_34_1496 ();
 sg13g2_decap_8 FILLER_34_1503 ();
 sg13g2_fill_1 FILLER_34_1510 ();
 sg13g2_decap_4 FILLER_34_1524 ();
 sg13g2_fill_2 FILLER_34_1528 ();
 sg13g2_decap_4 FILLER_34_1540 ();
 sg13g2_fill_1 FILLER_34_1565 ();
 sg13g2_fill_1 FILLER_34_1575 ();
 sg13g2_decap_4 FILLER_34_1584 ();
 sg13g2_fill_1 FILLER_34_1588 ();
 sg13g2_decap_8 FILLER_34_1622 ();
 sg13g2_fill_2 FILLER_34_1638 ();
 sg13g2_decap_4 FILLER_34_1658 ();
 sg13g2_fill_2 FILLER_34_1667 ();
 sg13g2_fill_1 FILLER_34_1676 ();
 sg13g2_fill_2 FILLER_34_1687 ();
 sg13g2_fill_1 FILLER_34_1694 ();
 sg13g2_fill_2 FILLER_34_1701 ();
 sg13g2_fill_1 FILLER_34_1703 ();
 sg13g2_decap_8 FILLER_34_1748 ();
 sg13g2_decap_8 FILLER_34_1755 ();
 sg13g2_decap_8 FILLER_34_1762 ();
 sg13g2_decap_4 FILLER_34_1769 ();
 sg13g2_fill_1 FILLER_34_1773 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_36 ();
 sg13g2_decap_8 FILLER_35_41 ();
 sg13g2_decap_8 FILLER_35_48 ();
 sg13g2_decap_8 FILLER_35_59 ();
 sg13g2_decap_8 FILLER_35_66 ();
 sg13g2_fill_2 FILLER_35_73 ();
 sg13g2_decap_4 FILLER_35_96 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_165 ();
 sg13g2_decap_4 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_174 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_decap_4 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_292 ();
 sg13g2_decap_4 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_303 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_4 FILLER_35_385 ();
 sg13g2_fill_1 FILLER_35_389 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_fill_1 FILLER_35_405 ();
 sg13g2_fill_1 FILLER_35_436 ();
 sg13g2_fill_2 FILLER_35_441 ();
 sg13g2_fill_1 FILLER_35_443 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_fill_1 FILLER_35_462 ();
 sg13g2_fill_1 FILLER_35_489 ();
 sg13g2_decap_8 FILLER_35_520 ();
 sg13g2_decap_4 FILLER_35_527 ();
 sg13g2_fill_1 FILLER_35_531 ();
 sg13g2_decap_4 FILLER_35_536 ();
 sg13g2_fill_1 FILLER_35_540 ();
 sg13g2_decap_8 FILLER_35_593 ();
 sg13g2_decap_8 FILLER_35_600 ();
 sg13g2_fill_2 FILLER_35_612 ();
 sg13g2_decap_8 FILLER_35_618 ();
 sg13g2_decap_8 FILLER_35_625 ();
 sg13g2_fill_2 FILLER_35_632 ();
 sg13g2_fill_1 FILLER_35_634 ();
 sg13g2_decap_8 FILLER_35_661 ();
 sg13g2_decap_8 FILLER_35_668 ();
 sg13g2_decap_4 FILLER_35_675 ();
 sg13g2_decap_8 FILLER_35_683 ();
 sg13g2_fill_2 FILLER_35_690 ();
 sg13g2_fill_1 FILLER_35_699 ();
 sg13g2_decap_4 FILLER_35_707 ();
 sg13g2_decap_4 FILLER_35_716 ();
 sg13g2_fill_2 FILLER_35_720 ();
 sg13g2_fill_1 FILLER_35_748 ();
 sg13g2_fill_2 FILLER_35_782 ();
 sg13g2_fill_1 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_789 ();
 sg13g2_decap_4 FILLER_35_796 ();
 sg13g2_fill_2 FILLER_35_800 ();
 sg13g2_fill_1 FILLER_35_828 ();
 sg13g2_fill_2 FILLER_35_855 ();
 sg13g2_decap_8 FILLER_35_887 ();
 sg13g2_decap_8 FILLER_35_894 ();
 sg13g2_decap_4 FILLER_35_901 ();
 sg13g2_fill_1 FILLER_35_905 ();
 sg13g2_fill_2 FILLER_35_936 ();
 sg13g2_fill_1 FILLER_35_950 ();
 sg13g2_fill_1 FILLER_35_977 ();
 sg13g2_decap_4 FILLER_35_1007 ();
 sg13g2_fill_1 FILLER_35_1011 ();
 sg13g2_decap_8 FILLER_35_1016 ();
 sg13g2_fill_2 FILLER_35_1023 ();
 sg13g2_fill_1 FILLER_35_1025 ();
 sg13g2_decap_8 FILLER_35_1030 ();
 sg13g2_decap_8 FILLER_35_1037 ();
 sg13g2_fill_1 FILLER_35_1044 ();
 sg13g2_fill_2 FILLER_35_1050 ();
 sg13g2_fill_2 FILLER_35_1078 ();
 sg13g2_fill_1 FILLER_35_1100 ();
 sg13g2_fill_2 FILLER_35_1127 ();
 sg13g2_fill_2 FILLER_35_1158 ();
 sg13g2_fill_1 FILLER_35_1160 ();
 sg13g2_decap_8 FILLER_35_1165 ();
 sg13g2_decap_8 FILLER_35_1176 ();
 sg13g2_decap_8 FILLER_35_1183 ();
 sg13g2_fill_2 FILLER_35_1190 ();
 sg13g2_fill_2 FILLER_35_1201 ();
 sg13g2_fill_1 FILLER_35_1203 ();
 sg13g2_decap_4 FILLER_35_1216 ();
 sg13g2_decap_4 FILLER_35_1224 ();
 sg13g2_decap_8 FILLER_35_1237 ();
 sg13g2_decap_4 FILLER_35_1244 ();
 sg13g2_decap_8 FILLER_35_1256 ();
 sg13g2_decap_8 FILLER_35_1263 ();
 sg13g2_decap_8 FILLER_35_1286 ();
 sg13g2_decap_8 FILLER_35_1293 ();
 sg13g2_decap_8 FILLER_35_1300 ();
 sg13g2_fill_2 FILLER_35_1307 ();
 sg13g2_decap_4 FILLER_35_1327 ();
 sg13g2_fill_1 FILLER_35_1331 ();
 sg13g2_decap_4 FILLER_35_1336 ();
 sg13g2_fill_1 FILLER_35_1340 ();
 sg13g2_decap_8 FILLER_35_1344 ();
 sg13g2_decap_8 FILLER_35_1351 ();
 sg13g2_decap_8 FILLER_35_1358 ();
 sg13g2_fill_1 FILLER_35_1365 ();
 sg13g2_decap_4 FILLER_35_1370 ();
 sg13g2_decap_8 FILLER_35_1387 ();
 sg13g2_decap_4 FILLER_35_1394 ();
 sg13g2_fill_2 FILLER_35_1398 ();
 sg13g2_fill_1 FILLER_35_1417 ();
 sg13g2_decap_4 FILLER_35_1422 ();
 sg13g2_decap_8 FILLER_35_1430 ();
 sg13g2_decap_4 FILLER_35_1437 ();
 sg13g2_fill_2 FILLER_35_1441 ();
 sg13g2_fill_1 FILLER_35_1477 ();
 sg13g2_fill_2 FILLER_35_1504 ();
 sg13g2_fill_1 FILLER_35_1506 ();
 sg13g2_fill_2 FILLER_35_1524 ();
 sg13g2_fill_1 FILLER_35_1526 ();
 sg13g2_fill_1 FILLER_35_1533 ();
 sg13g2_decap_8 FILLER_35_1565 ();
 sg13g2_fill_1 FILLER_35_1572 ();
 sg13g2_fill_1 FILLER_35_1577 ();
 sg13g2_fill_1 FILLER_35_1582 ();
 sg13g2_fill_2 FILLER_35_1592 ();
 sg13g2_fill_1 FILLER_35_1594 ();
 sg13g2_fill_1 FILLER_35_1619 ();
 sg13g2_decap_8 FILLER_35_1627 ();
 sg13g2_fill_1 FILLER_35_1634 ();
 sg13g2_decap_8 FILLER_35_1640 ();
 sg13g2_decap_4 FILLER_35_1647 ();
 sg13g2_decap_8 FILLER_35_1656 ();
 sg13g2_decap_8 FILLER_35_1663 ();
 sg13g2_fill_2 FILLER_35_1670 ();
 sg13g2_decap_4 FILLER_35_1676 ();
 sg13g2_fill_1 FILLER_35_1685 ();
 sg13g2_fill_1 FILLER_35_1694 ();
 sg13g2_fill_1 FILLER_35_1711 ();
 sg13g2_decap_8 FILLER_35_1717 ();
 sg13g2_decap_4 FILLER_35_1724 ();
 sg13g2_fill_2 FILLER_35_1728 ();
 sg13g2_decap_8 FILLER_35_1760 ();
 sg13g2_decap_8 FILLER_35_1767 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_74 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_decap_8 FILLER_36_136 ();
 sg13g2_decap_4 FILLER_36_143 ();
 sg13g2_fill_2 FILLER_36_173 ();
 sg13g2_fill_1 FILLER_36_175 ();
 sg13g2_decap_4 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_201 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_decap_4 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_decap_4 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_320 ();
 sg13g2_decap_8 FILLER_36_327 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_decap_4 FILLER_36_340 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_404 ();
 sg13g2_fill_2 FILLER_36_435 ();
 sg13g2_decap_4 FILLER_36_467 ();
 sg13g2_fill_2 FILLER_36_471 ();
 sg13g2_fill_2 FILLER_36_482 ();
 sg13g2_fill_2 FILLER_36_518 ();
 sg13g2_fill_1 FILLER_36_551 ();
 sg13g2_fill_2 FILLER_36_578 ();
 sg13g2_fill_1 FILLER_36_606 ();
 sg13g2_fill_2 FILLER_36_633 ();
 sg13g2_fill_2 FILLER_36_639 ();
 sg13g2_fill_1 FILLER_36_641 ();
 sg13g2_decap_8 FILLER_36_646 ();
 sg13g2_decap_8 FILLER_36_653 ();
 sg13g2_decap_4 FILLER_36_660 ();
 sg13g2_fill_1 FILLER_36_694 ();
 sg13g2_fill_2 FILLER_36_726 ();
 sg13g2_decap_8 FILLER_36_732 ();
 sg13g2_decap_4 FILLER_36_739 ();
 sg13g2_decap_4 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_813 ();
 sg13g2_decap_4 FILLER_36_820 ();
 sg13g2_fill_1 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_829 ();
 sg13g2_fill_1 FILLER_36_836 ();
 sg13g2_fill_1 FILLER_36_841 ();
 sg13g2_fill_1 FILLER_36_868 ();
 sg13g2_fill_1 FILLER_36_882 ();
 sg13g2_fill_2 FILLER_36_891 ();
 sg13g2_decap_4 FILLER_36_897 ();
 sg13g2_decap_8 FILLER_36_922 ();
 sg13g2_fill_1 FILLER_36_929 ();
 sg13g2_fill_2 FILLER_36_935 ();
 sg13g2_fill_2 FILLER_36_964 ();
 sg13g2_decap_8 FILLER_36_975 ();
 sg13g2_decap_8 FILLER_36_982 ();
 sg13g2_decap_8 FILLER_36_989 ();
 sg13g2_decap_4 FILLER_36_996 ();
 sg13g2_fill_1 FILLER_36_1000 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_fill_2 FILLER_36_1048 ();
 sg13g2_fill_1 FILLER_36_1050 ();
 sg13g2_fill_2 FILLER_36_1077 ();
 sg13g2_fill_2 FILLER_36_1107 ();
 sg13g2_fill_1 FILLER_36_1128 ();
 sg13g2_fill_2 FILLER_36_1180 ();
 sg13g2_fill_1 FILLER_36_1182 ();
 sg13g2_decap_8 FILLER_36_1201 ();
 sg13g2_decap_8 FILLER_36_1208 ();
 sg13g2_decap_4 FILLER_36_1215 ();
 sg13g2_fill_1 FILLER_36_1219 ();
 sg13g2_fill_2 FILLER_36_1224 ();
 sg13g2_fill_1 FILLER_36_1240 ();
 sg13g2_fill_1 FILLER_36_1267 ();
 sg13g2_fill_1 FILLER_36_1297 ();
 sg13g2_decap_4 FILLER_36_1302 ();
 sg13g2_decap_8 FILLER_36_1310 ();
 sg13g2_decap_4 FILLER_36_1317 ();
 sg13g2_fill_1 FILLER_36_1321 ();
 sg13g2_decap_8 FILLER_36_1387 ();
 sg13g2_decap_8 FILLER_36_1394 ();
 sg13g2_fill_1 FILLER_36_1401 ();
 sg13g2_decap_4 FILLER_36_1445 ();
 sg13g2_fill_2 FILLER_36_1461 ();
 sg13g2_decap_4 FILLER_36_1471 ();
 sg13g2_fill_1 FILLER_36_1499 ();
 sg13g2_decap_8 FILLER_36_1504 ();
 sg13g2_decap_4 FILLER_36_1511 ();
 sg13g2_fill_1 FILLER_36_1515 ();
 sg13g2_fill_1 FILLER_36_1525 ();
 sg13g2_fill_1 FILLER_36_1557 ();
 sg13g2_fill_1 FILLER_36_1563 ();
 sg13g2_fill_2 FILLER_36_1568 ();
 sg13g2_fill_1 FILLER_36_1575 ();
 sg13g2_decap_4 FILLER_36_1581 ();
 sg13g2_fill_2 FILLER_36_1585 ();
 sg13g2_decap_8 FILLER_36_1613 ();
 sg13g2_fill_1 FILLER_36_1620 ();
 sg13g2_decap_4 FILLER_36_1651 ();
 sg13g2_fill_1 FILLER_36_1655 ();
 sg13g2_decap_4 FILLER_36_1671 ();
 sg13g2_fill_2 FILLER_36_1675 ();
 sg13g2_decap_8 FILLER_36_1682 ();
 sg13g2_fill_1 FILLER_36_1689 ();
 sg13g2_decap_8 FILLER_36_1715 ();
 sg13g2_decap_8 FILLER_36_1727 ();
 sg13g2_fill_1 FILLER_36_1734 ();
 sg13g2_decap_8 FILLER_36_1740 ();
 sg13g2_decap_4 FILLER_36_1747 ();
 sg13g2_fill_1 FILLER_36_1751 ();
 sg13g2_decap_8 FILLER_36_1756 ();
 sg13g2_decap_8 FILLER_36_1763 ();
 sg13g2_decap_4 FILLER_36_1770 ();
 sg13g2_decap_8 FILLER_37_30 ();
 sg13g2_decap_8 FILLER_37_37 ();
 sg13g2_fill_2 FILLER_37_53 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_decap_8 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_73 ();
 sg13g2_decap_4 FILLER_37_80 ();
 sg13g2_decap_8 FILLER_37_88 ();
 sg13g2_decap_8 FILLER_37_95 ();
 sg13g2_decap_8 FILLER_37_106 ();
 sg13g2_decap_4 FILLER_37_113 ();
 sg13g2_fill_1 FILLER_37_117 ();
 sg13g2_fill_2 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_153 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_172 ();
 sg13g2_fill_1 FILLER_37_174 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_decap_4 FILLER_37_204 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_decap_8 FILLER_37_213 ();
 sg13g2_decap_4 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_224 ();
 sg13g2_decap_4 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_264 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_decap_4 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_342 ();
 sg13g2_decap_4 FILLER_37_349 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_4 FILLER_37_364 ();
 sg13g2_decap_4 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_375 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_400 ();
 sg13g2_fill_1 FILLER_37_409 ();
 sg13g2_fill_1 FILLER_37_416 ();
 sg13g2_fill_1 FILLER_37_451 ();
 sg13g2_decap_8 FILLER_37_456 ();
 sg13g2_fill_1 FILLER_37_463 ();
 sg13g2_fill_1 FILLER_37_497 ();
 sg13g2_decap_4 FILLER_37_524 ();
 sg13g2_fill_2 FILLER_37_528 ();
 sg13g2_fill_1 FILLER_37_534 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_fill_1 FILLER_37_553 ();
 sg13g2_fill_1 FILLER_37_558 ();
 sg13g2_fill_2 FILLER_37_563 ();
 sg13g2_fill_1 FILLER_37_570 ();
 sg13g2_fill_2 FILLER_37_575 ();
 sg13g2_fill_2 FILLER_37_586 ();
 sg13g2_fill_2 FILLER_37_592 ();
 sg13g2_decap_8 FILLER_37_626 ();
 sg13g2_fill_1 FILLER_37_633 ();
 sg13g2_decap_8 FILLER_37_639 ();
 sg13g2_fill_2 FILLER_37_656 ();
 sg13g2_fill_2 FILLER_37_668 ();
 sg13g2_fill_2 FILLER_37_679 ();
 sg13g2_fill_1 FILLER_37_681 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_fill_2 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_699 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_fill_1 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_753 ();
 sg13g2_decap_4 FILLER_37_760 ();
 sg13g2_fill_2 FILLER_37_764 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_4 FILLER_37_784 ();
 sg13g2_fill_1 FILLER_37_788 ();
 sg13g2_decap_4 FILLER_37_793 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_fill_1 FILLER_37_819 ();
 sg13g2_fill_2 FILLER_37_830 ();
 sg13g2_fill_1 FILLER_37_832 ();
 sg13g2_fill_2 FILLER_37_859 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_fill_1 FILLER_37_908 ();
 sg13g2_fill_1 FILLER_37_968 ();
 sg13g2_fill_1 FILLER_37_995 ();
 sg13g2_decap_4 FILLER_37_1000 ();
 sg13g2_fill_2 FILLER_37_1004 ();
 sg13g2_decap_8 FILLER_37_1036 ();
 sg13g2_decap_4 FILLER_37_1043 ();
 sg13g2_decap_4 FILLER_37_1051 ();
 sg13g2_fill_1 FILLER_37_1055 ();
 sg13g2_decap_8 FILLER_37_1060 ();
 sg13g2_decap_8 FILLER_37_1067 ();
 sg13g2_fill_2 FILLER_37_1074 ();
 sg13g2_decap_8 FILLER_37_1110 ();
 sg13g2_decap_4 FILLER_37_1117 ();
 sg13g2_fill_1 FILLER_37_1121 ();
 sg13g2_decap_4 FILLER_37_1125 ();
 sg13g2_fill_1 FILLER_37_1129 ();
 sg13g2_fill_2 FILLER_37_1136 ();
 sg13g2_decap_8 FILLER_37_1150 ();
 sg13g2_fill_1 FILLER_37_1157 ();
 sg13g2_decap_8 FILLER_37_1163 ();
 sg13g2_decap_8 FILLER_37_1170 ();
 sg13g2_decap_8 FILLER_37_1177 ();
 sg13g2_decap_4 FILLER_37_1184 ();
 sg13g2_fill_1 FILLER_37_1188 ();
 sg13g2_fill_1 FILLER_37_1201 ();
 sg13g2_fill_1 FILLER_37_1210 ();
 sg13g2_fill_2 FILLER_37_1237 ();
 sg13g2_fill_2 FILLER_37_1243 ();
 sg13g2_fill_2 FILLER_37_1248 ();
 sg13g2_fill_1 FILLER_37_1250 ();
 sg13g2_decap_8 FILLER_37_1255 ();
 sg13g2_decap_8 FILLER_37_1262 ();
 sg13g2_decap_4 FILLER_37_1269 ();
 sg13g2_decap_8 FILLER_37_1277 ();
 sg13g2_decap_4 FILLER_37_1284 ();
 sg13g2_fill_1 FILLER_37_1288 ();
 sg13g2_fill_2 FILLER_37_1293 ();
 sg13g2_fill_1 FILLER_37_1295 ();
 sg13g2_decap_8 FILLER_37_1327 ();
 sg13g2_decap_8 FILLER_37_1334 ();
 sg13g2_decap_8 FILLER_37_1341 ();
 sg13g2_decap_8 FILLER_37_1348 ();
 sg13g2_fill_2 FILLER_37_1355 ();
 sg13g2_fill_1 FILLER_37_1357 ();
 sg13g2_decap_4 FILLER_37_1362 ();
 sg13g2_fill_2 FILLER_37_1366 ();
 sg13g2_fill_1 FILLER_37_1402 ();
 sg13g2_decap_4 FILLER_37_1423 ();
 sg13g2_fill_1 FILLER_37_1427 ();
 sg13g2_decap_4 FILLER_37_1432 ();
 sg13g2_fill_2 FILLER_37_1436 ();
 sg13g2_decap_8 FILLER_37_1442 ();
 sg13g2_decap_8 FILLER_37_1453 ();
 sg13g2_fill_1 FILLER_37_1460 ();
 sg13g2_decap_8 FILLER_37_1465 ();
 sg13g2_fill_2 FILLER_37_1482 ();
 sg13g2_fill_1 FILLER_37_1502 ();
 sg13g2_fill_2 FILLER_37_1529 ();
 sg13g2_decap_4 FILLER_37_1540 ();
 sg13g2_decap_4 FILLER_37_1570 ();
 sg13g2_fill_1 FILLER_37_1574 ();
 sg13g2_decap_4 FILLER_37_1579 ();
 sg13g2_decap_4 FILLER_37_1587 ();
 sg13g2_fill_2 FILLER_37_1591 ();
 sg13g2_decap_8 FILLER_37_1597 ();
 sg13g2_decap_8 FILLER_37_1604 ();
 sg13g2_decap_8 FILLER_37_1615 ();
 sg13g2_decap_4 FILLER_37_1622 ();
 sg13g2_fill_2 FILLER_37_1626 ();
 sg13g2_fill_2 FILLER_37_1632 ();
 sg13g2_decap_8 FILLER_37_1650 ();
 sg13g2_decap_4 FILLER_37_1657 ();
 sg13g2_fill_1 FILLER_37_1661 ();
 sg13g2_fill_2 FILLER_37_1666 ();
 sg13g2_decap_4 FILLER_37_1673 ();
 sg13g2_fill_2 FILLER_37_1677 ();
 sg13g2_decap_8 FILLER_37_1683 ();
 sg13g2_decap_8 FILLER_37_1694 ();
 sg13g2_decap_4 FILLER_37_1701 ();
 sg13g2_fill_1 FILLER_37_1705 ();
 sg13g2_fill_1 FILLER_37_1733 ();
 sg13g2_fill_2 FILLER_37_1740 ();
 sg13g2_fill_1 FILLER_37_1742 ();
 sg13g2_decap_4 FILLER_37_1769 ();
 sg13g2_fill_1 FILLER_37_1773 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_11 ();
 sg13g2_decap_4 FILLER_38_18 ();
 sg13g2_fill_2 FILLER_38_22 ();
 sg13g2_decap_4 FILLER_38_29 ();
 sg13g2_fill_1 FILLER_38_33 ();
 sg13g2_decap_4 FILLER_38_64 ();
 sg13g2_decap_4 FILLER_38_86 ();
 sg13g2_fill_2 FILLER_38_90 ();
 sg13g2_decap_8 FILLER_38_97 ();
 sg13g2_fill_2 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_decap_4 FILLER_38_130 ();
 sg13g2_fill_1 FILLER_38_134 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_165 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_fill_1 FILLER_38_198 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_302 ();
 sg13g2_fill_1 FILLER_38_309 ();
 sg13g2_decap_8 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_fill_1 FILLER_38_336 ();
 sg13g2_fill_1 FILLER_38_363 ();
 sg13g2_fill_2 FILLER_38_371 ();
 sg13g2_fill_2 FILLER_38_403 ();
 sg13g2_fill_1 FILLER_38_412 ();
 sg13g2_fill_1 FILLER_38_417 ();
 sg13g2_fill_1 FILLER_38_422 ();
 sg13g2_decap_8 FILLER_38_433 ();
 sg13g2_decap_8 FILLER_38_440 ();
 sg13g2_fill_1 FILLER_38_447 ();
 sg13g2_fill_2 FILLER_38_474 ();
 sg13g2_fill_2 FILLER_38_502 ();
 sg13g2_fill_1 FILLER_38_509 ();
 sg13g2_decap_8 FILLER_38_514 ();
 sg13g2_fill_2 FILLER_38_521 ();
 sg13g2_fill_1 FILLER_38_523 ();
 sg13g2_decap_8 FILLER_38_558 ();
 sg13g2_fill_2 FILLER_38_565 ();
 sg13g2_fill_1 FILLER_38_571 ();
 sg13g2_fill_1 FILLER_38_580 ();
 sg13g2_decap_8 FILLER_38_595 ();
 sg13g2_fill_1 FILLER_38_602 ();
 sg13g2_fill_1 FILLER_38_612 ();
 sg13g2_decap_8 FILLER_38_621 ();
 sg13g2_fill_2 FILLER_38_628 ();
 sg13g2_decap_8 FILLER_38_651 ();
 sg13g2_fill_2 FILLER_38_658 ();
 sg13g2_fill_1 FILLER_38_660 ();
 sg13g2_fill_1 FILLER_38_683 ();
 sg13g2_fill_2 FILLER_38_724 ();
 sg13g2_decap_4 FILLER_38_774 ();
 sg13g2_fill_2 FILLER_38_778 ();
 sg13g2_decap_4 FILLER_38_790 ();
 sg13g2_decap_8 FILLER_38_824 ();
 sg13g2_decap_4 FILLER_38_831 ();
 sg13g2_fill_1 FILLER_38_835 ();
 sg13g2_decap_8 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_fill_2 FILLER_38_858 ();
 sg13g2_fill_1 FILLER_38_860 ();
 sg13g2_decap_8 FILLER_38_879 ();
 sg13g2_decap_8 FILLER_38_886 ();
 sg13g2_decap_4 FILLER_38_897 ();
 sg13g2_fill_2 FILLER_38_964 ();
 sg13g2_fill_2 FILLER_38_991 ();
 sg13g2_fill_1 FILLER_38_993 ();
 sg13g2_fill_1 FILLER_38_1004 ();
 sg13g2_decap_8 FILLER_38_1009 ();
 sg13g2_fill_2 FILLER_38_1020 ();
 sg13g2_decap_8 FILLER_38_1026 ();
 sg13g2_decap_4 FILLER_38_1033 ();
 sg13g2_decap_4 FILLER_38_1063 ();
 sg13g2_fill_2 FILLER_38_1067 ();
 sg13g2_decap_8 FILLER_38_1158 ();
 sg13g2_fill_1 FILLER_38_1165 ();
 sg13g2_fill_2 FILLER_38_1170 ();
 sg13g2_fill_1 FILLER_38_1201 ();
 sg13g2_decap_8 FILLER_38_1215 ();
 sg13g2_decap_4 FILLER_38_1222 ();
 sg13g2_fill_1 FILLER_38_1256 ();
 sg13g2_fill_1 FILLER_38_1283 ();
 sg13g2_fill_1 FILLER_38_1310 ();
 sg13g2_fill_1 FILLER_38_1315 ();
 sg13g2_fill_2 FILLER_38_1342 ();
 sg13g2_fill_2 FILLER_38_1370 ();
 sg13g2_fill_2 FILLER_38_1393 ();
 sg13g2_fill_1 FILLER_38_1395 ();
 sg13g2_fill_2 FILLER_38_1407 ();
 sg13g2_fill_1 FILLER_38_1409 ();
 sg13g2_decap_8 FILLER_38_1415 ();
 sg13g2_decap_4 FILLER_38_1448 ();
 sg13g2_decap_8 FILLER_38_1516 ();
 sg13g2_decap_8 FILLER_38_1523 ();
 sg13g2_decap_8 FILLER_38_1530 ();
 sg13g2_decap_8 FILLER_38_1537 ();
 sg13g2_decap_8 FILLER_38_1544 ();
 sg13g2_fill_2 FILLER_38_1551 ();
 sg13g2_fill_1 FILLER_38_1553 ();
 sg13g2_decap_8 FILLER_38_1558 ();
 sg13g2_decap_8 FILLER_38_1573 ();
 sg13g2_decap_4 FILLER_38_1580 ();
 sg13g2_fill_1 FILLER_38_1584 ();
 sg13g2_fill_1 FILLER_38_1594 ();
 sg13g2_fill_1 FILLER_38_1600 ();
 sg13g2_fill_2 FILLER_38_1624 ();
 sg13g2_fill_1 FILLER_38_1626 ();
 sg13g2_fill_2 FILLER_38_1630 ();
 sg13g2_fill_1 FILLER_38_1632 ();
 sg13g2_fill_1 FILLER_38_1638 ();
 sg13g2_decap_8 FILLER_38_1652 ();
 sg13g2_fill_2 FILLER_38_1659 ();
 sg13g2_fill_1 FILLER_38_1691 ();
 sg13g2_decap_8 FILLER_38_1705 ();
 sg13g2_fill_2 FILLER_38_1727 ();
 sg13g2_decap_4 FILLER_38_1733 ();
 sg13g2_fill_1 FILLER_38_1767 ();
 sg13g2_fill_2 FILLER_38_1772 ();
 sg13g2_fill_1 FILLER_39_26 ();
 sg13g2_fill_2 FILLER_39_32 ();
 sg13g2_fill_1 FILLER_39_34 ();
 sg13g2_decap_8 FILLER_39_39 ();
 sg13g2_decap_4 FILLER_39_46 ();
 sg13g2_fill_1 FILLER_39_55 ();
 sg13g2_fill_1 FILLER_39_60 ();
 sg13g2_fill_2 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_180 ();
 sg13g2_decap_8 FILLER_39_187 ();
 sg13g2_decap_8 FILLER_39_194 ();
 sg13g2_decap_4 FILLER_39_201 ();
 sg13g2_decap_4 FILLER_39_214 ();
 sg13g2_fill_2 FILLER_39_218 ();
 sg13g2_decap_4 FILLER_39_272 ();
 sg13g2_fill_1 FILLER_39_293 ();
 sg13g2_decap_8 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_331 ();
 sg13g2_fill_2 FILLER_39_342 ();
 sg13g2_decap_4 FILLER_39_348 ();
 sg13g2_fill_2 FILLER_39_352 ();
 sg13g2_decap_4 FILLER_39_380 ();
 sg13g2_decap_8 FILLER_39_398 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_decap_4 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_421 ();
 sg13g2_decap_8 FILLER_39_428 ();
 sg13g2_fill_1 FILLER_39_435 ();
 sg13g2_fill_2 FILLER_39_441 ();
 sg13g2_fill_2 FILLER_39_448 ();
 sg13g2_fill_1 FILLER_39_450 ();
 sg13g2_fill_2 FILLER_39_456 ();
 sg13g2_decap_4 FILLER_39_462 ();
 sg13g2_decap_4 FILLER_39_526 ();
 sg13g2_decap_8 FILLER_39_539 ();
 sg13g2_decap_4 FILLER_39_546 ();
 sg13g2_fill_2 FILLER_39_563 ();
 sg13g2_decap_4 FILLER_39_599 ();
 sg13g2_fill_1 FILLER_39_603 ();
 sg13g2_fill_1 FILLER_39_634 ();
 sg13g2_fill_2 FILLER_39_680 ();
 sg13g2_fill_1 FILLER_39_690 ();
 sg13g2_decap_4 FILLER_39_701 ();
 sg13g2_decap_4 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_722 ();
 sg13g2_fill_2 FILLER_39_729 ();
 sg13g2_fill_1 FILLER_39_731 ();
 sg13g2_fill_2 FILLER_39_747 ();
 sg13g2_fill_1 FILLER_39_749 ();
 sg13g2_decap_4 FILLER_39_761 ();
 sg13g2_fill_2 FILLER_39_765 ();
 sg13g2_fill_2 FILLER_39_770 ();
 sg13g2_fill_2 FILLER_39_787 ();
 sg13g2_decap_4 FILLER_39_819 ();
 sg13g2_fill_1 FILLER_39_823 ();
 sg13g2_fill_2 FILLER_39_863 ();
 sg13g2_decap_4 FILLER_39_895 ();
 sg13g2_fill_1 FILLER_39_899 ();
 sg13g2_fill_2 FILLER_39_909 ();
 sg13g2_decap_8 FILLER_39_915 ();
 sg13g2_decap_4 FILLER_39_922 ();
 sg13g2_fill_1 FILLER_39_926 ();
 sg13g2_decap_8 FILLER_39_932 ();
 sg13g2_fill_1 FILLER_39_939 ();
 sg13g2_fill_1 FILLER_39_962 ();
 sg13g2_fill_1 FILLER_39_970 ();
 sg13g2_decap_4 FILLER_39_988 ();
 sg13g2_fill_1 FILLER_39_992 ();
 sg13g2_decap_8 FILLER_39_996 ();
 sg13g2_decap_8 FILLER_39_1003 ();
 sg13g2_decap_4 FILLER_39_1010 ();
 sg13g2_fill_2 FILLER_39_1018 ();
 sg13g2_fill_1 FILLER_39_1020 ();
 sg13g2_decap_8 FILLER_39_1036 ();
 sg13g2_fill_1 FILLER_39_1043 ();
 sg13g2_decap_8 FILLER_39_1048 ();
 sg13g2_decap_4 FILLER_39_1101 ();
 sg13g2_fill_2 FILLER_39_1105 ();
 sg13g2_decap_8 FILLER_39_1111 ();
 sg13g2_decap_8 FILLER_39_1118 ();
 sg13g2_decap_8 FILLER_39_1125 ();
 sg13g2_fill_1 FILLER_39_1132 ();
 sg13g2_fill_2 FILLER_39_1138 ();
 sg13g2_fill_1 FILLER_39_1140 ();
 sg13g2_decap_8 FILLER_39_1151 ();
 sg13g2_fill_1 FILLER_39_1158 ();
 sg13g2_fill_1 FILLER_39_1185 ();
 sg13g2_fill_2 FILLER_39_1192 ();
 sg13g2_fill_1 FILLER_39_1194 ();
 sg13g2_fill_1 FILLER_39_1231 ();
 sg13g2_decap_4 FILLER_39_1245 ();
 sg13g2_fill_1 FILLER_39_1255 ();
 sg13g2_fill_2 FILLER_39_1261 ();
 sg13g2_decap_8 FILLER_39_1267 ();
 sg13g2_decap_4 FILLER_39_1279 ();
 sg13g2_fill_1 FILLER_39_1288 ();
 sg13g2_fill_1 FILLER_39_1294 ();
 sg13g2_fill_1 FILLER_39_1299 ();
 sg13g2_fill_1 FILLER_39_1311 ();
 sg13g2_fill_1 FILLER_39_1318 ();
 sg13g2_fill_1 FILLER_39_1324 ();
 sg13g2_fill_1 FILLER_39_1330 ();
 sg13g2_decap_8 FILLER_39_1335 ();
 sg13g2_fill_2 FILLER_39_1342 ();
 sg13g2_fill_1 FILLER_39_1349 ();
 sg13g2_fill_1 FILLER_39_1354 ();
 sg13g2_fill_1 FILLER_39_1360 ();
 sg13g2_fill_2 FILLER_39_1367 ();
 sg13g2_decap_4 FILLER_39_1433 ();
 sg13g2_fill_2 FILLER_39_1437 ();
 sg13g2_decap_4 FILLER_39_1465 ();
 sg13g2_fill_1 FILLER_39_1469 ();
 sg13g2_decap_4 FILLER_39_1486 ();
 sg13g2_fill_1 FILLER_39_1498 ();
 sg13g2_decap_8 FILLER_39_1503 ();
 sg13g2_fill_2 FILLER_39_1510 ();
 sg13g2_fill_2 FILLER_39_1517 ();
 sg13g2_fill_1 FILLER_39_1519 ();
 sg13g2_decap_8 FILLER_39_1546 ();
 sg13g2_decap_8 FILLER_39_1553 ();
 sg13g2_decap_4 FILLER_39_1560 ();
 sg13g2_fill_1 FILLER_39_1603 ();
 sg13g2_fill_2 FILLER_39_1609 ();
 sg13g2_fill_2 FILLER_39_1617 ();
 sg13g2_fill_1 FILLER_39_1619 ();
 sg13g2_fill_2 FILLER_39_1624 ();
 sg13g2_fill_1 FILLER_39_1626 ();
 sg13g2_fill_2 FILLER_39_1632 ();
 sg13g2_fill_1 FILLER_39_1634 ();
 sg13g2_decap_4 FILLER_39_1661 ();
 sg13g2_fill_2 FILLER_39_1675 ();
 sg13g2_fill_1 FILLER_39_1677 ();
 sg13g2_decap_8 FILLER_39_1684 ();
 sg13g2_decap_8 FILLER_39_1691 ();
 sg13g2_fill_1 FILLER_39_1704 ();
 sg13g2_fill_1 FILLER_39_1711 ();
 sg13g2_fill_1 FILLER_39_1716 ();
 sg13g2_fill_1 FILLER_39_1722 ();
 sg13g2_fill_1 FILLER_39_1729 ();
 sg13g2_decap_8 FILLER_39_1760 ();
 sg13g2_decap_8 FILLER_39_1767 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_9 ();
 sg13g2_decap_8 FILLER_40_40 ();
 sg13g2_fill_2 FILLER_40_73 ();
 sg13g2_fill_1 FILLER_40_75 ();
 sg13g2_decap_8 FILLER_40_80 ();
 sg13g2_decap_4 FILLER_40_87 ();
 sg13g2_decap_8 FILLER_40_95 ();
 sg13g2_decap_8 FILLER_40_102 ();
 sg13g2_fill_2 FILLER_40_109 ();
 sg13g2_decap_8 FILLER_40_116 ();
 sg13g2_decap_8 FILLER_40_123 ();
 sg13g2_fill_1 FILLER_40_130 ();
 sg13g2_decap_8 FILLER_40_139 ();
 sg13g2_fill_1 FILLER_40_146 ();
 sg13g2_decap_4 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_167 ();
 sg13g2_decap_8 FILLER_40_174 ();
 sg13g2_decap_8 FILLER_40_181 ();
 sg13g2_decap_8 FILLER_40_192 ();
 sg13g2_fill_2 FILLER_40_199 ();
 sg13g2_decap_8 FILLER_40_227 ();
 sg13g2_decap_8 FILLER_40_260 ();
 sg13g2_decap_8 FILLER_40_267 ();
 sg13g2_fill_2 FILLER_40_308 ();
 sg13g2_fill_1 FILLER_40_326 ();
 sg13g2_fill_1 FILLER_40_357 ();
 sg13g2_fill_2 FILLER_40_363 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_40_385 ();
 sg13g2_fill_1 FILLER_40_394 ();
 sg13g2_decap_4 FILLER_40_436 ();
 sg13g2_fill_1 FILLER_40_479 ();
 sg13g2_fill_2 FILLER_40_494 ();
 sg13g2_fill_1 FILLER_40_507 ();
 sg13g2_decap_8 FILLER_40_518 ();
 sg13g2_fill_2 FILLER_40_525 ();
 sg13g2_fill_1 FILLER_40_527 ();
 sg13g2_decap_8 FILLER_40_533 ();
 sg13g2_fill_2 FILLER_40_540 ();
 sg13g2_fill_1 FILLER_40_542 ();
 sg13g2_decap_4 FILLER_40_580 ();
 sg13g2_fill_1 FILLER_40_584 ();
 sg13g2_decap_4 FILLER_40_604 ();
 sg13g2_fill_1 FILLER_40_608 ();
 sg13g2_decap_4 FILLER_40_634 ();
 sg13g2_fill_2 FILLER_40_647 ();
 sg13g2_fill_1 FILLER_40_649 ();
 sg13g2_decap_8 FILLER_40_663 ();
 sg13g2_fill_1 FILLER_40_670 ();
 sg13g2_decap_8 FILLER_40_677 ();
 sg13g2_decap_4 FILLER_40_684 ();
 sg13g2_fill_1 FILLER_40_688 ();
 sg13g2_decap_8 FILLER_40_699 ();
 sg13g2_fill_1 FILLER_40_706 ();
 sg13g2_fill_2 FILLER_40_742 ();
 sg13g2_fill_2 FILLER_40_748 ();
 sg13g2_fill_1 FILLER_40_750 ();
 sg13g2_decap_8 FILLER_40_755 ();
 sg13g2_decap_4 FILLER_40_762 ();
 sg13g2_fill_2 FILLER_40_766 ();
 sg13g2_fill_2 FILLER_40_777 ();
 sg13g2_fill_1 FILLER_40_779 ();
 sg13g2_fill_2 FILLER_40_785 ();
 sg13g2_fill_1 FILLER_40_791 ();
 sg13g2_fill_1 FILLER_40_814 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_decap_4 FILLER_40_840 ();
 sg13g2_fill_1 FILLER_40_844 ();
 sg13g2_fill_1 FILLER_40_856 ();
 sg13g2_fill_1 FILLER_40_887 ();
 sg13g2_fill_1 FILLER_40_892 ();
 sg13g2_fill_2 FILLER_40_896 ();
 sg13g2_fill_1 FILLER_40_898 ();
 sg13g2_decap_4 FILLER_40_922 ();
 sg13g2_fill_2 FILLER_40_959 ();
 sg13g2_fill_2 FILLER_40_1004 ();
 sg13g2_decap_4 FILLER_40_1032 ();
 sg13g2_fill_2 FILLER_40_1040 ();
 sg13g2_fill_1 FILLER_40_1042 ();
 sg13g2_fill_1 FILLER_40_1048 ();
 sg13g2_fill_2 FILLER_40_1064 ();
 sg13g2_fill_2 FILLER_40_1097 ();
 sg13g2_fill_1 FILLER_40_1099 ();
 sg13g2_fill_2 FILLER_40_1126 ();
 sg13g2_fill_2 FILLER_40_1132 ();
 sg13g2_decap_4 FILLER_40_1144 ();
 sg13g2_decap_4 FILLER_40_1156 ();
 sg13g2_fill_1 FILLER_40_1160 ();
 sg13g2_fill_2 FILLER_40_1180 ();
 sg13g2_decap_8 FILLER_40_1188 ();
 sg13g2_decap_4 FILLER_40_1195 ();
 sg13g2_fill_2 FILLER_40_1199 ();
 sg13g2_decap_4 FILLER_40_1211 ();
 sg13g2_fill_1 FILLER_40_1215 ();
 sg13g2_decap_8 FILLER_40_1248 ();
 sg13g2_decap_8 FILLER_40_1255 ();
 sg13g2_decap_4 FILLER_40_1267 ();
 sg13g2_fill_1 FILLER_40_1271 ();
 sg13g2_fill_2 FILLER_40_1277 ();
 sg13g2_fill_1 FILLER_40_1298 ();
 sg13g2_decap_4 FILLER_40_1307 ();
 sg13g2_fill_1 FILLER_40_1324 ();
 sg13g2_fill_2 FILLER_40_1330 ();
 sg13g2_fill_1 FILLER_40_1338 ();
 sg13g2_fill_2 FILLER_40_1343 ();
 sg13g2_decap_8 FILLER_40_1355 ();
 sg13g2_decap_4 FILLER_40_1362 ();
 sg13g2_fill_1 FILLER_40_1366 ();
 sg13g2_decap_8 FILLER_40_1382 ();
 sg13g2_decap_4 FILLER_40_1389 ();
 sg13g2_fill_1 FILLER_40_1393 ();
 sg13g2_fill_2 FILLER_40_1397 ();
 sg13g2_decap_8 FILLER_40_1407 ();
 sg13g2_decap_8 FILLER_40_1418 ();
 sg13g2_decap_8 FILLER_40_1425 ();
 sg13g2_fill_2 FILLER_40_1432 ();
 sg13g2_fill_1 FILLER_40_1434 ();
 sg13g2_decap_8 FILLER_40_1447 ();
 sg13g2_decap_8 FILLER_40_1454 ();
 sg13g2_fill_2 FILLER_40_1461 ();
 sg13g2_fill_2 FILLER_40_1471 ();
 sg13g2_fill_1 FILLER_40_1478 ();
 sg13g2_decap_4 FILLER_40_1517 ();
 sg13g2_fill_2 FILLER_40_1521 ();
 sg13g2_fill_1 FILLER_40_1526 ();
 sg13g2_decap_8 FILLER_40_1548 ();
 sg13g2_decap_8 FILLER_40_1555 ();
 sg13g2_decap_8 FILLER_40_1562 ();
 sg13g2_decap_8 FILLER_40_1569 ();
 sg13g2_decap_8 FILLER_40_1576 ();
 sg13g2_decap_8 FILLER_40_1583 ();
 sg13g2_fill_1 FILLER_40_1590 ();
 sg13g2_fill_1 FILLER_40_1597 ();
 sg13g2_decap_4 FILLER_40_1604 ();
 sg13g2_fill_1 FILLER_40_1612 ();
 sg13g2_fill_2 FILLER_40_1647 ();
 sg13g2_fill_1 FILLER_40_1649 ();
 sg13g2_decap_8 FILLER_40_1662 ();
 sg13g2_decap_4 FILLER_40_1669 ();
 sg13g2_fill_1 FILLER_40_1696 ();
 sg13g2_decap_8 FILLER_40_1703 ();
 sg13g2_fill_1 FILLER_40_1710 ();
 sg13g2_decap_8 FILLER_40_1715 ();
 sg13g2_decap_4 FILLER_40_1722 ();
 sg13g2_decap_4 FILLER_40_1730 ();
 sg13g2_fill_2 FILLER_40_1734 ();
 sg13g2_decap_8 FILLER_40_1740 ();
 sg13g2_decap_8 FILLER_40_1747 ();
 sg13g2_decap_8 FILLER_40_1754 ();
 sg13g2_decap_8 FILLER_40_1761 ();
 sg13g2_decap_4 FILLER_40_1768 ();
 sg13g2_fill_2 FILLER_40_1772 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_4 FILLER_41_28 ();
 sg13g2_fill_2 FILLER_41_32 ();
 sg13g2_decap_8 FILLER_41_38 ();
 sg13g2_decap_8 FILLER_41_45 ();
 sg13g2_fill_2 FILLER_41_52 ();
 sg13g2_decap_4 FILLER_41_80 ();
 sg13g2_decap_8 FILLER_41_110 ();
 sg13g2_decap_8 FILLER_41_117 ();
 sg13g2_decap_4 FILLER_41_124 ();
 sg13g2_fill_2 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_212 ();
 sg13g2_decap_8 FILLER_41_219 ();
 sg13g2_fill_1 FILLER_41_226 ();
 sg13g2_decap_4 FILLER_41_239 ();
 sg13g2_decap_8 FILLER_41_247 ();
 sg13g2_fill_2 FILLER_41_254 ();
 sg13g2_fill_1 FILLER_41_256 ();
 sg13g2_decap_8 FILLER_41_261 ();
 sg13g2_decap_8 FILLER_41_268 ();
 sg13g2_decap_4 FILLER_41_275 ();
 sg13g2_fill_2 FILLER_41_318 ();
 sg13g2_fill_1 FILLER_41_325 ();
 sg13g2_fill_2 FILLER_41_334 ();
 sg13g2_fill_2 FILLER_41_341 ();
 sg13g2_fill_1 FILLER_41_343 ();
 sg13g2_fill_2 FILLER_41_349 ();
 sg13g2_fill_1 FILLER_41_351 ();
 sg13g2_fill_2 FILLER_41_356 ();
 sg13g2_fill_1 FILLER_41_374 ();
 sg13g2_decap_8 FILLER_41_405 ();
 sg13g2_fill_2 FILLER_41_430 ();
 sg13g2_decap_8 FILLER_41_438 ();
 sg13g2_fill_2 FILLER_41_445 ();
 sg13g2_fill_1 FILLER_41_447 ();
 sg13g2_decap_8 FILLER_41_452 ();
 sg13g2_decap_4 FILLER_41_463 ();
 sg13g2_fill_1 FILLER_41_467 ();
 sg13g2_decap_8 FILLER_41_473 ();
 sg13g2_decap_4 FILLER_41_480 ();
 sg13g2_fill_2 FILLER_41_484 ();
 sg13g2_decap_4 FILLER_41_501 ();
 sg13g2_fill_2 FILLER_41_505 ();
 sg13g2_decap_8 FILLER_41_519 ();
 sg13g2_decap_4 FILLER_41_526 ();
 sg13g2_fill_1 FILLER_41_530 ();
 sg13g2_decap_8 FILLER_41_536 ();
 sg13g2_decap_8 FILLER_41_543 ();
 sg13g2_decap_4 FILLER_41_550 ();
 sg13g2_fill_2 FILLER_41_554 ();
 sg13g2_fill_2 FILLER_41_564 ();
 sg13g2_fill_1 FILLER_41_571 ();
 sg13g2_decap_8 FILLER_41_576 ();
 sg13g2_decap_4 FILLER_41_583 ();
 sg13g2_fill_2 FILLER_41_587 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_fill_1 FILLER_41_602 ();
 sg13g2_fill_1 FILLER_41_629 ();
 sg13g2_fill_1 FILLER_41_634 ();
 sg13g2_fill_2 FILLER_41_640 ();
 sg13g2_fill_2 FILLER_41_646 ();
 sg13g2_fill_1 FILLER_41_648 ();
 sg13g2_fill_1 FILLER_41_653 ();
 sg13g2_fill_2 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_682 ();
 sg13g2_decap_4 FILLER_41_687 ();
 sg13g2_fill_1 FILLER_41_691 ();
 sg13g2_decap_8 FILLER_41_696 ();
 sg13g2_decap_8 FILLER_41_703 ();
 sg13g2_decap_8 FILLER_41_710 ();
 sg13g2_decap_8 FILLER_41_717 ();
 sg13g2_fill_2 FILLER_41_724 ();
 sg13g2_fill_1 FILLER_41_726 ();
 sg13g2_decap_8 FILLER_41_811 ();
 sg13g2_decap_8 FILLER_41_818 ();
 sg13g2_decap_4 FILLER_41_825 ();
 sg13g2_fill_2 FILLER_41_829 ();
 sg13g2_decap_4 FILLER_41_835 ();
 sg13g2_fill_2 FILLER_41_844 ();
 sg13g2_decap_4 FILLER_41_850 ();
 sg13g2_fill_1 FILLER_41_859 ();
 sg13g2_fill_2 FILLER_41_864 ();
 sg13g2_decap_4 FILLER_41_911 ();
 sg13g2_fill_1 FILLER_41_915 ();
 sg13g2_decap_8 FILLER_41_920 ();
 sg13g2_decap_8 FILLER_41_927 ();
 sg13g2_decap_8 FILLER_41_934 ();
 sg13g2_decap_8 FILLER_41_941 ();
 sg13g2_decap_4 FILLER_41_971 ();
 sg13g2_fill_2 FILLER_41_980 ();
 sg13g2_fill_1 FILLER_41_982 ();
 sg13g2_decap_4 FILLER_41_1018 ();
 sg13g2_fill_2 FILLER_41_1022 ();
 sg13g2_decap_8 FILLER_41_1054 ();
 sg13g2_decap_4 FILLER_41_1061 ();
 sg13g2_fill_1 FILLER_41_1065 ();
 sg13g2_decap_4 FILLER_41_1071 ();
 sg13g2_fill_1 FILLER_41_1075 ();
 sg13g2_fill_2 FILLER_41_1080 ();
 sg13g2_fill_1 FILLER_41_1082 ();
 sg13g2_decap_8 FILLER_41_1087 ();
 sg13g2_decap_4 FILLER_41_1094 ();
 sg13g2_fill_1 FILLER_41_1098 ();
 sg13g2_decap_8 FILLER_41_1104 ();
 sg13g2_fill_2 FILLER_41_1111 ();
 sg13g2_fill_1 FILLER_41_1113 ();
 sg13g2_fill_2 FILLER_41_1117 ();
 sg13g2_decap_4 FILLER_41_1123 ();
 sg13g2_fill_2 FILLER_41_1127 ();
 sg13g2_fill_2 FILLER_41_1141 ();
 sg13g2_fill_2 FILLER_41_1252 ();
 sg13g2_fill_2 FILLER_41_1294 ();
 sg13g2_fill_2 FILLER_41_1322 ();
 sg13g2_fill_2 FILLER_41_1355 ();
 sg13g2_fill_1 FILLER_41_1357 ();
 sg13g2_decap_8 FILLER_41_1389 ();
 sg13g2_fill_2 FILLER_41_1396 ();
 sg13g2_fill_1 FILLER_41_1398 ();
 sg13g2_decap_4 FILLER_41_1407 ();
 sg13g2_fill_1 FILLER_41_1411 ();
 sg13g2_decap_8 FILLER_41_1417 ();
 sg13g2_decap_8 FILLER_41_1424 ();
 sg13g2_fill_1 FILLER_41_1431 ();
 sg13g2_decap_8 FILLER_41_1457 ();
 sg13g2_decap_8 FILLER_41_1464 ();
 sg13g2_fill_2 FILLER_41_1471 ();
 sg13g2_decap_8 FILLER_41_1481 ();
 sg13g2_decap_8 FILLER_41_1488 ();
 sg13g2_decap_4 FILLER_41_1495 ();
 sg13g2_fill_1 FILLER_41_1499 ();
 sg13g2_fill_2 FILLER_41_1508 ();
 sg13g2_fill_1 FILLER_41_1526 ();
 sg13g2_fill_2 FILLER_41_1562 ();
 sg13g2_fill_1 FILLER_41_1564 ();
 sg13g2_decap_4 FILLER_41_1595 ();
 sg13g2_fill_1 FILLER_41_1599 ();
 sg13g2_decap_8 FILLER_41_1606 ();
 sg13g2_decap_4 FILLER_41_1613 ();
 sg13g2_fill_2 FILLER_41_1617 ();
 sg13g2_decap_8 FILLER_41_1623 ();
 sg13g2_decap_8 FILLER_41_1630 ();
 sg13g2_fill_1 FILLER_41_1637 ();
 sg13g2_decap_8 FILLER_41_1668 ();
 sg13g2_decap_8 FILLER_41_1675 ();
 sg13g2_decap_4 FILLER_41_1682 ();
 sg13g2_fill_1 FILLER_41_1686 ();
 sg13g2_decap_8 FILLER_41_1697 ();
 sg13g2_decap_8 FILLER_41_1734 ();
 sg13g2_decap_4 FILLER_41_1741 ();
 sg13g2_fill_1 FILLER_41_1745 ();
 sg13g2_fill_2 FILLER_41_1772 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_4 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_25 ();
 sg13g2_fill_2 FILLER_42_57 ();
 sg13g2_fill_1 FILLER_42_59 ();
 sg13g2_decap_8 FILLER_42_64 ();
 sg13g2_fill_2 FILLER_42_71 ();
 sg13g2_fill_1 FILLER_42_73 ();
 sg13g2_fill_2 FILLER_42_105 ();
 sg13g2_fill_1 FILLER_42_107 ();
 sg13g2_decap_8 FILLER_42_157 ();
 sg13g2_decap_8 FILLER_42_164 ();
 sg13g2_decap_8 FILLER_42_171 ();
 sg13g2_decap_4 FILLER_42_178 ();
 sg13g2_fill_1 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_188 ();
 sg13g2_decap_4 FILLER_42_200 ();
 sg13g2_fill_2 FILLER_42_209 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_decap_8 FILLER_42_232 ();
 sg13g2_fill_2 FILLER_42_239 ();
 sg13g2_fill_1 FILLER_42_256 ();
 sg13g2_decap_8 FILLER_42_270 ();
 sg13g2_decap_8 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_299 ();
 sg13g2_fill_2 FILLER_42_305 ();
 sg13g2_fill_1 FILLER_42_307 ();
 sg13g2_decap_4 FILLER_42_321 ();
 sg13g2_fill_1 FILLER_42_335 ();
 sg13g2_fill_2 FILLER_42_349 ();
 sg13g2_fill_1 FILLER_42_351 ();
 sg13g2_fill_2 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_370 ();
 sg13g2_decap_8 FILLER_42_377 ();
 sg13g2_fill_2 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_fill_2 FILLER_42_413 ();
 sg13g2_fill_2 FILLER_42_445 ();
 sg13g2_fill_2 FILLER_42_452 ();
 sg13g2_fill_1 FILLER_42_454 ();
 sg13g2_decap_8 FILLER_42_465 ();
 sg13g2_fill_1 FILLER_42_472 ();
 sg13g2_fill_1 FILLER_42_480 ();
 sg13g2_fill_2 FILLER_42_486 ();
 sg13g2_fill_2 FILLER_42_493 ();
 sg13g2_fill_2 FILLER_42_500 ();
 sg13g2_decap_4 FILLER_42_514 ();
 sg13g2_fill_1 FILLER_42_518 ();
 sg13g2_decap_4 FILLER_42_523 ();
 sg13g2_fill_1 FILLER_42_527 ();
 sg13g2_decap_8 FILLER_42_533 ();
 sg13g2_decap_4 FILLER_42_540 ();
 sg13g2_fill_1 FILLER_42_592 ();
 sg13g2_fill_2 FILLER_42_598 ();
 sg13g2_fill_1 FILLER_42_600 ();
 sg13g2_fill_2 FILLER_42_645 ();
 sg13g2_fill_1 FILLER_42_647 ();
 sg13g2_decap_8 FILLER_42_671 ();
 sg13g2_fill_1 FILLER_42_678 ();
 sg13g2_fill_2 FILLER_42_714 ();
 sg13g2_decap_8 FILLER_42_747 ();
 sg13g2_decap_4 FILLER_42_754 ();
 sg13g2_decap_8 FILLER_42_761 ();
 sg13g2_fill_2 FILLER_42_775 ();
 sg13g2_fill_1 FILLER_42_777 ();
 sg13g2_fill_1 FILLER_42_782 ();
 sg13g2_decap_8 FILLER_42_813 ();
 sg13g2_decap_4 FILLER_42_820 ();
 sg13g2_fill_2 FILLER_42_850 ();
 sg13g2_fill_1 FILLER_42_852 ();
 sg13g2_fill_1 FILLER_42_879 ();
 sg13g2_fill_2 FILLER_42_897 ();
 sg13g2_fill_1 FILLER_42_899 ();
 sg13g2_decap_4 FILLER_42_920 ();
 sg13g2_fill_1 FILLER_42_924 ();
 sg13g2_fill_1 FILLER_42_929 ();
 sg13g2_decap_4 FILLER_42_942 ();
 sg13g2_fill_1 FILLER_42_946 ();
 sg13g2_fill_2 FILLER_42_952 ();
 sg13g2_fill_1 FILLER_42_998 ();
 sg13g2_decap_4 FILLER_42_1035 ();
 sg13g2_fill_2 FILLER_42_1039 ();
 sg13g2_fill_1 FILLER_42_1044 ();
 sg13g2_decap_4 FILLER_42_1058 ();
 sg13g2_fill_2 FILLER_42_1062 ();
 sg13g2_fill_1 FILLER_42_1099 ();
 sg13g2_fill_2 FILLER_42_1135 ();
 sg13g2_fill_1 FILLER_42_1137 ();
 sg13g2_decap_8 FILLER_42_1155 ();
 sg13g2_fill_2 FILLER_42_1162 ();
 sg13g2_fill_1 FILLER_42_1164 ();
 sg13g2_decap_8 FILLER_42_1182 ();
 sg13g2_decap_8 FILLER_42_1189 ();
 sg13g2_decap_8 FILLER_42_1200 ();
 sg13g2_decap_8 FILLER_42_1211 ();
 sg13g2_fill_2 FILLER_42_1227 ();
 sg13g2_fill_1 FILLER_42_1229 ();
 sg13g2_fill_2 FILLER_42_1235 ();
 sg13g2_decap_4 FILLER_42_1242 ();
 sg13g2_decap_4 FILLER_42_1252 ();
 sg13g2_decap_4 FILLER_42_1260 ();
 sg13g2_decap_8 FILLER_42_1268 ();
 sg13g2_fill_2 FILLER_42_1275 ();
 sg13g2_decap_8 FILLER_42_1287 ();
 sg13g2_fill_2 FILLER_42_1299 ();
 sg13g2_decap_8 FILLER_42_1306 ();
 sg13g2_fill_1 FILLER_42_1322 ();
 sg13g2_fill_1 FILLER_42_1327 ();
 sg13g2_decap_8 FILLER_42_1332 ();
 sg13g2_decap_4 FILLER_42_1339 ();
 sg13g2_fill_1 FILLER_42_1343 ();
 sg13g2_decap_8 FILLER_42_1348 ();
 sg13g2_fill_2 FILLER_42_1355 ();
 sg13g2_decap_8 FILLER_42_1361 ();
 sg13g2_fill_2 FILLER_42_1368 ();
 sg13g2_decap_8 FILLER_42_1374 ();
 sg13g2_decap_8 FILLER_42_1381 ();
 sg13g2_fill_2 FILLER_42_1388 ();
 sg13g2_fill_2 FILLER_42_1420 ();
 sg13g2_fill_1 FILLER_42_1422 ();
 sg13g2_decap_4 FILLER_42_1428 ();
 sg13g2_fill_1 FILLER_42_1432 ();
 sg13g2_fill_1 FILLER_42_1441 ();
 sg13g2_decap_4 FILLER_42_1468 ();
 sg13g2_fill_2 FILLER_42_1480 ();
 sg13g2_fill_1 FILLER_42_1482 ();
 sg13g2_decap_8 FILLER_42_1486 ();
 sg13g2_decap_8 FILLER_42_1493 ();
 sg13g2_fill_2 FILLER_42_1500 ();
 sg13g2_fill_2 FILLER_42_1510 ();
 sg13g2_fill_1 FILLER_42_1512 ();
 sg13g2_decap_4 FILLER_42_1519 ();
 sg13g2_decap_8 FILLER_42_1554 ();
 sg13g2_decap_8 FILLER_42_1561 ();
 sg13g2_fill_2 FILLER_42_1568 ();
 sg13g2_fill_1 FILLER_42_1570 ();
 sg13g2_decap_8 FILLER_42_1576 ();
 sg13g2_decap_4 FILLER_42_1583 ();
 sg13g2_fill_1 FILLER_42_1587 ();
 sg13g2_decap_8 FILLER_42_1593 ();
 sg13g2_fill_2 FILLER_42_1600 ();
 sg13g2_fill_1 FILLER_42_1602 ();
 sg13g2_decap_8 FILLER_42_1639 ();
 sg13g2_decap_8 FILLER_42_1655 ();
 sg13g2_decap_4 FILLER_42_1662 ();
 sg13g2_fill_2 FILLER_42_1666 ();
 sg13g2_fill_2 FILLER_42_1673 ();
 sg13g2_decap_8 FILLER_42_1690 ();
 sg13g2_fill_2 FILLER_42_1697 ();
 sg13g2_fill_1 FILLER_42_1717 ();
 sg13g2_fill_1 FILLER_42_1731 ();
 sg13g2_fill_1 FILLER_42_1736 ();
 sg13g2_decap_4 FILLER_42_1747 ();
 sg13g2_fill_1 FILLER_42_1751 ();
 sg13g2_decap_4 FILLER_42_1756 ();
 sg13g2_fill_2 FILLER_42_1760 ();
 sg13g2_decap_8 FILLER_42_1766 ();
 sg13g2_fill_1 FILLER_42_1773 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_fill_1 FILLER_43_49 ();
 sg13g2_decap_4 FILLER_43_60 ();
 sg13g2_fill_2 FILLER_43_64 ();
 sg13g2_decap_8 FILLER_43_78 ();
 sg13g2_decap_8 FILLER_43_89 ();
 sg13g2_decap_8 FILLER_43_96 ();
 sg13g2_fill_1 FILLER_43_103 ();
 sg13g2_decap_4 FILLER_43_122 ();
 sg13g2_fill_1 FILLER_43_126 ();
 sg13g2_decap_4 FILLER_43_135 ();
 sg13g2_fill_1 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_149 ();
 sg13g2_decap_8 FILLER_43_163 ();
 sg13g2_fill_2 FILLER_43_170 ();
 sg13g2_fill_1 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_178 ();
 sg13g2_fill_2 FILLER_43_186 ();
 sg13g2_fill_1 FILLER_43_188 ();
 sg13g2_fill_2 FILLER_43_194 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_fill_2 FILLER_43_217 ();
 sg13g2_fill_1 FILLER_43_219 ();
 sg13g2_decap_8 FILLER_43_225 ();
 sg13g2_fill_2 FILLER_43_232 ();
 sg13g2_fill_1 FILLER_43_234 ();
 sg13g2_decap_4 FILLER_43_239 ();
 sg13g2_fill_2 FILLER_43_247 ();
 sg13g2_decap_4 FILLER_43_254 ();
 sg13g2_decap_4 FILLER_43_278 ();
 sg13g2_fill_2 FILLER_43_282 ();
 sg13g2_decap_8 FILLER_43_289 ();
 sg13g2_fill_1 FILLER_43_296 ();
 sg13g2_decap_8 FILLER_43_302 ();
 sg13g2_decap_8 FILLER_43_309 ();
 sg13g2_fill_2 FILLER_43_316 ();
 sg13g2_fill_1 FILLER_43_318 ();
 sg13g2_fill_2 FILLER_43_323 ();
 sg13g2_fill_1 FILLER_43_325 ();
 sg13g2_fill_2 FILLER_43_331 ();
 sg13g2_fill_2 FILLER_43_352 ();
 sg13g2_decap_4 FILLER_43_374 ();
 sg13g2_fill_2 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_390 ();
 sg13g2_decap_4 FILLER_43_397 ();
 sg13g2_fill_1 FILLER_43_401 ();
 sg13g2_decap_4 FILLER_43_414 ();
 sg13g2_fill_1 FILLER_43_430 ();
 sg13g2_decap_8 FILLER_43_443 ();
 sg13g2_decap_8 FILLER_43_450 ();
 sg13g2_decap_4 FILLER_43_457 ();
 sg13g2_fill_2 FILLER_43_471 ();
 sg13g2_decap_4 FILLER_43_477 ();
 sg13g2_decap_8 FILLER_43_486 ();
 sg13g2_decap_8 FILLER_43_493 ();
 sg13g2_decap_4 FILLER_43_500 ();
 sg13g2_fill_2 FILLER_43_504 ();
 sg13g2_decap_4 FILLER_43_525 ();
 sg13g2_fill_1 FILLER_43_529 ();
 sg13g2_fill_1 FILLER_43_549 ();
 sg13g2_decap_4 FILLER_43_554 ();
 sg13g2_fill_2 FILLER_43_567 ();
 sg13g2_fill_1 FILLER_43_573 ();
 sg13g2_decap_4 FILLER_43_578 ();
 sg13g2_decap_8 FILLER_43_586 ();
 sg13g2_fill_1 FILLER_43_593 ();
 sg13g2_fill_1 FILLER_43_609 ();
 sg13g2_decap_4 FILLER_43_641 ();
 sg13g2_fill_1 FILLER_43_645 ();
 sg13g2_decap_8 FILLER_43_655 ();
 sg13g2_decap_8 FILLER_43_662 ();
 sg13g2_fill_1 FILLER_43_727 ();
 sg13g2_decap_4 FILLER_43_787 ();
 sg13g2_fill_2 FILLER_43_791 ();
 sg13g2_fill_1 FILLER_43_797 ();
 sg13g2_fill_2 FILLER_43_824 ();
 sg13g2_decap_4 FILLER_43_830 ();
 sg13g2_fill_2 FILLER_43_834 ();
 sg13g2_fill_2 FILLER_43_845 ();
 sg13g2_fill_1 FILLER_43_847 ();
 sg13g2_fill_1 FILLER_43_853 ();
 sg13g2_fill_1 FILLER_43_859 ();
 sg13g2_fill_2 FILLER_43_865 ();
 sg13g2_fill_2 FILLER_43_872 ();
 sg13g2_fill_2 FILLER_43_879 ();
 sg13g2_fill_1 FILLER_43_881 ();
 sg13g2_fill_1 FILLER_43_887 ();
 sg13g2_decap_8 FILLER_43_892 ();
 sg13g2_decap_4 FILLER_43_899 ();
 sg13g2_fill_1 FILLER_43_907 ();
 sg13g2_fill_2 FILLER_43_963 ();
 sg13g2_fill_1 FILLER_43_978 ();
 sg13g2_decap_4 FILLER_43_988 ();
 sg13g2_fill_1 FILLER_43_997 ();
 sg13g2_decap_4 FILLER_43_1016 ();
 sg13g2_fill_1 FILLER_43_1020 ();
 sg13g2_fill_1 FILLER_43_1025 ();
 sg13g2_fill_1 FILLER_43_1048 ();
 sg13g2_fill_1 FILLER_43_1068 ();
 sg13g2_fill_2 FILLER_43_1083 ();
 sg13g2_decap_4 FILLER_43_1108 ();
 sg13g2_decap_8 FILLER_43_1116 ();
 sg13g2_decap_4 FILLER_43_1123 ();
 sg13g2_fill_1 FILLER_43_1146 ();
 sg13g2_fill_1 FILLER_43_1152 ();
 sg13g2_fill_2 FILLER_43_1157 ();
 sg13g2_fill_1 FILLER_43_1159 ();
 sg13g2_decap_4 FILLER_43_1170 ();
 sg13g2_fill_1 FILLER_43_1174 ();
 sg13g2_decap_8 FILLER_43_1180 ();
 sg13g2_decap_4 FILLER_43_1187 ();
 sg13g2_fill_2 FILLER_43_1191 ();
 sg13g2_decap_4 FILLER_43_1198 ();
 sg13g2_fill_1 FILLER_43_1215 ();
 sg13g2_decap_4 FILLER_43_1224 ();
 sg13g2_fill_1 FILLER_43_1228 ();
 sg13g2_fill_1 FILLER_43_1233 ();
 sg13g2_decap_8 FILLER_43_1238 ();
 sg13g2_decap_8 FILLER_43_1258 ();
 sg13g2_decap_4 FILLER_43_1265 ();
 sg13g2_fill_2 FILLER_43_1274 ();
 sg13g2_fill_1 FILLER_43_1276 ();
 sg13g2_decap_4 FILLER_43_1281 ();
 sg13g2_fill_1 FILLER_43_1285 ();
 sg13g2_decap_8 FILLER_43_1295 ();
 sg13g2_decap_8 FILLER_43_1302 ();
 sg13g2_fill_2 FILLER_43_1309 ();
 sg13g2_fill_1 FILLER_43_1311 ();
 sg13g2_fill_2 FILLER_43_1347 ();
 sg13g2_fill_1 FILLER_43_1349 ();
 sg13g2_fill_2 FILLER_43_1395 ();
 sg13g2_fill_2 FILLER_43_1402 ();
 sg13g2_fill_1 FILLER_43_1404 ();
 sg13g2_fill_1 FILLER_43_1409 ();
 sg13g2_fill_2 FILLER_43_1416 ();
 sg13g2_fill_1 FILLER_43_1418 ();
 sg13g2_fill_1 FILLER_43_1424 ();
 sg13g2_fill_1 FILLER_43_1512 ();
 sg13g2_decap_8 FILLER_43_1526 ();
 sg13g2_fill_2 FILLER_43_1533 ();
 sg13g2_decap_8 FILLER_43_1539 ();
 sg13g2_decap_8 FILLER_43_1546 ();
 sg13g2_decap_4 FILLER_43_1553 ();
 sg13g2_fill_1 FILLER_43_1557 ();
 sg13g2_decap_4 FILLER_43_1604 ();
 sg13g2_fill_1 FILLER_43_1608 ();
 sg13g2_fill_1 FILLER_43_1621 ();
 sg13g2_decap_8 FILLER_43_1631 ();
 sg13g2_decap_4 FILLER_43_1638 ();
 sg13g2_fill_2 FILLER_43_1642 ();
 sg13g2_fill_1 FILLER_43_1653 ();
 sg13g2_fill_2 FILLER_43_1664 ();
 sg13g2_fill_1 FILLER_43_1666 ();
 sg13g2_fill_2 FILLER_43_1672 ();
 sg13g2_fill_1 FILLER_43_1674 ();
 sg13g2_decap_4 FILLER_43_1698 ();
 sg13g2_fill_1 FILLER_43_1707 ();
 sg13g2_decap_8 FILLER_43_1713 ();
 sg13g2_fill_1 FILLER_43_1724 ();
 sg13g2_fill_1 FILLER_43_1730 ();
 sg13g2_fill_2 FILLER_43_1739 ();
 sg13g2_decap_8 FILLER_43_1746 ();
 sg13g2_fill_2 FILLER_43_1753 ();
 sg13g2_decap_8 FILLER_43_1759 ();
 sg13g2_decap_8 FILLER_43_1766 ();
 sg13g2_fill_1 FILLER_43_1773 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_fill_2 FILLER_44_49 ();
 sg13g2_fill_1 FILLER_44_51 ();
 sg13g2_fill_1 FILLER_44_61 ();
 sg13g2_fill_1 FILLER_44_72 ();
 sg13g2_decap_4 FILLER_44_77 ();
 sg13g2_fill_1 FILLER_44_81 ();
 sg13g2_decap_8 FILLER_44_86 ();
 sg13g2_decap_8 FILLER_44_93 ();
 sg13g2_fill_2 FILLER_44_100 ();
 sg13g2_fill_1 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_115 ();
 sg13g2_decap_8 FILLER_44_122 ();
 sg13g2_decap_4 FILLER_44_129 ();
 sg13g2_fill_1 FILLER_44_138 ();
 sg13g2_decap_8 FILLER_44_170 ();
 sg13g2_decap_4 FILLER_44_177 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_4 FILLER_44_200 ();
 sg13g2_fill_2 FILLER_44_204 ();
 sg13g2_decap_8 FILLER_44_242 ();
 sg13g2_decap_8 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_256 ();
 sg13g2_decap_8 FILLER_44_263 ();
 sg13g2_fill_2 FILLER_44_270 ();
 sg13g2_fill_1 FILLER_44_272 ();
 sg13g2_fill_1 FILLER_44_278 ();
 sg13g2_decap_4 FILLER_44_286 ();
 sg13g2_fill_2 FILLER_44_290 ();
 sg13g2_fill_1 FILLER_44_302 ();
 sg13g2_decap_4 FILLER_44_318 ();
 sg13g2_fill_1 FILLER_44_322 ();
 sg13g2_fill_2 FILLER_44_339 ();
 sg13g2_fill_2 FILLER_44_375 ();
 sg13g2_fill_1 FILLER_44_377 ();
 sg13g2_decap_4 FILLER_44_381 ();
 sg13g2_decap_4 FILLER_44_389 ();
 sg13g2_fill_1 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_4 FILLER_44_413 ();
 sg13g2_fill_2 FILLER_44_417 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_451 ();
 sg13g2_decap_8 FILLER_44_458 ();
 sg13g2_decap_8 FILLER_44_465 ();
 sg13g2_decap_4 FILLER_44_484 ();
 sg13g2_fill_1 FILLER_44_488 ();
 sg13g2_decap_8 FILLER_44_499 ();
 sg13g2_fill_2 FILLER_44_509 ();
 sg13g2_fill_2 FILLER_44_523 ();
 sg13g2_decap_4 FILLER_44_532 ();
 sg13g2_fill_2 FILLER_44_536 ();
 sg13g2_decap_8 FILLER_44_543 ();
 sg13g2_decap_4 FILLER_44_550 ();
 sg13g2_decap_8 FILLER_44_566 ();
 sg13g2_fill_2 FILLER_44_573 ();
 sg13g2_decap_4 FILLER_44_588 ();
 sg13g2_fill_2 FILLER_44_601 ();
 sg13g2_decap_8 FILLER_44_614 ();
 sg13g2_decap_8 FILLER_44_625 ();
 sg13g2_decap_4 FILLER_44_632 ();
 sg13g2_fill_2 FILLER_44_636 ();
 sg13g2_fill_2 FILLER_44_668 ();
 sg13g2_fill_1 FILLER_44_701 ();
 sg13g2_decap_8 FILLER_44_715 ();
 sg13g2_decap_8 FILLER_44_722 ();
 sg13g2_decap_8 FILLER_44_729 ();
 sg13g2_decap_8 FILLER_44_736 ();
 sg13g2_decap_8 FILLER_44_743 ();
 sg13g2_decap_4 FILLER_44_750 ();
 sg13g2_fill_1 FILLER_44_754 ();
 sg13g2_fill_2 FILLER_44_764 ();
 sg13g2_decap_8 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_4 FILLER_44_784 ();
 sg13g2_fill_2 FILLER_44_802 ();
 sg13g2_decap_4 FILLER_44_809 ();
 sg13g2_fill_2 FILLER_44_813 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_fill_1 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_832 ();
 sg13g2_fill_2 FILLER_44_839 ();
 sg13g2_fill_1 FILLER_44_841 ();
 sg13g2_fill_1 FILLER_44_876 ();
 sg13g2_decap_8 FILLER_44_907 ();
 sg13g2_decap_8 FILLER_44_914 ();
 sg13g2_fill_2 FILLER_44_921 ();
 sg13g2_fill_2 FILLER_44_927 ();
 sg13g2_fill_2 FILLER_44_946 ();
 sg13g2_decap_4 FILLER_44_987 ();
 sg13g2_fill_2 FILLER_44_1017 ();
 sg13g2_fill_1 FILLER_44_1044 ();
 sg13g2_fill_2 FILLER_44_1054 ();
 sg13g2_fill_1 FILLER_44_1060 ();
 sg13g2_fill_1 FILLER_44_1069 ();
 sg13g2_fill_1 FILLER_44_1085 ();
 sg13g2_decap_4 FILLER_44_1121 ();
 sg13g2_fill_1 FILLER_44_1169 ();
 sg13g2_fill_2 FILLER_44_1174 ();
 sg13g2_fill_1 FILLER_44_1176 ();
 sg13g2_fill_1 FILLER_44_1221 ();
 sg13g2_fill_2 FILLER_44_1313 ();
 sg13g2_fill_1 FILLER_44_1315 ();
 sg13g2_decap_4 FILLER_44_1326 ();
 sg13g2_fill_1 FILLER_44_1330 ();
 sg13g2_decap_8 FILLER_44_1335 ();
 sg13g2_decap_8 FILLER_44_1342 ();
 sg13g2_fill_2 FILLER_44_1349 ();
 sg13g2_decap_4 FILLER_44_1355 ();
 sg13g2_fill_2 FILLER_44_1359 ();
 sg13g2_fill_1 FILLER_44_1366 ();
 sg13g2_fill_1 FILLER_44_1381 ();
 sg13g2_fill_1 FILLER_44_1386 ();
 sg13g2_decap_4 FILLER_44_1395 ();
 sg13g2_fill_2 FILLER_44_1399 ();
 sg13g2_decap_4 FILLER_44_1410 ();
 sg13g2_fill_2 FILLER_44_1414 ();
 sg13g2_fill_1 FILLER_44_1420 ();
 sg13g2_decap_8 FILLER_44_1426 ();
 sg13g2_decap_8 FILLER_44_1433 ();
 sg13g2_decap_4 FILLER_44_1440 ();
 sg13g2_fill_2 FILLER_44_1449 ();
 sg13g2_decap_8 FILLER_44_1468 ();
 sg13g2_fill_1 FILLER_44_1475 ();
 sg13g2_decap_8 FILLER_44_1480 ();
 sg13g2_fill_2 FILLER_44_1487 ();
 sg13g2_fill_2 FILLER_44_1497 ();
 sg13g2_fill_1 FILLER_44_1499 ();
 sg13g2_decap_8 FILLER_44_1516 ();
 sg13g2_decap_4 FILLER_44_1523 ();
 sg13g2_fill_1 FILLER_44_1527 ();
 sg13g2_fill_2 FILLER_44_1554 ();
 sg13g2_decap_4 FILLER_44_1572 ();
 sg13g2_fill_1 FILLER_44_1576 ();
 sg13g2_decap_8 FILLER_44_1594 ();
 sg13g2_decap_8 FILLER_44_1601 ();
 sg13g2_fill_2 FILLER_44_1624 ();
 sg13g2_fill_1 FILLER_44_1662 ();
 sg13g2_decap_8 FILLER_44_1668 ();
 sg13g2_fill_2 FILLER_44_1675 ();
 sg13g2_fill_2 FILLER_44_1700 ();
 sg13g2_fill_2 FILLER_44_1707 ();
 sg13g2_fill_1 FILLER_44_1709 ();
 sg13g2_fill_2 FILLER_44_1714 ();
 sg13g2_fill_1 FILLER_44_1716 ();
 sg13g2_fill_1 FILLER_44_1747 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_9 ();
 sg13g2_fill_2 FILLER_45_20 ();
 sg13g2_decap_8 FILLER_45_32 ();
 sg13g2_fill_2 FILLER_45_39 ();
 sg13g2_decap_8 FILLER_45_54 ();
 sg13g2_decap_8 FILLER_45_61 ();
 sg13g2_decap_8 FILLER_45_68 ();
 sg13g2_fill_2 FILLER_45_75 ();
 sg13g2_decap_8 FILLER_45_93 ();
 sg13g2_decap_4 FILLER_45_104 ();
 sg13g2_decap_8 FILLER_45_113 ();
 sg13g2_decap_4 FILLER_45_120 ();
 sg13g2_fill_1 FILLER_45_124 ();
 sg13g2_fill_1 FILLER_45_130 ();
 sg13g2_decap_4 FILLER_45_147 ();
 sg13g2_fill_2 FILLER_45_151 ();
 sg13g2_decap_4 FILLER_45_156 ();
 sg13g2_decap_8 FILLER_45_167 ();
 sg13g2_fill_2 FILLER_45_174 ();
 sg13g2_fill_1 FILLER_45_176 ();
 sg13g2_decap_4 FILLER_45_187 ();
 sg13g2_fill_1 FILLER_45_205 ();
 sg13g2_decap_4 FILLER_45_211 ();
 sg13g2_fill_2 FILLER_45_215 ();
 sg13g2_decap_4 FILLER_45_225 ();
 sg13g2_fill_1 FILLER_45_229 ();
 sg13g2_fill_2 FILLER_45_257 ();
 sg13g2_fill_2 FILLER_45_296 ();
 sg13g2_decap_4 FILLER_45_323 ();
 sg13g2_fill_1 FILLER_45_327 ();
 sg13g2_fill_1 FILLER_45_333 ();
 sg13g2_fill_2 FILLER_45_339 ();
 sg13g2_fill_1 FILLER_45_346 ();
 sg13g2_fill_1 FILLER_45_360 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_372 ();
 sg13g2_fill_2 FILLER_45_379 ();
 sg13g2_fill_2 FILLER_45_400 ();
 sg13g2_decap_8 FILLER_45_416 ();
 sg13g2_fill_1 FILLER_45_423 ();
 sg13g2_fill_2 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_45_435 ();
 sg13g2_fill_2 FILLER_45_442 ();
 sg13g2_decap_8 FILLER_45_454 ();
 sg13g2_fill_2 FILLER_45_484 ();
 sg13g2_fill_1 FILLER_45_486 ();
 sg13g2_fill_2 FILLER_45_506 ();
 sg13g2_fill_1 FILLER_45_508 ();
 sg13g2_decap_8 FILLER_45_513 ();
 sg13g2_fill_2 FILLER_45_520 ();
 sg13g2_fill_2 FILLER_45_527 ();
 sg13g2_fill_1 FILLER_45_529 ();
 sg13g2_fill_1 FILLER_45_537 ();
 sg13g2_fill_2 FILLER_45_543 ();
 sg13g2_fill_1 FILLER_45_545 ();
 sg13g2_decap_8 FILLER_45_561 ();
 sg13g2_fill_2 FILLER_45_568 ();
 sg13g2_fill_1 FILLER_45_570 ();
 sg13g2_decap_8 FILLER_45_605 ();
 sg13g2_decap_8 FILLER_45_612 ();
 sg13g2_fill_1 FILLER_45_619 ();
 sg13g2_decap_8 FILLER_45_650 ();
 sg13g2_decap_8 FILLER_45_657 ();
 sg13g2_decap_4 FILLER_45_664 ();
 sg13g2_fill_2 FILLER_45_668 ();
 sg13g2_decap_4 FILLER_45_674 ();
 sg13g2_fill_1 FILLER_45_678 ();
 sg13g2_fill_1 FILLER_45_683 ();
 sg13g2_decap_8 FILLER_45_688 ();
 sg13g2_decap_4 FILLER_45_695 ();
 sg13g2_fill_1 FILLER_45_699 ();
 sg13g2_decap_8 FILLER_45_713 ();
 sg13g2_decap_4 FILLER_45_720 ();
 sg13g2_fill_2 FILLER_45_724 ();
 sg13g2_decap_8 FILLER_45_735 ();
 sg13g2_decap_8 FILLER_45_742 ();
 sg13g2_fill_2 FILLER_45_749 ();
 sg13g2_fill_1 FILLER_45_751 ();
 sg13g2_decap_8 FILLER_45_761 ();
 sg13g2_decap_8 FILLER_45_768 ();
 sg13g2_decap_8 FILLER_45_779 ();
 sg13g2_decap_4 FILLER_45_786 ();
 sg13g2_fill_2 FILLER_45_805 ();
 sg13g2_fill_1 FILLER_45_807 ();
 sg13g2_decap_4 FILLER_45_834 ();
 sg13g2_decap_4 FILLER_45_843 ();
 sg13g2_fill_1 FILLER_45_852 ();
 sg13g2_decap_8 FILLER_45_857 ();
 sg13g2_decap_8 FILLER_45_864 ();
 sg13g2_decap_8 FILLER_45_871 ();
 sg13g2_decap_8 FILLER_45_878 ();
 sg13g2_decap_4 FILLER_45_934 ();
 sg13g2_fill_1 FILLER_45_947 ();
 sg13g2_fill_2 FILLER_45_954 ();
 sg13g2_fill_1 FILLER_45_966 ();
 sg13g2_decap_8 FILLER_45_976 ();
 sg13g2_decap_8 FILLER_45_983 ();
 sg13g2_decap_4 FILLER_45_990 ();
 sg13g2_fill_2 FILLER_45_994 ();
 sg13g2_fill_1 FILLER_45_1021 ();
 sg13g2_fill_2 FILLER_45_1027 ();
 sg13g2_fill_1 FILLER_45_1039 ();
 sg13g2_fill_1 FILLER_45_1045 ();
 sg13g2_fill_2 FILLER_45_1082 ();
 sg13g2_fill_1 FILLER_45_1098 ();
 sg13g2_fill_1 FILLER_45_1115 ();
 sg13g2_decap_4 FILLER_45_1124 ();
 sg13g2_fill_2 FILLER_45_1128 ();
 sg13g2_decap_8 FILLER_45_1145 ();
 sg13g2_fill_1 FILLER_45_1152 ();
 sg13g2_decap_8 FILLER_45_1157 ();
 sg13g2_decap_4 FILLER_45_1164 ();
 sg13g2_decap_4 FILLER_45_1173 ();
 sg13g2_fill_1 FILLER_45_1177 ();
 sg13g2_decap_8 FILLER_45_1183 ();
 sg13g2_fill_2 FILLER_45_1190 ();
 sg13g2_decap_4 FILLER_45_1206 ();
 sg13g2_fill_2 FILLER_45_1210 ();
 sg13g2_decap_8 FILLER_45_1217 ();
 sg13g2_fill_2 FILLER_45_1229 ();
 sg13g2_fill_1 FILLER_45_1235 ();
 sg13g2_decap_8 FILLER_45_1240 ();
 sg13g2_fill_2 FILLER_45_1247 ();
 sg13g2_fill_1 FILLER_45_1249 ();
 sg13g2_decap_4 FILLER_45_1259 ();
 sg13g2_fill_2 FILLER_45_1272 ();
 sg13g2_fill_1 FILLER_45_1274 ();
 sg13g2_fill_2 FILLER_45_1293 ();
 sg13g2_fill_2 FILLER_45_1300 ();
 sg13g2_decap_4 FILLER_45_1307 ();
 sg13g2_fill_1 FILLER_45_1311 ();
 sg13g2_decap_8 FILLER_45_1316 ();
 sg13g2_fill_1 FILLER_45_1323 ();
 sg13g2_decap_8 FILLER_45_1329 ();
 sg13g2_fill_2 FILLER_45_1336 ();
 sg13g2_fill_2 FILLER_45_1396 ();
 sg13g2_fill_1 FILLER_45_1398 ();
 sg13g2_fill_2 FILLER_45_1408 ();
 sg13g2_fill_2 FILLER_45_1416 ();
 sg13g2_fill_1 FILLER_45_1418 ();
 sg13g2_fill_1 FILLER_45_1424 ();
 sg13g2_fill_2 FILLER_45_1451 ();
 sg13g2_fill_1 FILLER_45_1453 ();
 sg13g2_fill_1 FILLER_45_1462 ();
 sg13g2_fill_1 FILLER_45_1471 ();
 sg13g2_fill_1 FILLER_45_1477 ();
 sg13g2_decap_4 FILLER_45_1487 ();
 sg13g2_fill_1 FILLER_45_1496 ();
 sg13g2_fill_2 FILLER_45_1515 ();
 sg13g2_decap_4 FILLER_45_1532 ();
 sg13g2_fill_2 FILLER_45_1536 ();
 sg13g2_fill_2 FILLER_45_1542 ();
 sg13g2_fill_2 FILLER_45_1554 ();
 sg13g2_fill_1 FILLER_45_1569 ();
 sg13g2_decap_4 FILLER_45_1601 ();
 sg13g2_fill_2 FILLER_45_1605 ();
 sg13g2_fill_2 FILLER_45_1611 ();
 sg13g2_fill_1 FILLER_45_1617 ();
 sg13g2_decap_8 FILLER_45_1630 ();
 sg13g2_decap_4 FILLER_45_1637 ();
 sg13g2_fill_2 FILLER_45_1641 ();
 sg13g2_decap_8 FILLER_45_1647 ();
 sg13g2_fill_2 FILLER_45_1654 ();
 sg13g2_decap_8 FILLER_45_1661 ();
 sg13g2_fill_2 FILLER_45_1668 ();
 sg13g2_decap_4 FILLER_45_1678 ();
 sg13g2_fill_1 FILLER_45_1682 ();
 sg13g2_fill_2 FILLER_45_1687 ();
 sg13g2_decap_4 FILLER_45_1704 ();
 sg13g2_fill_2 FILLER_45_1708 ();
 sg13g2_fill_2 FILLER_45_1735 ();
 sg13g2_fill_2 FILLER_45_1750 ();
 sg13g2_fill_1 FILLER_45_1752 ();
 sg13g2_decap_4 FILLER_45_1757 ();
 sg13g2_fill_1 FILLER_45_1761 ();
 sg13g2_decap_8 FILLER_45_1766 ();
 sg13g2_fill_1 FILLER_45_1773 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_19 ();
 sg13g2_fill_2 FILLER_46_39 ();
 sg13g2_fill_1 FILLER_46_41 ();
 sg13g2_decap_8 FILLER_46_58 ();
 sg13g2_fill_2 FILLER_46_65 ();
 sg13g2_decap_4 FILLER_46_75 ();
 sg13g2_fill_2 FILLER_46_79 ();
 sg13g2_fill_2 FILLER_46_89 ();
 sg13g2_fill_2 FILLER_46_96 ();
 sg13g2_decap_8 FILLER_46_113 ();
 sg13g2_fill_2 FILLER_46_120 ();
 sg13g2_fill_1 FILLER_46_122 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_fill_1 FILLER_46_137 ();
 sg13g2_fill_1 FILLER_46_163 ();
 sg13g2_fill_1 FILLER_46_177 ();
 sg13g2_decap_4 FILLER_46_188 ();
 sg13g2_fill_2 FILLER_46_192 ();
 sg13g2_fill_2 FILLER_46_226 ();
 sg13g2_decap_8 FILLER_46_240 ();
 sg13g2_decap_8 FILLER_46_247 ();
 sg13g2_decap_4 FILLER_46_254 ();
 sg13g2_fill_1 FILLER_46_258 ();
 sg13g2_fill_2 FILLER_46_310 ();
 sg13g2_decap_8 FILLER_46_317 ();
 sg13g2_fill_2 FILLER_46_324 ();
 sg13g2_decap_4 FILLER_46_330 ();
 sg13g2_fill_1 FILLER_46_334 ();
 sg13g2_decap_4 FILLER_46_347 ();
 sg13g2_fill_1 FILLER_46_362 ();
 sg13g2_fill_1 FILLER_46_367 ();
 sg13g2_fill_2 FILLER_46_381 ();
 sg13g2_fill_2 FILLER_46_402 ();
 sg13g2_fill_2 FILLER_46_409 ();
 sg13g2_decap_8 FILLER_46_415 ();
 sg13g2_decap_8 FILLER_46_422 ();
 sg13g2_fill_2 FILLER_46_429 ();
 sg13g2_fill_1 FILLER_46_444 ();
 sg13g2_decap_8 FILLER_46_450 ();
 sg13g2_fill_2 FILLER_46_457 ();
 sg13g2_fill_1 FILLER_46_459 ();
 sg13g2_decap_4 FILLER_46_465 ();
 sg13g2_fill_1 FILLER_46_469 ();
 sg13g2_decap_4 FILLER_46_475 ();
 sg13g2_fill_2 FILLER_46_479 ();
 sg13g2_fill_1 FILLER_46_487 ();
 sg13g2_decap_8 FILLER_46_506 ();
 sg13g2_fill_1 FILLER_46_513 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_fill_1 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_559 ();
 sg13g2_decap_8 FILLER_46_580 ();
 sg13g2_decap_4 FILLER_46_587 ();
 sg13g2_decap_8 FILLER_46_596 ();
 sg13g2_decap_4 FILLER_46_612 ();
 sg13g2_fill_2 FILLER_46_622 ();
 sg13g2_decap_8 FILLER_46_628 ();
 sg13g2_fill_1 FILLER_46_635 ();
 sg13g2_decap_4 FILLER_46_647 ();
 sg13g2_fill_2 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_661 ();
 sg13g2_fill_2 FILLER_46_668 ();
 sg13g2_fill_1 FILLER_46_670 ();
 sg13g2_fill_2 FILLER_46_707 ();
 sg13g2_fill_1 FILLER_46_709 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_4 FILLER_46_721 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_fill_2 FILLER_46_749 ();
 sg13g2_fill_2 FILLER_46_765 ();
 sg13g2_fill_1 FILLER_46_767 ();
 sg13g2_decap_8 FILLER_46_804 ();
 sg13g2_decap_4 FILLER_46_811 ();
 sg13g2_fill_1 FILLER_46_815 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_8 FILLER_46_836 ();
 sg13g2_fill_1 FILLER_46_843 ();
 sg13g2_fill_2 FILLER_46_848 ();
 sg13g2_fill_1 FILLER_46_850 ();
 sg13g2_decap_4 FILLER_46_862 ();
 sg13g2_fill_2 FILLER_46_870 ();
 sg13g2_fill_1 FILLER_46_872 ();
 sg13g2_decap_8 FILLER_46_888 ();
 sg13g2_decap_8 FILLER_46_895 ();
 sg13g2_fill_2 FILLER_46_902 ();
 sg13g2_fill_1 FILLER_46_914 ();
 sg13g2_fill_2 FILLER_46_919 ();
 sg13g2_fill_1 FILLER_46_921 ();
 sg13g2_fill_1 FILLER_46_935 ();
 sg13g2_fill_2 FILLER_46_941 ();
 sg13g2_fill_1 FILLER_46_958 ();
 sg13g2_fill_1 FILLER_46_969 ();
 sg13g2_decap_4 FILLER_46_984 ();
 sg13g2_fill_1 FILLER_46_993 ();
 sg13g2_fill_2 FILLER_46_998 ();
 sg13g2_decap_4 FILLER_46_1004 ();
 sg13g2_fill_2 FILLER_46_1008 ();
 sg13g2_fill_2 FILLER_46_1026 ();
 sg13g2_fill_2 FILLER_46_1032 ();
 sg13g2_fill_1 FILLER_46_1058 ();
 sg13g2_fill_2 FILLER_46_1075 ();
 sg13g2_fill_1 FILLER_46_1077 ();
 sg13g2_fill_2 FILLER_46_1083 ();
 sg13g2_fill_2 FILLER_46_1110 ();
 sg13g2_decap_4 FILLER_46_1129 ();
 sg13g2_fill_2 FILLER_46_1138 ();
 sg13g2_fill_1 FILLER_46_1140 ();
 sg13g2_fill_2 FILLER_46_1176 ();
 sg13g2_decap_4 FILLER_46_1212 ();
 sg13g2_fill_1 FILLER_46_1216 ();
 sg13g2_fill_2 FILLER_46_1222 ();
 sg13g2_fill_1 FILLER_46_1224 ();
 sg13g2_decap_8 FILLER_46_1229 ();
 sg13g2_fill_1 FILLER_46_1240 ();
 sg13g2_decap_8 FILLER_46_1255 ();
 sg13g2_decap_8 FILLER_46_1297 ();
 sg13g2_fill_2 FILLER_46_1304 ();
 sg13g2_fill_1 FILLER_46_1320 ();
 sg13g2_decap_8 FILLER_46_1325 ();
 sg13g2_decap_4 FILLER_46_1332 ();
 sg13g2_fill_2 FILLER_46_1336 ();
 sg13g2_fill_1 FILLER_46_1352 ();
 sg13g2_decap_8 FILLER_46_1357 ();
 sg13g2_decap_8 FILLER_46_1364 ();
 sg13g2_decap_4 FILLER_46_1371 ();
 sg13g2_fill_2 FILLER_46_1410 ();
 sg13g2_fill_1 FILLER_46_1412 ();
 sg13g2_fill_1 FILLER_46_1431 ();
 sg13g2_decap_8 FILLER_46_1436 ();
 sg13g2_fill_2 FILLER_46_1443 ();
 sg13g2_fill_1 FILLER_46_1445 ();
 sg13g2_decap_4 FILLER_46_1491 ();
 sg13g2_fill_2 FILLER_46_1495 ();
 sg13g2_decap_8 FILLER_46_1515 ();
 sg13g2_fill_1 FILLER_46_1522 ();
 sg13g2_fill_1 FILLER_46_1552 ();
 sg13g2_decap_8 FILLER_46_1589 ();
 sg13g2_decap_8 FILLER_46_1596 ();
 sg13g2_fill_2 FILLER_46_1603 ();
 sg13g2_decap_8 FILLER_46_1625 ();
 sg13g2_fill_1 FILLER_46_1632 ();
 sg13g2_fill_2 FILLER_46_1650 ();
 sg13g2_fill_1 FILLER_46_1657 ();
 sg13g2_decap_4 FILLER_46_1663 ();
 sg13g2_decap_8 FILLER_46_1679 ();
 sg13g2_decap_8 FILLER_46_1686 ();
 sg13g2_fill_2 FILLER_46_1693 ();
 sg13g2_fill_1 FILLER_46_1695 ();
 sg13g2_fill_2 FILLER_46_1709 ();
 sg13g2_fill_2 FILLER_46_1772 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_fill_2 FILLER_47_21 ();
 sg13g2_fill_2 FILLER_47_36 ();
 sg13g2_fill_1 FILLER_47_38 ();
 sg13g2_fill_2 FILLER_47_60 ();
 sg13g2_decap_4 FILLER_47_89 ();
 sg13g2_fill_2 FILLER_47_93 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_fill_2 FILLER_47_112 ();
 sg13g2_fill_1 FILLER_47_114 ();
 sg13g2_decap_4 FILLER_47_133 ();
 sg13g2_decap_4 FILLER_47_141 ();
 sg13g2_fill_2 FILLER_47_151 ();
 sg13g2_fill_1 FILLER_47_169 ();
 sg13g2_decap_4 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_200 ();
 sg13g2_decap_4 FILLER_47_205 ();
 sg13g2_decap_4 FILLER_47_214 ();
 sg13g2_fill_1 FILLER_47_218 ();
 sg13g2_fill_2 FILLER_47_223 ();
 sg13g2_decap_4 FILLER_47_241 ();
 sg13g2_fill_2 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_262 ();
 sg13g2_decap_4 FILLER_47_274 ();
 sg13g2_fill_2 FILLER_47_287 ();
 sg13g2_fill_1 FILLER_47_294 ();
 sg13g2_decap_4 FILLER_47_300 ();
 sg13g2_fill_2 FILLER_47_304 ();
 sg13g2_decap_8 FILLER_47_314 ();
 sg13g2_fill_2 FILLER_47_321 ();
 sg13g2_fill_2 FILLER_47_332 ();
 sg13g2_fill_2 FILLER_47_339 ();
 sg13g2_fill_2 FILLER_47_347 ();
 sg13g2_fill_1 FILLER_47_349 ();
 sg13g2_decap_8 FILLER_47_355 ();
 sg13g2_fill_2 FILLER_47_362 ();
 sg13g2_fill_1 FILLER_47_364 ();
 sg13g2_decap_4 FILLER_47_376 ();
 sg13g2_fill_1 FILLER_47_380 ();
 sg13g2_fill_2 FILLER_47_386 ();
 sg13g2_decap_4 FILLER_47_393 ();
 sg13g2_fill_2 FILLER_47_403 ();
 sg13g2_fill_1 FILLER_47_405 ();
 sg13g2_fill_1 FILLER_47_411 ();
 sg13g2_fill_2 FILLER_47_429 ();
 sg13g2_fill_1 FILLER_47_431 ();
 sg13g2_fill_1 FILLER_47_436 ();
 sg13g2_fill_1 FILLER_47_442 ();
 sg13g2_fill_1 FILLER_47_447 ();
 sg13g2_fill_2 FILLER_47_458 ();
 sg13g2_fill_2 FILLER_47_479 ();
 sg13g2_fill_1 FILLER_47_481 ();
 sg13g2_decap_4 FILLER_47_505 ();
 sg13g2_fill_1 FILLER_47_509 ();
 sg13g2_fill_2 FILLER_47_521 ();
 sg13g2_fill_1 FILLER_47_523 ();
 sg13g2_decap_8 FILLER_47_529 ();
 sg13g2_decap_8 FILLER_47_536 ();
 sg13g2_decap_8 FILLER_47_543 ();
 sg13g2_fill_2 FILLER_47_550 ();
 sg13g2_fill_1 FILLER_47_566 ();
 sg13g2_fill_1 FILLER_47_574 ();
 sg13g2_fill_1 FILLER_47_586 ();
 sg13g2_fill_2 FILLER_47_592 ();
 sg13g2_fill_1 FILLER_47_594 ();
 sg13g2_fill_1 FILLER_47_607 ();
 sg13g2_fill_2 FILLER_47_636 ();
 sg13g2_fill_2 FILLER_47_648 ();
 sg13g2_decap_8 FILLER_47_662 ();
 sg13g2_decap_8 FILLER_47_669 ();
 sg13g2_fill_2 FILLER_47_685 ();
 sg13g2_decap_4 FILLER_47_696 ();
 sg13g2_fill_2 FILLER_47_700 ();
 sg13g2_fill_2 FILLER_47_741 ();
 sg13g2_fill_1 FILLER_47_743 ();
 sg13g2_decap_4 FILLER_47_774 ();
 sg13g2_decap_8 FILLER_47_804 ();
 sg13g2_decap_8 FILLER_47_811 ();
 sg13g2_fill_1 FILLER_47_862 ();
 sg13g2_decap_8 FILLER_47_881 ();
 sg13g2_fill_1 FILLER_47_893 ();
 sg13g2_decap_8 FILLER_47_898 ();
 sg13g2_decap_8 FILLER_47_905 ();
 sg13g2_decap_4 FILLER_47_912 ();
 sg13g2_fill_1 FILLER_47_916 ();
 sg13g2_decap_8 FILLER_47_921 ();
 sg13g2_fill_2 FILLER_47_928 ();
 sg13g2_fill_2 FILLER_47_934 ();
 sg13g2_fill_1 FILLER_47_936 ();
 sg13g2_fill_1 FILLER_47_982 ();
 sg13g2_decap_4 FILLER_47_987 ();
 sg13g2_fill_2 FILLER_47_991 ();
 sg13g2_fill_1 FILLER_47_998 ();
 sg13g2_fill_1 FILLER_47_1004 ();
 sg13g2_fill_1 FILLER_47_1047 ();
 sg13g2_fill_1 FILLER_47_1058 ();
 sg13g2_decap_4 FILLER_47_1067 ();
 sg13g2_fill_1 FILLER_47_1102 ();
 sg13g2_fill_2 FILLER_47_1112 ();
 sg13g2_fill_2 FILLER_47_1128 ();
 sg13g2_decap_8 FILLER_47_1135 ();
 sg13g2_fill_2 FILLER_47_1142 ();
 sg13g2_fill_1 FILLER_47_1149 ();
 sg13g2_decap_8 FILLER_47_1155 ();
 sg13g2_decap_8 FILLER_47_1162 ();
 sg13g2_decap_8 FILLER_47_1169 ();
 sg13g2_decap_4 FILLER_47_1176 ();
 sg13g2_fill_1 FILLER_47_1180 ();
 sg13g2_decap_8 FILLER_47_1189 ();
 sg13g2_decap_4 FILLER_47_1196 ();
 sg13g2_fill_1 FILLER_47_1200 ();
 sg13g2_decap_8 FILLER_47_1206 ();
 sg13g2_decap_8 FILLER_47_1213 ();
 sg13g2_decap_4 FILLER_47_1220 ();
 sg13g2_decap_8 FILLER_47_1260 ();
 sg13g2_fill_2 FILLER_47_1267 ();
 sg13g2_fill_1 FILLER_47_1269 ();
 sg13g2_fill_2 FILLER_47_1275 ();
 sg13g2_fill_1 FILLER_47_1277 ();
 sg13g2_decap_4 FILLER_47_1282 ();
 sg13g2_fill_1 FILLER_47_1286 ();
 sg13g2_fill_1 FILLER_47_1308 ();
 sg13g2_decap_8 FILLER_47_1340 ();
 sg13g2_fill_1 FILLER_47_1347 ();
 sg13g2_decap_4 FILLER_47_1352 ();
 sg13g2_fill_1 FILLER_47_1356 ();
 sg13g2_fill_1 FILLER_47_1360 ();
 sg13g2_fill_2 FILLER_47_1372 ();
 sg13g2_fill_1 FILLER_47_1378 ();
 sg13g2_fill_2 FILLER_47_1383 ();
 sg13g2_fill_2 FILLER_47_1403 ();
 sg13g2_fill_1 FILLER_47_1422 ();
 sg13g2_fill_1 FILLER_47_1431 ();
 sg13g2_decap_8 FILLER_47_1463 ();
 sg13g2_fill_2 FILLER_47_1470 ();
 sg13g2_fill_1 FILLER_47_1472 ();
 sg13g2_fill_2 FILLER_47_1477 ();
 sg13g2_decap_4 FILLER_47_1529 ();
 sg13g2_fill_2 FILLER_47_1533 ();
 sg13g2_decap_8 FILLER_47_1539 ();
 sg13g2_fill_2 FILLER_47_1546 ();
 sg13g2_fill_1 FILLER_47_1548 ();
 sg13g2_fill_2 FILLER_47_1594 ();
 sg13g2_decap_8 FILLER_47_1600 ();
 sg13g2_fill_1 FILLER_47_1607 ();
 sg13g2_decap_4 FILLER_47_1626 ();
 sg13g2_fill_1 FILLER_47_1630 ();
 sg13g2_decap_4 FILLER_47_1661 ();
 sg13g2_fill_2 FILLER_47_1665 ();
 sg13g2_decap_8 FILLER_47_1672 ();
 sg13g2_decap_8 FILLER_47_1679 ();
 sg13g2_decap_8 FILLER_47_1686 ();
 sg13g2_fill_2 FILLER_47_1693 ();
 sg13g2_fill_1 FILLER_47_1695 ();
 sg13g2_fill_1 FILLER_47_1706 ();
 sg13g2_fill_2 FILLER_47_1720 ();
 sg13g2_decap_8 FILLER_47_1740 ();
 sg13g2_decap_4 FILLER_47_1747 ();
 sg13g2_decap_8 FILLER_47_1755 ();
 sg13g2_decap_8 FILLER_47_1762 ();
 sg13g2_decap_4 FILLER_47_1769 ();
 sg13g2_fill_1 FILLER_47_1773 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_4 FILLER_48_14 ();
 sg13g2_fill_1 FILLER_48_18 ();
 sg13g2_fill_2 FILLER_48_31 ();
 sg13g2_fill_1 FILLER_48_37 ();
 sg13g2_fill_2 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_50 ();
 sg13g2_decap_4 FILLER_48_57 ();
 sg13g2_fill_1 FILLER_48_61 ();
 sg13g2_decap_8 FILLER_48_67 ();
 sg13g2_decap_8 FILLER_48_74 ();
 sg13g2_fill_1 FILLER_48_89 ();
 sg13g2_decap_4 FILLER_48_117 ();
 sg13g2_fill_2 FILLER_48_121 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_fill_2 FILLER_48_140 ();
 sg13g2_fill_1 FILLER_48_142 ();
 sg13g2_fill_1 FILLER_48_156 ();
 sg13g2_fill_2 FILLER_48_162 ();
 sg13g2_fill_1 FILLER_48_164 ();
 sg13g2_decap_8 FILLER_48_206 ();
 sg13g2_fill_2 FILLER_48_217 ();
 sg13g2_fill_1 FILLER_48_224 ();
 sg13g2_fill_2 FILLER_48_237 ();
 sg13g2_fill_1 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_fill_1 FILLER_48_259 ();
 sg13g2_fill_1 FILLER_48_265 ();
 sg13g2_fill_2 FILLER_48_273 ();
 sg13g2_fill_1 FILLER_48_275 ();
 sg13g2_fill_1 FILLER_48_286 ();
 sg13g2_fill_2 FILLER_48_294 ();
 sg13g2_fill_1 FILLER_48_296 ();
 sg13g2_decap_4 FILLER_48_302 ();
 sg13g2_fill_2 FILLER_48_306 ();
 sg13g2_fill_2 FILLER_48_318 ();
 sg13g2_decap_8 FILLER_48_327 ();
 sg13g2_decap_4 FILLER_48_334 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_354 ();
 sg13g2_decap_8 FILLER_48_361 ();
 sg13g2_fill_1 FILLER_48_368 ();
 sg13g2_decap_4 FILLER_48_373 ();
 sg13g2_fill_1 FILLER_48_382 ();
 sg13g2_fill_2 FILLER_48_393 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_415 ();
 sg13g2_fill_1 FILLER_48_417 ();
 sg13g2_fill_2 FILLER_48_443 ();
 sg13g2_decap_4 FILLER_48_449 ();
 sg13g2_fill_2 FILLER_48_458 ();
 sg13g2_decap_4 FILLER_48_477 ();
 sg13g2_fill_1 FILLER_48_481 ();
 sg13g2_decap_8 FILLER_48_486 ();
 sg13g2_fill_2 FILLER_48_493 ();
 sg13g2_decap_4 FILLER_48_500 ();
 sg13g2_decap_4 FILLER_48_509 ();
 sg13g2_fill_2 FILLER_48_513 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_fill_1 FILLER_48_532 ();
 sg13g2_fill_2 FILLER_48_540 ();
 sg13g2_fill_2 FILLER_48_561 ();
 sg13g2_fill_2 FILLER_48_568 ();
 sg13g2_fill_2 FILLER_48_586 ();
 sg13g2_fill_1 FILLER_48_596 ();
 sg13g2_fill_1 FILLER_48_607 ();
 sg13g2_fill_2 FILLER_48_622 ();
 sg13g2_fill_1 FILLER_48_643 ();
 sg13g2_decap_8 FILLER_48_648 ();
 sg13g2_decap_4 FILLER_48_655 ();
 sg13g2_fill_2 FILLER_48_674 ();
 sg13g2_fill_1 FILLER_48_676 ();
 sg13g2_fill_1 FILLER_48_681 ();
 sg13g2_fill_1 FILLER_48_689 ();
 sg13g2_decap_8 FILLER_48_702 ();
 sg13g2_fill_1 FILLER_48_721 ();
 sg13g2_decap_4 FILLER_48_745 ();
 sg13g2_decap_4 FILLER_48_753 ();
 sg13g2_fill_1 FILLER_48_757 ();
 sg13g2_fill_2 FILLER_48_771 ();
 sg13g2_decap_8 FILLER_48_778 ();
 sg13g2_fill_1 FILLER_48_785 ();
 sg13g2_decap_4 FILLER_48_790 ();
 sg13g2_fill_1 FILLER_48_794 ();
 sg13g2_decap_4 FILLER_48_825 ();
 sg13g2_fill_2 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_4 FILLER_48_875 ();
 sg13g2_fill_1 FILLER_48_883 ();
 sg13g2_fill_2 FILLER_48_889 ();
 sg13g2_decap_4 FILLER_48_895 ();
 sg13g2_fill_1 FILLER_48_899 ();
 sg13g2_fill_2 FILLER_48_905 ();
 sg13g2_decap_4 FILLER_48_912 ();
 sg13g2_fill_2 FILLER_48_916 ();
 sg13g2_decap_8 FILLER_48_923 ();
 sg13g2_fill_2 FILLER_48_930 ();
 sg13g2_fill_2 FILLER_48_941 ();
 sg13g2_fill_1 FILLER_48_943 ();
 sg13g2_fill_2 FILLER_48_966 ();
 sg13g2_decap_8 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_987 ();
 sg13g2_fill_2 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1009 ();
 sg13g2_decap_4 FILLER_48_1020 ();
 sg13g2_fill_2 FILLER_48_1024 ();
 sg13g2_decap_8 FILLER_48_1052 ();
 sg13g2_fill_2 FILLER_48_1059 ();
 sg13g2_fill_1 FILLER_48_1061 ();
 sg13g2_decap_8 FILLER_48_1066 ();
 sg13g2_decap_8 FILLER_48_1073 ();
 sg13g2_fill_2 FILLER_48_1080 ();
 sg13g2_fill_2 FILLER_48_1105 ();
 sg13g2_fill_2 FILLER_48_1140 ();
 sg13g2_fill_1 FILLER_48_1142 ();
 sg13g2_decap_8 FILLER_48_1148 ();
 sg13g2_decap_4 FILLER_48_1155 ();
 sg13g2_decap_4 FILLER_48_1196 ();
 sg13g2_fill_1 FILLER_48_1200 ();
 sg13g2_fill_1 FILLER_48_1210 ();
 sg13g2_decap_4 FILLER_48_1221 ();
 sg13g2_fill_1 FILLER_48_1225 ();
 sg13g2_fill_1 FILLER_48_1230 ();
 sg13g2_fill_1 FILLER_48_1235 ();
 sg13g2_fill_1 FILLER_48_1240 ();
 sg13g2_fill_1 FILLER_48_1246 ();
 sg13g2_fill_1 FILLER_48_1252 ();
 sg13g2_fill_2 FILLER_48_1257 ();
 sg13g2_fill_2 FILLER_48_1281 ();
 sg13g2_fill_1 FILLER_48_1283 ();
 sg13g2_fill_2 FILLER_48_1292 ();
 sg13g2_fill_2 FILLER_48_1299 ();
 sg13g2_fill_1 FILLER_48_1306 ();
 sg13g2_decap_8 FILLER_48_1338 ();
 sg13g2_fill_2 FILLER_48_1345 ();
 sg13g2_fill_1 FILLER_48_1356 ();
 sg13g2_decap_4 FILLER_48_1402 ();
 sg13g2_fill_1 FILLER_48_1406 ();
 sg13g2_fill_2 FILLER_48_1411 ();
 sg13g2_decap_8 FILLER_48_1434 ();
 sg13g2_fill_1 FILLER_48_1441 ();
 sg13g2_decap_8 FILLER_48_1446 ();
 sg13g2_decap_4 FILLER_48_1453 ();
 sg13g2_fill_1 FILLER_48_1457 ();
 sg13g2_decap_8 FILLER_48_1462 ();
 sg13g2_fill_1 FILLER_48_1469 ();
 sg13g2_fill_1 FILLER_48_1490 ();
 sg13g2_fill_2 FILLER_48_1513 ();
 sg13g2_fill_1 FILLER_48_1515 ();
 sg13g2_decap_8 FILLER_48_1525 ();
 sg13g2_decap_8 FILLER_48_1532 ();
 sg13g2_fill_2 FILLER_48_1539 ();
 sg13g2_decap_4 FILLER_48_1551 ();
 sg13g2_fill_1 FILLER_48_1555 ();
 sg13g2_fill_2 FILLER_48_1562 ();
 sg13g2_decap_8 FILLER_48_1574 ();
 sg13g2_decap_4 FILLER_48_1581 ();
 sg13g2_decap_8 FILLER_48_1615 ();
 sg13g2_decap_8 FILLER_48_1622 ();
 sg13g2_fill_1 FILLER_48_1629 ();
 sg13g2_decap_8 FILLER_48_1640 ();
 sg13g2_fill_2 FILLER_48_1647 ();
 sg13g2_fill_1 FILLER_48_1649 ();
 sg13g2_decap_8 FILLER_48_1668 ();
 sg13g2_decap_8 FILLER_48_1675 ();
 sg13g2_decap_8 FILLER_48_1682 ();
 sg13g2_decap_4 FILLER_48_1689 ();
 sg13g2_fill_1 FILLER_48_1693 ();
 sg13g2_fill_2 FILLER_48_1704 ();
 sg13g2_decap_8 FILLER_48_1711 ();
 sg13g2_decap_4 FILLER_48_1718 ();
 sg13g2_fill_2 FILLER_48_1722 ();
 sg13g2_decap_4 FILLER_48_1733 ();
 sg13g2_fill_1 FILLER_48_1737 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_19 ();
 sg13g2_fill_1 FILLER_49_26 ();
 sg13g2_fill_1 FILLER_49_32 ();
 sg13g2_decap_4 FILLER_49_37 ();
 sg13g2_fill_2 FILLER_49_45 ();
 sg13g2_fill_1 FILLER_49_47 ();
 sg13g2_decap_4 FILLER_49_53 ();
 sg13g2_fill_2 FILLER_49_57 ();
 sg13g2_fill_2 FILLER_49_66 ();
 sg13g2_decap_4 FILLER_49_72 ();
 sg13g2_fill_2 FILLER_49_76 ();
 sg13g2_decap_8 FILLER_49_82 ();
 sg13g2_decap_4 FILLER_49_89 ();
 sg13g2_fill_1 FILLER_49_93 ();
 sg13g2_decap_4 FILLER_49_103 ();
 sg13g2_fill_1 FILLER_49_107 ();
 sg13g2_decap_4 FILLER_49_113 ();
 sg13g2_decap_8 FILLER_49_121 ();
 sg13g2_fill_2 FILLER_49_128 ();
 sg13g2_fill_2 FILLER_49_138 ();
 sg13g2_decap_8 FILLER_49_152 ();
 sg13g2_decap_8 FILLER_49_159 ();
 sg13g2_fill_2 FILLER_49_166 ();
 sg13g2_fill_1 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_184 ();
 sg13g2_fill_2 FILLER_49_191 ();
 sg13g2_fill_2 FILLER_49_205 ();
 sg13g2_decap_8 FILLER_49_211 ();
 sg13g2_decap_8 FILLER_49_218 ();
 sg13g2_decap_4 FILLER_49_225 ();
 sg13g2_decap_4 FILLER_49_233 ();
 sg13g2_fill_1 FILLER_49_237 ();
 sg13g2_fill_1 FILLER_49_255 ();
 sg13g2_fill_2 FILLER_49_260 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_fill_1 FILLER_49_294 ();
 sg13g2_fill_1 FILLER_49_310 ();
 sg13g2_decap_8 FILLER_49_317 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_fill_1 FILLER_49_337 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_fill_1 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_360 ();
 sg13g2_decap_8 FILLER_49_367 ();
 sg13g2_decap_8 FILLER_49_374 ();
 sg13g2_fill_1 FILLER_49_381 ();
 sg13g2_fill_2 FILLER_49_401 ();
 sg13g2_fill_2 FILLER_49_408 ();
 sg13g2_fill_1 FILLER_49_410 ();
 sg13g2_decap_8 FILLER_49_415 ();
 sg13g2_decap_8 FILLER_49_422 ();
 sg13g2_decap_4 FILLER_49_429 ();
 sg13g2_fill_2 FILLER_49_438 ();
 sg13g2_fill_2 FILLER_49_445 ();
 sg13g2_fill_1 FILLER_49_447 ();
 sg13g2_decap_4 FILLER_49_466 ();
 sg13g2_fill_1 FILLER_49_480 ();
 sg13g2_decap_4 FILLER_49_491 ();
 sg13g2_fill_1 FILLER_49_495 ();
 sg13g2_decap_4 FILLER_49_500 ();
 sg13g2_decap_4 FILLER_49_527 ();
 sg13g2_decap_4 FILLER_49_542 ();
 sg13g2_decap_4 FILLER_49_550 ();
 sg13g2_fill_1 FILLER_49_554 ();
 sg13g2_decap_8 FILLER_49_606 ();
 sg13g2_decap_8 FILLER_49_645 ();
 sg13g2_fill_2 FILLER_49_666 ();
 sg13g2_fill_2 FILLER_49_674 ();
 sg13g2_fill_2 FILLER_49_681 ();
 sg13g2_decap_8 FILLER_49_688 ();
 sg13g2_fill_2 FILLER_49_695 ();
 sg13g2_fill_1 FILLER_49_702 ();
 sg13g2_fill_1 FILLER_49_710 ();
 sg13g2_fill_1 FILLER_49_720 ();
 sg13g2_decap_8 FILLER_49_739 ();
 sg13g2_fill_1 FILLER_49_746 ();
 sg13g2_decap_8 FILLER_49_760 ();
 sg13g2_fill_1 FILLER_49_767 ();
 sg13g2_fill_2 FILLER_49_773 ();
 sg13g2_fill_1 FILLER_49_775 ();
 sg13g2_decap_4 FILLER_49_781 ();
 sg13g2_fill_2 FILLER_49_803 ();
 sg13g2_decap_4 FILLER_49_809 ();
 sg13g2_fill_2 FILLER_49_813 ();
 sg13g2_decap_4 FILLER_49_820 ();
 sg13g2_fill_1 FILLER_49_824 ();
 sg13g2_fill_1 FILLER_49_830 ();
 sg13g2_fill_2 FILLER_49_836 ();
 sg13g2_decap_8 FILLER_49_846 ();
 sg13g2_fill_2 FILLER_49_853 ();
 sg13g2_fill_1 FILLER_49_855 ();
 sg13g2_fill_1 FILLER_49_864 ();
 sg13g2_fill_1 FILLER_49_869 ();
 sg13g2_fill_1 FILLER_49_901 ();
 sg13g2_fill_2 FILLER_49_932 ();
 sg13g2_fill_1 FILLER_49_934 ();
 sg13g2_fill_2 FILLER_49_939 ();
 sg13g2_fill_1 FILLER_49_945 ();
 sg13g2_fill_1 FILLER_49_1045 ();
 sg13g2_fill_1 FILLER_49_1050 ();
 sg13g2_fill_1 FILLER_49_1056 ();
 sg13g2_decap_4 FILLER_49_1080 ();
 sg13g2_fill_2 FILLER_49_1088 ();
 sg13g2_fill_1 FILLER_49_1095 ();
 sg13g2_decap_8 FILLER_49_1101 ();
 sg13g2_fill_2 FILLER_49_1108 ();
 sg13g2_fill_2 FILLER_49_1116 ();
 sg13g2_fill_1 FILLER_49_1118 ();
 sg13g2_decap_8 FILLER_49_1124 ();
 sg13g2_decap_4 FILLER_49_1131 ();
 sg13g2_fill_1 FILLER_49_1135 ();
 sg13g2_decap_8 FILLER_49_1164 ();
 sg13g2_decap_4 FILLER_49_1171 ();
 sg13g2_fill_1 FILLER_49_1175 ();
 sg13g2_decap_8 FILLER_49_1180 ();
 sg13g2_fill_1 FILLER_49_1187 ();
 sg13g2_fill_2 FILLER_49_1193 ();
 sg13g2_fill_1 FILLER_49_1195 ();
 sg13g2_decap_4 FILLER_49_1205 ();
 sg13g2_decap_8 FILLER_49_1269 ();
 sg13g2_decap_8 FILLER_49_1276 ();
 sg13g2_fill_1 FILLER_49_1296 ();
 sg13g2_fill_1 FILLER_49_1302 ();
 sg13g2_fill_1 FILLER_49_1313 ();
 sg13g2_fill_1 FILLER_49_1318 ();
 sg13g2_fill_2 FILLER_49_1322 ();
 sg13g2_decap_8 FILLER_49_1350 ();
 sg13g2_decap_8 FILLER_49_1357 ();
 sg13g2_fill_2 FILLER_49_1364 ();
 sg13g2_fill_1 FILLER_49_1374 ();
 sg13g2_fill_1 FILLER_49_1390 ();
 sg13g2_fill_2 FILLER_49_1407 ();
 sg13g2_decap_4 FILLER_49_1413 ();
 sg13g2_decap_4 FILLER_49_1421 ();
 sg13g2_fill_1 FILLER_49_1425 ();
 sg13g2_fill_1 FILLER_49_1431 ();
 sg13g2_fill_2 FILLER_49_1458 ();
 sg13g2_fill_1 FILLER_49_1460 ();
 sg13g2_decap_8 FILLER_49_1469 ();
 sg13g2_fill_2 FILLER_49_1476 ();
 sg13g2_fill_2 FILLER_49_1491 ();
 sg13g2_fill_1 FILLER_49_1493 ();
 sg13g2_decap_4 FILLER_49_1543 ();
 sg13g2_fill_2 FILLER_49_1583 ();
 sg13g2_fill_1 FILLER_49_1585 ();
 sg13g2_decap_8 FILLER_49_1590 ();
 sg13g2_decap_8 FILLER_49_1597 ();
 sg13g2_decap_8 FILLER_49_1604 ();
 sg13g2_decap_4 FILLER_49_1611 ();
 sg13g2_fill_2 FILLER_49_1627 ();
 sg13g2_decap_8 FILLER_49_1648 ();
 sg13g2_decap_4 FILLER_49_1689 ();
 sg13g2_fill_1 FILLER_49_1714 ();
 sg13g2_decap_4 FILLER_49_1720 ();
 sg13g2_fill_1 FILLER_49_1724 ();
 sg13g2_decap_4 FILLER_49_1737 ();
 sg13g2_decap_4 FILLER_49_1751 ();
 sg13g2_fill_2 FILLER_49_1755 ();
 sg13g2_fill_1 FILLER_49_1761 ();
 sg13g2_decap_8 FILLER_49_1766 ();
 sg13g2_fill_1 FILLER_49_1773 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_31 ();
 sg13g2_fill_1 FILLER_50_46 ();
 sg13g2_decap_4 FILLER_50_51 ();
 sg13g2_decap_4 FILLER_50_81 ();
 sg13g2_fill_2 FILLER_50_85 ();
 sg13g2_decap_8 FILLER_50_97 ();
 sg13g2_fill_1 FILLER_50_124 ();
 sg13g2_fill_1 FILLER_50_135 ();
 sg13g2_fill_1 FILLER_50_141 ();
 sg13g2_fill_1 FILLER_50_146 ();
 sg13g2_fill_1 FILLER_50_151 ();
 sg13g2_decap_8 FILLER_50_159 ();
 sg13g2_fill_2 FILLER_50_166 ();
 sg13g2_fill_1 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_183 ();
 sg13g2_decap_4 FILLER_50_190 ();
 sg13g2_fill_2 FILLER_50_194 ();
 sg13g2_decap_8 FILLER_50_218 ();
 sg13g2_fill_2 FILLER_50_225 ();
 sg13g2_fill_1 FILLER_50_227 ();
 sg13g2_fill_1 FILLER_50_233 ();
 sg13g2_fill_2 FILLER_50_240 ();
 sg13g2_decap_8 FILLER_50_247 ();
 sg13g2_decap_8 FILLER_50_254 ();
 sg13g2_decap_8 FILLER_50_261 ();
 sg13g2_fill_1 FILLER_50_268 ();
 sg13g2_decap_8 FILLER_50_281 ();
 sg13g2_decap_8 FILLER_50_301 ();
 sg13g2_decap_8 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_315 ();
 sg13g2_decap_4 FILLER_50_322 ();
 sg13g2_fill_1 FILLER_50_342 ();
 sg13g2_decap_4 FILLER_50_348 ();
 sg13g2_fill_2 FILLER_50_352 ();
 sg13g2_decap_8 FILLER_50_359 ();
 sg13g2_decap_4 FILLER_50_366 ();
 sg13g2_fill_2 FILLER_50_370 ();
 sg13g2_decap_8 FILLER_50_381 ();
 sg13g2_decap_4 FILLER_50_388 ();
 sg13g2_decap_4 FILLER_50_396 ();
 sg13g2_fill_1 FILLER_50_400 ();
 sg13g2_decap_8 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_50_412 ();
 sg13g2_fill_2 FILLER_50_419 ();
 sg13g2_decap_8 FILLER_50_426 ();
 sg13g2_decap_8 FILLER_50_433 ();
 sg13g2_decap_8 FILLER_50_440 ();
 sg13g2_decap_8 FILLER_50_447 ();
 sg13g2_decap_8 FILLER_50_454 ();
 sg13g2_decap_4 FILLER_50_461 ();
 sg13g2_fill_1 FILLER_50_465 ();
 sg13g2_decap_4 FILLER_50_471 ();
 sg13g2_decap_8 FILLER_50_485 ();
 sg13g2_fill_2 FILLER_50_492 ();
 sg13g2_decap_4 FILLER_50_518 ();
 sg13g2_decap_4 FILLER_50_526 ();
 sg13g2_decap_4 FILLER_50_535 ();
 sg13g2_decap_8 FILLER_50_547 ();
 sg13g2_fill_2 FILLER_50_554 ();
 sg13g2_fill_2 FILLER_50_579 ();
 sg13g2_decap_8 FILLER_50_605 ();
 sg13g2_decap_8 FILLER_50_612 ();
 sg13g2_decap_8 FILLER_50_619 ();
 sg13g2_fill_2 FILLER_50_626 ();
 sg13g2_fill_1 FILLER_50_628 ();
 sg13g2_fill_2 FILLER_50_657 ();
 sg13g2_decap_4 FILLER_50_666 ();
 sg13g2_decap_8 FILLER_50_675 ();
 sg13g2_decap_8 FILLER_50_682 ();
 sg13g2_decap_8 FILLER_50_689 ();
 sg13g2_fill_1 FILLER_50_706 ();
 sg13g2_fill_2 FILLER_50_744 ();
 sg13g2_fill_1 FILLER_50_746 ();
 sg13g2_fill_1 FILLER_50_773 ();
 sg13g2_decap_8 FILLER_50_812 ();
 sg13g2_decap_8 FILLER_50_864 ();
 sg13g2_fill_1 FILLER_50_899 ();
 sg13g2_fill_2 FILLER_50_910 ();
 sg13g2_decap_8 FILLER_50_927 ();
 sg13g2_fill_2 FILLER_50_934 ();
 sg13g2_fill_1 FILLER_50_936 ();
 sg13g2_fill_1 FILLER_50_946 ();
 sg13g2_fill_2 FILLER_50_961 ();
 sg13g2_fill_2 FILLER_50_979 ();
 sg13g2_fill_2 FILLER_50_990 ();
 sg13g2_fill_2 FILLER_50_996 ();
 sg13g2_decap_4 FILLER_50_1002 ();
 sg13g2_decap_8 FILLER_50_1011 ();
 sg13g2_decap_4 FILLER_50_1018 ();
 sg13g2_fill_1 FILLER_50_1031 ();
 sg13g2_fill_2 FILLER_50_1036 ();
 sg13g2_decap_4 FILLER_50_1102 ();
 sg13g2_fill_1 FILLER_50_1106 ();
 sg13g2_decap_8 FILLER_50_1112 ();
 sg13g2_decap_8 FILLER_50_1119 ();
 sg13g2_decap_4 FILLER_50_1126 ();
 sg13g2_fill_1 FILLER_50_1130 ();
 sg13g2_fill_2 FILLER_50_1141 ();
 sg13g2_fill_1 FILLER_50_1143 ();
 sg13g2_decap_4 FILLER_50_1148 ();
 sg13g2_decap_8 FILLER_50_1160 ();
 sg13g2_decap_4 FILLER_50_1167 ();
 sg13g2_fill_2 FILLER_50_1175 ();
 sg13g2_decap_8 FILLER_50_1185 ();
 sg13g2_decap_4 FILLER_50_1192 ();
 sg13g2_decap_4 FILLER_50_1201 ();
 sg13g2_decap_8 FILLER_50_1209 ();
 sg13g2_fill_2 FILLER_50_1216 ();
 sg13g2_decap_4 FILLER_50_1226 ();
 sg13g2_fill_1 FILLER_50_1230 ();
 sg13g2_decap_8 FILLER_50_1235 ();
 sg13g2_decap_4 FILLER_50_1242 ();
 sg13g2_fill_1 FILLER_50_1250 ();
 sg13g2_decap_8 FILLER_50_1256 ();
 sg13g2_decap_4 FILLER_50_1263 ();
 sg13g2_fill_1 FILLER_50_1267 ();
 sg13g2_fill_2 FILLER_50_1281 ();
 sg13g2_fill_1 FILLER_50_1283 ();
 sg13g2_fill_1 FILLER_50_1318 ();
 sg13g2_decap_8 FILLER_50_1336 ();
 sg13g2_fill_1 FILLER_50_1348 ();
 sg13g2_fill_1 FILLER_50_1362 ();
 sg13g2_decap_4 FILLER_50_1381 ();
 sg13g2_fill_1 FILLER_50_1385 ();
 sg13g2_fill_1 FILLER_50_1396 ();
 sg13g2_decap_4 FILLER_50_1402 ();
 sg13g2_fill_1 FILLER_50_1414 ();
 sg13g2_fill_2 FILLER_50_1420 ();
 sg13g2_decap_4 FILLER_50_1427 ();
 sg13g2_decap_8 FILLER_50_1461 ();
 sg13g2_decap_4 FILLER_50_1468 ();
 sg13g2_decap_8 FILLER_50_1498 ();
 sg13g2_decap_8 FILLER_50_1505 ();
 sg13g2_fill_2 FILLER_50_1512 ();
 sg13g2_fill_1 FILLER_50_1530 ();
 sg13g2_decap_4 FILLER_50_1536 ();
 sg13g2_fill_1 FILLER_50_1545 ();
 sg13g2_fill_2 FILLER_50_1551 ();
 sg13g2_fill_1 FILLER_50_1553 ();
 sg13g2_decap_8 FILLER_50_1558 ();
 sg13g2_decap_8 FILLER_50_1565 ();
 sg13g2_fill_2 FILLER_50_1572 ();
 sg13g2_fill_1 FILLER_50_1574 ();
 sg13g2_decap_8 FILLER_50_1606 ();
 sg13g2_fill_2 FILLER_50_1613 ();
 sg13g2_decap_8 FILLER_50_1620 ();
 sg13g2_decap_8 FILLER_50_1627 ();
 sg13g2_decap_4 FILLER_50_1634 ();
 sg13g2_fill_1 FILLER_50_1638 ();
 sg13g2_decap_8 FILLER_50_1644 ();
 sg13g2_decap_8 FILLER_50_1670 ();
 sg13g2_decap_8 FILLER_50_1677 ();
 sg13g2_decap_4 FILLER_50_1684 ();
 sg13g2_fill_1 FILLER_50_1688 ();
 sg13g2_fill_1 FILLER_50_1712 ();
 sg13g2_fill_2 FILLER_50_1740 ();
 sg13g2_fill_1 FILLER_50_1742 ();
 sg13g2_fill_1 FILLER_50_1773 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_11 ();
 sg13g2_decap_4 FILLER_51_18 ();
 sg13g2_fill_1 FILLER_51_22 ();
 sg13g2_fill_1 FILLER_51_27 ();
 sg13g2_fill_1 FILLER_51_46 ();
 sg13g2_decap_4 FILLER_51_57 ();
 sg13g2_fill_2 FILLER_51_94 ();
 sg13g2_fill_1 FILLER_51_96 ();
 sg13g2_decap_8 FILLER_51_109 ();
 sg13g2_decap_8 FILLER_51_121 ();
 sg13g2_fill_1 FILLER_51_128 ();
 sg13g2_fill_1 FILLER_51_152 ();
 sg13g2_fill_2 FILLER_51_157 ();
 sg13g2_decap_4 FILLER_51_164 ();
 sg13g2_fill_1 FILLER_51_177 ();
 sg13g2_fill_1 FILLER_51_189 ();
 sg13g2_fill_1 FILLER_51_194 ();
 sg13g2_decap_4 FILLER_51_215 ();
 sg13g2_fill_2 FILLER_51_219 ();
 sg13g2_decap_8 FILLER_51_250 ();
 sg13g2_decap_8 FILLER_51_257 ();
 sg13g2_fill_1 FILLER_51_276 ();
 sg13g2_fill_2 FILLER_51_292 ();
 sg13g2_decap_8 FILLER_51_298 ();
 sg13g2_fill_2 FILLER_51_305 ();
 sg13g2_fill_2 FILLER_51_317 ();
 sg13g2_fill_1 FILLER_51_319 ();
 sg13g2_decap_4 FILLER_51_324 ();
 sg13g2_fill_2 FILLER_51_328 ();
 sg13g2_fill_1 FILLER_51_352 ();
 sg13g2_decap_4 FILLER_51_360 ();
 sg13g2_fill_2 FILLER_51_364 ();
 sg13g2_fill_2 FILLER_51_376 ();
 sg13g2_fill_1 FILLER_51_378 ();
 sg13g2_fill_1 FILLER_51_393 ();
 sg13g2_decap_4 FILLER_51_406 ();
 sg13g2_fill_2 FILLER_51_415 ();
 sg13g2_fill_1 FILLER_51_417 ();
 sg13g2_decap_4 FILLER_51_425 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_decap_4 FILLER_51_434 ();
 sg13g2_decap_4 FILLER_51_458 ();
 sg13g2_fill_2 FILLER_51_462 ();
 sg13g2_fill_1 FILLER_51_469 ();
 sg13g2_decap_4 FILLER_51_485 ();
 sg13g2_fill_1 FILLER_51_489 ();
 sg13g2_decap_8 FILLER_51_495 ();
 sg13g2_decap_8 FILLER_51_502 ();
 sg13g2_decap_4 FILLER_51_509 ();
 sg13g2_fill_1 FILLER_51_513 ();
 sg13g2_decap_4 FILLER_51_519 ();
 sg13g2_fill_2 FILLER_51_529 ();
 sg13g2_fill_1 FILLER_51_531 ();
 sg13g2_fill_2 FILLER_51_538 ();
 sg13g2_decap_4 FILLER_51_544 ();
 sg13g2_fill_1 FILLER_51_548 ();
 sg13g2_decap_4 FILLER_51_554 ();
 sg13g2_fill_1 FILLER_51_558 ();
 sg13g2_fill_1 FILLER_51_564 ();
 sg13g2_fill_1 FILLER_51_583 ();
 sg13g2_decap_8 FILLER_51_592 ();
 sg13g2_decap_4 FILLER_51_599 ();
 sg13g2_fill_2 FILLER_51_603 ();
 sg13g2_fill_2 FILLER_51_617 ();
 sg13g2_decap_4 FILLER_51_622 ();
 sg13g2_fill_1 FILLER_51_626 ();
 sg13g2_decap_8 FILLER_51_632 ();
 sg13g2_decap_8 FILLER_51_639 ();
 sg13g2_decap_8 FILLER_51_646 ();
 sg13g2_decap_8 FILLER_51_657 ();
 sg13g2_decap_8 FILLER_51_664 ();
 sg13g2_decap_8 FILLER_51_671 ();
 sg13g2_fill_1 FILLER_51_678 ();
 sg13g2_fill_1 FILLER_51_738 ();
 sg13g2_decap_8 FILLER_51_748 ();
 sg13g2_decap_8 FILLER_51_755 ();
 sg13g2_fill_2 FILLER_51_762 ();
 sg13g2_fill_2 FILLER_51_778 ();
 sg13g2_fill_1 FILLER_51_780 ();
 sg13g2_decap_4 FILLER_51_786 ();
 sg13g2_decap_4 FILLER_51_795 ();
 sg13g2_decap_4 FILLER_51_813 ();
 sg13g2_fill_1 FILLER_51_817 ();
 sg13g2_fill_1 FILLER_51_832 ();
 sg13g2_fill_1 FILLER_51_842 ();
 sg13g2_decap_8 FILLER_51_848 ();
 sg13g2_fill_2 FILLER_51_855 ();
 sg13g2_decap_4 FILLER_51_865 ();
 sg13g2_fill_2 FILLER_51_869 ();
 sg13g2_fill_1 FILLER_51_905 ();
 sg13g2_fill_2 FILLER_51_910 ();
 sg13g2_fill_2 FILLER_51_917 ();
 sg13g2_decap_8 FILLER_51_926 ();
 sg13g2_decap_4 FILLER_51_938 ();
 sg13g2_fill_1 FILLER_51_951 ();
 sg13g2_fill_1 FILLER_51_957 ();
 sg13g2_fill_2 FILLER_51_1023 ();
 sg13g2_decap_4 FILLER_51_1030 ();
 sg13g2_decap_4 FILLER_51_1085 ();
 sg13g2_decap_8 FILLER_51_1095 ();
 sg13g2_fill_1 FILLER_51_1102 ();
 sg13g2_decap_8 FILLER_51_1108 ();
 sg13g2_fill_1 FILLER_51_1115 ();
 sg13g2_decap_4 FILLER_51_1126 ();
 sg13g2_fill_2 FILLER_51_1130 ();
 sg13g2_decap_8 FILLER_51_1151 ();
 sg13g2_fill_1 FILLER_51_1158 ();
 sg13g2_decap_4 FILLER_51_1194 ();
 sg13g2_decap_8 FILLER_51_1227 ();
 sg13g2_fill_2 FILLER_51_1247 ();
 sg13g2_fill_1 FILLER_51_1249 ();
 sg13g2_fill_2 FILLER_51_1260 ();
 sg13g2_fill_1 FILLER_51_1262 ();
 sg13g2_fill_1 FILLER_51_1273 ();
 sg13g2_decap_4 FILLER_51_1279 ();
 sg13g2_fill_2 FILLER_51_1283 ();
 sg13g2_decap_4 FILLER_51_1290 ();
 sg13g2_fill_2 FILLER_51_1294 ();
 sg13g2_fill_1 FILLER_51_1300 ();
 sg13g2_fill_2 FILLER_51_1320 ();
 sg13g2_decap_8 FILLER_51_1329 ();
 sg13g2_decap_4 FILLER_51_1336 ();
 sg13g2_fill_1 FILLER_51_1353 ();
 sg13g2_decap_4 FILLER_51_1369 ();
 sg13g2_fill_1 FILLER_51_1373 ();
 sg13g2_fill_1 FILLER_51_1387 ();
 sg13g2_decap_8 FILLER_51_1392 ();
 sg13g2_decap_8 FILLER_51_1399 ();
 sg13g2_decap_8 FILLER_51_1415 ();
 sg13g2_fill_2 FILLER_51_1422 ();
 sg13g2_decap_4 FILLER_51_1450 ();
 sg13g2_decap_8 FILLER_51_1458 ();
 sg13g2_decap_8 FILLER_51_1484 ();
 sg13g2_decap_4 FILLER_51_1491 ();
 sg13g2_fill_1 FILLER_51_1502 ();
 sg13g2_decap_8 FILLER_51_1507 ();
 sg13g2_decap_4 FILLER_51_1514 ();
 sg13g2_decap_8 FILLER_51_1536 ();
 sg13g2_fill_1 FILLER_51_1573 ();
 sg13g2_decap_8 FILLER_51_1578 ();
 sg13g2_fill_1 FILLER_51_1585 ();
 sg13g2_decap_8 FILLER_51_1590 ();
 sg13g2_decap_4 FILLER_51_1597 ();
 sg13g2_fill_2 FILLER_51_1627 ();
 sg13g2_fill_1 FILLER_51_1629 ();
 sg13g2_decap_8 FILLER_51_1669 ();
 sg13g2_decap_8 FILLER_51_1676 ();
 sg13g2_decap_4 FILLER_51_1683 ();
 sg13g2_fill_2 FILLER_51_1721 ();
 sg13g2_fill_2 FILLER_51_1729 ();
 sg13g2_fill_1 FILLER_51_1731 ();
 sg13g2_decap_4 FILLER_51_1737 ();
 sg13g2_decap_4 FILLER_51_1750 ();
 sg13g2_fill_2 FILLER_51_1758 ();
 sg13g2_fill_1 FILLER_51_1760 ();
 sg13g2_decap_8 FILLER_51_1765 ();
 sg13g2_fill_2 FILLER_51_1772 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_46 ();
 sg13g2_decap_8 FILLER_52_58 ();
 sg13g2_decap_4 FILLER_52_65 ();
 sg13g2_fill_1 FILLER_52_78 ();
 sg13g2_fill_1 FILLER_52_83 ();
 sg13g2_decap_4 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_95 ();
 sg13g2_decap_8 FILLER_52_116 ();
 sg13g2_fill_2 FILLER_52_123 ();
 sg13g2_fill_1 FILLER_52_125 ();
 sg13g2_fill_1 FILLER_52_131 ();
 sg13g2_decap_4 FILLER_52_137 ();
 sg13g2_fill_2 FILLER_52_145 ();
 sg13g2_fill_1 FILLER_52_151 ();
 sg13g2_decap_4 FILLER_52_161 ();
 sg13g2_fill_2 FILLER_52_170 ();
 sg13g2_fill_1 FILLER_52_183 ();
 sg13g2_decap_8 FILLER_52_188 ();
 sg13g2_decap_8 FILLER_52_195 ();
 sg13g2_fill_1 FILLER_52_202 ();
 sg13g2_fill_2 FILLER_52_215 ();
 sg13g2_fill_1 FILLER_52_229 ();
 sg13g2_fill_1 FILLER_52_251 ();
 sg13g2_fill_1 FILLER_52_256 ();
 sg13g2_fill_2 FILLER_52_276 ();
 sg13g2_fill_1 FILLER_52_278 ();
 sg13g2_decap_8 FILLER_52_287 ();
 sg13g2_decap_4 FILLER_52_294 ();
 sg13g2_decap_4 FILLER_52_303 ();
 sg13g2_fill_1 FILLER_52_307 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_decap_8 FILLER_52_336 ();
 sg13g2_decap_4 FILLER_52_343 ();
 sg13g2_fill_2 FILLER_52_361 ();
 sg13g2_decap_8 FILLER_52_368 ();
 sg13g2_decap_4 FILLER_52_375 ();
 sg13g2_fill_2 FILLER_52_379 ();
 sg13g2_fill_1 FILLER_52_392 ();
 sg13g2_decap_4 FILLER_52_406 ();
 sg13g2_fill_1 FILLER_52_410 ();
 sg13g2_fill_2 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_52_436 ();
 sg13g2_decap_8 FILLER_52_443 ();
 sg13g2_decap_8 FILLER_52_450 ();
 sg13g2_decap_8 FILLER_52_457 ();
 sg13g2_decap_4 FILLER_52_464 ();
 sg13g2_fill_2 FILLER_52_472 ();
 sg13g2_fill_1 FILLER_52_474 ();
 sg13g2_decap_4 FILLER_52_480 ();
 sg13g2_fill_1 FILLER_52_484 ();
 sg13g2_decap_8 FILLER_52_491 ();
 sg13g2_decap_8 FILLER_52_498 ();
 sg13g2_decap_4 FILLER_52_505 ();
 sg13g2_fill_1 FILLER_52_509 ();
 sg13g2_decap_8 FILLER_52_514 ();
 sg13g2_decap_4 FILLER_52_521 ();
 sg13g2_fill_2 FILLER_52_529 ();
 sg13g2_fill_1 FILLER_52_531 ();
 sg13g2_fill_2 FILLER_52_537 ();
 sg13g2_fill_2 FILLER_52_565 ();
 sg13g2_decap_4 FILLER_52_618 ();
 sg13g2_decap_4 FILLER_52_649 ();
 sg13g2_fill_1 FILLER_52_659 ();
 sg13g2_fill_1 FILLER_52_664 ();
 sg13g2_fill_2 FILLER_52_671 ();
 sg13g2_fill_1 FILLER_52_688 ();
 sg13g2_fill_2 FILLER_52_700 ();
 sg13g2_fill_2 FILLER_52_732 ();
 sg13g2_decap_8 FILLER_52_739 ();
 sg13g2_fill_2 FILLER_52_746 ();
 sg13g2_fill_2 FILLER_52_752 ();
 sg13g2_fill_2 FILLER_52_780 ();
 sg13g2_fill_1 FILLER_52_782 ();
 sg13g2_fill_2 FILLER_52_788 ();
 sg13g2_fill_1 FILLER_52_790 ();
 sg13g2_decap_8 FILLER_52_821 ();
 sg13g2_fill_1 FILLER_52_828 ();
 sg13g2_fill_2 FILLER_52_833 ();
 sg13g2_fill_1 FILLER_52_842 ();
 sg13g2_fill_2 FILLER_52_848 ();
 sg13g2_fill_1 FILLER_52_881 ();
 sg13g2_fill_2 FILLER_52_887 ();
 sg13g2_fill_2 FILLER_52_892 ();
 sg13g2_fill_2 FILLER_52_898 ();
 sg13g2_fill_2 FILLER_52_921 ();
 sg13g2_fill_1 FILLER_52_923 ();
 sg13g2_fill_2 FILLER_52_956 ();
 sg13g2_decap_8 FILLER_52_982 ();
 sg13g2_fill_2 FILLER_52_989 ();
 sg13g2_fill_2 FILLER_52_996 ();
 sg13g2_decap_8 FILLER_52_1002 ();
 sg13g2_decap_8 FILLER_52_1009 ();
 sg13g2_decap_8 FILLER_52_1016 ();
 sg13g2_decap_8 FILLER_52_1023 ();
 sg13g2_decap_8 FILLER_52_1030 ();
 sg13g2_decap_4 FILLER_52_1037 ();
 sg13g2_decap_4 FILLER_52_1080 ();
 sg13g2_decap_4 FILLER_52_1091 ();
 sg13g2_fill_1 FILLER_52_1095 ();
 sg13g2_fill_2 FILLER_52_1124 ();
 sg13g2_decap_4 FILLER_52_1135 ();
 sg13g2_fill_1 FILLER_52_1139 ();
 sg13g2_fill_2 FILLER_52_1149 ();
 sg13g2_decap_8 FILLER_52_1163 ();
 sg13g2_decap_8 FILLER_52_1170 ();
 sg13g2_decap_4 FILLER_52_1177 ();
 sg13g2_fill_2 FILLER_52_1181 ();
 sg13g2_fill_2 FILLER_52_1203 ();
 sg13g2_fill_1 FILLER_52_1205 ();
 sg13g2_decap_8 FILLER_52_1222 ();
 sg13g2_decap_4 FILLER_52_1229 ();
 sg13g2_fill_1 FILLER_52_1233 ();
 sg13g2_decap_8 FILLER_52_1242 ();
 sg13g2_fill_2 FILLER_52_1249 ();
 sg13g2_decap_4 FILLER_52_1256 ();
 sg13g2_fill_2 FILLER_52_1260 ();
 sg13g2_decap_8 FILLER_52_1266 ();
 sg13g2_fill_1 FILLER_52_1273 ();
 sg13g2_fill_2 FILLER_52_1279 ();
 sg13g2_decap_4 FILLER_52_1286 ();
 sg13g2_fill_2 FILLER_52_1294 ();
 sg13g2_fill_2 FILLER_52_1314 ();
 sg13g2_fill_1 FILLER_52_1316 ();
 sg13g2_decap_8 FILLER_52_1322 ();
 sg13g2_decap_8 FILLER_52_1329 ();
 sg13g2_decap_4 FILLER_52_1336 ();
 sg13g2_decap_8 FILLER_52_1349 ();
 sg13g2_fill_2 FILLER_52_1356 ();
 sg13g2_decap_4 FILLER_52_1366 ();
 sg13g2_decap_4 FILLER_52_1382 ();
 sg13g2_fill_2 FILLER_52_1386 ();
 sg13g2_fill_2 FILLER_52_1393 ();
 sg13g2_fill_2 FILLER_52_1444 ();
 sg13g2_fill_1 FILLER_52_1446 ();
 sg13g2_decap_8 FILLER_52_1454 ();
 sg13g2_fill_1 FILLER_52_1461 ();
 sg13g2_fill_2 FILLER_52_1472 ();
 sg13g2_decap_8 FILLER_52_1508 ();
 sg13g2_fill_1 FILLER_52_1515 ();
 sg13g2_decap_8 FILLER_52_1539 ();
 sg13g2_fill_1 FILLER_52_1546 ();
 sg13g2_fill_2 FILLER_52_1559 ();
 sg13g2_fill_1 FILLER_52_1561 ();
 sg13g2_decap_4 FILLER_52_1609 ();
 sg13g2_fill_1 FILLER_52_1613 ();
 sg13g2_decap_8 FILLER_52_1623 ();
 sg13g2_decap_8 FILLER_52_1657 ();
 sg13g2_decap_4 FILLER_52_1664 ();
 sg13g2_fill_2 FILLER_52_1668 ();
 sg13g2_decap_8 FILLER_52_1679 ();
 sg13g2_decap_8 FILLER_52_1686 ();
 sg13g2_decap_4 FILLER_52_1698 ();
 sg13g2_decap_8 FILLER_52_1706 ();
 sg13g2_decap_4 FILLER_52_1713 ();
 sg13g2_decap_4 FILLER_52_1720 ();
 sg13g2_fill_1 FILLER_52_1724 ();
 sg13g2_fill_1 FILLER_52_1729 ();
 sg13g2_decap_4 FILLER_52_1770 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_2 ();
 sg13g2_decap_8 FILLER_53_8 ();
 sg13g2_fill_2 FILLER_53_15 ();
 sg13g2_fill_1 FILLER_53_17 ();
 sg13g2_decap_8 FILLER_53_55 ();
 sg13g2_fill_1 FILLER_53_75 ();
 sg13g2_fill_2 FILLER_53_89 ();
 sg13g2_fill_1 FILLER_53_102 ();
 sg13g2_fill_2 FILLER_53_109 ();
 sg13g2_decap_8 FILLER_53_120 ();
 sg13g2_fill_1 FILLER_53_127 ();
 sg13g2_fill_2 FILLER_53_140 ();
 sg13g2_decap_4 FILLER_53_150 ();
 sg13g2_fill_2 FILLER_53_173 ();
 sg13g2_fill_1 FILLER_53_175 ();
 sg13g2_decap_4 FILLER_53_188 ();
 sg13g2_fill_2 FILLER_53_192 ();
 sg13g2_fill_2 FILLER_53_202 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_4 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_236 ();
 sg13g2_decap_8 FILLER_53_243 ();
 sg13g2_fill_1 FILLER_53_255 ();
 sg13g2_decap_4 FILLER_53_269 ();
 sg13g2_fill_2 FILLER_53_273 ();
 sg13g2_fill_1 FILLER_53_302 ();
 sg13g2_fill_1 FILLER_53_307 ();
 sg13g2_fill_1 FILLER_53_313 ();
 sg13g2_fill_1 FILLER_53_319 ();
 sg13g2_fill_1 FILLER_53_326 ();
 sg13g2_fill_2 FILLER_53_335 ();
 sg13g2_fill_2 FILLER_53_341 ();
 sg13g2_fill_2 FILLER_53_348 ();
 sg13g2_fill_1 FILLER_53_350 ();
 sg13g2_decap_8 FILLER_53_357 ();
 sg13g2_decap_4 FILLER_53_364 ();
 sg13g2_fill_1 FILLER_53_368 ();
 sg13g2_decap_4 FILLER_53_397 ();
 sg13g2_fill_2 FILLER_53_401 ();
 sg13g2_decap_8 FILLER_53_414 ();
 sg13g2_decap_4 FILLER_53_421 ();
 sg13g2_decap_8 FILLER_53_439 ();
 sg13g2_decap_8 FILLER_53_446 ();
 sg13g2_decap_8 FILLER_53_453 ();
 sg13g2_decap_4 FILLER_53_460 ();
 sg13g2_fill_2 FILLER_53_464 ();
 sg13g2_fill_2 FILLER_53_476 ();
 sg13g2_fill_1 FILLER_53_482 ();
 sg13g2_fill_2 FILLER_53_493 ();
 sg13g2_decap_4 FILLER_53_499 ();
 sg13g2_fill_1 FILLER_53_513 ();
 sg13g2_decap_4 FILLER_53_518 ();
 sg13g2_decap_8 FILLER_53_534 ();
 sg13g2_decap_4 FILLER_53_541 ();
 sg13g2_fill_1 FILLER_53_545 ();
 sg13g2_decap_4 FILLER_53_550 ();
 sg13g2_fill_1 FILLER_53_554 ();
 sg13g2_fill_1 FILLER_53_565 ();
 sg13g2_fill_2 FILLER_53_575 ();
 sg13g2_fill_1 FILLER_53_577 ();
 sg13g2_decap_8 FILLER_53_583 ();
 sg13g2_decap_8 FILLER_53_590 ();
 sg13g2_decap_4 FILLER_53_597 ();
 sg13g2_decap_8 FILLER_53_620 ();
 sg13g2_fill_1 FILLER_53_627 ();
 sg13g2_decap_8 FILLER_53_664 ();
 sg13g2_decap_8 FILLER_53_671 ();
 sg13g2_decap_4 FILLER_53_678 ();
 sg13g2_fill_1 FILLER_53_685 ();
 sg13g2_decap_8 FILLER_53_696 ();
 sg13g2_decap_8 FILLER_53_708 ();
 sg13g2_fill_1 FILLER_53_722 ();
 sg13g2_decap_8 FILLER_53_732 ();
 sg13g2_decap_4 FILLER_53_739 ();
 sg13g2_fill_2 FILLER_53_743 ();
 sg13g2_decap_8 FILLER_53_749 ();
 sg13g2_decap_4 FILLER_53_756 ();
 sg13g2_decap_8 FILLER_53_764 ();
 sg13g2_fill_1 FILLER_53_771 ();
 sg13g2_decap_8 FILLER_53_777 ();
 sg13g2_decap_8 FILLER_53_784 ();
 sg13g2_fill_2 FILLER_53_791 ();
 sg13g2_fill_1 FILLER_53_803 ();
 sg13g2_decap_8 FILLER_53_808 ();
 sg13g2_decap_4 FILLER_53_815 ();
 sg13g2_fill_1 FILLER_53_819 ();
 sg13g2_fill_2 FILLER_53_851 ();
 sg13g2_fill_1 FILLER_53_853 ();
 sg13g2_decap_8 FILLER_53_861 ();
 sg13g2_fill_2 FILLER_53_868 ();
 sg13g2_fill_1 FILLER_53_870 ();
 sg13g2_fill_1 FILLER_53_879 ();
 sg13g2_fill_1 FILLER_53_885 ();
 sg13g2_decap_4 FILLER_53_916 ();
 sg13g2_fill_2 FILLER_53_920 ();
 sg13g2_decap_8 FILLER_53_927 ();
 sg13g2_decap_8 FILLER_53_934 ();
 sg13g2_decap_4 FILLER_53_941 ();
 sg13g2_fill_1 FILLER_53_945 ();
 sg13g2_fill_2 FILLER_53_951 ();
 sg13g2_decap_8 FILLER_53_970 ();
 sg13g2_fill_2 FILLER_53_977 ();
 sg13g2_decap_4 FILLER_53_992 ();
 sg13g2_fill_1 FILLER_53_996 ();
 sg13g2_decap_8 FILLER_53_1015 ();
 sg13g2_fill_1 FILLER_53_1022 ();
 sg13g2_fill_1 FILLER_53_1026 ();
 sg13g2_decap_4 FILLER_53_1035 ();
 sg13g2_fill_2 FILLER_53_1049 ();
 sg13g2_fill_1 FILLER_53_1051 ();
 sg13g2_fill_1 FILLER_53_1056 ();
 sg13g2_fill_1 FILLER_53_1075 ();
 sg13g2_fill_2 FILLER_53_1081 ();
 sg13g2_fill_2 FILLER_53_1101 ();
 sg13g2_fill_1 FILLER_53_1103 ();
 sg13g2_decap_8 FILLER_53_1130 ();
 sg13g2_fill_1 FILLER_53_1137 ();
 sg13g2_decap_4 FILLER_53_1142 ();
 sg13g2_decap_8 FILLER_53_1172 ();
 sg13g2_decap_8 FILLER_53_1189 ();
 sg13g2_decap_4 FILLER_53_1196 ();
 sg13g2_fill_1 FILLER_53_1200 ();
 sg13g2_decap_4 FILLER_53_1206 ();
 sg13g2_fill_1 FILLER_53_1210 ();
 sg13g2_fill_2 FILLER_53_1216 ();
 sg13g2_decap_4 FILLER_53_1222 ();
 sg13g2_decap_8 FILLER_53_1229 ();
 sg13g2_fill_2 FILLER_53_1236 ();
 sg13g2_fill_1 FILLER_53_1238 ();
 sg13g2_decap_4 FILLER_53_1286 ();
 sg13g2_decap_4 FILLER_53_1299 ();
 sg13g2_fill_2 FILLER_53_1303 ();
 sg13g2_decap_4 FILLER_53_1309 ();
 sg13g2_decap_4 FILLER_53_1325 ();
 sg13g2_fill_1 FILLER_53_1346 ();
 sg13g2_fill_2 FILLER_53_1352 ();
 sg13g2_fill_1 FILLER_53_1354 ();
 sg13g2_fill_2 FILLER_53_1406 ();
 sg13g2_fill_1 FILLER_53_1408 ();
 sg13g2_fill_2 FILLER_53_1414 ();
 sg13g2_fill_1 FILLER_53_1416 ();
 sg13g2_decap_8 FILLER_53_1425 ();
 sg13g2_decap_8 FILLER_53_1436 ();
 sg13g2_decap_8 FILLER_53_1443 ();
 sg13g2_fill_2 FILLER_53_1458 ();
 sg13g2_fill_2 FILLER_53_1468 ();
 sg13g2_fill_2 FILLER_53_1479 ();
 sg13g2_decap_8 FILLER_53_1485 ();
 sg13g2_decap_8 FILLER_53_1492 ();
 sg13g2_decap_4 FILLER_53_1499 ();
 sg13g2_decap_4 FILLER_53_1508 ();
 sg13g2_fill_1 FILLER_53_1512 ();
 sg13g2_fill_2 FILLER_53_1518 ();
 sg13g2_decap_8 FILLER_53_1525 ();
 sg13g2_decap_4 FILLER_53_1532 ();
 sg13g2_fill_1 FILLER_53_1544 ();
 sg13g2_decap_8 FILLER_53_1551 ();
 sg13g2_decap_8 FILLER_53_1558 ();
 sg13g2_fill_2 FILLER_53_1565 ();
 sg13g2_fill_1 FILLER_53_1567 ();
 sg13g2_decap_8 FILLER_53_1581 ();
 sg13g2_decap_4 FILLER_53_1588 ();
 sg13g2_fill_1 FILLER_53_1592 ();
 sg13g2_decap_8 FILLER_53_1597 ();
 sg13g2_decap_4 FILLER_53_1609 ();
 sg13g2_decap_4 FILLER_53_1639 ();
 sg13g2_decap_4 FILLER_53_1660 ();
 sg13g2_fill_1 FILLER_53_1694 ();
 sg13g2_decap_4 FILLER_53_1744 ();
 sg13g2_fill_1 FILLER_53_1748 ();
 sg13g2_decap_8 FILLER_53_1753 ();
 sg13g2_decap_8 FILLER_53_1760 ();
 sg13g2_decap_8 FILLER_53_1767 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_4 FILLER_54_21 ();
 sg13g2_fill_1 FILLER_54_25 ();
 sg13g2_fill_2 FILLER_54_31 ();
 sg13g2_fill_1 FILLER_54_33 ();
 sg13g2_decap_8 FILLER_54_53 ();
 sg13g2_fill_1 FILLER_54_60 ();
 sg13g2_decap_8 FILLER_54_66 ();
 sg13g2_fill_1 FILLER_54_73 ();
 sg13g2_decap_8 FILLER_54_78 ();
 sg13g2_decap_8 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_97 ();
 sg13g2_decap_8 FILLER_54_102 ();
 sg13g2_decap_4 FILLER_54_109 ();
 sg13g2_fill_1 FILLER_54_113 ();
 sg13g2_fill_2 FILLER_54_119 ();
 sg13g2_fill_1 FILLER_54_121 ();
 sg13g2_fill_2 FILLER_54_126 ();
 sg13g2_decap_4 FILLER_54_143 ();
 sg13g2_decap_8 FILLER_54_153 ();
 sg13g2_decap_8 FILLER_54_160 ();
 sg13g2_decap_4 FILLER_54_167 ();
 sg13g2_fill_1 FILLER_54_171 ();
 sg13g2_fill_2 FILLER_54_182 ();
 sg13g2_fill_2 FILLER_54_189 ();
 sg13g2_fill_1 FILLER_54_191 ();
 sg13g2_fill_1 FILLER_54_196 ();
 sg13g2_fill_2 FILLER_54_205 ();
 sg13g2_fill_1 FILLER_54_207 ();
 sg13g2_decap_8 FILLER_54_213 ();
 sg13g2_fill_2 FILLER_54_220 ();
 sg13g2_decap_4 FILLER_54_227 ();
 sg13g2_fill_1 FILLER_54_231 ();
 sg13g2_fill_2 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_241 ();
 sg13g2_fill_1 FILLER_54_263 ();
 sg13g2_decap_8 FILLER_54_269 ();
 sg13g2_decap_4 FILLER_54_276 ();
 sg13g2_fill_1 FILLER_54_280 ();
 sg13g2_fill_1 FILLER_54_291 ();
 sg13g2_decap_8 FILLER_54_297 ();
 sg13g2_fill_1 FILLER_54_304 ();
 sg13g2_fill_1 FILLER_54_311 ();
 sg13g2_fill_2 FILLER_54_316 ();
 sg13g2_fill_1 FILLER_54_318 ();
 sg13g2_decap_8 FILLER_54_323 ();
 sg13g2_fill_2 FILLER_54_335 ();
 sg13g2_decap_4 FILLER_54_348 ();
 sg13g2_fill_1 FILLER_54_352 ();
 sg13g2_decap_8 FILLER_54_362 ();
 sg13g2_decap_8 FILLER_54_369 ();
 sg13g2_decap_4 FILLER_54_376 ();
 sg13g2_fill_2 FILLER_54_380 ();
 sg13g2_decap_4 FILLER_54_393 ();
 sg13g2_fill_2 FILLER_54_397 ();
 sg13g2_decap_4 FILLER_54_404 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_fill_2 FILLER_54_417 ();
 sg13g2_decap_8 FILLER_54_427 ();
 sg13g2_decap_4 FILLER_54_434 ();
 sg13g2_fill_2 FILLER_54_438 ();
 sg13g2_decap_4 FILLER_54_452 ();
 sg13g2_decap_8 FILLER_54_460 ();
 sg13g2_fill_2 FILLER_54_472 ();
 sg13g2_decap_8 FILLER_54_478 ();
 sg13g2_decap_8 FILLER_54_485 ();
 sg13g2_fill_2 FILLER_54_492 ();
 sg13g2_decap_8 FILLER_54_499 ();
 sg13g2_decap_8 FILLER_54_510 ();
 sg13g2_decap_8 FILLER_54_517 ();
 sg13g2_fill_1 FILLER_54_524 ();
 sg13g2_decap_4 FILLER_54_530 ();
 sg13g2_fill_1 FILLER_54_534 ();
 sg13g2_decap_8 FILLER_54_539 ();
 sg13g2_decap_8 FILLER_54_546 ();
 sg13g2_fill_2 FILLER_54_553 ();
 sg13g2_fill_1 FILLER_54_559 ();
 sg13g2_fill_1 FILLER_54_591 ();
 sg13g2_fill_1 FILLER_54_595 ();
 sg13g2_decap_4 FILLER_54_600 ();
 sg13g2_decap_8 FILLER_54_628 ();
 sg13g2_fill_2 FILLER_54_635 ();
 sg13g2_fill_1 FILLER_54_637 ();
 sg13g2_decap_8 FILLER_54_642 ();
 sg13g2_decap_4 FILLER_54_649 ();
 sg13g2_fill_1 FILLER_54_653 ();
 sg13g2_fill_2 FILLER_54_658 ();
 sg13g2_fill_1 FILLER_54_660 ();
 sg13g2_decap_4 FILLER_54_676 ();
 sg13g2_fill_2 FILLER_54_680 ();
 sg13g2_fill_2 FILLER_54_726 ();
 sg13g2_fill_1 FILLER_54_728 ();
 sg13g2_fill_2 FILLER_54_765 ();
 sg13g2_fill_2 FILLER_54_793 ();
 sg13g2_fill_1 FILLER_54_795 ();
 sg13g2_fill_1 FILLER_54_799 ();
 sg13g2_decap_8 FILLER_54_803 ();
 sg13g2_decap_8 FILLER_54_810 ();
 sg13g2_decap_8 FILLER_54_817 ();
 sg13g2_fill_2 FILLER_54_824 ();
 sg13g2_fill_2 FILLER_54_830 ();
 sg13g2_fill_1 FILLER_54_832 ();
 sg13g2_decap_4 FILLER_54_839 ();
 sg13g2_fill_1 FILLER_54_843 ();
 sg13g2_decap_8 FILLER_54_849 ();
 sg13g2_fill_1 FILLER_54_856 ();
 sg13g2_fill_1 FILLER_54_867 ();
 sg13g2_fill_1 FILLER_54_873 ();
 sg13g2_fill_1 FILLER_54_879 ();
 sg13g2_fill_2 FILLER_54_884 ();
 sg13g2_decap_4 FILLER_54_891 ();
 sg13g2_fill_2 FILLER_54_895 ();
 sg13g2_decap_4 FILLER_54_901 ();
 sg13g2_decap_8 FILLER_54_915 ();
 sg13g2_decap_8 FILLER_54_922 ();
 sg13g2_decap_8 FILLER_54_929 ();
 sg13g2_decap_8 FILLER_54_936 ();
 sg13g2_fill_2 FILLER_54_943 ();
 sg13g2_fill_1 FILLER_54_956 ();
 sg13g2_fill_1 FILLER_54_968 ();
 sg13g2_decap_4 FILLER_54_975 ();
 sg13g2_decap_8 FILLER_54_1000 ();
 sg13g2_fill_1 FILLER_54_1026 ();
 sg13g2_decap_4 FILLER_54_1032 ();
 sg13g2_fill_1 FILLER_54_1036 ();
 sg13g2_decap_8 FILLER_54_1049 ();
 sg13g2_fill_2 FILLER_54_1056 ();
 sg13g2_decap_8 FILLER_54_1061 ();
 sg13g2_decap_4 FILLER_54_1068 ();
 sg13g2_fill_2 FILLER_54_1072 ();
 sg13g2_decap_8 FILLER_54_1097 ();
 sg13g2_decap_4 FILLER_54_1104 ();
 sg13g2_fill_2 FILLER_54_1108 ();
 sg13g2_decap_8 FILLER_54_1114 ();
 sg13g2_fill_1 FILLER_54_1121 ();
 sg13g2_decap_4 FILLER_54_1128 ();
 sg13g2_fill_2 FILLER_54_1132 ();
 sg13g2_fill_2 FILLER_54_1189 ();
 sg13g2_decap_8 FILLER_54_1203 ();
 sg13g2_decap_8 FILLER_54_1210 ();
 sg13g2_fill_1 FILLER_54_1217 ();
 sg13g2_fill_2 FILLER_54_1264 ();
 sg13g2_fill_1 FILLER_54_1266 ();
 sg13g2_fill_2 FILLER_54_1293 ();
 sg13g2_fill_2 FILLER_54_1301 ();
 sg13g2_fill_2 FILLER_54_1312 ();
 sg13g2_decap_8 FILLER_54_1329 ();
 sg13g2_fill_1 FILLER_54_1336 ();
 sg13g2_decap_8 FILLER_54_1341 ();
 sg13g2_decap_4 FILLER_54_1348 ();
 sg13g2_decap_8 FILLER_54_1356 ();
 sg13g2_decap_8 FILLER_54_1363 ();
 sg13g2_fill_2 FILLER_54_1370 ();
 sg13g2_decap_8 FILLER_54_1389 ();
 sg13g2_decap_4 FILLER_54_1396 ();
 sg13g2_fill_1 FILLER_54_1400 ();
 sg13g2_fill_2 FILLER_54_1405 ();
 sg13g2_fill_2 FILLER_54_1412 ();
 sg13g2_fill_2 FILLER_54_1423 ();
 sg13g2_decap_8 FILLER_54_1435 ();
 sg13g2_fill_1 FILLER_54_1452 ();
 sg13g2_decap_4 FILLER_54_1483 ();
 sg13g2_decap_4 FILLER_54_1541 ();
 sg13g2_decap_4 FILLER_54_1571 ();
 sg13g2_fill_2 FILLER_54_1575 ();
 sg13g2_fill_1 FILLER_54_1585 ();
 sg13g2_decap_8 FILLER_54_1612 ();
 sg13g2_decap_8 FILLER_54_1623 ();
 sg13g2_fill_2 FILLER_54_1630 ();
 sg13g2_fill_1 FILLER_54_1632 ();
 sg13g2_decap_8 FILLER_54_1636 ();
 sg13g2_decap_8 FILLER_54_1669 ();
 sg13g2_decap_8 FILLER_54_1684 ();
 sg13g2_fill_2 FILLER_54_1691 ();
 sg13g2_fill_2 FILLER_54_1707 ();
 sg13g2_fill_2 FILLER_54_1721 ();
 sg13g2_fill_1 FILLER_54_1723 ();
 sg13g2_decap_8 FILLER_54_1728 ();
 sg13g2_fill_2 FILLER_54_1739 ();
 sg13g2_decap_8 FILLER_54_1746 ();
 sg13g2_decap_8 FILLER_54_1753 ();
 sg13g2_decap_8 FILLER_54_1760 ();
 sg13g2_decap_8 FILLER_54_1767 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_4 FILLER_55_52 ();
 sg13g2_fill_2 FILLER_55_56 ();
 sg13g2_decap_4 FILLER_55_70 ();
 sg13g2_fill_2 FILLER_55_74 ();
 sg13g2_fill_2 FILLER_55_91 ();
 sg13g2_fill_1 FILLER_55_102 ();
 sg13g2_decap_8 FILLER_55_108 ();
 sg13g2_decap_8 FILLER_55_121 ();
 sg13g2_fill_2 FILLER_55_128 ();
 sg13g2_decap_4 FILLER_55_140 ();
 sg13g2_decap_4 FILLER_55_148 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_decap_4 FILLER_55_168 ();
 sg13g2_decap_4 FILLER_55_190 ();
 sg13g2_fill_2 FILLER_55_194 ();
 sg13g2_decap_8 FILLER_55_204 ();
 sg13g2_decap_8 FILLER_55_211 ();
 sg13g2_decap_8 FILLER_55_218 ();
 sg13g2_decap_8 FILLER_55_225 ();
 sg13g2_fill_2 FILLER_55_232 ();
 sg13g2_fill_1 FILLER_55_234 ();
 sg13g2_decap_4 FILLER_55_239 ();
 sg13g2_decap_8 FILLER_55_250 ();
 sg13g2_decap_8 FILLER_55_257 ();
 sg13g2_fill_2 FILLER_55_264 ();
 sg13g2_decap_8 FILLER_55_284 ();
 sg13g2_fill_2 FILLER_55_291 ();
 sg13g2_fill_1 FILLER_55_298 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_fill_2 FILLER_55_311 ();
 sg13g2_fill_2 FILLER_55_318 ();
 sg13g2_fill_1 FILLER_55_327 ();
 sg13g2_fill_1 FILLER_55_338 ();
 sg13g2_decap_8 FILLER_55_349 ();
 sg13g2_fill_2 FILLER_55_356 ();
 sg13g2_fill_1 FILLER_55_358 ();
 sg13g2_fill_1 FILLER_55_368 ();
 sg13g2_fill_2 FILLER_55_374 ();
 sg13g2_fill_1 FILLER_55_376 ();
 sg13g2_fill_2 FILLER_55_398 ();
 sg13g2_fill_2 FILLER_55_405 ();
 sg13g2_decap_8 FILLER_55_411 ();
 sg13g2_decap_8 FILLER_55_430 ();
 sg13g2_fill_2 FILLER_55_437 ();
 sg13g2_fill_1 FILLER_55_439 ();
 sg13g2_fill_1 FILLER_55_449 ();
 sg13g2_fill_1 FILLER_55_458 ();
 sg13g2_fill_2 FILLER_55_467 ();
 sg13g2_fill_1 FILLER_55_469 ();
 sg13g2_decap_8 FILLER_55_473 ();
 sg13g2_decap_8 FILLER_55_480 ();
 sg13g2_fill_1 FILLER_55_487 ();
 sg13g2_decap_4 FILLER_55_500 ();
 sg13g2_fill_2 FILLER_55_532 ();
 sg13g2_fill_2 FILLER_55_549 ();
 sg13g2_fill_1 FILLER_55_556 ();
 sg13g2_decap_8 FILLER_55_572 ();
 sg13g2_fill_1 FILLER_55_579 ();
 sg13g2_fill_2 FILLER_55_591 ();
 sg13g2_decap_4 FILLER_55_598 ();
 sg13g2_decap_8 FILLER_55_611 ();
 sg13g2_decap_8 FILLER_55_618 ();
 sg13g2_fill_2 FILLER_55_625 ();
 sg13g2_fill_1 FILLER_55_627 ();
 sg13g2_decap_8 FILLER_55_631 ();
 sg13g2_decap_8 FILLER_55_638 ();
 sg13g2_decap_8 FILLER_55_675 ();
 sg13g2_decap_8 FILLER_55_682 ();
 sg13g2_fill_1 FILLER_55_689 ();
 sg13g2_decap_8 FILLER_55_694 ();
 sg13g2_decap_8 FILLER_55_705 ();
 sg13g2_fill_2 FILLER_55_712 ();
 sg13g2_decap_8 FILLER_55_717 ();
 sg13g2_decap_8 FILLER_55_724 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_fill_2 FILLER_55_737 ();
 sg13g2_fill_1 FILLER_55_739 ();
 sg13g2_decap_8 FILLER_55_754 ();
 sg13g2_fill_2 FILLER_55_778 ();
 sg13g2_decap_4 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_792 ();
 sg13g2_fill_2 FILLER_55_799 ();
 sg13g2_decap_8 FILLER_55_804 ();
 sg13g2_decap_4 FILLER_55_811 ();
 sg13g2_fill_1 FILLER_55_815 ();
 sg13g2_fill_1 FILLER_55_821 ();
 sg13g2_decap_4 FILLER_55_827 ();
 sg13g2_fill_1 FILLER_55_831 ();
 sg13g2_decap_8 FILLER_55_843 ();
 sg13g2_decap_8 FILLER_55_850 ();
 sg13g2_decap_8 FILLER_55_857 ();
 sg13g2_decap_8 FILLER_55_864 ();
 sg13g2_fill_2 FILLER_55_871 ();
 sg13g2_fill_1 FILLER_55_877 ();
 sg13g2_decap_8 FILLER_55_883 ();
 sg13g2_decap_8 FILLER_55_890 ();
 sg13g2_decap_4 FILLER_55_897 ();
 sg13g2_fill_2 FILLER_55_901 ();
 sg13g2_fill_2 FILLER_55_923 ();
 sg13g2_decap_8 FILLER_55_937 ();
 sg13g2_decap_4 FILLER_55_944 ();
 sg13g2_fill_1 FILLER_55_948 ();
 sg13g2_decap_8 FILLER_55_953 ();
 sg13g2_decap_4 FILLER_55_960 ();
 sg13g2_fill_1 FILLER_55_964 ();
 sg13g2_fill_2 FILLER_55_977 ();
 sg13g2_fill_1 FILLER_55_979 ();
 sg13g2_fill_1 FILLER_55_985 ();
 sg13g2_decap_8 FILLER_55_994 ();
 sg13g2_decap_4 FILLER_55_1009 ();
 sg13g2_fill_1 FILLER_55_1013 ();
 sg13g2_fill_1 FILLER_55_1021 ();
 sg13g2_fill_1 FILLER_55_1033 ();
 sg13g2_fill_1 FILLER_55_1044 ();
 sg13g2_fill_2 FILLER_55_1050 ();
 sg13g2_fill_1 FILLER_55_1052 ();
 sg13g2_fill_1 FILLER_55_1069 ();
 sg13g2_fill_2 FILLER_55_1078 ();
 sg13g2_fill_2 FILLER_55_1088 ();
 sg13g2_fill_2 FILLER_55_1094 ();
 sg13g2_decap_8 FILLER_55_1100 ();
 sg13g2_decap_8 FILLER_55_1107 ();
 sg13g2_decap_4 FILLER_55_1114 ();
 sg13g2_fill_1 FILLER_55_1118 ();
 sg13g2_decap_8 FILLER_55_1124 ();
 sg13g2_decap_4 FILLER_55_1131 ();
 sg13g2_fill_2 FILLER_55_1135 ();
 sg13g2_fill_1 FILLER_55_1164 ();
 sg13g2_decap_8 FILLER_55_1174 ();
 sg13g2_fill_2 FILLER_55_1181 ();
 sg13g2_fill_1 FILLER_55_1183 ();
 sg13g2_fill_2 FILLER_55_1196 ();
 sg13g2_fill_1 FILLER_55_1198 ();
 sg13g2_decap_8 FILLER_55_1204 ();
 sg13g2_decap_4 FILLER_55_1211 ();
 sg13g2_decap_4 FILLER_55_1232 ();
 sg13g2_fill_2 FILLER_55_1240 ();
 sg13g2_fill_1 FILLER_55_1242 ();
 sg13g2_fill_2 FILLER_55_1248 ();
 sg13g2_fill_1 FILLER_55_1250 ();
 sg13g2_decap_4 FILLER_55_1261 ();
 sg13g2_decap_4 FILLER_55_1299 ();
 sg13g2_fill_1 FILLER_55_1303 ();
 sg13g2_fill_1 FILLER_55_1310 ();
 sg13g2_decap_4 FILLER_55_1321 ();
 sg13g2_decap_4 FILLER_55_1362 ();
 sg13g2_fill_1 FILLER_55_1418 ();
 sg13g2_fill_2 FILLER_55_1423 ();
 sg13g2_fill_2 FILLER_55_1430 ();
 sg13g2_fill_1 FILLER_55_1437 ();
 sg13g2_decap_4 FILLER_55_1446 ();
 sg13g2_fill_2 FILLER_55_1450 ();
 sg13g2_decap_4 FILLER_55_1473 ();
 sg13g2_decap_8 FILLER_55_1486 ();
 sg13g2_decap_8 FILLER_55_1493 ();
 sg13g2_fill_1 FILLER_55_1500 ();
 sg13g2_decap_4 FILLER_55_1537 ();
 sg13g2_fill_1 FILLER_55_1541 ();
 sg13g2_decap_4 FILLER_55_1558 ();
 sg13g2_fill_1 FILLER_55_1562 ();
 sg13g2_decap_8 FILLER_55_1606 ();
 sg13g2_fill_2 FILLER_55_1613 ();
 sg13g2_fill_1 FILLER_55_1615 ();
 sg13g2_fill_2 FILLER_55_1646 ();
 sg13g2_fill_2 FILLER_55_1652 ();
 sg13g2_fill_1 FILLER_55_1654 ();
 sg13g2_fill_2 FILLER_55_1659 ();
 sg13g2_fill_1 FILLER_55_1661 ();
 sg13g2_decap_8 FILLER_55_1672 ();
 sg13g2_decap_8 FILLER_55_1679 ();
 sg13g2_decap_8 FILLER_55_1686 ();
 sg13g2_decap_4 FILLER_55_1693 ();
 sg13g2_fill_2 FILLER_55_1697 ();
 sg13g2_decap_8 FILLER_55_1749 ();
 sg13g2_decap_8 FILLER_55_1756 ();
 sg13g2_decap_8 FILLER_55_1763 ();
 sg13g2_decap_4 FILLER_55_1770 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_23 ();
 sg13g2_fill_2 FILLER_56_30 ();
 sg13g2_fill_2 FILLER_56_41 ();
 sg13g2_decap_4 FILLER_56_49 ();
 sg13g2_fill_2 FILLER_56_58 ();
 sg13g2_fill_1 FILLER_56_76 ();
 sg13g2_fill_1 FILLER_56_91 ();
 sg13g2_fill_1 FILLER_56_100 ();
 sg13g2_fill_2 FILLER_56_114 ();
 sg13g2_fill_1 FILLER_56_116 ();
 sg13g2_decap_4 FILLER_56_125 ();
 sg13g2_fill_2 FILLER_56_133 ();
 sg13g2_fill_1 FILLER_56_140 ();
 sg13g2_fill_2 FILLER_56_146 ();
 sg13g2_fill_1 FILLER_56_148 ();
 sg13g2_decap_8 FILLER_56_159 ();
 sg13g2_decap_8 FILLER_56_166 ();
 sg13g2_fill_1 FILLER_56_173 ();
 sg13g2_fill_1 FILLER_56_180 ();
 sg13g2_decap_8 FILLER_56_185 ();
 sg13g2_fill_1 FILLER_56_192 ();
 sg13g2_decap_4 FILLER_56_209 ();
 sg13g2_fill_2 FILLER_56_229 ();
 sg13g2_fill_1 FILLER_56_231 ();
 sg13g2_decap_4 FILLER_56_239 ();
 sg13g2_fill_1 FILLER_56_243 ();
 sg13g2_decap_4 FILLER_56_252 ();
 sg13g2_fill_1 FILLER_56_256 ();
 sg13g2_fill_2 FILLER_56_262 ();
 sg13g2_fill_1 FILLER_56_264 ();
 sg13g2_decap_8 FILLER_56_273 ();
 sg13g2_fill_2 FILLER_56_280 ();
 sg13g2_fill_1 FILLER_56_282 ();
 sg13g2_decap_4 FILLER_56_300 ();
 sg13g2_decap_8 FILLER_56_310 ();
 sg13g2_decap_8 FILLER_56_317 ();
 sg13g2_decap_8 FILLER_56_324 ();
 sg13g2_decap_8 FILLER_56_331 ();
 sg13g2_decap_8 FILLER_56_338 ();
 sg13g2_fill_2 FILLER_56_345 ();
 sg13g2_fill_1 FILLER_56_347 ();
 sg13g2_fill_2 FILLER_56_367 ();
 sg13g2_decap_8 FILLER_56_374 ();
 sg13g2_decap_8 FILLER_56_381 ();
 sg13g2_decap_8 FILLER_56_388 ();
 sg13g2_fill_2 FILLER_56_408 ();
 sg13g2_fill_1 FILLER_56_410 ();
 sg13g2_decap_8 FILLER_56_416 ();
 sg13g2_fill_1 FILLER_56_423 ();
 sg13g2_fill_2 FILLER_56_442 ();
 sg13g2_fill_1 FILLER_56_452 ();
 sg13g2_decap_4 FILLER_56_458 ();
 sg13g2_fill_2 FILLER_56_467 ();
 sg13g2_fill_1 FILLER_56_469 ();
 sg13g2_fill_2 FILLER_56_479 ();
 sg13g2_fill_1 FILLER_56_481 ();
 sg13g2_decap_4 FILLER_56_495 ();
 sg13g2_fill_1 FILLER_56_499 ();
 sg13g2_decap_8 FILLER_56_504 ();
 sg13g2_decap_4 FILLER_56_511 ();
 sg13g2_fill_2 FILLER_56_519 ();
 sg13g2_fill_2 FILLER_56_526 ();
 sg13g2_fill_1 FILLER_56_528 ();
 sg13g2_decap_8 FILLER_56_533 ();
 sg13g2_fill_1 FILLER_56_540 ();
 sg13g2_fill_2 FILLER_56_556 ();
 sg13g2_decap_4 FILLER_56_575 ();
 sg13g2_fill_1 FILLER_56_583 ();
 sg13g2_decap_8 FILLER_56_593 ();
 sg13g2_fill_1 FILLER_56_600 ();
 sg13g2_fill_1 FILLER_56_608 ();
 sg13g2_fill_2 FILLER_56_626 ();
 sg13g2_fill_2 FILLER_56_640 ();
 sg13g2_decap_4 FILLER_56_656 ();
 sg13g2_fill_2 FILLER_56_660 ();
 sg13g2_decap_8 FILLER_56_666 ();
 sg13g2_decap_8 FILLER_56_673 ();
 sg13g2_decap_4 FILLER_56_680 ();
 sg13g2_fill_2 FILLER_56_684 ();
 sg13g2_fill_2 FILLER_56_696 ();
 sg13g2_fill_1 FILLER_56_698 ();
 sg13g2_fill_2 FILLER_56_712 ();
 sg13g2_decap_4 FILLER_56_720 ();
 sg13g2_fill_2 FILLER_56_724 ();
 sg13g2_decap_4 FILLER_56_734 ();
 sg13g2_fill_1 FILLER_56_738 ();
 sg13g2_decap_4 FILLER_56_748 ();
 sg13g2_decap_4 FILLER_56_758 ();
 sg13g2_fill_2 FILLER_56_762 ();
 sg13g2_decap_4 FILLER_56_803 ();
 sg13g2_fill_1 FILLER_56_807 ();
 sg13g2_fill_1 FILLER_56_821 ();
 sg13g2_fill_2 FILLER_56_827 ();
 sg13g2_decap_4 FILLER_56_834 ();
 sg13g2_fill_1 FILLER_56_838 ();
 sg13g2_fill_2 FILLER_56_869 ();
 sg13g2_fill_1 FILLER_56_871 ();
 sg13g2_decap_8 FILLER_56_891 ();
 sg13g2_decap_8 FILLER_56_898 ();
 sg13g2_fill_1 FILLER_56_905 ();
 sg13g2_decap_4 FILLER_56_911 ();
 sg13g2_decap_4 FILLER_56_931 ();
 sg13g2_decap_4 FILLER_56_950 ();
 sg13g2_fill_1 FILLER_56_954 ();
 sg13g2_decap_8 FILLER_56_964 ();
 sg13g2_fill_1 FILLER_56_971 ();
 sg13g2_decap_4 FILLER_56_981 ();
 sg13g2_fill_2 FILLER_56_985 ();
 sg13g2_decap_8 FILLER_56_1013 ();
 sg13g2_decap_4 FILLER_56_1020 ();
 sg13g2_decap_8 FILLER_56_1028 ();
 sg13g2_decap_8 FILLER_56_1056 ();
 sg13g2_fill_1 FILLER_56_1063 ();
 sg13g2_decap_8 FILLER_56_1081 ();
 sg13g2_fill_1 FILLER_56_1088 ();
 sg13g2_decap_4 FILLER_56_1115 ();
 sg13g2_fill_2 FILLER_56_1142 ();
 sg13g2_fill_1 FILLER_56_1149 ();
 sg13g2_decap_4 FILLER_56_1155 ();
 sg13g2_fill_1 FILLER_56_1167 ();
 sg13g2_decap_4 FILLER_56_1173 ();
 sg13g2_fill_1 FILLER_56_1177 ();
 sg13g2_decap_8 FILLER_56_1190 ();
 sg13g2_fill_1 FILLER_56_1208 ();
 sg13g2_decap_4 FILLER_56_1214 ();
 sg13g2_fill_1 FILLER_56_1245 ();
 sg13g2_fill_2 FILLER_56_1251 ();
 sg13g2_fill_1 FILLER_56_1258 ();
 sg13g2_decap_8 FILLER_56_1272 ();
 sg13g2_decap_8 FILLER_56_1279 ();
 sg13g2_decap_8 FILLER_56_1286 ();
 sg13g2_decap_8 FILLER_56_1293 ();
 sg13g2_fill_2 FILLER_56_1300 ();
 sg13g2_decap_8 FILLER_56_1314 ();
 sg13g2_decap_8 FILLER_56_1321 ();
 sg13g2_decap_4 FILLER_56_1328 ();
 sg13g2_decap_8 FILLER_56_1340 ();
 sg13g2_decap_8 FILLER_56_1347 ();
 sg13g2_fill_2 FILLER_56_1354 ();
 sg13g2_fill_1 FILLER_56_1356 ();
 sg13g2_decap_8 FILLER_56_1381 ();
 sg13g2_decap_8 FILLER_56_1392 ();
 sg13g2_fill_2 FILLER_56_1404 ();
 sg13g2_fill_1 FILLER_56_1406 ();
 sg13g2_fill_1 FILLER_56_1411 ();
 sg13g2_fill_2 FILLER_56_1423 ();
 sg13g2_decap_8 FILLER_56_1430 ();
 sg13g2_fill_1 FILLER_56_1437 ();
 sg13g2_fill_1 FILLER_56_1505 ();
 sg13g2_decap_4 FILLER_56_1536 ();
 sg13g2_fill_2 FILLER_56_1540 ();
 sg13g2_decap_8 FILLER_56_1562 ();
 sg13g2_decap_8 FILLER_56_1569 ();
 sg13g2_decap_8 FILLER_56_1576 ();
 sg13g2_fill_2 FILLER_56_1583 ();
 sg13g2_fill_1 FILLER_56_1585 ();
 sg13g2_decap_8 FILLER_56_1595 ();
 sg13g2_decap_8 FILLER_56_1602 ();
 sg13g2_decap_4 FILLER_56_1609 ();
 sg13g2_fill_2 FILLER_56_1613 ();
 sg13g2_fill_2 FILLER_56_1620 ();
 sg13g2_fill_2 FILLER_56_1630 ();
 sg13g2_fill_1 FILLER_56_1632 ();
 sg13g2_decap_8 FILLER_56_1637 ();
 sg13g2_fill_2 FILLER_56_1644 ();
 sg13g2_fill_1 FILLER_56_1646 ();
 sg13g2_fill_2 FILLER_56_1652 ();
 sg13g2_decap_4 FILLER_56_1659 ();
 sg13g2_decap_8 FILLER_56_1711 ();
 sg13g2_decap_8 FILLER_56_1718 ();
 sg13g2_fill_1 FILLER_56_1725 ();
 sg13g2_decap_8 FILLER_56_1730 ();
 sg13g2_decap_8 FILLER_56_1737 ();
 sg13g2_decap_8 FILLER_56_1744 ();
 sg13g2_decap_8 FILLER_56_1751 ();
 sg13g2_decap_8 FILLER_56_1758 ();
 sg13g2_decap_8 FILLER_56_1765 ();
 sg13g2_fill_2 FILLER_56_1772 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_19 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_4 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_50 ();
 sg13g2_fill_1 FILLER_57_63 ();
 sg13g2_decap_4 FILLER_57_87 ();
 sg13g2_decap_4 FILLER_57_98 ();
 sg13g2_fill_2 FILLER_57_102 ();
 sg13g2_decap_8 FILLER_57_146 ();
 sg13g2_fill_1 FILLER_57_153 ();
 sg13g2_fill_2 FILLER_57_169 ();
 sg13g2_fill_1 FILLER_57_171 ();
 sg13g2_decap_8 FILLER_57_190 ();
 sg13g2_fill_2 FILLER_57_207 ();
 sg13g2_fill_2 FILLER_57_213 ();
 sg13g2_fill_1 FILLER_57_215 ();
 sg13g2_fill_2 FILLER_57_222 ();
 sg13g2_fill_1 FILLER_57_253 ();
 sg13g2_decap_4 FILLER_57_262 ();
 sg13g2_fill_1 FILLER_57_266 ();
 sg13g2_decap_8 FILLER_57_277 ();
 sg13g2_fill_1 FILLER_57_284 ();
 sg13g2_fill_2 FILLER_57_312 ();
 sg13g2_fill_1 FILLER_57_314 ();
 sg13g2_decap_8 FILLER_57_320 ();
 sg13g2_decap_4 FILLER_57_327 ();
 sg13g2_fill_2 FILLER_57_331 ();
 sg13g2_decap_8 FILLER_57_343 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_decap_4 FILLER_57_355 ();
 sg13g2_decap_8 FILLER_57_368 ();
 sg13g2_decap_4 FILLER_57_375 ();
 sg13g2_fill_1 FILLER_57_379 ();
 sg13g2_decap_4 FILLER_57_386 ();
 sg13g2_decap_8 FILLER_57_397 ();
 sg13g2_fill_2 FILLER_57_424 ();
 sg13g2_fill_1 FILLER_57_426 ();
 sg13g2_fill_2 FILLER_57_431 ();
 sg13g2_decap_8 FILLER_57_437 ();
 sg13g2_decap_4 FILLER_57_444 ();
 sg13g2_fill_2 FILLER_57_448 ();
 sg13g2_fill_2 FILLER_57_458 ();
 sg13g2_fill_2 FILLER_57_465 ();
 sg13g2_fill_2 FILLER_57_471 ();
 sg13g2_fill_2 FILLER_57_490 ();
 sg13g2_fill_1 FILLER_57_504 ();
 sg13g2_fill_2 FILLER_57_514 ();
 sg13g2_fill_1 FILLER_57_516 ();
 sg13g2_decap_8 FILLER_57_536 ();
 sg13g2_fill_1 FILLER_57_560 ();
 sg13g2_decap_8 FILLER_57_571 ();
 sg13g2_fill_2 FILLER_57_578 ();
 sg13g2_fill_1 FILLER_57_580 ();
 sg13g2_fill_2 FILLER_57_596 ();
 sg13g2_fill_1 FILLER_57_613 ();
 sg13g2_fill_1 FILLER_57_618 ();
 sg13g2_decap_8 FILLER_57_651 ();
 sg13g2_fill_2 FILLER_57_658 ();
 sg13g2_decap_8 FILLER_57_665 ();
 sg13g2_decap_8 FILLER_57_676 ();
 sg13g2_fill_2 FILLER_57_686 ();
 sg13g2_fill_2 FILLER_57_728 ();
 sg13g2_decap_8 FILLER_57_765 ();
 sg13g2_decap_8 FILLER_57_772 ();
 sg13g2_decap_8 FILLER_57_779 ();
 sg13g2_fill_1 FILLER_57_786 ();
 sg13g2_decap_4 FILLER_57_820 ();
 sg13g2_fill_1 FILLER_57_824 ();
 sg13g2_fill_1 FILLER_57_830 ();
 sg13g2_decap_4 FILLER_57_835 ();
 sg13g2_fill_2 FILLER_57_847 ();
 sg13g2_fill_1 FILLER_57_849 ();
 sg13g2_decap_4 FILLER_57_854 ();
 sg13g2_fill_2 FILLER_57_858 ();
 sg13g2_fill_1 FILLER_57_864 ();
 sg13g2_decap_4 FILLER_57_870 ();
 sg13g2_decap_4 FILLER_57_878 ();
 sg13g2_fill_1 FILLER_57_882 ();
 sg13g2_decap_4 FILLER_57_891 ();
 sg13g2_fill_1 FILLER_57_895 ();
 sg13g2_decap_4 FILLER_57_901 ();
 sg13g2_fill_1 FILLER_57_905 ();
 sg13g2_fill_2 FILLER_57_913 ();
 sg13g2_fill_1 FILLER_57_915 ();
 sg13g2_fill_1 FILLER_57_921 ();
 sg13g2_fill_2 FILLER_57_926 ();
 sg13g2_fill_1 FILLER_57_933 ();
 sg13g2_decap_4 FILLER_57_952 ();
 sg13g2_fill_1 FILLER_57_961 ();
 sg13g2_decap_4 FILLER_57_967 ();
 sg13g2_fill_1 FILLER_57_971 ();
 sg13g2_decap_8 FILLER_57_977 ();
 sg13g2_fill_2 FILLER_57_984 ();
 sg13g2_fill_1 FILLER_57_986 ();
 sg13g2_decap_4 FILLER_57_991 ();
 sg13g2_decap_8 FILLER_57_1000 ();
 sg13g2_decap_4 FILLER_57_1027 ();
 sg13g2_decap_8 FILLER_57_1035 ();
 sg13g2_decap_4 FILLER_57_1042 ();
 sg13g2_decap_8 FILLER_57_1051 ();
 sg13g2_decap_4 FILLER_57_1058 ();
 sg13g2_fill_1 FILLER_57_1062 ();
 sg13g2_decap_8 FILLER_57_1067 ();
 sg13g2_fill_1 FILLER_57_1074 ();
 sg13g2_decap_8 FILLER_57_1080 ();
 sg13g2_decap_4 FILLER_57_1087 ();
 sg13g2_fill_2 FILLER_57_1094 ();
 sg13g2_fill_1 FILLER_57_1096 ();
 sg13g2_decap_8 FILLER_57_1117 ();
 sg13g2_fill_2 FILLER_57_1124 ();
 sg13g2_decap_4 FILLER_57_1132 ();
 sg13g2_fill_1 FILLER_57_1144 ();
 sg13g2_fill_1 FILLER_57_1152 ();
 sg13g2_fill_1 FILLER_57_1166 ();
 sg13g2_fill_1 FILLER_57_1171 ();
 sg13g2_fill_2 FILLER_57_1193 ();
 sg13g2_fill_2 FILLER_57_1202 ();
 sg13g2_fill_1 FILLER_57_1215 ();
 sg13g2_decap_4 FILLER_57_1243 ();
 sg13g2_fill_2 FILLER_57_1247 ();
 sg13g2_fill_2 FILLER_57_1262 ();
 sg13g2_decap_8 FILLER_57_1268 ();
 sg13g2_decap_8 FILLER_57_1281 ();
 sg13g2_decap_8 FILLER_57_1288 ();
 sg13g2_decap_8 FILLER_57_1295 ();
 sg13g2_decap_4 FILLER_57_1302 ();
 sg13g2_fill_1 FILLER_57_1306 ();
 sg13g2_decap_8 FILLER_57_1311 ();
 sg13g2_decap_8 FILLER_57_1318 ();
 sg13g2_fill_1 FILLER_57_1325 ();
 sg13g2_fill_1 FILLER_57_1356 ();
 sg13g2_decap_4 FILLER_57_1361 ();
 sg13g2_fill_1 FILLER_57_1365 ();
 sg13g2_fill_2 FILLER_57_1392 ();
 sg13g2_fill_1 FILLER_57_1394 ();
 sg13g2_fill_1 FILLER_57_1423 ();
 sg13g2_decap_8 FILLER_57_1432 ();
 sg13g2_decap_4 FILLER_57_1439 ();
 sg13g2_fill_1 FILLER_57_1443 ();
 sg13g2_fill_2 FILLER_57_1448 ();
 sg13g2_fill_1 FILLER_57_1450 ();
 sg13g2_decap_8 FILLER_57_1467 ();
 sg13g2_decap_4 FILLER_57_1474 ();
 sg13g2_decap_4 FILLER_57_1482 ();
 sg13g2_decap_8 FILLER_57_1490 ();
 sg13g2_decap_8 FILLER_57_1497 ();
 sg13g2_decap_8 FILLER_57_1504 ();
 sg13g2_decap_4 FILLER_57_1511 ();
 sg13g2_fill_2 FILLER_57_1515 ();
 sg13g2_decap_8 FILLER_57_1521 ();
 sg13g2_decap_8 FILLER_57_1528 ();
 sg13g2_decap_8 FILLER_57_1535 ();
 sg13g2_decap_4 FILLER_57_1542 ();
 sg13g2_decap_8 FILLER_57_1561 ();
 sg13g2_fill_1 FILLER_57_1573 ();
 sg13g2_fill_1 FILLER_57_1590 ();
 sg13g2_fill_1 FILLER_57_1621 ();
 sg13g2_decap_8 FILLER_57_1627 ();
 sg13g2_fill_2 FILLER_57_1634 ();
 sg13g2_fill_1 FILLER_57_1636 ();
 sg13g2_fill_2 FILLER_57_1658 ();
 sg13g2_fill_2 FILLER_57_1701 ();
 sg13g2_decap_8 FILLER_57_1707 ();
 sg13g2_decap_8 FILLER_57_1714 ();
 sg13g2_decap_8 FILLER_57_1721 ();
 sg13g2_decap_8 FILLER_57_1728 ();
 sg13g2_decap_8 FILLER_57_1735 ();
 sg13g2_decap_8 FILLER_57_1742 ();
 sg13g2_decap_8 FILLER_57_1749 ();
 sg13g2_decap_8 FILLER_57_1756 ();
 sg13g2_decap_8 FILLER_57_1763 ();
 sg13g2_decap_4 FILLER_57_1770 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_2 ();
 sg13g2_fill_2 FILLER_58_8 ();
 sg13g2_decap_4 FILLER_58_14 ();
 sg13g2_fill_2 FILLER_58_37 ();
 sg13g2_fill_1 FILLER_58_39 ();
 sg13g2_fill_2 FILLER_58_44 ();
 sg13g2_fill_1 FILLER_58_46 ();
 sg13g2_decap_4 FILLER_58_71 ();
 sg13g2_fill_1 FILLER_58_75 ();
 sg13g2_decap_8 FILLER_58_85 ();
 sg13g2_decap_4 FILLER_58_92 ();
 sg13g2_fill_2 FILLER_58_96 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_4 FILLER_58_126 ();
 sg13g2_fill_2 FILLER_58_130 ();
 sg13g2_fill_1 FILLER_58_146 ();
 sg13g2_decap_4 FILLER_58_157 ();
 sg13g2_decap_4 FILLER_58_186 ();
 sg13g2_fill_2 FILLER_58_190 ();
 sg13g2_fill_1 FILLER_58_196 ();
 sg13g2_fill_2 FILLER_58_217 ();
 sg13g2_decap_4 FILLER_58_224 ();
 sg13g2_decap_4 FILLER_58_233 ();
 sg13g2_decap_8 FILLER_58_246 ();
 sg13g2_decap_8 FILLER_58_261 ();
 sg13g2_decap_8 FILLER_58_268 ();
 sg13g2_decap_4 FILLER_58_275 ();
 sg13g2_fill_1 FILLER_58_279 ();
 sg13g2_decap_8 FILLER_58_285 ();
 sg13g2_decap_4 FILLER_58_292 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_323 ();
 sg13g2_fill_1 FILLER_58_325 ();
 sg13g2_decap_8 FILLER_58_339 ();
 sg13g2_decap_4 FILLER_58_346 ();
 sg13g2_fill_2 FILLER_58_350 ();
 sg13g2_decap_4 FILLER_58_357 ();
 sg13g2_fill_2 FILLER_58_361 ();
 sg13g2_fill_2 FILLER_58_371 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_1 FILLER_58_379 ();
 sg13g2_decap_4 FILLER_58_387 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_2 FILLER_58_414 ();
 sg13g2_fill_1 FILLER_58_416 ();
 sg13g2_fill_1 FILLER_58_432 ();
 sg13g2_fill_2 FILLER_58_438 ();
 sg13g2_fill_2 FILLER_58_448 ();
 sg13g2_fill_2 FILLER_58_457 ();
 sg13g2_fill_2 FILLER_58_464 ();
 sg13g2_fill_1 FILLER_58_483 ();
 sg13g2_fill_2 FILLER_58_489 ();
 sg13g2_fill_2 FILLER_58_504 ();
 sg13g2_decap_4 FILLER_58_515 ();
 sg13g2_fill_2 FILLER_58_519 ();
 sg13g2_fill_1 FILLER_58_526 ();
 sg13g2_fill_1 FILLER_58_532 ();
 sg13g2_fill_1 FILLER_58_541 ();
 sg13g2_fill_2 FILLER_58_548 ();
 sg13g2_decap_4 FILLER_58_554 ();
 sg13g2_decap_8 FILLER_58_562 ();
 sg13g2_decap_8 FILLER_58_569 ();
 sg13g2_decap_4 FILLER_58_576 ();
 sg13g2_fill_1 FILLER_58_585 ();
 sg13g2_fill_1 FILLER_58_591 ();
 sg13g2_decap_4 FILLER_58_642 ();
 sg13g2_decap_4 FILLER_58_651 ();
 sg13g2_fill_2 FILLER_58_655 ();
 sg13g2_fill_2 FILLER_58_668 ();
 sg13g2_fill_2 FILLER_58_686 ();
 sg13g2_fill_2 FILLER_58_692 ();
 sg13g2_fill_2 FILLER_58_699 ();
 sg13g2_fill_1 FILLER_58_706 ();
 sg13g2_decap_8 FILLER_58_728 ();
 sg13g2_fill_2 FILLER_58_735 ();
 sg13g2_fill_1 FILLER_58_737 ();
 sg13g2_decap_4 FILLER_58_743 ();
 sg13g2_fill_2 FILLER_58_747 ();
 sg13g2_fill_2 FILLER_58_755 ();
 sg13g2_decap_8 FILLER_58_761 ();
 sg13g2_fill_2 FILLER_58_768 ();
 sg13g2_fill_1 FILLER_58_779 ();
 sg13g2_fill_2 FILLER_58_798 ();
 sg13g2_fill_2 FILLER_58_824 ();
 sg13g2_fill_1 FILLER_58_826 ();
 sg13g2_decap_8 FILLER_58_865 ();
 sg13g2_fill_1 FILLER_58_880 ();
 sg13g2_fill_1 FILLER_58_885 ();
 sg13g2_decap_4 FILLER_58_895 ();
 sg13g2_decap_4 FILLER_58_904 ();
 sg13g2_fill_2 FILLER_58_908 ();
 sg13g2_decap_4 FILLER_58_929 ();
 sg13g2_decap_4 FILLER_58_942 ();
 sg13g2_fill_2 FILLER_58_946 ();
 sg13g2_decap_8 FILLER_58_952 ();
 sg13g2_fill_1 FILLER_58_964 ();
 sg13g2_decap_8 FILLER_58_979 ();
 sg13g2_fill_2 FILLER_58_986 ();
 sg13g2_fill_2 FILLER_58_991 ();
 sg13g2_fill_1 FILLER_58_993 ();
 sg13g2_fill_2 FILLER_58_1002 ();
 sg13g2_fill_1 FILLER_58_1033 ();
 sg13g2_fill_2 FILLER_58_1041 ();
 sg13g2_fill_2 FILLER_58_1063 ();
 sg13g2_fill_1 FILLER_58_1065 ();
 sg13g2_fill_2 FILLER_58_1089 ();
 sg13g2_fill_1 FILLER_58_1091 ();
 sg13g2_fill_1 FILLER_58_1097 ();
 sg13g2_decap_8 FILLER_58_1102 ();
 sg13g2_decap_4 FILLER_58_1109 ();
 sg13g2_decap_8 FILLER_58_1118 ();
 sg13g2_fill_2 FILLER_58_1125 ();
 sg13g2_fill_1 FILLER_58_1131 ();
 sg13g2_decap_4 FILLER_58_1135 ();
 sg13g2_decap_4 FILLER_58_1160 ();
 sg13g2_fill_1 FILLER_58_1164 ();
 sg13g2_fill_2 FILLER_58_1181 ();
 sg13g2_fill_1 FILLER_58_1183 ();
 sg13g2_decap_4 FILLER_58_1188 ();
 sg13g2_fill_2 FILLER_58_1192 ();
 sg13g2_fill_1 FILLER_58_1199 ();
 sg13g2_fill_1 FILLER_58_1204 ();
 sg13g2_fill_1 FILLER_58_1210 ();
 sg13g2_fill_1 FILLER_58_1216 ();
 sg13g2_decap_4 FILLER_58_1232 ();
 sg13g2_fill_2 FILLER_58_1236 ();
 sg13g2_fill_2 FILLER_58_1254 ();
 sg13g2_fill_2 FILLER_58_1270 ();
 sg13g2_fill_1 FILLER_58_1332 ();
 sg13g2_fill_1 FILLER_58_1337 ();
 sg13g2_fill_1 FILLER_58_1364 ();
 sg13g2_fill_2 FILLER_58_1369 ();
 sg13g2_decap_8 FILLER_58_1375 ();
 sg13g2_decap_4 FILLER_58_1382 ();
 sg13g2_fill_2 FILLER_58_1386 ();
 sg13g2_decap_8 FILLER_58_1392 ();
 sg13g2_decap_8 FILLER_58_1399 ();
 sg13g2_fill_2 FILLER_58_1413 ();
 sg13g2_fill_1 FILLER_58_1415 ();
 sg13g2_fill_1 FILLER_58_1427 ();
 sg13g2_decap_8 FILLER_58_1440 ();
 sg13g2_fill_2 FILLER_58_1447 ();
 sg13g2_fill_1 FILLER_58_1449 ();
 sg13g2_decap_8 FILLER_58_1467 ();
 sg13g2_fill_2 FILLER_58_1474 ();
 sg13g2_fill_1 FILLER_58_1476 ();
 sg13g2_decap_8 FILLER_58_1485 ();
 sg13g2_decap_4 FILLER_58_1492 ();
 sg13g2_decap_8 FILLER_58_1500 ();
 sg13g2_decap_4 FILLER_58_1511 ();
 sg13g2_fill_2 FILLER_58_1515 ();
 sg13g2_fill_2 FILLER_58_1533 ();
 sg13g2_fill_2 FILLER_58_1539 ();
 sg13g2_fill_2 FILLER_58_1547 ();
 sg13g2_fill_1 FILLER_58_1549 ();
 sg13g2_fill_2 FILLER_58_1556 ();
 sg13g2_fill_1 FILLER_58_1558 ();
 sg13g2_fill_2 FILLER_58_1567 ();
 sg13g2_fill_1 FILLER_58_1569 ();
 sg13g2_decap_8 FILLER_58_1578 ();
 sg13g2_fill_2 FILLER_58_1585 ();
 sg13g2_decap_8 FILLER_58_1591 ();
 sg13g2_decap_8 FILLER_58_1602 ();
 sg13g2_decap_8 FILLER_58_1609 ();
 sg13g2_decap_4 FILLER_58_1652 ();
 sg13g2_decap_4 FILLER_58_1660 ();
 sg13g2_fill_1 FILLER_58_1664 ();
 sg13g2_fill_1 FILLER_58_1669 ();
 sg13g2_decap_4 FILLER_58_1675 ();
 sg13g2_fill_1 FILLER_58_1679 ();
 sg13g2_decap_8 FILLER_58_1684 ();
 sg13g2_decap_8 FILLER_58_1691 ();
 sg13g2_decap_8 FILLER_58_1698 ();
 sg13g2_decap_8 FILLER_58_1705 ();
 sg13g2_decap_8 FILLER_58_1712 ();
 sg13g2_decap_8 FILLER_58_1719 ();
 sg13g2_decap_8 FILLER_58_1726 ();
 sg13g2_decap_8 FILLER_58_1733 ();
 sg13g2_decap_8 FILLER_58_1740 ();
 sg13g2_decap_8 FILLER_58_1747 ();
 sg13g2_decap_8 FILLER_58_1754 ();
 sg13g2_decap_8 FILLER_58_1761 ();
 sg13g2_decap_4 FILLER_58_1768 ();
 sg13g2_fill_2 FILLER_58_1772 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_11 ();
 sg13g2_fill_2 FILLER_59_25 ();
 sg13g2_fill_1 FILLER_59_27 ();
 sg13g2_fill_2 FILLER_59_33 ();
 sg13g2_fill_2 FILLER_59_43 ();
 sg13g2_fill_1 FILLER_59_45 ();
 sg13g2_decap_4 FILLER_59_51 ();
 sg13g2_fill_2 FILLER_59_55 ();
 sg13g2_fill_2 FILLER_59_63 ();
 sg13g2_fill_2 FILLER_59_71 ();
 sg13g2_decap_8 FILLER_59_78 ();
 sg13g2_decap_4 FILLER_59_85 ();
 sg13g2_fill_2 FILLER_59_89 ();
 sg13g2_fill_2 FILLER_59_99 ();
 sg13g2_fill_1 FILLER_59_101 ();
 sg13g2_fill_2 FILLER_59_107 ();
 sg13g2_fill_1 FILLER_59_109 ();
 sg13g2_decap_8 FILLER_59_115 ();
 sg13g2_fill_2 FILLER_59_131 ();
 sg13g2_decap_8 FILLER_59_160 ();
 sg13g2_decap_8 FILLER_59_167 ();
 sg13g2_decap_8 FILLER_59_174 ();
 sg13g2_fill_2 FILLER_59_185 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_fill_2 FILLER_59_216 ();
 sg13g2_decap_4 FILLER_59_250 ();
 sg13g2_fill_1 FILLER_59_254 ();
 sg13g2_decap_4 FILLER_59_261 ();
 sg13g2_decap_8 FILLER_59_270 ();
 sg13g2_fill_2 FILLER_59_277 ();
 sg13g2_fill_1 FILLER_59_279 ();
 sg13g2_decap_8 FILLER_59_288 ();
 sg13g2_decap_4 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_299 ();
 sg13g2_fill_1 FILLER_59_316 ();
 sg13g2_decap_4 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_337 ();
 sg13g2_decap_4 FILLER_59_344 ();
 sg13g2_fill_2 FILLER_59_348 ();
 sg13g2_decap_8 FILLER_59_359 ();
 sg13g2_decap_8 FILLER_59_366 ();
 sg13g2_fill_2 FILLER_59_373 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_fill_2 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_439 ();
 sg13g2_decap_8 FILLER_59_446 ();
 sg13g2_decap_8 FILLER_59_453 ();
 sg13g2_decap_8 FILLER_59_460 ();
 sg13g2_decap_8 FILLER_59_467 ();
 sg13g2_fill_2 FILLER_59_489 ();
 sg13g2_fill_1 FILLER_59_491 ();
 sg13g2_fill_2 FILLER_59_508 ();
 sg13g2_fill_1 FILLER_59_510 ();
 sg13g2_decap_4 FILLER_59_542 ();
 sg13g2_fill_2 FILLER_59_546 ();
 sg13g2_decap_8 FILLER_59_560 ();
 sg13g2_decap_8 FILLER_59_567 ();
 sg13g2_decap_4 FILLER_59_574 ();
 sg13g2_fill_2 FILLER_59_578 ();
 sg13g2_fill_2 FILLER_59_598 ();
 sg13g2_fill_2 FILLER_59_617 ();
 sg13g2_decap_8 FILLER_59_629 ();
 sg13g2_fill_2 FILLER_59_636 ();
 sg13g2_fill_1 FILLER_59_638 ();
 sg13g2_decap_8 FILLER_59_644 ();
 sg13g2_decap_8 FILLER_59_651 ();
 sg13g2_fill_1 FILLER_59_658 ();
 sg13g2_fill_1 FILLER_59_737 ();
 sg13g2_fill_1 FILLER_59_743 ();
 sg13g2_fill_2 FILLER_59_779 ();
 sg13g2_fill_1 FILLER_59_781 ();
 sg13g2_decap_8 FILLER_59_787 ();
 sg13g2_decap_4 FILLER_59_794 ();
 sg13g2_decap_8 FILLER_59_805 ();
 sg13g2_decap_4 FILLER_59_812 ();
 sg13g2_fill_2 FILLER_59_816 ();
 sg13g2_decap_8 FILLER_59_823 ();
 sg13g2_decap_4 FILLER_59_834 ();
 sg13g2_decap_8 FILLER_59_849 ();
 sg13g2_decap_8 FILLER_59_856 ();
 sg13g2_fill_2 FILLER_59_863 ();
 sg13g2_fill_1 FILLER_59_865 ();
 sg13g2_decap_8 FILLER_59_886 ();
 sg13g2_decap_8 FILLER_59_893 ();
 sg13g2_decap_8 FILLER_59_900 ();
 sg13g2_decap_8 FILLER_59_907 ();
 sg13g2_fill_2 FILLER_59_914 ();
 sg13g2_decap_4 FILLER_59_930 ();
 sg13g2_fill_2 FILLER_59_934 ();
 sg13g2_fill_1 FILLER_59_941 ();
 sg13g2_fill_2 FILLER_59_947 ();
 sg13g2_fill_1 FILLER_59_949 ();
 sg13g2_decap_8 FILLER_59_954 ();
 sg13g2_fill_2 FILLER_59_970 ();
 sg13g2_decap_4 FILLER_59_981 ();
 sg13g2_fill_1 FILLER_59_985 ();
 sg13g2_decap_8 FILLER_59_989 ();
 sg13g2_fill_1 FILLER_59_996 ();
 sg13g2_fill_2 FILLER_59_1002 ();
 sg13g2_fill_1 FILLER_59_1004 ();
 sg13g2_fill_1 FILLER_59_1030 ();
 sg13g2_fill_2 FILLER_59_1054 ();
 sg13g2_decap_8 FILLER_59_1060 ();
 sg13g2_fill_1 FILLER_59_1067 ();
 sg13g2_decap_4 FILLER_59_1072 ();
 sg13g2_fill_1 FILLER_59_1088 ();
 sg13g2_fill_2 FILLER_59_1093 ();
 sg13g2_fill_1 FILLER_59_1095 ();
 sg13g2_fill_1 FILLER_59_1113 ();
 sg13g2_fill_1 FILLER_59_1118 ();
 sg13g2_fill_1 FILLER_59_1127 ();
 sg13g2_fill_1 FILLER_59_1134 ();
 sg13g2_fill_1 FILLER_59_1146 ();
 sg13g2_decap_8 FILLER_59_1163 ();
 sg13g2_decap_4 FILLER_59_1170 ();
 sg13g2_fill_1 FILLER_59_1174 ();
 sg13g2_fill_1 FILLER_59_1184 ();
 sg13g2_decap_8 FILLER_59_1194 ();
 sg13g2_decap_4 FILLER_59_1201 ();
 sg13g2_fill_1 FILLER_59_1205 ();
 sg13g2_fill_2 FILLER_59_1224 ();
 sg13g2_decap_4 FILLER_59_1234 ();
 sg13g2_fill_2 FILLER_59_1248 ();
 sg13g2_decap_4 FILLER_59_1256 ();
 sg13g2_decap_8 FILLER_59_1266 ();
 sg13g2_fill_1 FILLER_59_1273 ();
 sg13g2_fill_2 FILLER_59_1279 ();
 sg13g2_fill_1 FILLER_59_1281 ();
 sg13g2_decap_8 FILLER_59_1290 ();
 sg13g2_decap_4 FILLER_59_1297 ();
 sg13g2_fill_2 FILLER_59_1301 ();
 sg13g2_decap_8 FILLER_59_1312 ();
 sg13g2_decap_8 FILLER_59_1319 ();
 sg13g2_fill_2 FILLER_59_1326 ();
 sg13g2_fill_1 FILLER_59_1328 ();
 sg13g2_fill_2 FILLER_59_1365 ();
 sg13g2_decap_8 FILLER_59_1373 ();
 sg13g2_decap_8 FILLER_59_1380 ();
 sg13g2_decap_8 FILLER_59_1387 ();
 sg13g2_decap_8 FILLER_59_1394 ();
 sg13g2_decap_4 FILLER_59_1401 ();
 sg13g2_fill_2 FILLER_59_1413 ();
 sg13g2_fill_1 FILLER_59_1415 ();
 sg13g2_fill_2 FILLER_59_1431 ();
 sg13g2_decap_8 FILLER_59_1441 ();
 sg13g2_decap_4 FILLER_59_1478 ();
 sg13g2_fill_2 FILLER_59_1486 ();
 sg13g2_decap_4 FILLER_59_1514 ();
 sg13g2_decap_8 FILLER_59_1558 ();
 sg13g2_decap_8 FILLER_59_1565 ();
 sg13g2_fill_2 FILLER_59_1572 ();
 sg13g2_fill_2 FILLER_59_1578 ();
 sg13g2_decap_8 FILLER_59_1610 ();
 sg13g2_decap_8 FILLER_59_1617 ();
 sg13g2_decap_8 FILLER_59_1684 ();
 sg13g2_decap_8 FILLER_59_1691 ();
 sg13g2_decap_8 FILLER_59_1698 ();
 sg13g2_decap_8 FILLER_59_1705 ();
 sg13g2_decap_8 FILLER_59_1712 ();
 sg13g2_decap_8 FILLER_59_1719 ();
 sg13g2_decap_8 FILLER_59_1726 ();
 sg13g2_decap_8 FILLER_59_1733 ();
 sg13g2_decap_8 FILLER_59_1740 ();
 sg13g2_decap_8 FILLER_59_1747 ();
 sg13g2_decap_8 FILLER_59_1754 ();
 sg13g2_decap_8 FILLER_59_1761 ();
 sg13g2_decap_4 FILLER_59_1768 ();
 sg13g2_fill_2 FILLER_59_1772 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_15 ();
 sg13g2_fill_2 FILLER_60_19 ();
 sg13g2_fill_2 FILLER_60_27 ();
 sg13g2_decap_8 FILLER_60_34 ();
 sg13g2_fill_1 FILLER_60_41 ();
 sg13g2_decap_8 FILLER_60_61 ();
 sg13g2_decap_8 FILLER_60_68 ();
 sg13g2_decap_4 FILLER_60_75 ();
 sg13g2_fill_1 FILLER_60_79 ();
 sg13g2_decap_8 FILLER_60_83 ();
 sg13g2_fill_2 FILLER_60_90 ();
 sg13g2_fill_1 FILLER_60_110 ();
 sg13g2_decap_8 FILLER_60_117 ();
 sg13g2_decap_8 FILLER_60_124 ();
 sg13g2_decap_4 FILLER_60_135 ();
 sg13g2_fill_2 FILLER_60_139 ();
 sg13g2_fill_1 FILLER_60_145 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_4 FILLER_60_168 ();
 sg13g2_fill_2 FILLER_60_172 ();
 sg13g2_decap_8 FILLER_60_186 ();
 sg13g2_decap_8 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_200 ();
 sg13g2_decap_4 FILLER_60_207 ();
 sg13g2_decap_4 FILLER_60_223 ();
 sg13g2_decap_4 FILLER_60_232 ();
 sg13g2_fill_1 FILLER_60_236 ();
 sg13g2_fill_1 FILLER_60_258 ();
 sg13g2_decap_8 FILLER_60_266 ();
 sg13g2_fill_1 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_286 ();
 sg13g2_decap_4 FILLER_60_293 ();
 sg13g2_fill_1 FILLER_60_297 ();
 sg13g2_decap_4 FILLER_60_314 ();
 sg13g2_fill_2 FILLER_60_318 ();
 sg13g2_decap_8 FILLER_60_323 ();
 sg13g2_fill_2 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_332 ();
 sg13g2_fill_1 FILLER_60_348 ();
 sg13g2_decap_4 FILLER_60_355 ();
 sg13g2_fill_1 FILLER_60_359 ();
 sg13g2_decap_4 FILLER_60_365 ();
 sg13g2_decap_8 FILLER_60_376 ();
 sg13g2_fill_2 FILLER_60_396 ();
 sg13g2_decap_8 FILLER_60_429 ();
 sg13g2_fill_2 FILLER_60_436 ();
 sg13g2_fill_1 FILLER_60_443 ();
 sg13g2_decap_8 FILLER_60_453 ();
 sg13g2_decap_4 FILLER_60_460 ();
 sg13g2_fill_2 FILLER_60_469 ();
 sg13g2_fill_1 FILLER_60_476 ();
 sg13g2_decap_8 FILLER_60_481 ();
 sg13g2_decap_4 FILLER_60_501 ();
 sg13g2_decap_4 FILLER_60_514 ();
 sg13g2_fill_1 FILLER_60_518 ();
 sg13g2_fill_1 FILLER_60_536 ();
 sg13g2_fill_1 FILLER_60_543 ();
 sg13g2_decap_8 FILLER_60_553 ();
 sg13g2_decap_8 FILLER_60_560 ();
 sg13g2_decap_4 FILLER_60_567 ();
 sg13g2_decap_8 FILLER_60_575 ();
 sg13g2_decap_8 FILLER_60_582 ();
 sg13g2_fill_1 FILLER_60_589 ();
 sg13g2_fill_1 FILLER_60_621 ();
 sg13g2_decap_4 FILLER_60_634 ();
 sg13g2_decap_8 FILLER_60_642 ();
 sg13g2_decap_4 FILLER_60_649 ();
 sg13g2_fill_2 FILLER_60_653 ();
 sg13g2_decap_8 FILLER_60_658 ();
 sg13g2_decap_4 FILLER_60_665 ();
 sg13g2_fill_2 FILLER_60_669 ();
 sg13g2_decap_8 FILLER_60_675 ();
 sg13g2_decap_8 FILLER_60_682 ();
 sg13g2_decap_4 FILLER_60_689 ();
 sg13g2_fill_1 FILLER_60_693 ();
 sg13g2_fill_1 FILLER_60_698 ();
 sg13g2_fill_1 FILLER_60_711 ();
 sg13g2_decap_4 FILLER_60_721 ();
 sg13g2_fill_2 FILLER_60_725 ();
 sg13g2_decap_8 FILLER_60_732 ();
 sg13g2_fill_1 FILLER_60_739 ();
 sg13g2_fill_2 FILLER_60_744 ();
 sg13g2_fill_1 FILLER_60_746 ();
 sg13g2_decap_4 FILLER_60_755 ();
 sg13g2_decap_4 FILLER_60_764 ();
 sg13g2_decap_4 FILLER_60_772 ();
 sg13g2_decap_4 FILLER_60_784 ();
 sg13g2_fill_2 FILLER_60_788 ();
 sg13g2_fill_1 FILLER_60_797 ();
 sg13g2_fill_1 FILLER_60_824 ();
 sg13g2_fill_1 FILLER_60_829 ();
 sg13g2_decap_4 FILLER_60_834 ();
 sg13g2_fill_1 FILLER_60_838 ();
 sg13g2_fill_2 FILLER_60_865 ();
 sg13g2_decap_8 FILLER_60_874 ();
 sg13g2_decap_8 FILLER_60_881 ();
 sg13g2_fill_2 FILLER_60_888 ();
 sg13g2_decap_8 FILLER_60_905 ();
 sg13g2_decap_8 FILLER_60_912 ();
 sg13g2_decap_8 FILLER_60_919 ();
 sg13g2_decap_8 FILLER_60_926 ();
 sg13g2_decap_8 FILLER_60_933 ();
 sg13g2_decap_4 FILLER_60_940 ();
 sg13g2_fill_1 FILLER_60_944 ();
 sg13g2_decap_4 FILLER_60_954 ();
 sg13g2_decap_8 FILLER_60_962 ();
 sg13g2_fill_2 FILLER_60_969 ();
 sg13g2_decap_8 FILLER_60_989 ();
 sg13g2_fill_2 FILLER_60_1014 ();
 sg13g2_fill_1 FILLER_60_1016 ();
 sg13g2_fill_2 FILLER_60_1038 ();
 sg13g2_fill_2 FILLER_60_1046 ();
 sg13g2_decap_8 FILLER_60_1053 ();
 sg13g2_decap_8 FILLER_60_1060 ();
 sg13g2_decap_4 FILLER_60_1067 ();
 sg13g2_fill_2 FILLER_60_1071 ();
 sg13g2_fill_1 FILLER_60_1077 ();
 sg13g2_fill_1 FILLER_60_1082 ();
 sg13g2_fill_2 FILLER_60_1094 ();
 sg13g2_decap_4 FILLER_60_1114 ();
 sg13g2_fill_1 FILLER_60_1118 ();
 sg13g2_fill_2 FILLER_60_1147 ();
 sg13g2_decap_8 FILLER_60_1162 ();
 sg13g2_decap_4 FILLER_60_1169 ();
 sg13g2_fill_2 FILLER_60_1173 ();
 sg13g2_decap_8 FILLER_60_1191 ();
 sg13g2_decap_8 FILLER_60_1198 ();
 sg13g2_decap_4 FILLER_60_1205 ();
 sg13g2_fill_1 FILLER_60_1209 ();
 sg13g2_fill_2 FILLER_60_1223 ();
 sg13g2_fill_1 FILLER_60_1225 ();
 sg13g2_fill_2 FILLER_60_1234 ();
 sg13g2_decap_8 FILLER_60_1246 ();
 sg13g2_decap_4 FILLER_60_1253 ();
 sg13g2_decap_8 FILLER_60_1261 ();
 sg13g2_decap_8 FILLER_60_1272 ();
 sg13g2_fill_2 FILLER_60_1279 ();
 sg13g2_decap_4 FILLER_60_1290 ();
 sg13g2_decap_8 FILLER_60_1320 ();
 sg13g2_fill_2 FILLER_60_1327 ();
 sg13g2_decap_4 FILLER_60_1338 ();
 sg13g2_fill_1 FILLER_60_1342 ();
 sg13g2_decap_4 FILLER_60_1347 ();
 sg13g2_fill_2 FILLER_60_1351 ();
 sg13g2_decap_8 FILLER_60_1357 ();
 sg13g2_fill_2 FILLER_60_1364 ();
 sg13g2_fill_1 FILLER_60_1366 ();
 sg13g2_decap_8 FILLER_60_1371 ();
 sg13g2_decap_8 FILLER_60_1378 ();
 sg13g2_decap_8 FILLER_60_1385 ();
 sg13g2_decap_4 FILLER_60_1392 ();
 sg13g2_fill_1 FILLER_60_1396 ();
 sg13g2_fill_2 FILLER_60_1401 ();
 sg13g2_fill_1 FILLER_60_1411 ();
 sg13g2_fill_2 FILLER_60_1426 ();
 sg13g2_fill_1 FILLER_60_1428 ();
 sg13g2_decap_4 FILLER_60_1447 ();
 sg13g2_fill_1 FILLER_60_1451 ();
 sg13g2_decap_4 FILLER_60_1463 ();
 sg13g2_fill_2 FILLER_60_1467 ();
 sg13g2_decap_8 FILLER_60_1480 ();
 sg13g2_decap_4 FILLER_60_1487 ();
 sg13g2_fill_1 FILLER_60_1495 ();
 sg13g2_decap_8 FILLER_60_1508 ();
 sg13g2_fill_1 FILLER_60_1515 ();
 sg13g2_fill_1 FILLER_60_1520 ();
 sg13g2_decap_8 FILLER_60_1530 ();
 sg13g2_decap_8 FILLER_60_1537 ();
 sg13g2_fill_1 FILLER_60_1544 ();
 sg13g2_decap_4 FILLER_60_1550 ();
 sg13g2_fill_2 FILLER_60_1554 ();
 sg13g2_decap_4 FILLER_60_1572 ();
 sg13g2_decap_4 FILLER_60_1580 ();
 sg13g2_decap_4 FILLER_60_1593 ();
 sg13g2_fill_2 FILLER_60_1597 ();
 sg13g2_decap_8 FILLER_60_1603 ();
 sg13g2_fill_1 FILLER_60_1610 ();
 sg13g2_fill_2 FILLER_60_1620 ();
 sg13g2_fill_2 FILLER_60_1631 ();
 sg13g2_fill_1 FILLER_60_1644 ();
 sg13g2_fill_2 FILLER_60_1652 ();
 sg13g2_fill_1 FILLER_60_1672 ();
 sg13g2_decap_8 FILLER_60_1683 ();
 sg13g2_decap_8 FILLER_60_1690 ();
 sg13g2_decap_8 FILLER_60_1697 ();
 sg13g2_decap_8 FILLER_60_1704 ();
 sg13g2_decap_8 FILLER_60_1711 ();
 sg13g2_decap_8 FILLER_60_1718 ();
 sg13g2_decap_8 FILLER_60_1725 ();
 sg13g2_decap_8 FILLER_60_1732 ();
 sg13g2_decap_8 FILLER_60_1739 ();
 sg13g2_decap_8 FILLER_60_1746 ();
 sg13g2_decap_8 FILLER_60_1753 ();
 sg13g2_decap_8 FILLER_60_1760 ();
 sg13g2_decap_8 FILLER_60_1767 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_17 ();
 sg13g2_fill_1 FILLER_61_19 ();
 sg13g2_fill_2 FILLER_61_25 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_fill_2 FILLER_61_42 ();
 sg13g2_fill_1 FILLER_61_44 ();
 sg13g2_fill_2 FILLER_61_57 ();
 sg13g2_fill_2 FILLER_61_64 ();
 sg13g2_fill_1 FILLER_61_66 ();
 sg13g2_fill_2 FILLER_61_75 ();
 sg13g2_fill_1 FILLER_61_77 ();
 sg13g2_fill_2 FILLER_61_88 ();
 sg13g2_fill_1 FILLER_61_95 ();
 sg13g2_decap_8 FILLER_61_116 ();
 sg13g2_decap_8 FILLER_61_123 ();
 sg13g2_decap_8 FILLER_61_141 ();
 sg13g2_decap_8 FILLER_61_148 ();
 sg13g2_decap_8 FILLER_61_155 ();
 sg13g2_decap_8 FILLER_61_162 ();
 sg13g2_fill_1 FILLER_61_169 ();
 sg13g2_decap_4 FILLER_61_194 ();
 sg13g2_fill_1 FILLER_61_198 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_fill_1 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_215 ();
 sg13g2_decap_4 FILLER_61_222 ();
 sg13g2_fill_2 FILLER_61_226 ();
 sg13g2_decap_4 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_242 ();
 sg13g2_fill_2 FILLER_61_248 ();
 sg13g2_decap_8 FILLER_61_254 ();
 sg13g2_decap_8 FILLER_61_261 ();
 sg13g2_decap_4 FILLER_61_268 ();
 sg13g2_fill_1 FILLER_61_285 ();
 sg13g2_decap_8 FILLER_61_296 ();
 sg13g2_decap_8 FILLER_61_303 ();
 sg13g2_fill_1 FILLER_61_310 ();
 sg13g2_decap_8 FILLER_61_330 ();
 sg13g2_fill_2 FILLER_61_337 ();
 sg13g2_fill_1 FILLER_61_339 ();
 sg13g2_fill_2 FILLER_61_354 ();
 sg13g2_decap_8 FILLER_61_360 ();
 sg13g2_fill_1 FILLER_61_367 ();
 sg13g2_decap_8 FILLER_61_376 ();
 sg13g2_fill_1 FILLER_61_383 ();
 sg13g2_decap_8 FILLER_61_390 ();
 sg13g2_decap_8 FILLER_61_397 ();
 sg13g2_decap_8 FILLER_61_404 ();
 sg13g2_decap_4 FILLER_61_411 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_decap_4 FILLER_61_428 ();
 sg13g2_fill_2 FILLER_61_432 ();
 sg13g2_fill_2 FILLER_61_442 ();
 sg13g2_fill_1 FILLER_61_444 ();
 sg13g2_decap_8 FILLER_61_450 ();
 sg13g2_decap_8 FILLER_61_457 ();
 sg13g2_fill_2 FILLER_61_464 ();
 sg13g2_decap_8 FILLER_61_490 ();
 sg13g2_decap_8 FILLER_61_501 ();
 sg13g2_fill_1 FILLER_61_508 ();
 sg13g2_decap_8 FILLER_61_519 ();
 sg13g2_decap_4 FILLER_61_526 ();
 sg13g2_fill_2 FILLER_61_530 ();
 sg13g2_decap_8 FILLER_61_561 ();
 sg13g2_decap_8 FILLER_61_568 ();
 sg13g2_decap_8 FILLER_61_575 ();
 sg13g2_fill_2 FILLER_61_582 ();
 sg13g2_fill_1 FILLER_61_584 ();
 sg13g2_fill_2 FILLER_61_590 ();
 sg13g2_fill_1 FILLER_61_592 ();
 sg13g2_decap_8 FILLER_61_598 ();
 sg13g2_fill_2 FILLER_61_605 ();
 sg13g2_fill_1 FILLER_61_607 ();
 sg13g2_decap_4 FILLER_61_613 ();
 sg13g2_decap_4 FILLER_61_626 ();
 sg13g2_decap_8 FILLER_61_635 ();
 sg13g2_fill_2 FILLER_61_642 ();
 sg13g2_fill_1 FILLER_61_644 ();
 sg13g2_decap_8 FILLER_61_654 ();
 sg13g2_decap_4 FILLER_61_661 ();
 sg13g2_fill_2 FILLER_61_665 ();
 sg13g2_decap_4 FILLER_61_686 ();
 sg13g2_fill_2 FILLER_61_694 ();
 sg13g2_decap_4 FILLER_61_708 ();
 sg13g2_fill_2 FILLER_61_712 ();
 sg13g2_fill_1 FILLER_61_740 ();
 sg13g2_decap_8 FILLER_61_745 ();
 sg13g2_decap_8 FILLER_61_752 ();
 sg13g2_fill_1 FILLER_61_759 ();
 sg13g2_fill_1 FILLER_61_800 ();
 sg13g2_decap_8 FILLER_61_812 ();
 sg13g2_decap_8 FILLER_61_819 ();
 sg13g2_decap_4 FILLER_61_826 ();
 sg13g2_fill_1 FILLER_61_839 ();
 sg13g2_decap_8 FILLER_61_848 ();
 sg13g2_decap_4 FILLER_61_855 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_decap_4 FILLER_61_868 ();
 sg13g2_fill_1 FILLER_61_886 ();
 sg13g2_decap_4 FILLER_61_891 ();
 sg13g2_decap_8 FILLER_61_921 ();
 sg13g2_decap_8 FILLER_61_928 ();
 sg13g2_fill_2 FILLER_61_935 ();
 sg13g2_decap_4 FILLER_61_946 ();
 sg13g2_fill_2 FILLER_61_950 ();
 sg13g2_fill_2 FILLER_61_961 ();
 sg13g2_fill_2 FILLER_61_970 ();
 sg13g2_decap_8 FILLER_61_978 ();
 sg13g2_decap_4 FILLER_61_985 ();
 sg13g2_fill_2 FILLER_61_1015 ();
 sg13g2_fill_2 FILLER_61_1035 ();
 sg13g2_decap_8 FILLER_61_1063 ();
 sg13g2_decap_8 FILLER_61_1070 ();
 sg13g2_decap_8 FILLER_61_1077 ();
 sg13g2_decap_4 FILLER_61_1084 ();
 sg13g2_fill_2 FILLER_61_1088 ();
 sg13g2_decap_8 FILLER_61_1095 ();
 sg13g2_decap_8 FILLER_61_1112 ();
 sg13g2_decap_8 FILLER_61_1119 ();
 sg13g2_decap_8 FILLER_61_1126 ();
 sg13g2_decap_4 FILLER_61_1144 ();
 sg13g2_fill_2 FILLER_61_1148 ();
 sg13g2_fill_2 FILLER_61_1180 ();
 sg13g2_fill_1 FILLER_61_1182 ();
 sg13g2_decap_8 FILLER_61_1213 ();
 sg13g2_decap_4 FILLER_61_1220 ();
 sg13g2_fill_2 FILLER_61_1224 ();
 sg13g2_fill_1 FILLER_61_1248 ();
 sg13g2_decap_4 FILLER_61_1253 ();
 sg13g2_decap_8 FILLER_61_1288 ();
 sg13g2_decap_4 FILLER_61_1295 ();
 sg13g2_decap_4 FILLER_61_1415 ();
 sg13g2_fill_1 FILLER_61_1419 ();
 sg13g2_decap_8 FILLER_61_1441 ();
 sg13g2_fill_2 FILLER_61_1453 ();
 sg13g2_fill_2 FILLER_61_1459 ();
 sg13g2_decap_4 FILLER_61_1469 ();
 sg13g2_decap_4 FILLER_61_1477 ();
 sg13g2_fill_2 FILLER_61_1481 ();
 sg13g2_decap_4 FILLER_61_1487 ();
 sg13g2_fill_2 FILLER_61_1491 ();
 sg13g2_fill_2 FILLER_61_1519 ();
 sg13g2_fill_1 FILLER_61_1521 ();
 sg13g2_decap_4 FILLER_61_1617 ();
 sg13g2_fill_2 FILLER_61_1621 ();
 sg13g2_fill_2 FILLER_61_1664 ();
 sg13g2_decap_8 FILLER_61_1692 ();
 sg13g2_decap_8 FILLER_61_1699 ();
 sg13g2_decap_8 FILLER_61_1706 ();
 sg13g2_decap_8 FILLER_61_1713 ();
 sg13g2_decap_8 FILLER_61_1720 ();
 sg13g2_decap_8 FILLER_61_1727 ();
 sg13g2_decap_8 FILLER_61_1734 ();
 sg13g2_decap_8 FILLER_61_1741 ();
 sg13g2_decap_8 FILLER_61_1748 ();
 sg13g2_decap_8 FILLER_61_1755 ();
 sg13g2_decap_8 FILLER_61_1762 ();
 sg13g2_decap_4 FILLER_61_1769 ();
 sg13g2_fill_1 FILLER_61_1773 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_29 ();
 sg13g2_decap_8 FILLER_62_36 ();
 sg13g2_fill_2 FILLER_62_43 ();
 sg13g2_fill_1 FILLER_62_45 ();
 sg13g2_decap_8 FILLER_62_55 ();
 sg13g2_fill_1 FILLER_62_62 ();
 sg13g2_decap_4 FILLER_62_76 ();
 sg13g2_fill_1 FILLER_62_80 ();
 sg13g2_decap_4 FILLER_62_116 ();
 sg13g2_fill_1 FILLER_62_120 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_4 FILLER_62_161 ();
 sg13g2_decap_4 FILLER_62_169 ();
 sg13g2_fill_2 FILLER_62_180 ();
 sg13g2_decap_4 FILLER_62_200 ();
 sg13g2_fill_1 FILLER_62_204 ();
 sg13g2_fill_1 FILLER_62_218 ();
 sg13g2_decap_8 FILLER_62_223 ();
 sg13g2_decap_8 FILLER_62_243 ();
 sg13g2_decap_4 FILLER_62_250 ();
 sg13g2_fill_1 FILLER_62_254 ();
 sg13g2_fill_2 FILLER_62_263 ();
 sg13g2_fill_2 FILLER_62_278 ();
 sg13g2_fill_1 FILLER_62_280 ();
 sg13g2_decap_8 FILLER_62_286 ();
 sg13g2_fill_2 FILLER_62_293 ();
 sg13g2_fill_2 FILLER_62_303 ();
 sg13g2_decap_4 FILLER_62_310 ();
 sg13g2_fill_2 FILLER_62_314 ();
 sg13g2_fill_2 FILLER_62_327 ();
 sg13g2_decap_8 FILLER_62_337 ();
 sg13g2_decap_4 FILLER_62_344 ();
 sg13g2_fill_2 FILLER_62_393 ();
 sg13g2_fill_1 FILLER_62_395 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_fill_1 FILLER_62_409 ();
 sg13g2_decap_4 FILLER_62_415 ();
 sg13g2_decap_4 FILLER_62_431 ();
 sg13g2_fill_1 FILLER_62_435 ();
 sg13g2_fill_2 FILLER_62_445 ();
 sg13g2_fill_2 FILLER_62_455 ();
 sg13g2_fill_1 FILLER_62_457 ();
 sg13g2_decap_8 FILLER_62_462 ();
 sg13g2_decap_4 FILLER_62_469 ();
 sg13g2_fill_1 FILLER_62_473 ();
 sg13g2_decap_8 FILLER_62_494 ();
 sg13g2_fill_2 FILLER_62_501 ();
 sg13g2_decap_8 FILLER_62_516 ();
 sg13g2_fill_2 FILLER_62_523 ();
 sg13g2_fill_2 FILLER_62_535 ();
 sg13g2_fill_2 FILLER_62_542 ();
 sg13g2_fill_1 FILLER_62_544 ();
 sg13g2_decap_8 FILLER_62_569 ();
 sg13g2_fill_2 FILLER_62_576 ();
 sg13g2_fill_1 FILLER_62_588 ();
 sg13g2_decap_8 FILLER_62_598 ();
 sg13g2_decap_8 FILLER_62_605 ();
 sg13g2_decap_4 FILLER_62_612 ();
 sg13g2_fill_2 FILLER_62_616 ();
 sg13g2_decap_4 FILLER_62_634 ();
 sg13g2_fill_2 FILLER_62_638 ();
 sg13g2_decap_8 FILLER_62_653 ();
 sg13g2_decap_8 FILLER_62_681 ();
 sg13g2_decap_4 FILLER_62_688 ();
 sg13g2_decap_4 FILLER_62_718 ();
 sg13g2_fill_1 FILLER_62_722 ();
 sg13g2_decap_4 FILLER_62_727 ();
 sg13g2_fill_1 FILLER_62_731 ();
 sg13g2_decap_4 FILLER_62_758 ();
 sg13g2_fill_1 FILLER_62_762 ();
 sg13g2_decap_8 FILLER_62_789 ();
 sg13g2_decap_4 FILLER_62_831 ();
 sg13g2_decap_8 FILLER_62_845 ();
 sg13g2_fill_1 FILLER_62_852 ();
 sg13g2_fill_1 FILLER_62_857 ();
 sg13g2_fill_1 FILLER_62_863 ();
 sg13g2_decap_4 FILLER_62_873 ();
 sg13g2_fill_1 FILLER_62_877 ();
 sg13g2_decap_8 FILLER_62_883 ();
 sg13g2_decap_8 FILLER_62_890 ();
 sg13g2_decap_8 FILLER_62_897 ();
 sg13g2_decap_4 FILLER_62_909 ();
 sg13g2_decap_4 FILLER_62_917 ();
 sg13g2_fill_1 FILLER_62_921 ();
 sg13g2_decap_8 FILLER_62_927 ();
 sg13g2_decap_8 FILLER_62_934 ();
 sg13g2_decap_8 FILLER_62_941 ();
 sg13g2_fill_1 FILLER_62_948 ();
 sg13g2_decap_8 FILLER_62_954 ();
 sg13g2_fill_2 FILLER_62_961 ();
 sg13g2_fill_1 FILLER_62_963 ();
 sg13g2_fill_1 FILLER_62_988 ();
 sg13g2_fill_2 FILLER_62_994 ();
 sg13g2_decap_8 FILLER_62_1001 ();
 sg13g2_fill_2 FILLER_62_1008 ();
 sg13g2_fill_2 FILLER_62_1017 ();
 sg13g2_fill_1 FILLER_62_1019 ();
 sg13g2_decap_4 FILLER_62_1027 ();
 sg13g2_fill_1 FILLER_62_1031 ();
 sg13g2_decap_8 FILLER_62_1035 ();
 sg13g2_fill_2 FILLER_62_1042 ();
 sg13g2_fill_1 FILLER_62_1044 ();
 sg13g2_decap_8 FILLER_62_1049 ();
 sg13g2_fill_1 FILLER_62_1056 ();
 sg13g2_decap_4 FILLER_62_1087 ();
 sg13g2_fill_2 FILLER_62_1091 ();
 sg13g2_decap_4 FILLER_62_1123 ();
 sg13g2_decap_8 FILLER_62_1131 ();
 sg13g2_decap_8 FILLER_62_1138 ();
 sg13g2_fill_2 FILLER_62_1145 ();
 sg13g2_fill_1 FILLER_62_1147 ();
 sg13g2_decap_8 FILLER_62_1152 ();
 sg13g2_decap_8 FILLER_62_1168 ();
 sg13g2_fill_2 FILLER_62_1175 ();
 sg13g2_fill_1 FILLER_62_1177 ();
 sg13g2_decap_8 FILLER_62_1182 ();
 sg13g2_fill_2 FILLER_62_1203 ();
 sg13g2_fill_1 FILLER_62_1205 ();
 sg13g2_decap_8 FILLER_62_1267 ();
 sg13g2_fill_2 FILLER_62_1274 ();
 sg13g2_decap_4 FILLER_62_1280 ();
 sg13g2_decap_4 FILLER_62_1288 ();
 sg13g2_fill_1 FILLER_62_1292 ();
 sg13g2_fill_1 FILLER_62_1298 ();
 sg13g2_decap_4 FILLER_62_1304 ();
 sg13g2_decap_4 FILLER_62_1313 ();
 sg13g2_decap_8 FILLER_62_1321 ();
 sg13g2_fill_2 FILLER_62_1332 ();
 sg13g2_fill_1 FILLER_62_1334 ();
 sg13g2_decap_8 FILLER_62_1340 ();
 sg13g2_decap_8 FILLER_62_1356 ();
 sg13g2_decap_8 FILLER_62_1363 ();
 sg13g2_fill_2 FILLER_62_1370 ();
 sg13g2_decap_8 FILLER_62_1376 ();
 sg13g2_decap_8 FILLER_62_1383 ();
 sg13g2_fill_2 FILLER_62_1390 ();
 sg13g2_fill_1 FILLER_62_1392 ();
 sg13g2_decap_4 FILLER_62_1397 ();
 sg13g2_decap_8 FILLER_62_1414 ();
 sg13g2_decap_4 FILLER_62_1421 ();
 sg13g2_fill_2 FILLER_62_1425 ();
 sg13g2_decap_4 FILLER_62_1457 ();
 sg13g2_fill_1 FILLER_62_1465 ();
 sg13g2_decap_4 FILLER_62_1497 ();
 sg13g2_fill_2 FILLER_62_1505 ();
 sg13g2_fill_1 FILLER_62_1507 ();
 sg13g2_decap_8 FILLER_62_1513 ();
 sg13g2_decap_8 FILLER_62_1520 ();
 sg13g2_fill_2 FILLER_62_1527 ();
 sg13g2_fill_2 FILLER_62_1547 ();
 sg13g2_fill_1 FILLER_62_1632 ();
 sg13g2_fill_1 FILLER_62_1636 ();
 sg13g2_fill_1 FILLER_62_1641 ();
 sg13g2_fill_1 FILLER_62_1650 ();
 sg13g2_fill_1 FILLER_62_1660 ();
 sg13g2_fill_2 FILLER_62_1665 ();
 sg13g2_fill_1 FILLER_62_1667 ();
 sg13g2_fill_2 FILLER_62_1672 ();
 sg13g2_fill_1 FILLER_62_1674 ();
 sg13g2_decap_8 FILLER_62_1679 ();
 sg13g2_decap_8 FILLER_62_1686 ();
 sg13g2_decap_8 FILLER_62_1693 ();
 sg13g2_decap_8 FILLER_62_1700 ();
 sg13g2_decap_8 FILLER_62_1707 ();
 sg13g2_decap_8 FILLER_62_1714 ();
 sg13g2_decap_8 FILLER_62_1721 ();
 sg13g2_decap_8 FILLER_62_1728 ();
 sg13g2_decap_8 FILLER_62_1735 ();
 sg13g2_decap_8 FILLER_62_1742 ();
 sg13g2_decap_8 FILLER_62_1749 ();
 sg13g2_decap_8 FILLER_62_1756 ();
 sg13g2_decap_8 FILLER_62_1763 ();
 sg13g2_decap_4 FILLER_62_1770 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_fill_2 FILLER_63_14 ();
 sg13g2_decap_4 FILLER_63_47 ();
 sg13g2_fill_1 FILLER_63_51 ();
 sg13g2_decap_4 FILLER_63_57 ();
 sg13g2_decap_4 FILLER_63_66 ();
 sg13g2_fill_1 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_76 ();
 sg13g2_decap_4 FILLER_63_96 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_fill_2 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_107 ();
 sg13g2_decap_4 FILLER_63_114 ();
 sg13g2_fill_1 FILLER_63_118 ();
 sg13g2_decap_4 FILLER_63_127 ();
 sg13g2_fill_1 FILLER_63_131 ();
 sg13g2_fill_2 FILLER_63_137 ();
 sg13g2_fill_1 FILLER_63_139 ();
 sg13g2_fill_2 FILLER_63_144 ();
 sg13g2_fill_1 FILLER_63_153 ();
 sg13g2_decap_8 FILLER_63_159 ();
 sg13g2_fill_1 FILLER_63_166 ();
 sg13g2_decap_4 FILLER_63_171 ();
 sg13g2_decap_4 FILLER_63_182 ();
 sg13g2_fill_2 FILLER_63_186 ();
 sg13g2_decap_4 FILLER_63_206 ();
 sg13g2_fill_1 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_231 ();
 sg13g2_decap_4 FILLER_63_236 ();
 sg13g2_fill_1 FILLER_63_240 ();
 sg13g2_fill_1 FILLER_63_259 ();
 sg13g2_fill_1 FILLER_63_275 ();
 sg13g2_decap_4 FILLER_63_280 ();
 sg13g2_decap_4 FILLER_63_296 ();
 sg13g2_fill_1 FILLER_63_300 ();
 sg13g2_fill_1 FILLER_63_306 ();
 sg13g2_fill_2 FILLER_63_311 ();
 sg13g2_fill_1 FILLER_63_313 ();
 sg13g2_decap_8 FILLER_63_321 ();
 sg13g2_decap_4 FILLER_63_328 ();
 sg13g2_decap_8 FILLER_63_337 ();
 sg13g2_decap_4 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_358 ();
 sg13g2_decap_8 FILLER_63_365 ();
 sg13g2_decap_8 FILLER_63_372 ();
 sg13g2_fill_1 FILLER_63_379 ();
 sg13g2_decap_8 FILLER_63_384 ();
 sg13g2_decap_4 FILLER_63_413 ();
 sg13g2_fill_2 FILLER_63_417 ();
 sg13g2_fill_2 FILLER_63_424 ();
 sg13g2_fill_1 FILLER_63_426 ();
 sg13g2_decap_4 FILLER_63_440 ();
 sg13g2_fill_2 FILLER_63_444 ();
 sg13g2_fill_1 FILLER_63_456 ();
 sg13g2_fill_2 FILLER_63_481 ();
 sg13g2_decap_4 FILLER_63_514 ();
 sg13g2_decap_8 FILLER_63_524 ();
 sg13g2_fill_2 FILLER_63_540 ();
 sg13g2_fill_1 FILLER_63_542 ();
 sg13g2_fill_1 FILLER_63_552 ();
 sg13g2_fill_1 FILLER_63_562 ();
 sg13g2_decap_4 FILLER_63_573 ();
 sg13g2_fill_2 FILLER_63_592 ();
 sg13g2_fill_2 FILLER_63_600 ();
 sg13g2_fill_1 FILLER_63_602 ();
 sg13g2_fill_2 FILLER_63_610 ();
 sg13g2_decap_4 FILLER_63_620 ();
 sg13g2_fill_2 FILLER_63_624 ();
 sg13g2_fill_1 FILLER_63_631 ();
 sg13g2_decap_8 FILLER_63_639 ();
 sg13g2_decap_8 FILLER_63_646 ();
 sg13g2_fill_2 FILLER_63_653 ();
 sg13g2_fill_1 FILLER_63_655 ();
 sg13g2_decap_8 FILLER_63_672 ();
 sg13g2_decap_8 FILLER_63_679 ();
 sg13g2_decap_8 FILLER_63_686 ();
 sg13g2_decap_4 FILLER_63_693 ();
 sg13g2_fill_2 FILLER_63_697 ();
 sg13g2_fill_2 FILLER_63_703 ();
 sg13g2_fill_2 FILLER_63_721 ();
 sg13g2_fill_1 FILLER_63_723 ();
 sg13g2_decap_8 FILLER_63_733 ();
 sg13g2_decap_8 FILLER_63_740 ();
 sg13g2_fill_1 FILLER_63_747 ();
 sg13g2_decap_8 FILLER_63_758 ();
 sg13g2_decap_4 FILLER_63_765 ();
 sg13g2_decap_8 FILLER_63_773 ();
 sg13g2_decap_8 FILLER_63_780 ();
 sg13g2_decap_8 FILLER_63_787 ();
 sg13g2_decap_8 FILLER_63_794 ();
 sg13g2_fill_2 FILLER_63_801 ();
 sg13g2_decap_8 FILLER_63_807 ();
 sg13g2_fill_1 FILLER_63_814 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_fill_2 FILLER_63_826 ();
 sg13g2_decap_4 FILLER_63_832 ();
 sg13g2_fill_1 FILLER_63_836 ();
 sg13g2_decap_8 FILLER_63_841 ();
 sg13g2_decap_4 FILLER_63_848 ();
 sg13g2_fill_2 FILLER_63_852 ();
 sg13g2_fill_2 FILLER_63_888 ();
 sg13g2_fill_2 FILLER_63_894 ();
 sg13g2_fill_1 FILLER_63_896 ();
 sg13g2_fill_2 FILLER_63_902 ();
 sg13g2_decap_8 FILLER_63_918 ();
 sg13g2_decap_8 FILLER_63_925 ();
 sg13g2_decap_8 FILLER_63_932 ();
 sg13g2_fill_1 FILLER_63_939 ();
 sg13g2_decap_8 FILLER_63_996 ();
 sg13g2_fill_2 FILLER_63_1020 ();
 sg13g2_decap_8 FILLER_63_1074 ();
 sg13g2_fill_2 FILLER_63_1081 ();
 sg13g2_fill_1 FILLER_63_1083 ();
 sg13g2_decap_4 FILLER_63_1114 ();
 sg13g2_fill_2 FILLER_63_1118 ();
 sg13g2_decap_4 FILLER_63_1146 ();
 sg13g2_fill_1 FILLER_63_1150 ();
 sg13g2_fill_2 FILLER_63_1156 ();
 sg13g2_fill_2 FILLER_63_1162 ();
 sg13g2_decap_8 FILLER_63_1190 ();
 sg13g2_decap_8 FILLER_63_1201 ();
 sg13g2_decap_8 FILLER_63_1208 ();
 sg13g2_fill_2 FILLER_63_1215 ();
 sg13g2_fill_1 FILLER_63_1222 ();
 sg13g2_fill_2 FILLER_63_1227 ();
 sg13g2_fill_1 FILLER_63_1229 ();
 sg13g2_decap_8 FILLER_63_1234 ();
 sg13g2_decap_4 FILLER_63_1241 ();
 sg13g2_fill_2 FILLER_63_1245 ();
 sg13g2_fill_1 FILLER_63_1278 ();
 sg13g2_fill_2 FILLER_63_1310 ();
 sg13g2_fill_2 FILLER_63_1356 ();
 sg13g2_decap_8 FILLER_63_1384 ();
 sg13g2_fill_2 FILLER_63_1391 ();
 sg13g2_fill_1 FILLER_63_1393 ();
 sg13g2_fill_2 FILLER_63_1424 ();
 sg13g2_fill_1 FILLER_63_1426 ();
 sg13g2_decap_4 FILLER_63_1432 ();
 sg13g2_fill_1 FILLER_63_1436 ();
 sg13g2_decap_4 FILLER_63_1447 ();
 sg13g2_fill_2 FILLER_63_1451 ();
 sg13g2_decap_4 FILLER_63_1483 ();
 sg13g2_decap_4 FILLER_63_1539 ();
 sg13g2_fill_2 FILLER_63_1569 ();
 sg13g2_decap_8 FILLER_63_1576 ();
 sg13g2_decap_4 FILLER_63_1583 ();
 sg13g2_decap_8 FILLER_63_1591 ();
 sg13g2_decap_8 FILLER_63_1598 ();
 sg13g2_decap_8 FILLER_63_1605 ();
 sg13g2_fill_1 FILLER_63_1612 ();
 sg13g2_fill_2 FILLER_63_1626 ();
 sg13g2_fill_2 FILLER_63_1658 ();
 sg13g2_decap_8 FILLER_63_1698 ();
 sg13g2_decap_8 FILLER_63_1705 ();
 sg13g2_decap_8 FILLER_63_1712 ();
 sg13g2_decap_8 FILLER_63_1719 ();
 sg13g2_decap_8 FILLER_63_1726 ();
 sg13g2_decap_8 FILLER_63_1733 ();
 sg13g2_decap_8 FILLER_63_1740 ();
 sg13g2_decap_8 FILLER_63_1747 ();
 sg13g2_decap_8 FILLER_63_1754 ();
 sg13g2_decap_8 FILLER_63_1761 ();
 sg13g2_decap_4 FILLER_63_1768 ();
 sg13g2_fill_2 FILLER_63_1772 ();
 sg13g2_decap_4 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_4 ();
 sg13g2_decap_8 FILLER_64_18 ();
 sg13g2_fill_1 FILLER_64_25 ();
 sg13g2_fill_2 FILLER_64_36 ();
 sg13g2_decap_4 FILLER_64_69 ();
 sg13g2_fill_2 FILLER_64_73 ();
 sg13g2_decap_8 FILLER_64_79 ();
 sg13g2_decap_8 FILLER_64_99 ();
 sg13g2_fill_2 FILLER_64_106 ();
 sg13g2_fill_2 FILLER_64_126 ();
 sg13g2_fill_1 FILLER_64_128 ();
 sg13g2_fill_2 FILLER_64_142 ();
 sg13g2_fill_2 FILLER_64_151 ();
 sg13g2_fill_2 FILLER_64_161 ();
 sg13g2_fill_1 FILLER_64_163 ();
 sg13g2_fill_1 FILLER_64_191 ();
 sg13g2_decap_8 FILLER_64_205 ();
 sg13g2_fill_2 FILLER_64_212 ();
 sg13g2_fill_1 FILLER_64_214 ();
 sg13g2_decap_8 FILLER_64_220 ();
 sg13g2_decap_4 FILLER_64_227 ();
 sg13g2_decap_8 FILLER_64_236 ();
 sg13g2_decap_8 FILLER_64_243 ();
 sg13g2_decap_4 FILLER_64_250 ();
 sg13g2_decap_8 FILLER_64_274 ();
 sg13g2_decap_8 FILLER_64_281 ();
 sg13g2_decap_8 FILLER_64_288 ();
 sg13g2_decap_4 FILLER_64_295 ();
 sg13g2_fill_1 FILLER_64_299 ();
 sg13g2_fill_1 FILLER_64_311 ();
 sg13g2_decap_8 FILLER_64_340 ();
 sg13g2_decap_4 FILLER_64_347 ();
 sg13g2_fill_1 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_357 ();
 sg13g2_decap_8 FILLER_64_364 ();
 sg13g2_decap_4 FILLER_64_371 ();
 sg13g2_fill_2 FILLER_64_385 ();
 sg13g2_fill_2 FILLER_64_414 ();
 sg13g2_decap_8 FILLER_64_422 ();
 sg13g2_fill_1 FILLER_64_429 ();
 sg13g2_decap_8 FILLER_64_435 ();
 sg13g2_decap_8 FILLER_64_442 ();
 sg13g2_decap_8 FILLER_64_449 ();
 sg13g2_fill_2 FILLER_64_456 ();
 sg13g2_fill_1 FILLER_64_458 ();
 sg13g2_fill_1 FILLER_64_464 ();
 sg13g2_decap_8 FILLER_64_485 ();
 sg13g2_decap_4 FILLER_64_492 ();
 sg13g2_fill_2 FILLER_64_496 ();
 sg13g2_fill_2 FILLER_64_506 ();
 sg13g2_fill_1 FILLER_64_508 ();
 sg13g2_decap_8 FILLER_64_518 ();
 sg13g2_decap_8 FILLER_64_525 ();
 sg13g2_fill_2 FILLER_64_532 ();
 sg13g2_fill_1 FILLER_64_534 ();
 sg13g2_decap_4 FILLER_64_539 ();
 sg13g2_fill_1 FILLER_64_560 ();
 sg13g2_fill_2 FILLER_64_567 ();
 sg13g2_fill_1 FILLER_64_569 ();
 sg13g2_fill_2 FILLER_64_575 ();
 sg13g2_fill_2 FILLER_64_584 ();
 sg13g2_decap_4 FILLER_64_593 ();
 sg13g2_decap_4 FILLER_64_602 ();
 sg13g2_fill_2 FILLER_64_611 ();
 sg13g2_decap_8 FILLER_64_618 ();
 sg13g2_decap_8 FILLER_64_625 ();
 sg13g2_decap_4 FILLER_64_632 ();
 sg13g2_fill_1 FILLER_64_636 ();
 sg13g2_fill_2 FILLER_64_642 ();
 sg13g2_fill_2 FILLER_64_648 ();
 sg13g2_fill_1 FILLER_64_650 ();
 sg13g2_fill_2 FILLER_64_673 ();
 sg13g2_fill_2 FILLER_64_679 ();
 sg13g2_fill_1 FILLER_64_681 ();
 sg13g2_fill_1 FILLER_64_723 ();
 sg13g2_decap_4 FILLER_64_759 ();
 sg13g2_fill_1 FILLER_64_772 ();
 sg13g2_fill_1 FILLER_64_783 ();
 sg13g2_fill_2 FILLER_64_804 ();
 sg13g2_fill_2 FILLER_64_821 ();
 sg13g2_fill_1 FILLER_64_833 ();
 sg13g2_fill_2 FILLER_64_841 ();
 sg13g2_decap_8 FILLER_64_848 ();
 sg13g2_decap_8 FILLER_64_859 ();
 sg13g2_decap_8 FILLER_64_866 ();
 sg13g2_decap_4 FILLER_64_873 ();
 sg13g2_fill_1 FILLER_64_877 ();
 sg13g2_fill_1 FILLER_64_888 ();
 sg13g2_fill_2 FILLER_64_899 ();
 sg13g2_fill_1 FILLER_64_901 ();
 sg13g2_fill_2 FILLER_64_912 ();
 sg13g2_fill_2 FILLER_64_924 ();
 sg13g2_fill_2 FILLER_64_930 ();
 sg13g2_fill_1 FILLER_64_932 ();
 sg13g2_fill_2 FILLER_64_946 ();
 sg13g2_decap_8 FILLER_64_952 ();
 sg13g2_decap_8 FILLER_64_959 ();
 sg13g2_decap_8 FILLER_64_966 ();
 sg13g2_decap_4 FILLER_64_973 ();
 sg13g2_decap_8 FILLER_64_981 ();
 sg13g2_decap_8 FILLER_64_988 ();
 sg13g2_decap_8 FILLER_64_995 ();
 sg13g2_fill_1 FILLER_64_1002 ();
 sg13g2_fill_2 FILLER_64_1029 ();
 sg13g2_decap_8 FILLER_64_1035 ();
 sg13g2_decap_8 FILLER_64_1042 ();
 sg13g2_decap_4 FILLER_64_1049 ();
 sg13g2_fill_2 FILLER_64_1053 ();
 sg13g2_decap_8 FILLER_64_1059 ();
 sg13g2_decap_8 FILLER_64_1066 ();
 sg13g2_decap_8 FILLER_64_1073 ();
 sg13g2_fill_1 FILLER_64_1080 ();
 sg13g2_decap_8 FILLER_64_1085 ();
 sg13g2_decap_8 FILLER_64_1092 ();
 sg13g2_decap_8 FILLER_64_1099 ();
 sg13g2_decap_4 FILLER_64_1106 ();
 sg13g2_fill_1 FILLER_64_1110 ();
 sg13g2_fill_1 FILLER_64_1159 ();
 sg13g2_fill_1 FILLER_64_1165 ();
 sg13g2_fill_1 FILLER_64_1170 ();
 sg13g2_fill_2 FILLER_64_1175 ();
 sg13g2_fill_2 FILLER_64_1186 ();
 sg13g2_fill_1 FILLER_64_1188 ();
 sg13g2_decap_8 FILLER_64_1246 ();
 sg13g2_decap_8 FILLER_64_1253 ();
 sg13g2_fill_2 FILLER_64_1260 ();
 sg13g2_fill_1 FILLER_64_1262 ();
 sg13g2_decap_8 FILLER_64_1267 ();
 sg13g2_decap_8 FILLER_64_1274 ();
 sg13g2_decap_8 FILLER_64_1281 ();
 sg13g2_fill_1 FILLER_64_1292 ();
 sg13g2_decap_8 FILLER_64_1305 ();
 sg13g2_decap_4 FILLER_64_1312 ();
 sg13g2_fill_2 FILLER_64_1316 ();
 sg13g2_fill_2 FILLER_64_1322 ();
 sg13g2_fill_1 FILLER_64_1324 ();
 sg13g2_fill_2 FILLER_64_1333 ();
 sg13g2_fill_1 FILLER_64_1335 ();
 sg13g2_fill_2 FILLER_64_1340 ();
 sg13g2_fill_1 FILLER_64_1342 ();
 sg13g2_decap_8 FILLER_64_1373 ();
 sg13g2_fill_1 FILLER_64_1380 ();
 sg13g2_decap_8 FILLER_64_1385 ();
 sg13g2_decap_8 FILLER_64_1392 ();
 sg13g2_fill_2 FILLER_64_1399 ();
 sg13g2_fill_1 FILLER_64_1401 ();
 sg13g2_decap_8 FILLER_64_1407 ();
 sg13g2_decap_4 FILLER_64_1414 ();
 sg13g2_decap_8 FILLER_64_1453 ();
 sg13g2_decap_8 FILLER_64_1460 ();
 sg13g2_fill_1 FILLER_64_1467 ();
 sg13g2_decap_8 FILLER_64_1472 ();
 sg13g2_decap_8 FILLER_64_1479 ();
 sg13g2_fill_2 FILLER_64_1508 ();
 sg13g2_decap_8 FILLER_64_1514 ();
 sg13g2_fill_1 FILLER_64_1521 ();
 sg13g2_decap_8 FILLER_64_1526 ();
 sg13g2_decap_8 FILLER_64_1533 ();
 sg13g2_fill_1 FILLER_64_1540 ();
 sg13g2_decap_4 FILLER_64_1546 ();
 sg13g2_decap_4 FILLER_64_1554 ();
 sg13g2_fill_1 FILLER_64_1558 ();
 sg13g2_decap_4 FILLER_64_1562 ();
 sg13g2_decap_4 FILLER_64_1576 ();
 sg13g2_decap_8 FILLER_64_1606 ();
 sg13g2_decap_8 FILLER_64_1613 ();
 sg13g2_decap_8 FILLER_64_1620 ();
 sg13g2_decap_8 FILLER_64_1627 ();
 sg13g2_decap_4 FILLER_64_1634 ();
 sg13g2_fill_1 FILLER_64_1638 ();
 sg13g2_decap_4 FILLER_64_1643 ();
 sg13g2_fill_2 FILLER_64_1647 ();
 sg13g2_decap_8 FILLER_64_1653 ();
 sg13g2_decap_8 FILLER_64_1660 ();
 sg13g2_decap_8 FILLER_64_1667 ();
 sg13g2_decap_8 FILLER_64_1674 ();
 sg13g2_decap_8 FILLER_64_1681 ();
 sg13g2_decap_8 FILLER_64_1688 ();
 sg13g2_decap_8 FILLER_64_1695 ();
 sg13g2_decap_8 FILLER_64_1702 ();
 sg13g2_decap_8 FILLER_64_1709 ();
 sg13g2_decap_8 FILLER_64_1716 ();
 sg13g2_decap_8 FILLER_64_1723 ();
 sg13g2_decap_8 FILLER_64_1730 ();
 sg13g2_decap_8 FILLER_64_1737 ();
 sg13g2_decap_8 FILLER_64_1744 ();
 sg13g2_decap_8 FILLER_64_1751 ();
 sg13g2_decap_8 FILLER_64_1758 ();
 sg13g2_decap_8 FILLER_64_1765 ();
 sg13g2_fill_2 FILLER_64_1772 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_11 ();
 sg13g2_decap_4 FILLER_65_25 ();
 sg13g2_fill_1 FILLER_65_29 ();
 sg13g2_fill_2 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_63 ();
 sg13g2_fill_1 FILLER_65_71 ();
 sg13g2_fill_1 FILLER_65_76 ();
 sg13g2_fill_1 FILLER_65_82 ();
 sg13g2_fill_2 FILLER_65_87 ();
 sg13g2_fill_1 FILLER_65_89 ();
 sg13g2_decap_8 FILLER_65_99 ();
 sg13g2_fill_2 FILLER_65_106 ();
 sg13g2_fill_1 FILLER_65_108 ();
 sg13g2_fill_1 FILLER_65_114 ();
 sg13g2_fill_2 FILLER_65_125 ();
 sg13g2_decap_8 FILLER_65_131 ();
 sg13g2_fill_1 FILLER_65_138 ();
 sg13g2_decap_8 FILLER_65_156 ();
 sg13g2_decap_8 FILLER_65_163 ();
 sg13g2_fill_2 FILLER_65_170 ();
 sg13g2_fill_1 FILLER_65_172 ();
 sg13g2_decap_8 FILLER_65_177 ();
 sg13g2_fill_1 FILLER_65_184 ();
 sg13g2_fill_1 FILLER_65_194 ();
 sg13g2_fill_1 FILLER_65_205 ();
 sg13g2_fill_2 FILLER_65_227 ();
 sg13g2_decap_4 FILLER_65_234 ();
 sg13g2_fill_1 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_249 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_decap_4 FILLER_65_295 ();
 sg13g2_fill_1 FILLER_65_299 ();
 sg13g2_decap_8 FILLER_65_305 ();
 sg13g2_decap_8 FILLER_65_312 ();
 sg13g2_fill_1 FILLER_65_319 ();
 sg13g2_fill_2 FILLER_65_336 ();
 sg13g2_fill_1 FILLER_65_338 ();
 sg13g2_decap_8 FILLER_65_351 ();
 sg13g2_decap_4 FILLER_65_358 ();
 sg13g2_fill_2 FILLER_65_362 ();
 sg13g2_fill_2 FILLER_65_386 ();
 sg13g2_fill_1 FILLER_65_388 ();
 sg13g2_decap_4 FILLER_65_394 ();
 sg13g2_fill_1 FILLER_65_398 ();
 sg13g2_decap_8 FILLER_65_413 ();
 sg13g2_fill_2 FILLER_65_420 ();
 sg13g2_decap_4 FILLER_65_432 ();
 sg13g2_fill_1 FILLER_65_436 ();
 sg13g2_fill_2 FILLER_65_443 ();
 sg13g2_decap_4 FILLER_65_450 ();
 sg13g2_fill_2 FILLER_65_454 ();
 sg13g2_fill_2 FILLER_65_469 ();
 sg13g2_fill_1 FILLER_65_471 ();
 sg13g2_fill_2 FILLER_65_478 ();
 sg13g2_fill_2 FILLER_65_484 ();
 sg13g2_fill_2 FILLER_65_501 ();
 sg13g2_fill_1 FILLER_65_512 ();
 sg13g2_fill_2 FILLER_65_518 ();
 sg13g2_fill_2 FILLER_65_546 ();
 sg13g2_fill_1 FILLER_65_548 ();
 sg13g2_fill_2 FILLER_65_557 ();
 sg13g2_fill_1 FILLER_65_559 ();
 sg13g2_fill_2 FILLER_65_573 ();
 sg13g2_fill_2 FILLER_65_582 ();
 sg13g2_fill_1 FILLER_65_584 ();
 sg13g2_fill_2 FILLER_65_593 ();
 sg13g2_fill_1 FILLER_65_595 ();
 sg13g2_fill_2 FILLER_65_602 ();
 sg13g2_fill_1 FILLER_65_604 ();
 sg13g2_decap_8 FILLER_65_622 ();
 sg13g2_decap_8 FILLER_65_629 ();
 sg13g2_decap_8 FILLER_65_636 ();
 sg13g2_fill_2 FILLER_65_643 ();
 sg13g2_fill_1 FILLER_65_645 ();
 sg13g2_decap_8 FILLER_65_651 ();
 sg13g2_decap_4 FILLER_65_658 ();
 sg13g2_decap_8 FILLER_65_670 ();
 sg13g2_decap_8 FILLER_65_677 ();
 sg13g2_decap_8 FILLER_65_684 ();
 sg13g2_decap_4 FILLER_65_691 ();
 sg13g2_fill_2 FILLER_65_695 ();
 sg13g2_fill_2 FILLER_65_701 ();
 sg13g2_fill_2 FILLER_65_707 ();
 sg13g2_fill_2 FILLER_65_714 ();
 sg13g2_fill_2 FILLER_65_721 ();
 sg13g2_fill_1 FILLER_65_723 ();
 sg13g2_fill_2 FILLER_65_728 ();
 sg13g2_fill_1 FILLER_65_730 ();
 sg13g2_fill_2 FILLER_65_741 ();
 sg13g2_decap_8 FILLER_65_747 ();
 sg13g2_decap_8 FILLER_65_754 ();
 sg13g2_decap_8 FILLER_65_761 ();
 sg13g2_fill_1 FILLER_65_773 ();
 sg13g2_decap_4 FILLER_65_778 ();
 sg13g2_fill_1 FILLER_65_782 ();
 sg13g2_decap_4 FILLER_65_787 ();
 sg13g2_fill_1 FILLER_65_800 ();
 sg13g2_fill_2 FILLER_65_806 ();
 sg13g2_fill_1 FILLER_65_812 ();
 sg13g2_fill_1 FILLER_65_823 ();
 sg13g2_decap_4 FILLER_65_833 ();
 sg13g2_fill_2 FILLER_65_837 ();
 sg13g2_fill_1 FILLER_65_853 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_fill_1 FILLER_65_870 ();
 sg13g2_fill_2 FILLER_65_875 ();
 sg13g2_decap_4 FILLER_65_881 ();
 sg13g2_fill_1 FILLER_65_885 ();
 sg13g2_fill_2 FILLER_65_905 ();
 sg13g2_fill_1 FILLER_65_917 ();
 sg13g2_fill_2 FILLER_65_930 ();
 sg13g2_fill_1 FILLER_65_932 ();
 sg13g2_fill_1 FILLER_65_940 ();
 sg13g2_decap_8 FILLER_65_967 ();
 sg13g2_fill_2 FILLER_65_974 ();
 sg13g2_decap_4 FILLER_65_980 ();
 sg13g2_fill_1 FILLER_65_984 ();
 sg13g2_fill_2 FILLER_65_993 ();
 sg13g2_fill_1 FILLER_65_995 ();
 sg13g2_fill_1 FILLER_65_1030 ();
 sg13g2_decap_8 FILLER_65_1035 ();
 sg13g2_fill_1 FILLER_65_1042 ();
 sg13g2_fill_2 FILLER_65_1100 ();
 sg13g2_fill_1 FILLER_65_1102 ();
 sg13g2_decap_8 FILLER_65_1111 ();
 sg13g2_decap_8 FILLER_65_1118 ();
 sg13g2_decap_8 FILLER_65_1125 ();
 sg13g2_decap_4 FILLER_65_1132 ();
 sg13g2_fill_2 FILLER_65_1136 ();
 sg13g2_fill_2 FILLER_65_1143 ();
 sg13g2_decap_8 FILLER_65_1189 ();
 sg13g2_decap_4 FILLER_65_1196 ();
 sg13g2_fill_1 FILLER_65_1200 ();
 sg13g2_decap_8 FILLER_65_1209 ();
 sg13g2_fill_1 FILLER_65_1216 ();
 sg13g2_decap_8 FILLER_65_1221 ();
 sg13g2_fill_2 FILLER_65_1228 ();
 sg13g2_fill_2 FILLER_65_1274 ();
 sg13g2_fill_1 FILLER_65_1276 ();
 sg13g2_fill_1 FILLER_65_1317 ();
 sg13g2_fill_2 FILLER_65_1349 ();
 sg13g2_fill_2 FILLER_65_1373 ();
 sg13g2_fill_2 FILLER_65_1409 ();
 sg13g2_decap_4 FILLER_65_1437 ();
 sg13g2_fill_2 FILLER_65_1441 ();
 sg13g2_decap_8 FILLER_65_1452 ();
 sg13g2_fill_2 FILLER_65_1459 ();
 sg13g2_fill_1 FILLER_65_1461 ();
 sg13g2_decap_4 FILLER_65_1497 ();
 sg13g2_fill_2 FILLER_65_1501 ();
 sg13g2_fill_2 FILLER_65_1507 ();
 sg13g2_fill_2 FILLER_65_1535 ();
 sg13g2_fill_2 FILLER_65_1547 ();
 sg13g2_fill_1 FILLER_65_1549 ();
 sg13g2_decap_4 FILLER_65_1554 ();
 sg13g2_fill_2 FILLER_65_1558 ();
 sg13g2_fill_2 FILLER_65_1572 ();
 sg13g2_decap_8 FILLER_65_1579 ();
 sg13g2_decap_8 FILLER_65_1590 ();
 sg13g2_decap_4 FILLER_65_1597 ();
 sg13g2_fill_2 FILLER_65_1601 ();
 sg13g2_decap_4 FILLER_65_1624 ();
 sg13g2_fill_1 FILLER_65_1628 ();
 sg13g2_decap_8 FILLER_65_1633 ();
 sg13g2_decap_8 FILLER_65_1640 ();
 sg13g2_decap_8 FILLER_65_1647 ();
 sg13g2_decap_8 FILLER_65_1654 ();
 sg13g2_decap_8 FILLER_65_1661 ();
 sg13g2_decap_8 FILLER_65_1668 ();
 sg13g2_decap_8 FILLER_65_1675 ();
 sg13g2_decap_8 FILLER_65_1682 ();
 sg13g2_decap_8 FILLER_65_1689 ();
 sg13g2_decap_8 FILLER_65_1696 ();
 sg13g2_decap_8 FILLER_65_1703 ();
 sg13g2_decap_8 FILLER_65_1710 ();
 sg13g2_decap_8 FILLER_65_1717 ();
 sg13g2_decap_8 FILLER_65_1724 ();
 sg13g2_decap_8 FILLER_65_1731 ();
 sg13g2_decap_8 FILLER_65_1738 ();
 sg13g2_decap_8 FILLER_65_1745 ();
 sg13g2_decap_8 FILLER_65_1752 ();
 sg13g2_decap_8 FILLER_65_1759 ();
 sg13g2_decap_8 FILLER_65_1766 ();
 sg13g2_fill_1 FILLER_65_1773 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_4 FILLER_66_14 ();
 sg13g2_fill_1 FILLER_66_18 ();
 sg13g2_fill_1 FILLER_66_65 ();
 sg13g2_fill_1 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_75 ();
 sg13g2_fill_1 FILLER_66_81 ();
 sg13g2_decap_4 FILLER_66_90 ();
 sg13g2_fill_2 FILLER_66_94 ();
 sg13g2_decap_4 FILLER_66_101 ();
 sg13g2_decap_8 FILLER_66_130 ();
 sg13g2_fill_1 FILLER_66_137 ();
 sg13g2_decap_4 FILLER_66_153 ();
 sg13g2_fill_1 FILLER_66_178 ();
 sg13g2_fill_1 FILLER_66_184 ();
 sg13g2_decap_8 FILLER_66_190 ();
 sg13g2_decap_4 FILLER_66_197 ();
 sg13g2_fill_1 FILLER_66_201 ();
 sg13g2_decap_4 FILLER_66_205 ();
 sg13g2_fill_1 FILLER_66_209 ();
 sg13g2_fill_2 FILLER_66_250 ();
 sg13g2_fill_1 FILLER_66_260 ();
 sg13g2_fill_1 FILLER_66_269 ();
 sg13g2_fill_1 FILLER_66_274 ();
 sg13g2_fill_1 FILLER_66_280 ();
 sg13g2_decap_4 FILLER_66_286 ();
 sg13g2_fill_1 FILLER_66_290 ();
 sg13g2_decap_4 FILLER_66_299 ();
 sg13g2_fill_1 FILLER_66_303 ();
 sg13g2_fill_1 FILLER_66_312 ();
 sg13g2_decap_8 FILLER_66_321 ();
 sg13g2_fill_2 FILLER_66_328 ();
 sg13g2_fill_2 FILLER_66_335 ();
 sg13g2_fill_2 FILLER_66_345 ();
 sg13g2_fill_1 FILLER_66_352 ();
 sg13g2_fill_1 FILLER_66_363 ();
 sg13g2_fill_1 FILLER_66_368 ();
 sg13g2_fill_1 FILLER_66_374 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_fill_2 FILLER_66_399 ();
 sg13g2_fill_2 FILLER_66_416 ();
 sg13g2_fill_1 FILLER_66_418 ();
 sg13g2_fill_2 FILLER_66_423 ();
 sg13g2_fill_1 FILLER_66_425 ();
 sg13g2_fill_2 FILLER_66_431 ();
 sg13g2_fill_1 FILLER_66_433 ();
 sg13g2_fill_1 FILLER_66_440 ();
 sg13g2_decap_4 FILLER_66_465 ();
 sg13g2_fill_2 FILLER_66_475 ();
 sg13g2_decap_8 FILLER_66_501 ();
 sg13g2_fill_2 FILLER_66_508 ();
 sg13g2_decap_8 FILLER_66_514 ();
 sg13g2_decap_8 FILLER_66_521 ();
 sg13g2_decap_4 FILLER_66_552 ();
 sg13g2_fill_2 FILLER_66_556 ();
 sg13g2_fill_2 FILLER_66_563 ();
 sg13g2_decap_8 FILLER_66_569 ();
 sg13g2_decap_4 FILLER_66_576 ();
 sg13g2_fill_1 FILLER_66_580 ();
 sg13g2_fill_2 FILLER_66_588 ();
 sg13g2_fill_1 FILLER_66_594 ();
 sg13g2_fill_1 FILLER_66_599 ();
 sg13g2_fill_1 FILLER_66_605 ();
 sg13g2_fill_1 FILLER_66_610 ();
 sg13g2_decap_8 FILLER_66_618 ();
 sg13g2_decap_8 FILLER_66_625 ();
 sg13g2_decap_4 FILLER_66_632 ();
 sg13g2_fill_1 FILLER_66_636 ();
 sg13g2_fill_1 FILLER_66_642 ();
 sg13g2_decap_8 FILLER_66_647 ();
 sg13g2_fill_2 FILLER_66_654 ();
 sg13g2_decap_8 FILLER_66_669 ();
 sg13g2_fill_2 FILLER_66_676 ();
 sg13g2_decap_8 FILLER_66_692 ();
 sg13g2_fill_2 FILLER_66_699 ();
 sg13g2_decap_8 FILLER_66_741 ();
 sg13g2_decap_8 FILLER_66_748 ();
 sg13g2_decap_4 FILLER_66_755 ();
 sg13g2_fill_1 FILLER_66_759 ();
 sg13g2_fill_1 FILLER_66_770 ();
 sg13g2_fill_1 FILLER_66_834 ();
 sg13g2_fill_2 FILLER_66_855 ();
 sg13g2_fill_1 FILLER_66_857 ();
 sg13g2_fill_2 FILLER_66_866 ();
 sg13g2_fill_1 FILLER_66_877 ();
 sg13g2_decap_8 FILLER_66_883 ();
 sg13g2_decap_8 FILLER_66_890 ();
 sg13g2_fill_1 FILLER_66_897 ();
 sg13g2_decap_4 FILLER_66_903 ();
 sg13g2_fill_2 FILLER_66_907 ();
 sg13g2_fill_2 FILLER_66_919 ();
 sg13g2_fill_1 FILLER_66_926 ();
 sg13g2_decap_4 FILLER_66_931 ();
 sg13g2_fill_1 FILLER_66_935 ();
 sg13g2_decap_8 FILLER_66_966 ();
 sg13g2_fill_2 FILLER_66_977 ();
 sg13g2_decap_4 FILLER_66_1009 ();
 sg13g2_fill_1 FILLER_66_1013 ();
 sg13g2_decap_4 FILLER_66_1044 ();
 sg13g2_fill_2 FILLER_66_1048 ();
 sg13g2_fill_2 FILLER_66_1054 ();
 sg13g2_fill_2 FILLER_66_1069 ();
 sg13g2_fill_1 FILLER_66_1071 ();
 sg13g2_decap_8 FILLER_66_1085 ();
 sg13g2_fill_2 FILLER_66_1092 ();
 sg13g2_fill_1 FILLER_66_1094 ();
 sg13g2_decap_4 FILLER_66_1130 ();
 sg13g2_decap_4 FILLER_66_1165 ();
 sg13g2_fill_2 FILLER_66_1169 ();
 sg13g2_decap_8 FILLER_66_1180 ();
 sg13g2_decap_4 FILLER_66_1187 ();
 sg13g2_fill_1 FILLER_66_1191 ();
 sg13g2_fill_1 FILLER_66_1196 ();
 sg13g2_decap_8 FILLER_66_1223 ();
 sg13g2_decap_8 FILLER_66_1230 ();
 sg13g2_decap_8 FILLER_66_1237 ();
 sg13g2_fill_2 FILLER_66_1244 ();
 sg13g2_fill_1 FILLER_66_1251 ();
 sg13g2_decap_8 FILLER_66_1261 ();
 sg13g2_fill_2 FILLER_66_1268 ();
 sg13g2_decap_8 FILLER_66_1300 ();
 sg13g2_fill_1 FILLER_66_1307 ();
 sg13g2_fill_2 FILLER_66_1318 ();
 sg13g2_fill_2 FILLER_66_1330 ();
 sg13g2_fill_1 FILLER_66_1332 ();
 sg13g2_fill_2 FILLER_66_1338 ();
 sg13g2_fill_1 FILLER_66_1340 ();
 sg13g2_decap_8 FILLER_66_1360 ();
 sg13g2_decap_8 FILLER_66_1367 ();
 sg13g2_decap_8 FILLER_66_1374 ();
 sg13g2_decap_8 FILLER_66_1381 ();
 sg13g2_fill_1 FILLER_66_1388 ();
 sg13g2_decap_8 FILLER_66_1393 ();
 sg13g2_fill_2 FILLER_66_1400 ();
 sg13g2_fill_1 FILLER_66_1402 ();
 sg13g2_fill_1 FILLER_66_1412 ();
 sg13g2_fill_1 FILLER_66_1418 ();
 sg13g2_fill_1 FILLER_66_1427 ();
 sg13g2_fill_2 FILLER_66_1438 ();
 sg13g2_fill_1 FILLER_66_1449 ();
 sg13g2_fill_1 FILLER_66_1480 ();
 sg13g2_fill_2 FILLER_66_1485 ();
 sg13g2_decap_4 FILLER_66_1496 ();
 sg13g2_fill_1 FILLER_66_1500 ();
 sg13g2_decap_8 FILLER_66_1506 ();
 sg13g2_fill_2 FILLER_66_1513 ();
 sg13g2_decap_8 FILLER_66_1519 ();
 sg13g2_decap_8 FILLER_66_1526 ();
 sg13g2_decap_4 FILLER_66_1533 ();
 sg13g2_fill_1 FILLER_66_1537 ();
 sg13g2_decap_4 FILLER_66_1605 ();
 sg13g2_fill_2 FILLER_66_1609 ();
 sg13g2_fill_2 FILLER_66_1621 ();
 sg13g2_decap_8 FILLER_66_1649 ();
 sg13g2_decap_8 FILLER_66_1656 ();
 sg13g2_decap_8 FILLER_66_1663 ();
 sg13g2_decap_8 FILLER_66_1670 ();
 sg13g2_decap_8 FILLER_66_1677 ();
 sg13g2_decap_8 FILLER_66_1684 ();
 sg13g2_decap_8 FILLER_66_1691 ();
 sg13g2_decap_8 FILLER_66_1698 ();
 sg13g2_decap_8 FILLER_66_1705 ();
 sg13g2_decap_8 FILLER_66_1712 ();
 sg13g2_decap_8 FILLER_66_1719 ();
 sg13g2_decap_8 FILLER_66_1726 ();
 sg13g2_decap_8 FILLER_66_1733 ();
 sg13g2_decap_8 FILLER_66_1740 ();
 sg13g2_decap_8 FILLER_66_1747 ();
 sg13g2_decap_8 FILLER_66_1754 ();
 sg13g2_decap_8 FILLER_66_1761 ();
 sg13g2_decap_4 FILLER_66_1768 ();
 sg13g2_fill_2 FILLER_66_1772 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_4 FILLER_67_28 ();
 sg13g2_fill_1 FILLER_67_32 ();
 sg13g2_decap_4 FILLER_67_72 ();
 sg13g2_decap_8 FILLER_67_85 ();
 sg13g2_decap_8 FILLER_67_92 ();
 sg13g2_decap_8 FILLER_67_99 ();
 sg13g2_fill_2 FILLER_67_106 ();
 sg13g2_fill_2 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_134 ();
 sg13g2_fill_1 FILLER_67_141 ();
 sg13g2_fill_1 FILLER_67_153 ();
 sg13g2_decap_8 FILLER_67_158 ();
 sg13g2_fill_1 FILLER_67_165 ();
 sg13g2_decap_4 FILLER_67_171 ();
 sg13g2_decap_8 FILLER_67_186 ();
 sg13g2_fill_1 FILLER_67_193 ();
 sg13g2_decap_4 FILLER_67_199 ();
 sg13g2_fill_1 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_216 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_decap_4 FILLER_67_237 ();
 sg13g2_fill_1 FILLER_67_241 ();
 sg13g2_decap_4 FILLER_67_249 ();
 sg13g2_decap_8 FILLER_67_265 ();
 sg13g2_decap_8 FILLER_67_272 ();
 sg13g2_fill_2 FILLER_67_294 ();
 sg13g2_fill_1 FILLER_67_296 ();
 sg13g2_decap_4 FILLER_67_302 ();
 sg13g2_fill_1 FILLER_67_314 ();
 sg13g2_decap_4 FILLER_67_331 ();
 sg13g2_decap_8 FILLER_67_352 ();
 sg13g2_decap_4 FILLER_67_359 ();
 sg13g2_fill_2 FILLER_67_363 ();
 sg13g2_decap_4 FILLER_67_381 ();
 sg13g2_fill_2 FILLER_67_394 ();
 sg13g2_fill_2 FILLER_67_400 ();
 sg13g2_decap_4 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_67_433 ();
 sg13g2_decap_4 FILLER_67_440 ();
 sg13g2_fill_2 FILLER_67_444 ();
 sg13g2_fill_1 FILLER_67_461 ();
 sg13g2_decap_8 FILLER_67_477 ();
 sg13g2_fill_1 FILLER_67_484 ();
 sg13g2_decap_4 FILLER_67_507 ();
 sg13g2_fill_2 FILLER_67_511 ();
 sg13g2_decap_8 FILLER_67_519 ();
 sg13g2_fill_2 FILLER_67_526 ();
 sg13g2_fill_1 FILLER_67_528 ();
 sg13g2_decap_4 FILLER_67_543 ();
 sg13g2_fill_1 FILLER_67_547 ();
 sg13g2_decap_4 FILLER_67_572 ();
 sg13g2_fill_1 FILLER_67_576 ();
 sg13g2_decap_8 FILLER_67_597 ();
 sg13g2_decap_8 FILLER_67_604 ();
 sg13g2_decap_8 FILLER_67_611 ();
 sg13g2_decap_8 FILLER_67_618 ();
 sg13g2_decap_8 FILLER_67_629 ();
 sg13g2_decap_8 FILLER_67_636 ();
 sg13g2_fill_2 FILLER_67_643 ();
 sg13g2_fill_1 FILLER_67_649 ();
 sg13g2_fill_2 FILLER_67_669 ();
 sg13g2_decap_4 FILLER_67_689 ();
 sg13g2_fill_1 FILLER_67_693 ();
 sg13g2_decap_4 FILLER_67_719 ();
 sg13g2_fill_2 FILLER_67_723 ();
 sg13g2_decap_8 FILLER_67_733 ();
 sg13g2_decap_8 FILLER_67_740 ();
 sg13g2_decap_4 FILLER_67_747 ();
 sg13g2_fill_1 FILLER_67_760 ();
 sg13g2_fill_2 FILLER_67_770 ();
 sg13g2_fill_2 FILLER_67_776 ();
 sg13g2_fill_1 FILLER_67_778 ();
 sg13g2_decap_8 FILLER_67_783 ();
 sg13g2_fill_2 FILLER_67_806 ();
 sg13g2_fill_1 FILLER_67_808 ();
 sg13g2_fill_2 FILLER_67_813 ();
 sg13g2_fill_1 FILLER_67_824 ();
 sg13g2_fill_1 FILLER_67_829 ();
 sg13g2_decap_8 FILLER_67_838 ();
 sg13g2_decap_8 FILLER_67_845 ();
 sg13g2_decap_4 FILLER_67_857 ();
 sg13g2_decap_4 FILLER_67_865 ();
 sg13g2_fill_2 FILLER_67_869 ();
 sg13g2_decap_8 FILLER_67_880 ();
 sg13g2_fill_2 FILLER_67_892 ();
 sg13g2_fill_1 FILLER_67_894 ();
 sg13g2_decap_4 FILLER_67_906 ();
 sg13g2_fill_2 FILLER_67_910 ();
 sg13g2_fill_2 FILLER_67_916 ();
 sg13g2_fill_1 FILLER_67_918 ();
 sg13g2_fill_2 FILLER_67_964 ();
 sg13g2_decap_8 FILLER_67_992 ();
 sg13g2_decap_8 FILLER_67_999 ();
 sg13g2_fill_2 FILLER_67_1006 ();
 sg13g2_fill_1 FILLER_67_1008 ();
 sg13g2_fill_1 FILLER_67_1018 ();
 sg13g2_decap_8 FILLER_67_1028 ();
 sg13g2_decap_4 FILLER_67_1035 ();
 sg13g2_fill_1 FILLER_67_1070 ();
 sg13g2_fill_1 FILLER_67_1101 ();
 sg13g2_decap_4 FILLER_67_1136 ();
 sg13g2_fill_1 FILLER_67_1140 ();
 sg13g2_fill_1 FILLER_67_1149 ();
 sg13g2_decap_8 FILLER_67_1154 ();
 sg13g2_decap_8 FILLER_67_1161 ();
 sg13g2_decap_4 FILLER_67_1199 ();
 sg13g2_decap_4 FILLER_67_1207 ();
 sg13g2_decap_8 FILLER_67_1216 ();
 sg13g2_decap_4 FILLER_67_1223 ();
 sg13g2_decap_8 FILLER_67_1252 ();
 sg13g2_decap_4 FILLER_67_1259 ();
 sg13g2_fill_1 FILLER_67_1263 ();
 sg13g2_decap_4 FILLER_67_1268 ();
 sg13g2_fill_2 FILLER_67_1272 ();
 sg13g2_fill_1 FILLER_67_1278 ();
 sg13g2_fill_1 FILLER_67_1303 ();
 sg13g2_decap_4 FILLER_67_1308 ();
 sg13g2_fill_1 FILLER_67_1312 ();
 sg13g2_fill_1 FILLER_67_1318 ();
 sg13g2_fill_2 FILLER_67_1339 ();
 sg13g2_fill_1 FILLER_67_1341 ();
 sg13g2_fill_1 FILLER_67_1357 ();
 sg13g2_decap_8 FILLER_67_1363 ();
 sg13g2_decap_8 FILLER_67_1370 ();
 sg13g2_decap_4 FILLER_67_1377 ();
 sg13g2_fill_1 FILLER_67_1381 ();
 sg13g2_decap_8 FILLER_67_1413 ();
 sg13g2_decap_8 FILLER_67_1420 ();
 sg13g2_fill_1 FILLER_67_1427 ();
 sg13g2_fill_1 FILLER_67_1433 ();
 sg13g2_decap_4 FILLER_67_1439 ();
 sg13g2_fill_1 FILLER_67_1452 ();
 sg13g2_fill_1 FILLER_67_1456 ();
 sg13g2_fill_1 FILLER_67_1466 ();
 sg13g2_fill_1 FILLER_67_1472 ();
 sg13g2_decap_8 FILLER_67_1508 ();
 sg13g2_decap_8 FILLER_67_1524 ();
 sg13g2_decap_8 FILLER_67_1531 ();
 sg13g2_decap_8 FILLER_67_1542 ();
 sg13g2_fill_2 FILLER_67_1549 ();
 sg13g2_fill_1 FILLER_67_1551 ();
 sg13g2_decap_8 FILLER_67_1556 ();
 sg13g2_decap_8 FILLER_67_1600 ();
 sg13g2_decap_8 FILLER_67_1607 ();
 sg13g2_decap_4 FILLER_67_1614 ();
 sg13g2_fill_1 FILLER_67_1618 ();
 sg13g2_decap_8 FILLER_67_1624 ();
 sg13g2_decap_8 FILLER_67_1631 ();
 sg13g2_decap_8 FILLER_67_1638 ();
 sg13g2_decap_8 FILLER_67_1645 ();
 sg13g2_decap_8 FILLER_67_1652 ();
 sg13g2_decap_8 FILLER_67_1659 ();
 sg13g2_decap_8 FILLER_67_1666 ();
 sg13g2_decap_8 FILLER_67_1673 ();
 sg13g2_decap_8 FILLER_67_1680 ();
 sg13g2_decap_8 FILLER_67_1687 ();
 sg13g2_decap_8 FILLER_67_1694 ();
 sg13g2_decap_8 FILLER_67_1701 ();
 sg13g2_decap_8 FILLER_67_1708 ();
 sg13g2_decap_8 FILLER_67_1715 ();
 sg13g2_decap_8 FILLER_67_1722 ();
 sg13g2_decap_8 FILLER_67_1729 ();
 sg13g2_decap_8 FILLER_67_1736 ();
 sg13g2_decap_8 FILLER_67_1743 ();
 sg13g2_decap_8 FILLER_67_1750 ();
 sg13g2_decap_8 FILLER_67_1757 ();
 sg13g2_decap_8 FILLER_67_1764 ();
 sg13g2_fill_2 FILLER_67_1771 ();
 sg13g2_fill_1 FILLER_67_1773 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_58 ();
 sg13g2_fill_1 FILLER_68_65 ();
 sg13g2_fill_1 FILLER_68_71 ();
 sg13g2_fill_2 FILLER_68_99 ();
 sg13g2_fill_1 FILLER_68_125 ();
 sg13g2_decap_4 FILLER_68_141 ();
 sg13g2_fill_2 FILLER_68_162 ();
 sg13g2_decap_4 FILLER_68_190 ();
 sg13g2_fill_2 FILLER_68_194 ();
 sg13g2_fill_2 FILLER_68_216 ();
 sg13g2_fill_2 FILLER_68_247 ();
 sg13g2_decap_8 FILLER_68_259 ();
 sg13g2_decap_8 FILLER_68_266 ();
 sg13g2_decap_8 FILLER_68_273 ();
 sg13g2_fill_1 FILLER_68_284 ();
 sg13g2_fill_2 FILLER_68_289 ();
 sg13g2_fill_1 FILLER_68_303 ();
 sg13g2_fill_2 FILLER_68_311 ();
 sg13g2_fill_2 FILLER_68_318 ();
 sg13g2_fill_1 FILLER_68_320 ();
 sg13g2_decap_8 FILLER_68_331 ();
 sg13g2_fill_1 FILLER_68_338 ();
 sg13g2_fill_2 FILLER_68_343 ();
 sg13g2_fill_1 FILLER_68_345 ();
 sg13g2_decap_8 FILLER_68_358 ();
 sg13g2_fill_1 FILLER_68_365 ();
 sg13g2_decap_4 FILLER_68_376 ();
 sg13g2_fill_1 FILLER_68_380 ();
 sg13g2_fill_1 FILLER_68_386 ();
 sg13g2_fill_2 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_68_402 ();
 sg13g2_decap_8 FILLER_68_409 ();
 sg13g2_fill_1 FILLER_68_416 ();
 sg13g2_decap_4 FILLER_68_433 ();
 sg13g2_fill_1 FILLER_68_437 ();
 sg13g2_decap_4 FILLER_68_443 ();
 sg13g2_decap_8 FILLER_68_455 ();
 sg13g2_decap_8 FILLER_68_462 ();
 sg13g2_decap_8 FILLER_68_469 ();
 sg13g2_fill_2 FILLER_68_476 ();
 sg13g2_fill_1 FILLER_68_478 ();
 sg13g2_fill_1 FILLER_68_483 ();
 sg13g2_decap_8 FILLER_68_505 ();
 sg13g2_decap_8 FILLER_68_512 ();
 sg13g2_decap_8 FILLER_68_519 ();
 sg13g2_fill_1 FILLER_68_526 ();
 sg13g2_decap_8 FILLER_68_546 ();
 sg13g2_decap_4 FILLER_68_553 ();
 sg13g2_fill_1 FILLER_68_557 ();
 sg13g2_fill_1 FILLER_68_563 ();
 sg13g2_fill_1 FILLER_68_576 ();
 sg13g2_fill_1 FILLER_68_584 ();
 sg13g2_fill_2 FILLER_68_593 ();
 sg13g2_fill_2 FILLER_68_632 ();
 sg13g2_decap_4 FILLER_68_641 ();
 sg13g2_fill_1 FILLER_68_645 ();
 sg13g2_fill_2 FILLER_68_650 ();
 sg13g2_fill_1 FILLER_68_652 ();
 sg13g2_fill_2 FILLER_68_668 ();
 sg13g2_fill_1 FILLER_68_670 ();
 sg13g2_decap_8 FILLER_68_675 ();
 sg13g2_decap_8 FILLER_68_682 ();
 sg13g2_fill_2 FILLER_68_689 ();
 sg13g2_decap_4 FILLER_68_695 ();
 sg13g2_fill_2 FILLER_68_699 ();
 sg13g2_fill_1 FILLER_68_711 ();
 sg13g2_decap_4 FILLER_68_748 ();
 sg13g2_fill_2 FILLER_68_752 ();
 sg13g2_decap_8 FILLER_68_759 ();
 sg13g2_fill_2 FILLER_68_770 ();
 sg13g2_decap_8 FILLER_68_777 ();
 sg13g2_decap_8 FILLER_68_784 ();
 sg13g2_fill_1 FILLER_68_791 ();
 sg13g2_fill_2 FILLER_68_811 ();
 sg13g2_fill_1 FILLER_68_813 ();
 sg13g2_decap_4 FILLER_68_856 ();
 sg13g2_fill_1 FILLER_68_860 ();
 sg13g2_decap_8 FILLER_68_871 ();
 sg13g2_decap_8 FILLER_68_878 ();
 sg13g2_decap_8 FILLER_68_885 ();
 sg13g2_fill_1 FILLER_68_892 ();
 sg13g2_fill_2 FILLER_68_900 ();
 sg13g2_fill_2 FILLER_68_933 ();
 sg13g2_fill_1 FILLER_68_935 ();
 sg13g2_fill_1 FILLER_68_943 ();
 sg13g2_decap_8 FILLER_68_995 ();
 sg13g2_decap_8 FILLER_68_1002 ();
 sg13g2_decap_4 FILLER_68_1009 ();
 sg13g2_fill_2 FILLER_68_1028 ();
 sg13g2_decap_4 FILLER_68_1038 ();
 sg13g2_fill_1 FILLER_68_1042 ();
 sg13g2_fill_2 FILLER_68_1056 ();
 sg13g2_decap_4 FILLER_68_1062 ();
 sg13g2_fill_2 FILLER_68_1066 ();
 sg13g2_decap_8 FILLER_68_1074 ();
 sg13g2_fill_2 FILLER_68_1081 ();
 sg13g2_decap_4 FILLER_68_1088 ();
 sg13g2_fill_1 FILLER_68_1092 ();
 sg13g2_fill_1 FILLER_68_1101 ();
 sg13g2_fill_1 FILLER_68_1109 ();
 sg13g2_fill_1 FILLER_68_1114 ();
 sg13g2_fill_1 FILLER_68_1120 ();
 sg13g2_decap_8 FILLER_68_1126 ();
 sg13g2_decap_8 FILLER_68_1137 ();
 sg13g2_fill_2 FILLER_68_1144 ();
 sg13g2_fill_1 FILLER_68_1146 ();
 sg13g2_fill_2 FILLER_68_1171 ();
 sg13g2_fill_1 FILLER_68_1177 ();
 sg13g2_fill_2 FILLER_68_1183 ();
 sg13g2_fill_1 FILLER_68_1185 ();
 sg13g2_decap_4 FILLER_68_1201 ();
 sg13g2_fill_2 FILLER_68_1205 ();
 sg13g2_fill_1 FILLER_68_1212 ();
 sg13g2_decap_4 FILLER_68_1218 ();
 sg13g2_decap_4 FILLER_68_1227 ();
 sg13g2_fill_1 FILLER_68_1231 ();
 sg13g2_decap_8 FILLER_68_1270 ();
 sg13g2_decap_8 FILLER_68_1277 ();
 sg13g2_decap_4 FILLER_68_1284 ();
 sg13g2_fill_1 FILLER_68_1288 ();
 sg13g2_decap_8 FILLER_68_1294 ();
 sg13g2_decap_8 FILLER_68_1321 ();
 sg13g2_fill_1 FILLER_68_1328 ();
 sg13g2_fill_1 FILLER_68_1344 ();
 sg13g2_decap_8 FILLER_68_1355 ();
 sg13g2_decap_8 FILLER_68_1362 ();
 sg13g2_decap_8 FILLER_68_1369 ();
 sg13g2_fill_2 FILLER_68_1376 ();
 sg13g2_fill_1 FILLER_68_1378 ();
 sg13g2_fill_1 FILLER_68_1405 ();
 sg13g2_fill_2 FILLER_68_1416 ();
 sg13g2_fill_1 FILLER_68_1418 ();
 sg13g2_decap_8 FILLER_68_1423 ();
 sg13g2_decap_8 FILLER_68_1430 ();
 sg13g2_fill_1 FILLER_68_1473 ();
 sg13g2_fill_1 FILLER_68_1507 ();
 sg13g2_decap_4 FILLER_68_1534 ();
 sg13g2_fill_2 FILLER_68_1538 ();
 sg13g2_decap_8 FILLER_68_1571 ();
 sg13g2_fill_1 FILLER_68_1578 ();
 sg13g2_decap_8 FILLER_68_1605 ();
 sg13g2_decap_8 FILLER_68_1612 ();
 sg13g2_decap_8 FILLER_68_1619 ();
 sg13g2_decap_8 FILLER_68_1626 ();
 sg13g2_decap_8 FILLER_68_1633 ();
 sg13g2_decap_8 FILLER_68_1640 ();
 sg13g2_decap_8 FILLER_68_1647 ();
 sg13g2_decap_8 FILLER_68_1654 ();
 sg13g2_decap_8 FILLER_68_1661 ();
 sg13g2_decap_8 FILLER_68_1668 ();
 sg13g2_decap_8 FILLER_68_1675 ();
 sg13g2_decap_8 FILLER_68_1682 ();
 sg13g2_decap_8 FILLER_68_1689 ();
 sg13g2_decap_8 FILLER_68_1696 ();
 sg13g2_decap_8 FILLER_68_1703 ();
 sg13g2_decap_8 FILLER_68_1710 ();
 sg13g2_decap_8 FILLER_68_1717 ();
 sg13g2_decap_8 FILLER_68_1724 ();
 sg13g2_decap_8 FILLER_68_1731 ();
 sg13g2_decap_8 FILLER_68_1738 ();
 sg13g2_decap_8 FILLER_68_1745 ();
 sg13g2_decap_8 FILLER_68_1752 ();
 sg13g2_decap_8 FILLER_68_1759 ();
 sg13g2_decap_8 FILLER_68_1766 ();
 sg13g2_fill_1 FILLER_68_1773 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_11 ();
 sg13g2_decap_8 FILLER_69_16 ();
 sg13g2_decap_8 FILLER_69_23 ();
 sg13g2_decap_8 FILLER_69_30 ();
 sg13g2_decap_8 FILLER_69_37 ();
 sg13g2_fill_1 FILLER_69_44 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_fill_2 FILLER_69_70 ();
 sg13g2_fill_1 FILLER_69_72 ();
 sg13g2_decap_8 FILLER_69_83 ();
 sg13g2_decap_8 FILLER_69_90 ();
 sg13g2_decap_4 FILLER_69_97 ();
 sg13g2_decap_8 FILLER_69_137 ();
 sg13g2_decap_8 FILLER_69_144 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_fill_1 FILLER_69_157 ();
 sg13g2_fill_1 FILLER_69_162 ();
 sg13g2_decap_4 FILLER_69_168 ();
 sg13g2_fill_2 FILLER_69_172 ();
 sg13g2_fill_2 FILLER_69_186 ();
 sg13g2_decap_8 FILLER_69_192 ();
 sg13g2_decap_4 FILLER_69_199 ();
 sg13g2_fill_1 FILLER_69_203 ();
 sg13g2_decap_4 FILLER_69_212 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_fill_2 FILLER_69_263 ();
 sg13g2_fill_2 FILLER_69_270 ();
 sg13g2_fill_1 FILLER_69_272 ();
 sg13g2_fill_1 FILLER_69_281 ();
 sg13g2_decap_8 FILLER_69_286 ();
 sg13g2_fill_1 FILLER_69_293 ();
 sg13g2_decap_8 FILLER_69_306 ();
 sg13g2_fill_2 FILLER_69_313 ();
 sg13g2_decap_8 FILLER_69_333 ();
 sg13g2_fill_2 FILLER_69_340 ();
 sg13g2_fill_1 FILLER_69_342 ();
 sg13g2_fill_2 FILLER_69_377 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_decap_4 FILLER_69_391 ();
 sg13g2_fill_2 FILLER_69_395 ();
 sg13g2_fill_2 FILLER_69_402 ();
 sg13g2_decap_8 FILLER_69_409 ();
 sg13g2_decap_4 FILLER_69_416 ();
 sg13g2_fill_2 FILLER_69_420 ();
 sg13g2_decap_8 FILLER_69_431 ();
 sg13g2_fill_1 FILLER_69_438 ();
 sg13g2_fill_1 FILLER_69_449 ();
 sg13g2_decap_8 FILLER_69_458 ();
 sg13g2_fill_2 FILLER_69_465 ();
 sg13g2_fill_1 FILLER_69_467 ();
 sg13g2_decap_4 FILLER_69_472 ();
 sg13g2_fill_1 FILLER_69_476 ();
 sg13g2_decap_8 FILLER_69_481 ();
 sg13g2_fill_2 FILLER_69_488 ();
 sg13g2_fill_1 FILLER_69_490 ();
 sg13g2_decap_4 FILLER_69_509 ();
 sg13g2_decap_8 FILLER_69_517 ();
 sg13g2_fill_2 FILLER_69_524 ();
 sg13g2_fill_1 FILLER_69_526 ();
 sg13g2_decap_8 FILLER_69_542 ();
 sg13g2_fill_2 FILLER_69_549 ();
 sg13g2_fill_2 FILLER_69_573 ();
 sg13g2_fill_1 FILLER_69_575 ();
 sg13g2_decap_8 FILLER_69_588 ();
 sg13g2_decap_8 FILLER_69_595 ();
 sg13g2_decap_8 FILLER_69_602 ();
 sg13g2_fill_2 FILLER_69_609 ();
 sg13g2_fill_2 FILLER_69_643 ();
 sg13g2_decap_8 FILLER_69_660 ();
 sg13g2_fill_2 FILLER_69_667 ();
 sg13g2_decap_4 FILLER_69_673 ();
 sg13g2_fill_2 FILLER_69_712 ();
 sg13g2_decap_8 FILLER_69_718 ();
 sg13g2_decap_8 FILLER_69_725 ();
 sg13g2_decap_8 FILLER_69_748 ();
 sg13g2_decap_8 FILLER_69_755 ();
 sg13g2_decap_8 FILLER_69_762 ();
 sg13g2_decap_4 FILLER_69_799 ();
 sg13g2_fill_1 FILLER_69_803 ();
 sg13g2_decap_8 FILLER_69_821 ();
 sg13g2_decap_8 FILLER_69_828 ();
 sg13g2_decap_8 FILLER_69_835 ();
 sg13g2_fill_1 FILLER_69_842 ();
 sg13g2_fill_1 FILLER_69_852 ();
 sg13g2_fill_2 FILLER_69_863 ();
 sg13g2_fill_1 FILLER_69_865 ();
 sg13g2_fill_1 FILLER_69_870 ();
 sg13g2_decap_4 FILLER_69_897 ();
 sg13g2_fill_2 FILLER_69_905 ();
 sg13g2_fill_1 FILLER_69_907 ();
 sg13g2_fill_1 FILLER_69_913 ();
 sg13g2_decap_8 FILLER_69_918 ();
 sg13g2_fill_2 FILLER_69_925 ();
 sg13g2_decap_4 FILLER_69_931 ();
 sg13g2_fill_2 FILLER_69_935 ();
 sg13g2_decap_8 FILLER_69_941 ();
 sg13g2_fill_1 FILLER_69_948 ();
 sg13g2_decap_4 FILLER_69_959 ();
 sg13g2_fill_1 FILLER_69_963 ();
 sg13g2_fill_1 FILLER_69_969 ();
 sg13g2_fill_2 FILLER_69_974 ();
 sg13g2_fill_2 FILLER_69_980 ();
 sg13g2_fill_2 FILLER_69_1008 ();
 sg13g2_fill_1 FILLER_69_1010 ();
 sg13g2_decap_8 FILLER_69_1015 ();
 sg13g2_fill_2 FILLER_69_1022 ();
 sg13g2_fill_1 FILLER_69_1028 ();
 sg13g2_fill_2 FILLER_69_1034 ();
 sg13g2_decap_8 FILLER_69_1041 ();
 sg13g2_decap_8 FILLER_69_1048 ();
 sg13g2_decap_4 FILLER_69_1055 ();
 sg13g2_fill_2 FILLER_69_1059 ();
 sg13g2_decap_8 FILLER_69_1065 ();
 sg13g2_fill_1 FILLER_69_1072 ();
 sg13g2_fill_2 FILLER_69_1085 ();
 sg13g2_fill_2 FILLER_69_1095 ();
 sg13g2_fill_1 FILLER_69_1097 ();
 sg13g2_decap_8 FILLER_69_1102 ();
 sg13g2_decap_4 FILLER_69_1109 ();
 sg13g2_fill_1 FILLER_69_1113 ();
 sg13g2_decap_8 FILLER_69_1119 ();
 sg13g2_decap_8 FILLER_69_1126 ();
 sg13g2_decap_4 FILLER_69_1133 ();
 sg13g2_fill_2 FILLER_69_1137 ();
 sg13g2_decap_8 FILLER_69_1144 ();
 sg13g2_fill_1 FILLER_69_1151 ();
 sg13g2_fill_2 FILLER_69_1176 ();
 sg13g2_fill_1 FILLER_69_1187 ();
 sg13g2_fill_1 FILLER_69_1203 ();
 sg13g2_fill_2 FILLER_69_1214 ();
 sg13g2_fill_1 FILLER_69_1216 ();
 sg13g2_fill_2 FILLER_69_1230 ();
 sg13g2_fill_2 FILLER_69_1237 ();
 sg13g2_fill_1 FILLER_69_1263 ();
 sg13g2_decap_4 FILLER_69_1282 ();
 sg13g2_fill_1 FILLER_69_1286 ();
 sg13g2_fill_2 FILLER_69_1300 ();
 sg13g2_fill_2 FILLER_69_1332 ();
 sg13g2_decap_8 FILLER_69_1338 ();
 sg13g2_decap_4 FILLER_69_1345 ();
 sg13g2_fill_1 FILLER_69_1383 ();
 sg13g2_decap_4 FILLER_69_1388 ();
 sg13g2_fill_1 FILLER_69_1392 ();
 sg13g2_decap_8 FILLER_69_1420 ();
 sg13g2_fill_2 FILLER_69_1435 ();
 sg13g2_fill_1 FILLER_69_1452 ();
 sg13g2_fill_1 FILLER_69_1471 ();
 sg13g2_fill_1 FILLER_69_1502 ();
 sg13g2_decap_4 FILLER_69_1508 ();
 sg13g2_decap_4 FILLER_69_1524 ();
 sg13g2_fill_2 FILLER_69_1528 ();
 sg13g2_fill_1 FILLER_69_1535 ();
 sg13g2_fill_2 FILLER_69_1543 ();
 sg13g2_fill_1 FILLER_69_1551 ();
 sg13g2_fill_2 FILLER_69_1560 ();
 sg13g2_decap_4 FILLER_69_1567 ();
 sg13g2_decap_4 FILLER_69_1585 ();
 sg13g2_fill_1 FILLER_69_1589 ();
 sg13g2_decap_8 FILLER_69_1594 ();
 sg13g2_decap_8 FILLER_69_1601 ();
 sg13g2_decap_8 FILLER_69_1608 ();
 sg13g2_decap_8 FILLER_69_1615 ();
 sg13g2_decap_8 FILLER_69_1622 ();
 sg13g2_decap_8 FILLER_69_1629 ();
 sg13g2_decap_8 FILLER_69_1636 ();
 sg13g2_decap_8 FILLER_69_1643 ();
 sg13g2_decap_8 FILLER_69_1650 ();
 sg13g2_decap_8 FILLER_69_1657 ();
 sg13g2_decap_8 FILLER_69_1664 ();
 sg13g2_decap_8 FILLER_69_1671 ();
 sg13g2_decap_8 FILLER_69_1678 ();
 sg13g2_decap_8 FILLER_69_1685 ();
 sg13g2_decap_8 FILLER_69_1692 ();
 sg13g2_decap_8 FILLER_69_1699 ();
 sg13g2_decap_8 FILLER_69_1706 ();
 sg13g2_decap_8 FILLER_69_1713 ();
 sg13g2_decap_8 FILLER_69_1720 ();
 sg13g2_decap_8 FILLER_69_1727 ();
 sg13g2_decap_8 FILLER_69_1734 ();
 sg13g2_decap_8 FILLER_69_1741 ();
 sg13g2_decap_8 FILLER_69_1748 ();
 sg13g2_decap_8 FILLER_69_1755 ();
 sg13g2_decap_8 FILLER_69_1762 ();
 sg13g2_decap_4 FILLER_69_1769 ();
 sg13g2_fill_1 FILLER_69_1773 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_4 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_42 ();
 sg13g2_fill_1 FILLER_70_57 ();
 sg13g2_decap_8 FILLER_70_66 ();
 sg13g2_fill_2 FILLER_70_77 ();
 sg13g2_fill_1 FILLER_70_79 ();
 sg13g2_decap_8 FILLER_70_90 ();
 sg13g2_fill_1 FILLER_70_97 ();
 sg13g2_decap_8 FILLER_70_108 ();
 sg13g2_decap_4 FILLER_70_115 ();
 sg13g2_fill_2 FILLER_70_119 ();
 sg13g2_decap_4 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_132 ();
 sg13g2_decap_8 FILLER_70_143 ();
 sg13g2_decap_4 FILLER_70_150 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_169 ();
 sg13g2_fill_2 FILLER_70_176 ();
 sg13g2_fill_1 FILLER_70_178 ();
 sg13g2_fill_1 FILLER_70_201 ();
 sg13g2_decap_4 FILLER_70_210 ();
 sg13g2_fill_2 FILLER_70_221 ();
 sg13g2_decap_8 FILLER_70_233 ();
 sg13g2_decap_4 FILLER_70_240 ();
 sg13g2_decap_8 FILLER_70_257 ();
 sg13g2_decap_4 FILLER_70_264 ();
 sg13g2_fill_2 FILLER_70_268 ();
 sg13g2_fill_2 FILLER_70_292 ();
 sg13g2_fill_1 FILLER_70_299 ();
 sg13g2_decap_4 FILLER_70_308 ();
 sg13g2_decap_8 FILLER_70_333 ();
 sg13g2_decap_4 FILLER_70_360 ();
 sg13g2_fill_2 FILLER_70_364 ();
 sg13g2_decap_4 FILLER_70_381 ();
 sg13g2_decap_8 FILLER_70_390 ();
 sg13g2_fill_2 FILLER_70_397 ();
 sg13g2_decap_8 FILLER_70_414 ();
 sg13g2_decap_8 FILLER_70_421 ();
 sg13g2_fill_2 FILLER_70_428 ();
 sg13g2_fill_2 FILLER_70_439 ();
 sg13g2_decap_4 FILLER_70_446 ();
 sg13g2_decap_4 FILLER_70_466 ();
 sg13g2_fill_1 FILLER_70_470 ();
 sg13g2_decap_8 FILLER_70_479 ();
 sg13g2_decap_8 FILLER_70_486 ();
 sg13g2_decap_8 FILLER_70_493 ();
 sg13g2_decap_4 FILLER_70_512 ();
 sg13g2_fill_1 FILLER_70_516 ();
 sg13g2_fill_2 FILLER_70_533 ();
 sg13g2_fill_1 FILLER_70_535 ();
 sg13g2_fill_2 FILLER_70_541 ();
 sg13g2_fill_2 FILLER_70_547 ();
 sg13g2_fill_1 FILLER_70_549 ();
 sg13g2_decap_4 FILLER_70_559 ();
 sg13g2_fill_1 FILLER_70_563 ();
 sg13g2_decap_8 FILLER_70_574 ();
 sg13g2_decap_8 FILLER_70_581 ();
 sg13g2_decap_8 FILLER_70_588 ();
 sg13g2_decap_4 FILLER_70_595 ();
 sg13g2_decap_8 FILLER_70_607 ();
 sg13g2_decap_4 FILLER_70_614 ();
 sg13g2_decap_4 FILLER_70_625 ();
 sg13g2_fill_2 FILLER_70_629 ();
 sg13g2_decap_8 FILLER_70_646 ();
 sg13g2_fill_2 FILLER_70_653 ();
 sg13g2_fill_1 FILLER_70_655 ();
 sg13g2_fill_2 FILLER_70_669 ();
 sg13g2_fill_1 FILLER_70_676 ();
 sg13g2_fill_2 FILLER_70_681 ();
 sg13g2_decap_4 FILLER_70_687 ();
 sg13g2_decap_8 FILLER_70_695 ();
 sg13g2_decap_4 FILLER_70_702 ();
 sg13g2_fill_2 FILLER_70_706 ();
 sg13g2_decap_4 FILLER_70_789 ();
 sg13g2_fill_1 FILLER_70_793 ();
 sg13g2_fill_2 FILLER_70_798 ();
 sg13g2_fill_2 FILLER_70_838 ();
 sg13g2_fill_1 FILLER_70_840 ();
 sg13g2_decap_4 FILLER_70_846 ();
 sg13g2_fill_1 FILLER_70_850 ();
 sg13g2_fill_2 FILLER_70_855 ();
 sg13g2_fill_1 FILLER_70_857 ();
 sg13g2_fill_2 FILLER_70_862 ();
 sg13g2_fill_1 FILLER_70_864 ();
 sg13g2_fill_1 FILLER_70_870 ();
 sg13g2_fill_2 FILLER_70_875 ();
 sg13g2_fill_1 FILLER_70_877 ();
 sg13g2_decap_8 FILLER_70_882 ();
 sg13g2_decap_8 FILLER_70_889 ();
 sg13g2_decap_8 FILLER_70_931 ();
 sg13g2_fill_1 FILLER_70_938 ();
 sg13g2_decap_4 FILLER_70_944 ();
 sg13g2_fill_1 FILLER_70_948 ();
 sg13g2_decap_8 FILLER_70_953 ();
 sg13g2_decap_4 FILLER_70_960 ();
 sg13g2_fill_1 FILLER_70_964 ();
 sg13g2_decap_8 FILLER_70_995 ();
 sg13g2_decap_8 FILLER_70_1002 ();
 sg13g2_fill_1 FILLER_70_1009 ();
 sg13g2_fill_2 FILLER_70_1025 ();
 sg13g2_fill_1 FILLER_70_1027 ();
 sg13g2_fill_1 FILLER_70_1033 ();
 sg13g2_fill_2 FILLER_70_1064 ();
 sg13g2_fill_1 FILLER_70_1066 ();
 sg13g2_fill_1 FILLER_70_1073 ();
 sg13g2_fill_1 FILLER_70_1110 ();
 sg13g2_fill_1 FILLER_70_1115 ();
 sg13g2_fill_1 FILLER_70_1121 ();
 sg13g2_fill_2 FILLER_70_1127 ();
 sg13g2_decap_4 FILLER_70_1134 ();
 sg13g2_fill_1 FILLER_70_1189 ();
 sg13g2_decap_8 FILLER_70_1195 ();
 sg13g2_decap_8 FILLER_70_1202 ();
 sg13g2_fill_2 FILLER_70_1209 ();
 sg13g2_decap_4 FILLER_70_1215 ();
 sg13g2_fill_2 FILLER_70_1219 ();
 sg13g2_decap_8 FILLER_70_1235 ();
 sg13g2_decap_4 FILLER_70_1242 ();
 sg13g2_fill_2 FILLER_70_1264 ();
 sg13g2_fill_1 FILLER_70_1266 ();
 sg13g2_fill_2 FILLER_70_1271 ();
 sg13g2_decap_4 FILLER_70_1278 ();
 sg13g2_fill_2 FILLER_70_1282 ();
 sg13g2_decap_8 FILLER_70_1292 ();
 sg13g2_decap_8 FILLER_70_1299 ();
 sg13g2_decap_4 FILLER_70_1306 ();
 sg13g2_decap_8 FILLER_70_1314 ();
 sg13g2_decap_4 FILLER_70_1321 ();
 sg13g2_fill_2 FILLER_70_1325 ();
 sg13g2_decap_4 FILLER_70_1353 ();
 sg13g2_fill_2 FILLER_70_1357 ();
 sg13g2_decap_4 FILLER_70_1363 ();
 sg13g2_fill_1 FILLER_70_1367 ();
 sg13g2_decap_4 FILLER_70_1372 ();
 sg13g2_fill_2 FILLER_70_1376 ();
 sg13g2_decap_8 FILLER_70_1382 ();
 sg13g2_decap_4 FILLER_70_1389 ();
 sg13g2_fill_2 FILLER_70_1450 ();
 sg13g2_fill_2 FILLER_70_1457 ();
 sg13g2_fill_2 FILLER_70_1468 ();
 sg13g2_fill_1 FILLER_70_1485 ();
 sg13g2_decap_4 FILLER_70_1494 ();
 sg13g2_fill_1 FILLER_70_1506 ();
 sg13g2_fill_2 FILLER_70_1512 ();
 sg13g2_fill_2 FILLER_70_1553 ();
 sg13g2_fill_1 FILLER_70_1555 ();
 sg13g2_decap_4 FILLER_70_1560 ();
 sg13g2_fill_1 FILLER_70_1564 ();
 sg13g2_decap_4 FILLER_70_1569 ();
 sg13g2_fill_1 FILLER_70_1573 ();
 sg13g2_decap_4 FILLER_70_1579 ();
 sg13g2_decap_8 FILLER_70_1609 ();
 sg13g2_decap_8 FILLER_70_1616 ();
 sg13g2_decap_8 FILLER_70_1623 ();
 sg13g2_decap_8 FILLER_70_1630 ();
 sg13g2_decap_8 FILLER_70_1637 ();
 sg13g2_decap_8 FILLER_70_1644 ();
 sg13g2_decap_8 FILLER_70_1651 ();
 sg13g2_decap_8 FILLER_70_1658 ();
 sg13g2_decap_8 FILLER_70_1665 ();
 sg13g2_decap_8 FILLER_70_1672 ();
 sg13g2_decap_8 FILLER_70_1679 ();
 sg13g2_decap_8 FILLER_70_1686 ();
 sg13g2_decap_8 FILLER_70_1693 ();
 sg13g2_decap_8 FILLER_70_1700 ();
 sg13g2_decap_8 FILLER_70_1707 ();
 sg13g2_decap_8 FILLER_70_1714 ();
 sg13g2_decap_8 FILLER_70_1721 ();
 sg13g2_decap_8 FILLER_70_1728 ();
 sg13g2_decap_8 FILLER_70_1735 ();
 sg13g2_decap_8 FILLER_70_1742 ();
 sg13g2_decap_8 FILLER_70_1749 ();
 sg13g2_decap_8 FILLER_70_1756 ();
 sg13g2_decap_8 FILLER_70_1763 ();
 sg13g2_decap_4 FILLER_70_1770 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_4 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_46 ();
 sg13g2_decap_8 FILLER_71_52 ();
 sg13g2_decap_8 FILLER_71_59 ();
 sg13g2_decap_8 FILLER_71_66 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_4 FILLER_71_98 ();
 sg13g2_fill_2 FILLER_71_107 ();
 sg13g2_fill_1 FILLER_71_128 ();
 sg13g2_decap_8 FILLER_71_144 ();
 sg13g2_fill_2 FILLER_71_151 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_fill_2 FILLER_71_189 ();
 sg13g2_fill_1 FILLER_71_191 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_208 ();
 sg13g2_fill_2 FILLER_71_215 ();
 sg13g2_fill_2 FILLER_71_263 ();
 sg13g2_decap_8 FILLER_71_291 ();
 sg13g2_fill_1 FILLER_71_298 ();
 sg13g2_fill_2 FILLER_71_304 ();
 sg13g2_decap_8 FILLER_71_314 ();
 sg13g2_decap_8 FILLER_71_321 ();
 sg13g2_decap_4 FILLER_71_328 ();
 sg13g2_fill_1 FILLER_71_341 ();
 sg13g2_fill_2 FILLER_71_346 ();
 sg13g2_fill_1 FILLER_71_348 ();
 sg13g2_decap_8 FILLER_71_360 ();
 sg13g2_decap_8 FILLER_71_393 ();
 sg13g2_fill_1 FILLER_71_400 ();
 sg13g2_decap_4 FILLER_71_415 ();
 sg13g2_fill_1 FILLER_71_419 ();
 sg13g2_fill_2 FILLER_71_439 ();
 sg13g2_fill_1 FILLER_71_448 ();
 sg13g2_fill_2 FILLER_71_454 ();
 sg13g2_decap_8 FILLER_71_460 ();
 sg13g2_fill_2 FILLER_71_467 ();
 sg13g2_fill_1 FILLER_71_469 ();
 sg13g2_fill_2 FILLER_71_475 ();
 sg13g2_fill_1 FILLER_71_477 ();
 sg13g2_fill_2 FILLER_71_483 ();
 sg13g2_fill_1 FILLER_71_485 ();
 sg13g2_decap_4 FILLER_71_492 ();
 sg13g2_fill_1 FILLER_71_496 ();
 sg13g2_fill_2 FILLER_71_512 ();
 sg13g2_decap_8 FILLER_71_535 ();
 sg13g2_fill_2 FILLER_71_542 ();
 sg13g2_fill_1 FILLER_71_544 ();
 sg13g2_fill_1 FILLER_71_549 ();
 sg13g2_fill_1 FILLER_71_554 ();
 sg13g2_fill_1 FILLER_71_562 ();
 sg13g2_fill_1 FILLER_71_568 ();
 sg13g2_fill_1 FILLER_71_579 ();
 sg13g2_fill_1 FILLER_71_585 ();
 sg13g2_decap_4 FILLER_71_596 ();
 sg13g2_fill_2 FILLER_71_620 ();
 sg13g2_decap_4 FILLER_71_641 ();
 sg13g2_fill_1 FILLER_71_645 ();
 sg13g2_decap_8 FILLER_71_706 ();
 sg13g2_decap_8 FILLER_71_713 ();
 sg13g2_decap_4 FILLER_71_720 ();
 sg13g2_decap_8 FILLER_71_728 ();
 sg13g2_decap_4 FILLER_71_735 ();
 sg13g2_fill_1 FILLER_71_739 ();
 sg13g2_decap_8 FILLER_71_745 ();
 sg13g2_fill_2 FILLER_71_752 ();
 sg13g2_fill_1 FILLER_71_754 ();
 sg13g2_fill_1 FILLER_71_759 ();
 sg13g2_fill_1 FILLER_71_783 ();
 sg13g2_fill_2 FILLER_71_788 ();
 sg13g2_fill_2 FILLER_71_794 ();
 sg13g2_fill_1 FILLER_71_796 ();
 sg13g2_fill_1 FILLER_71_802 ();
 sg13g2_fill_2 FILLER_71_816 ();
 sg13g2_decap_4 FILLER_71_822 ();
 sg13g2_fill_1 FILLER_71_826 ();
 sg13g2_decap_4 FILLER_71_832 ();
 sg13g2_fill_2 FILLER_71_836 ();
 sg13g2_fill_1 FILLER_71_869 ();
 sg13g2_fill_1 FILLER_71_874 ();
 sg13g2_fill_1 FILLER_71_880 ();
 sg13g2_fill_1 FILLER_71_886 ();
 sg13g2_fill_1 FILLER_71_896 ();
 sg13g2_decap_8 FILLER_71_905 ();
 sg13g2_decap_4 FILLER_71_912 ();
 sg13g2_decap_8 FILLER_71_920 ();
 sg13g2_fill_1 FILLER_71_927 ();
 sg13g2_decap_4 FILLER_71_932 ();
 sg13g2_fill_1 FILLER_71_936 ();
 sg13g2_fill_2 FILLER_71_966 ();
 sg13g2_decap_8 FILLER_71_985 ();
 sg13g2_decap_8 FILLER_71_992 ();
 sg13g2_fill_1 FILLER_71_999 ();
 sg13g2_decap_8 FILLER_71_1005 ();
 sg13g2_decap_8 FILLER_71_1012 ();
 sg13g2_decap_4 FILLER_71_1019 ();
 sg13g2_fill_1 FILLER_71_1023 ();
 sg13g2_decap_4 FILLER_71_1036 ();
 sg13g2_fill_1 FILLER_71_1044 ();
 sg13g2_fill_2 FILLER_71_1053 ();
 sg13g2_fill_1 FILLER_71_1055 ();
 sg13g2_decap_8 FILLER_71_1069 ();
 sg13g2_decap_4 FILLER_71_1076 ();
 sg13g2_decap_4 FILLER_71_1084 ();
 sg13g2_fill_2 FILLER_71_1088 ();
 sg13g2_decap_8 FILLER_71_1097 ();
 sg13g2_decap_8 FILLER_71_1104 ();
 sg13g2_decap_4 FILLER_71_1111 ();
 sg13g2_decap_4 FILLER_71_1120 ();
 sg13g2_fill_2 FILLER_71_1129 ();
 sg13g2_fill_1 FILLER_71_1131 ();
 sg13g2_decap_8 FILLER_71_1137 ();
 sg13g2_decap_4 FILLER_71_1144 ();
 sg13g2_fill_2 FILLER_71_1148 ();
 sg13g2_fill_2 FILLER_71_1158 ();
 sg13g2_fill_1 FILLER_71_1164 ();
 sg13g2_fill_2 FILLER_71_1174 ();
 sg13g2_fill_1 FILLER_71_1176 ();
 sg13g2_decap_4 FILLER_71_1187 ();
 sg13g2_fill_1 FILLER_71_1191 ();
 sg13g2_decap_8 FILLER_71_1196 ();
 sg13g2_fill_1 FILLER_71_1203 ();
 sg13g2_decap_4 FILLER_71_1208 ();
 sg13g2_fill_1 FILLER_71_1225 ();
 sg13g2_decap_8 FILLER_71_1244 ();
 sg13g2_decap_8 FILLER_71_1251 ();
 sg13g2_fill_2 FILLER_71_1267 ();
 sg13g2_fill_1 FILLER_71_1279 ();
 sg13g2_fill_1 FILLER_71_1284 ();
 sg13g2_fill_1 FILLER_71_1290 ();
 sg13g2_fill_1 FILLER_71_1295 ();
 sg13g2_decap_4 FILLER_71_1300 ();
 sg13g2_fill_2 FILLER_71_1304 ();
 sg13g2_decap_4 FILLER_71_1315 ();
 sg13g2_fill_1 FILLER_71_1319 ();
 sg13g2_decap_8 FILLER_71_1324 ();
 sg13g2_decap_8 FILLER_71_1331 ();
 sg13g2_fill_2 FILLER_71_1342 ();
 sg13g2_fill_1 FILLER_71_1344 ();
 sg13g2_decap_4 FILLER_71_1353 ();
 sg13g2_fill_1 FILLER_71_1357 ();
 sg13g2_fill_1 FILLER_71_1399 ();
 sg13g2_fill_1 FILLER_71_1416 ();
 sg13g2_fill_2 FILLER_71_1454 ();
 sg13g2_decap_4 FILLER_71_1473 ();
 sg13g2_fill_2 FILLER_71_1477 ();
 sg13g2_decap_8 FILLER_71_1505 ();
 sg13g2_decap_8 FILLER_71_1512 ();
 sg13g2_fill_2 FILLER_71_1519 ();
 sg13g2_fill_1 FILLER_71_1525 ();
 sg13g2_decap_8 FILLER_71_1530 ();
 sg13g2_decap_8 FILLER_71_1545 ();
 sg13g2_fill_1 FILLER_71_1552 ();
 sg13g2_decap_8 FILLER_71_1557 ();
 sg13g2_fill_1 FILLER_71_1564 ();
 sg13g2_fill_2 FILLER_71_1594 ();
 sg13g2_decap_8 FILLER_71_1600 ();
 sg13g2_decap_8 FILLER_71_1607 ();
 sg13g2_decap_8 FILLER_71_1614 ();
 sg13g2_decap_8 FILLER_71_1621 ();
 sg13g2_decap_8 FILLER_71_1628 ();
 sg13g2_decap_8 FILLER_71_1635 ();
 sg13g2_decap_8 FILLER_71_1642 ();
 sg13g2_decap_8 FILLER_71_1649 ();
 sg13g2_decap_8 FILLER_71_1656 ();
 sg13g2_decap_8 FILLER_71_1663 ();
 sg13g2_decap_8 FILLER_71_1670 ();
 sg13g2_decap_8 FILLER_71_1677 ();
 sg13g2_decap_8 FILLER_71_1684 ();
 sg13g2_decap_8 FILLER_71_1691 ();
 sg13g2_decap_8 FILLER_71_1698 ();
 sg13g2_decap_8 FILLER_71_1705 ();
 sg13g2_decap_8 FILLER_71_1712 ();
 sg13g2_decap_8 FILLER_71_1719 ();
 sg13g2_decap_8 FILLER_71_1726 ();
 sg13g2_decap_8 FILLER_71_1733 ();
 sg13g2_decap_8 FILLER_71_1740 ();
 sg13g2_decap_8 FILLER_71_1747 ();
 sg13g2_decap_8 FILLER_71_1754 ();
 sg13g2_decap_8 FILLER_71_1761 ();
 sg13g2_decap_4 FILLER_71_1768 ();
 sg13g2_fill_2 FILLER_71_1772 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_11 ();
 sg13g2_decap_8 FILLER_72_17 ();
 sg13g2_fill_2 FILLER_72_24 ();
 sg13g2_fill_1 FILLER_72_26 ();
 sg13g2_fill_1 FILLER_72_40 ();
 sg13g2_fill_2 FILLER_72_50 ();
 sg13g2_fill_1 FILLER_72_52 ();
 sg13g2_decap_8 FILLER_72_58 ();
 sg13g2_fill_2 FILLER_72_65 ();
 sg13g2_decap_4 FILLER_72_72 ();
 sg13g2_fill_2 FILLER_72_76 ();
 sg13g2_decap_4 FILLER_72_86 ();
 sg13g2_fill_1 FILLER_72_94 ();
 sg13g2_fill_1 FILLER_72_99 ();
 sg13g2_decap_8 FILLER_72_106 ();
 sg13g2_decap_4 FILLER_72_113 ();
 sg13g2_fill_2 FILLER_72_154 ();
 sg13g2_fill_1 FILLER_72_156 ();
 sg13g2_fill_2 FILLER_72_175 ();
 sg13g2_fill_2 FILLER_72_182 ();
 sg13g2_fill_1 FILLER_72_213 ();
 sg13g2_decap_4 FILLER_72_217 ();
 sg13g2_fill_1 FILLER_72_221 ();
 sg13g2_decap_4 FILLER_72_227 ();
 sg13g2_decap_8 FILLER_72_236 ();
 sg13g2_decap_8 FILLER_72_253 ();
 sg13g2_decap_8 FILLER_72_265 ();
 sg13g2_decap_8 FILLER_72_272 ();
 sg13g2_decap_8 FILLER_72_279 ();
 sg13g2_decap_8 FILLER_72_286 ();
 sg13g2_fill_2 FILLER_72_305 ();
 sg13g2_decap_4 FILLER_72_318 ();
 sg13g2_fill_2 FILLER_72_322 ();
 sg13g2_fill_2 FILLER_72_329 ();
 sg13g2_fill_1 FILLER_72_339 ();
 sg13g2_fill_1 FILLER_72_345 ();
 sg13g2_decap_4 FILLER_72_355 ();
 sg13g2_fill_2 FILLER_72_359 ();
 sg13g2_decap_4 FILLER_72_371 ();
 sg13g2_fill_2 FILLER_72_375 ();
 sg13g2_decap_8 FILLER_72_386 ();
 sg13g2_fill_1 FILLER_72_406 ();
 sg13g2_decap_4 FILLER_72_412 ();
 sg13g2_decap_8 FILLER_72_425 ();
 sg13g2_decap_4 FILLER_72_432 ();
 sg13g2_fill_1 FILLER_72_436 ();
 sg13g2_fill_1 FILLER_72_470 ();
 sg13g2_fill_2 FILLER_72_486 ();
 sg13g2_decap_8 FILLER_72_498 ();
 sg13g2_decap_8 FILLER_72_505 ();
 sg13g2_fill_2 FILLER_72_512 ();
 sg13g2_fill_2 FILLER_72_519 ();
 sg13g2_fill_1 FILLER_72_521 ();
 sg13g2_decap_8 FILLER_72_526 ();
 sg13g2_decap_8 FILLER_72_558 ();
 sg13g2_decap_8 FILLER_72_565 ();
 sg13g2_decap_8 FILLER_72_572 ();
 sg13g2_decap_4 FILLER_72_579 ();
 sg13g2_fill_1 FILLER_72_601 ();
 sg13g2_decap_8 FILLER_72_607 ();
 sg13g2_fill_2 FILLER_72_614 ();
 sg13g2_fill_1 FILLER_72_616 ();
 sg13g2_fill_2 FILLER_72_628 ();
 sg13g2_fill_1 FILLER_72_630 ();
 sg13g2_fill_1 FILLER_72_652 ();
 sg13g2_fill_2 FILLER_72_694 ();
 sg13g2_fill_2 FILLER_72_701 ();
 sg13g2_decap_8 FILLER_72_711 ();
 sg13g2_decap_8 FILLER_72_718 ();
 sg13g2_decap_4 FILLER_72_725 ();
 sg13g2_fill_1 FILLER_72_748 ();
 sg13g2_fill_2 FILLER_72_758 ();
 sg13g2_decap_4 FILLER_72_768 ();
 sg13g2_decap_8 FILLER_72_816 ();
 sg13g2_decap_8 FILLER_72_823 ();
 sg13g2_fill_2 FILLER_72_830 ();
 sg13g2_fill_1 FILLER_72_842 ();
 sg13g2_fill_2 FILLER_72_847 ();
 sg13g2_fill_2 FILLER_72_853 ();
 sg13g2_fill_2 FILLER_72_859 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_fill_2 FILLER_72_882 ();
 sg13g2_decap_8 FILLER_72_915 ();
 sg13g2_decap_4 FILLER_72_987 ();
 sg13g2_fill_1 FILLER_72_991 ();
 sg13g2_decap_8 FILLER_72_996 ();
 sg13g2_fill_2 FILLER_72_1027 ();
 sg13g2_fill_1 FILLER_72_1049 ();
 sg13g2_fill_2 FILLER_72_1055 ();
 sg13g2_fill_1 FILLER_72_1057 ();
 sg13g2_fill_1 FILLER_72_1089 ();
 sg13g2_fill_1 FILLER_72_1116 ();
 sg13g2_fill_2 FILLER_72_1126 ();
 sg13g2_decap_8 FILLER_72_1133 ();
 sg13g2_decap_8 FILLER_72_1140 ();
 sg13g2_fill_2 FILLER_72_1147 ();
 sg13g2_fill_1 FILLER_72_1149 ();
 sg13g2_decap_4 FILLER_72_1155 ();
 sg13g2_fill_1 FILLER_72_1168 ();
 sg13g2_fill_1 FILLER_72_1174 ();
 sg13g2_decap_8 FILLER_72_1205 ();
 sg13g2_decap_4 FILLER_72_1212 ();
 sg13g2_decap_4 FILLER_72_1221 ();
 sg13g2_fill_1 FILLER_72_1225 ();
 sg13g2_fill_1 FILLER_72_1241 ();
 sg13g2_fill_2 FILLER_72_1260 ();
 sg13g2_fill_2 FILLER_72_1267 ();
 sg13g2_fill_1 FILLER_72_1269 ();
 sg13g2_fill_1 FILLER_72_1275 ();
 sg13g2_decap_4 FILLER_72_1281 ();
 sg13g2_fill_2 FILLER_72_1298 ();
 sg13g2_fill_1 FILLER_72_1326 ();
 sg13g2_fill_1 FILLER_72_1331 ();
 sg13g2_fill_2 FILLER_72_1362 ();
 sg13g2_fill_1 FILLER_72_1364 ();
 sg13g2_fill_2 FILLER_72_1391 ();
 sg13g2_fill_1 FILLER_72_1424 ();
 sg13g2_fill_2 FILLER_72_1439 ();
 sg13g2_fill_2 FILLER_72_1485 ();
 sg13g2_fill_1 FILLER_72_1487 ();
 sg13g2_decap_4 FILLER_72_1493 ();
 sg13g2_fill_2 FILLER_72_1497 ();
 sg13g2_decap_8 FILLER_72_1503 ();
 sg13g2_decap_8 FILLER_72_1510 ();
 sg13g2_decap_8 FILLER_72_1517 ();
 sg13g2_decap_8 FILLER_72_1524 ();
 sg13g2_fill_1 FILLER_72_1531 ();
 sg13g2_fill_2 FILLER_72_1536 ();
 sg13g2_fill_1 FILLER_72_1542 ();
 sg13g2_fill_2 FILLER_72_1556 ();
 sg13g2_fill_1 FILLER_72_1558 ();
 sg13g2_decap_8 FILLER_72_1615 ();
 sg13g2_decap_8 FILLER_72_1622 ();
 sg13g2_decap_8 FILLER_72_1629 ();
 sg13g2_decap_8 FILLER_72_1636 ();
 sg13g2_decap_8 FILLER_72_1643 ();
 sg13g2_decap_8 FILLER_72_1650 ();
 sg13g2_decap_8 FILLER_72_1657 ();
 sg13g2_decap_8 FILLER_72_1664 ();
 sg13g2_decap_8 FILLER_72_1671 ();
 sg13g2_decap_8 FILLER_72_1678 ();
 sg13g2_decap_8 FILLER_72_1685 ();
 sg13g2_decap_8 FILLER_72_1692 ();
 sg13g2_decap_8 FILLER_72_1699 ();
 sg13g2_decap_8 FILLER_72_1706 ();
 sg13g2_decap_8 FILLER_72_1713 ();
 sg13g2_decap_8 FILLER_72_1720 ();
 sg13g2_decap_8 FILLER_72_1727 ();
 sg13g2_decap_8 FILLER_72_1734 ();
 sg13g2_decap_8 FILLER_72_1741 ();
 sg13g2_decap_8 FILLER_72_1748 ();
 sg13g2_decap_8 FILLER_72_1755 ();
 sg13g2_decap_8 FILLER_72_1762 ();
 sg13g2_decap_4 FILLER_72_1769 ();
 sg13g2_fill_1 FILLER_72_1773 ();
 sg13g2_fill_2 FILLER_73_26 ();
 sg13g2_fill_2 FILLER_73_32 ();
 sg13g2_fill_1 FILLER_73_34 ();
 sg13g2_fill_2 FILLER_73_44 ();
 sg13g2_fill_1 FILLER_73_60 ();
 sg13g2_decap_8 FILLER_73_71 ();
 sg13g2_fill_2 FILLER_73_78 ();
 sg13g2_fill_1 FILLER_73_80 ();
 sg13g2_decap_8 FILLER_73_96 ();
 sg13g2_decap_8 FILLER_73_103 ();
 sg13g2_decap_8 FILLER_73_110 ();
 sg13g2_decap_8 FILLER_73_117 ();
 sg13g2_decap_8 FILLER_73_124 ();
 sg13g2_fill_1 FILLER_73_131 ();
 sg13g2_decap_4 FILLER_73_136 ();
 sg13g2_decap_4 FILLER_73_145 ();
 sg13g2_fill_2 FILLER_73_149 ();
 sg13g2_fill_2 FILLER_73_172 ();
 sg13g2_fill_2 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_180 ();
 sg13g2_fill_2 FILLER_73_191 ();
 sg13g2_fill_1 FILLER_73_193 ();
 sg13g2_fill_1 FILLER_73_199 ();
 sg13g2_decap_8 FILLER_73_205 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_fill_1 FILLER_73_224 ();
 sg13g2_fill_2 FILLER_73_232 ();
 sg13g2_fill_1 FILLER_73_234 ();
 sg13g2_fill_1 FILLER_73_240 ();
 sg13g2_fill_1 FILLER_73_245 ();
 sg13g2_fill_1 FILLER_73_256 ();
 sg13g2_fill_1 FILLER_73_263 ();
 sg13g2_fill_1 FILLER_73_269 ();
 sg13g2_fill_1 FILLER_73_275 ();
 sg13g2_decap_4 FILLER_73_281 ();
 sg13g2_fill_2 FILLER_73_285 ();
 sg13g2_fill_2 FILLER_73_291 ();
 sg13g2_fill_1 FILLER_73_293 ();
 sg13g2_fill_2 FILLER_73_345 ();
 sg13g2_decap_4 FILLER_73_362 ();
 sg13g2_fill_2 FILLER_73_366 ();
 sg13g2_decap_8 FILLER_73_376 ();
 sg13g2_decap_8 FILLER_73_383 ();
 sg13g2_fill_2 FILLER_73_390 ();
 sg13g2_fill_1 FILLER_73_397 ();
 sg13g2_fill_2 FILLER_73_403 ();
 sg13g2_decap_8 FILLER_73_425 ();
 sg13g2_decap_8 FILLER_73_432 ();
 sg13g2_decap_4 FILLER_73_439 ();
 sg13g2_decap_8 FILLER_73_448 ();
 sg13g2_decap_4 FILLER_73_455 ();
 sg13g2_decap_8 FILLER_73_463 ();
 sg13g2_fill_2 FILLER_73_484 ();
 sg13g2_fill_2 FILLER_73_491 ();
 sg13g2_fill_1 FILLER_73_493 ();
 sg13g2_fill_2 FILLER_73_499 ();
 sg13g2_fill_1 FILLER_73_501 ();
 sg13g2_fill_2 FILLER_73_507 ();
 sg13g2_decap_8 FILLER_73_516 ();
 sg13g2_fill_2 FILLER_73_523 ();
 sg13g2_fill_1 FILLER_73_525 ();
 sg13g2_fill_1 FILLER_73_531 ();
 sg13g2_fill_2 FILLER_73_537 ();
 sg13g2_fill_1 FILLER_73_539 ();
 sg13g2_fill_1 FILLER_73_549 ();
 sg13g2_decap_4 FILLER_73_554 ();
 sg13g2_fill_1 FILLER_73_558 ();
 sg13g2_decap_4 FILLER_73_571 ();
 sg13g2_fill_1 FILLER_73_575 ();
 sg13g2_decap_8 FILLER_73_586 ();
 sg13g2_decap_4 FILLER_73_593 ();
 sg13g2_fill_1 FILLER_73_597 ();
 sg13g2_decap_8 FILLER_73_602 ();
 sg13g2_decap_8 FILLER_73_609 ();
 sg13g2_decap_4 FILLER_73_616 ();
 sg13g2_decap_8 FILLER_73_623 ();
 sg13g2_decap_8 FILLER_73_630 ();
 sg13g2_fill_1 FILLER_73_637 ();
 sg13g2_decap_8 FILLER_73_641 ();
 sg13g2_decap_8 FILLER_73_648 ();
 sg13g2_fill_1 FILLER_73_655 ();
 sg13g2_decap_8 FILLER_73_678 ();
 sg13g2_decap_4 FILLER_73_715 ();
 sg13g2_fill_1 FILLER_73_719 ();
 sg13g2_decap_8 FILLER_73_725 ();
 sg13g2_fill_2 FILLER_73_736 ();
 sg13g2_fill_1 FILLER_73_738 ();
 sg13g2_decap_8 FILLER_73_744 ();
 sg13g2_decap_8 FILLER_73_751 ();
 sg13g2_fill_2 FILLER_73_758 ();
 sg13g2_fill_1 FILLER_73_760 ();
 sg13g2_fill_2 FILLER_73_775 ();
 sg13g2_fill_1 FILLER_73_777 ();
 sg13g2_decap_8 FILLER_73_783 ();
 sg13g2_decap_4 FILLER_73_795 ();
 sg13g2_fill_2 FILLER_73_799 ();
 sg13g2_fill_2 FILLER_73_831 ();
 sg13g2_fill_1 FILLER_73_841 ();
 sg13g2_fill_1 FILLER_73_847 ();
 sg13g2_decap_8 FILLER_73_851 ();
 sg13g2_fill_2 FILLER_73_858 ();
 sg13g2_fill_1 FILLER_73_860 ();
 sg13g2_fill_2 FILLER_73_866 ();
 sg13g2_fill_1 FILLER_73_868 ();
 sg13g2_fill_2 FILLER_73_874 ();
 sg13g2_fill_2 FILLER_73_885 ();
 sg13g2_fill_1 FILLER_73_887 ();
 sg13g2_decap_8 FILLER_73_892 ();
 sg13g2_fill_2 FILLER_73_899 ();
 sg13g2_fill_1 FILLER_73_901 ();
 sg13g2_decap_8 FILLER_73_928 ();
 sg13g2_decap_8 FILLER_73_935 ();
 sg13g2_fill_2 FILLER_73_942 ();
 sg13g2_fill_1 FILLER_73_944 ();
 sg13g2_decap_4 FILLER_73_949 ();
 sg13g2_decap_8 FILLER_73_956 ();
 sg13g2_decap_8 FILLER_73_963 ();
 sg13g2_decap_8 FILLER_73_970 ();
 sg13g2_fill_2 FILLER_73_977 ();
 sg13g2_fill_1 FILLER_73_984 ();
 sg13g2_decap_8 FILLER_73_1011 ();
 sg13g2_fill_1 FILLER_73_1040 ();
 sg13g2_fill_1 FILLER_73_1046 ();
 sg13g2_fill_2 FILLER_73_1067 ();
 sg13g2_fill_1 FILLER_73_1069 ();
 sg13g2_fill_2 FILLER_73_1074 ();
 sg13g2_fill_1 FILLER_73_1076 ();
 sg13g2_fill_2 FILLER_73_1085 ();
 sg13g2_fill_1 FILLER_73_1087 ();
 sg13g2_decap_4 FILLER_73_1092 ();
 sg13g2_fill_1 FILLER_73_1096 ();
 sg13g2_fill_1 FILLER_73_1101 ();
 sg13g2_decap_8 FILLER_73_1106 ();
 sg13g2_fill_1 FILLER_73_1113 ();
 sg13g2_decap_4 FILLER_73_1124 ();
 sg13g2_decap_8 FILLER_73_1132 ();
 sg13g2_decap_8 FILLER_73_1139 ();
 sg13g2_decap_8 FILLER_73_1146 ();
 sg13g2_fill_2 FILLER_73_1153 ();
 sg13g2_fill_1 FILLER_73_1155 ();
 sg13g2_decap_8 FILLER_73_1176 ();
 sg13g2_fill_2 FILLER_73_1183 ();
 sg13g2_decap_4 FILLER_73_1194 ();
 sg13g2_fill_1 FILLER_73_1198 ();
 sg13g2_fill_2 FILLER_73_1208 ();
 sg13g2_decap_8 FILLER_73_1219 ();
 sg13g2_decap_8 FILLER_73_1226 ();
 sg13g2_decap_4 FILLER_73_1233 ();
 sg13g2_fill_2 FILLER_73_1247 ();
 sg13g2_fill_2 FILLER_73_1257 ();
 sg13g2_fill_1 FILLER_73_1259 ();
 sg13g2_fill_2 FILLER_73_1265 ();
 sg13g2_fill_1 FILLER_73_1267 ();
 sg13g2_fill_2 FILLER_73_1272 ();
 sg13g2_decap_4 FILLER_73_1304 ();
 sg13g2_fill_1 FILLER_73_1308 ();
 sg13g2_decap_4 FILLER_73_1314 ();
 sg13g2_fill_1 FILLER_73_1322 ();
 sg13g2_fill_1 FILLER_73_1349 ();
 sg13g2_decap_4 FILLER_73_1367 ();
 sg13g2_fill_1 FILLER_73_1371 ();
 sg13g2_fill_2 FILLER_73_1376 ();
 sg13g2_fill_1 FILLER_73_1408 ();
 sg13g2_fill_2 FILLER_73_1431 ();
 sg13g2_fill_1 FILLER_73_1450 ();
 sg13g2_fill_2 FILLER_73_1490 ();
 sg13g2_decap_8 FILLER_73_1522 ();
 sg13g2_fill_2 FILLER_73_1529 ();
 sg13g2_decap_8 FILLER_73_1557 ();
 sg13g2_fill_2 FILLER_73_1564 ();
 sg13g2_decap_8 FILLER_73_1570 ();
 sg13g2_decap_8 FILLER_73_1577 ();
 sg13g2_decap_8 FILLER_73_1584 ();
 sg13g2_decap_8 FILLER_73_1591 ();
 sg13g2_decap_8 FILLER_73_1598 ();
 sg13g2_decap_8 FILLER_73_1605 ();
 sg13g2_decap_8 FILLER_73_1612 ();
 sg13g2_decap_8 FILLER_73_1619 ();
 sg13g2_decap_8 FILLER_73_1626 ();
 sg13g2_decap_8 FILLER_73_1633 ();
 sg13g2_decap_8 FILLER_73_1640 ();
 sg13g2_decap_8 FILLER_73_1647 ();
 sg13g2_decap_8 FILLER_73_1654 ();
 sg13g2_decap_8 FILLER_73_1661 ();
 sg13g2_decap_8 FILLER_73_1668 ();
 sg13g2_decap_8 FILLER_73_1675 ();
 sg13g2_decap_8 FILLER_73_1682 ();
 sg13g2_decap_8 FILLER_73_1689 ();
 sg13g2_decap_8 FILLER_73_1696 ();
 sg13g2_decap_8 FILLER_73_1703 ();
 sg13g2_decap_8 FILLER_73_1710 ();
 sg13g2_decap_8 FILLER_73_1717 ();
 sg13g2_decap_8 FILLER_73_1724 ();
 sg13g2_decap_8 FILLER_73_1731 ();
 sg13g2_decap_8 FILLER_73_1738 ();
 sg13g2_decap_8 FILLER_73_1745 ();
 sg13g2_decap_8 FILLER_73_1752 ();
 sg13g2_decap_8 FILLER_73_1759 ();
 sg13g2_decap_8 FILLER_73_1766 ();
 sg13g2_fill_1 FILLER_73_1773 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_28 ();
 sg13g2_fill_1 FILLER_74_30 ();
 sg13g2_fill_1 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_40 ();
 sg13g2_decap_4 FILLER_74_51 ();
 sg13g2_fill_2 FILLER_74_55 ();
 sg13g2_decap_4 FILLER_74_72 ();
 sg13g2_fill_1 FILLER_74_76 ();
 sg13g2_fill_2 FILLER_74_111 ();
 sg13g2_fill_1 FILLER_74_113 ();
 sg13g2_decap_4 FILLER_74_128 ();
 sg13g2_decap_8 FILLER_74_137 ();
 sg13g2_decap_8 FILLER_74_144 ();
 sg13g2_decap_8 FILLER_74_151 ();
 sg13g2_decap_8 FILLER_74_163 ();
 sg13g2_decap_8 FILLER_74_170 ();
 sg13g2_decap_4 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_195 ();
 sg13g2_fill_1 FILLER_74_201 ();
 sg13g2_fill_2 FILLER_74_206 ();
 sg13g2_fill_1 FILLER_74_212 ();
 sg13g2_fill_2 FILLER_74_221 ();
 sg13g2_fill_2 FILLER_74_228 ();
 sg13g2_fill_1 FILLER_74_235 ();
 sg13g2_fill_2 FILLER_74_244 ();
 sg13g2_fill_2 FILLER_74_250 ();
 sg13g2_fill_1 FILLER_74_252 ();
 sg13g2_fill_1 FILLER_74_257 ();
 sg13g2_fill_2 FILLER_74_285 ();
 sg13g2_decap_4 FILLER_74_292 ();
 sg13g2_decap_4 FILLER_74_301 ();
 sg13g2_fill_2 FILLER_74_305 ();
 sg13g2_decap_8 FILLER_74_328 ();
 sg13g2_decap_8 FILLER_74_335 ();
 sg13g2_fill_2 FILLER_74_342 ();
 sg13g2_fill_1 FILLER_74_349 ();
 sg13g2_decap_4 FILLER_74_354 ();
 sg13g2_fill_2 FILLER_74_358 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_2 FILLER_74_397 ();
 sg13g2_fill_1 FILLER_74_399 ();
 sg13g2_fill_1 FILLER_74_414 ();
 sg13g2_fill_2 FILLER_74_418 ();
 sg13g2_fill_1 FILLER_74_433 ();
 sg13g2_fill_1 FILLER_74_442 ();
 sg13g2_fill_1 FILLER_74_453 ();
 sg13g2_fill_2 FILLER_74_459 ();
 sg13g2_fill_1 FILLER_74_461 ();
 sg13g2_fill_1 FILLER_74_474 ();
 sg13g2_fill_2 FILLER_74_480 ();
 sg13g2_fill_1 FILLER_74_482 ();
 sg13g2_fill_2 FILLER_74_487 ();
 sg13g2_fill_1 FILLER_74_494 ();
 sg13g2_fill_1 FILLER_74_503 ();
 sg13g2_fill_1 FILLER_74_509 ();
 sg13g2_fill_2 FILLER_74_515 ();
 sg13g2_fill_1 FILLER_74_549 ();
 sg13g2_fill_1 FILLER_74_554 ();
 sg13g2_decap_4 FILLER_74_564 ();
 sg13g2_fill_1 FILLER_74_568 ();
 sg13g2_fill_2 FILLER_74_575 ();
 sg13g2_fill_2 FILLER_74_582 ();
 sg13g2_decap_8 FILLER_74_588 ();
 sg13g2_decap_4 FILLER_74_595 ();
 sg13g2_fill_2 FILLER_74_599 ();
 sg13g2_decap_4 FILLER_74_606 ();
 sg13g2_fill_2 FILLER_74_610 ();
 sg13g2_fill_1 FILLER_74_638 ();
 sg13g2_decap_8 FILLER_74_675 ();
 sg13g2_decap_8 FILLER_74_682 ();
 sg13g2_fill_2 FILLER_74_689 ();
 sg13g2_decap_4 FILLER_74_695 ();
 sg13g2_decap_8 FILLER_74_703 ();
 sg13g2_decap_4 FILLER_74_710 ();
 sg13g2_decap_4 FILLER_74_719 ();
 sg13g2_fill_2 FILLER_74_727 ();
 sg13g2_fill_2 FILLER_74_769 ();
 sg13g2_decap_8 FILLER_74_802 ();
 sg13g2_decap_8 FILLER_74_813 ();
 sg13g2_decap_4 FILLER_74_820 ();
 sg13g2_fill_2 FILLER_74_824 ();
 sg13g2_fill_1 FILLER_74_907 ();
 sg13g2_decap_8 FILLER_74_912 ();
 sg13g2_fill_2 FILLER_74_919 ();
 sg13g2_fill_2 FILLER_74_925 ();
 sg13g2_fill_1 FILLER_74_927 ();
 sg13g2_fill_2 FILLER_74_968 ();
 sg13g2_fill_2 FILLER_74_987 ();
 sg13g2_fill_1 FILLER_74_989 ();
 sg13g2_decap_4 FILLER_74_1003 ();
 sg13g2_fill_1 FILLER_74_1007 ();
 sg13g2_decap_4 FILLER_74_1013 ();
 sg13g2_decap_4 FILLER_74_1027 ();
 sg13g2_decap_8 FILLER_74_1036 ();
 sg13g2_fill_1 FILLER_74_1073 ();
 sg13g2_decap_4 FILLER_74_1117 ();
 sg13g2_decap_8 FILLER_74_1151 ();
 sg13g2_fill_1 FILLER_74_1158 ();
 sg13g2_decap_4 FILLER_74_1169 ();
 sg13g2_decap_8 FILLER_74_1177 ();
 sg13g2_fill_1 FILLER_74_1184 ();
 sg13g2_decap_8 FILLER_74_1195 ();
 sg13g2_decap_4 FILLER_74_1221 ();
 sg13g2_fill_1 FILLER_74_1225 ();
 sg13g2_fill_1 FILLER_74_1239 ();
 sg13g2_fill_1 FILLER_74_1245 ();
 sg13g2_fill_1 FILLER_74_1251 ();
 sg13g2_fill_1 FILLER_74_1257 ();
 sg13g2_fill_1 FILLER_74_1262 ();
 sg13g2_fill_2 FILLER_74_1271 ();
 sg13g2_decap_4 FILLER_74_1278 ();
 sg13g2_fill_2 FILLER_74_1286 ();
 sg13g2_fill_1 FILLER_74_1288 ();
 sg13g2_fill_1 FILLER_74_1293 ();
 sg13g2_decap_8 FILLER_74_1304 ();
 sg13g2_fill_1 FILLER_74_1311 ();
 sg13g2_decap_8 FILLER_74_1316 ();
 sg13g2_fill_1 FILLER_74_1323 ();
 sg13g2_fill_2 FILLER_74_1329 ();
 sg13g2_decap_8 FILLER_74_1391 ();
 sg13g2_fill_2 FILLER_74_1398 ();
 sg13g2_fill_1 FILLER_74_1400 ();
 sg13g2_decap_4 FILLER_74_1407 ();
 sg13g2_fill_2 FILLER_74_1411 ();
 sg13g2_fill_1 FILLER_74_1478 ();
 sg13g2_fill_2 FILLER_74_1508 ();
 sg13g2_fill_1 FILLER_74_1510 ();
 sg13g2_decap_8 FILLER_74_1527 ();
 sg13g2_decap_4 FILLER_74_1538 ();
 sg13g2_fill_1 FILLER_74_1542 ();
 sg13g2_decap_8 FILLER_74_1546 ();
 sg13g2_decap_8 FILLER_74_1553 ();
 sg13g2_decap_8 FILLER_74_1560 ();
 sg13g2_decap_8 FILLER_74_1567 ();
 sg13g2_decap_8 FILLER_74_1574 ();
 sg13g2_decap_8 FILLER_74_1581 ();
 sg13g2_decap_8 FILLER_74_1588 ();
 sg13g2_decap_8 FILLER_74_1595 ();
 sg13g2_decap_8 FILLER_74_1602 ();
 sg13g2_decap_8 FILLER_74_1609 ();
 sg13g2_decap_8 FILLER_74_1616 ();
 sg13g2_decap_8 FILLER_74_1623 ();
 sg13g2_decap_8 FILLER_74_1630 ();
 sg13g2_decap_8 FILLER_74_1637 ();
 sg13g2_decap_8 FILLER_74_1644 ();
 sg13g2_decap_8 FILLER_74_1651 ();
 sg13g2_decap_8 FILLER_74_1658 ();
 sg13g2_decap_8 FILLER_74_1665 ();
 sg13g2_decap_8 FILLER_74_1672 ();
 sg13g2_decap_8 FILLER_74_1679 ();
 sg13g2_decap_8 FILLER_74_1686 ();
 sg13g2_decap_8 FILLER_74_1693 ();
 sg13g2_decap_8 FILLER_74_1700 ();
 sg13g2_decap_8 FILLER_74_1707 ();
 sg13g2_decap_8 FILLER_74_1714 ();
 sg13g2_decap_8 FILLER_74_1721 ();
 sg13g2_decap_8 FILLER_74_1728 ();
 sg13g2_decap_8 FILLER_74_1735 ();
 sg13g2_decap_8 FILLER_74_1742 ();
 sg13g2_decap_8 FILLER_74_1749 ();
 sg13g2_decap_8 FILLER_74_1756 ();
 sg13g2_decap_8 FILLER_74_1763 ();
 sg13g2_decap_4 FILLER_74_1770 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_7 ();
 sg13g2_decap_4 FILLER_75_13 ();
 sg13g2_fill_1 FILLER_75_17 ();
 sg13g2_decap_8 FILLER_75_22 ();
 sg13g2_fill_2 FILLER_75_29 ();
 sg13g2_decap_8 FILLER_75_53 ();
 sg13g2_decap_8 FILLER_75_60 ();
 sg13g2_decap_8 FILLER_75_67 ();
 sg13g2_decap_4 FILLER_75_74 ();
 sg13g2_fill_1 FILLER_75_87 ();
 sg13g2_decap_8 FILLER_75_92 ();
 sg13g2_decap_8 FILLER_75_99 ();
 sg13g2_fill_2 FILLER_75_106 ();
 sg13g2_fill_2 FILLER_75_117 ();
 sg13g2_decap_8 FILLER_75_136 ();
 sg13g2_fill_1 FILLER_75_143 ();
 sg13g2_decap_8 FILLER_75_148 ();
 sg13g2_fill_1 FILLER_75_155 ();
 sg13g2_decap_8 FILLER_75_170 ();
 sg13g2_fill_1 FILLER_75_177 ();
 sg13g2_decap_4 FILLER_75_187 ();
 sg13g2_fill_1 FILLER_75_191 ();
 sg13g2_fill_2 FILLER_75_196 ();
 sg13g2_decap_4 FILLER_75_212 ();
 sg13g2_fill_2 FILLER_75_216 ();
 sg13g2_fill_2 FILLER_75_227 ();
 sg13g2_fill_1 FILLER_75_244 ();
 sg13g2_fill_1 FILLER_75_253 ();
 sg13g2_fill_2 FILLER_75_265 ();
 sg13g2_decap_8 FILLER_75_272 ();
 sg13g2_decap_8 FILLER_75_279 ();
 sg13g2_decap_8 FILLER_75_286 ();
 sg13g2_decap_8 FILLER_75_293 ();
 sg13g2_decap_8 FILLER_75_300 ();
 sg13g2_decap_8 FILLER_75_307 ();
 sg13g2_decap_8 FILLER_75_314 ();
 sg13g2_decap_8 FILLER_75_321 ();
 sg13g2_decap_8 FILLER_75_328 ();
 sg13g2_decap_4 FILLER_75_335 ();
 sg13g2_fill_2 FILLER_75_339 ();
 sg13g2_fill_2 FILLER_75_349 ();
 sg13g2_fill_1 FILLER_75_351 ();
 sg13g2_decap_4 FILLER_75_356 ();
 sg13g2_fill_1 FILLER_75_360 ();
 sg13g2_fill_1 FILLER_75_368 ();
 sg13g2_fill_2 FILLER_75_383 ();
 sg13g2_decap_8 FILLER_75_390 ();
 sg13g2_decap_4 FILLER_75_397 ();
 sg13g2_fill_2 FILLER_75_401 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_fill_1 FILLER_75_409 ();
 sg13g2_fill_2 FILLER_75_415 ();
 sg13g2_fill_1 FILLER_75_432 ();
 sg13g2_decap_4 FILLER_75_439 ();
 sg13g2_fill_2 FILLER_75_448 ();
 sg13g2_fill_2 FILLER_75_456 ();
 sg13g2_fill_2 FILLER_75_468 ();
 sg13g2_fill_1 FILLER_75_470 ();
 sg13g2_fill_1 FILLER_75_479 ();
 sg13g2_decap_8 FILLER_75_484 ();
 sg13g2_decap_8 FILLER_75_500 ();
 sg13g2_decap_8 FILLER_75_507 ();
 sg13g2_decap_8 FILLER_75_514 ();
 sg13g2_fill_2 FILLER_75_521 ();
 sg13g2_fill_1 FILLER_75_523 ();
 sg13g2_decap_8 FILLER_75_529 ();
 sg13g2_fill_2 FILLER_75_536 ();
 sg13g2_fill_1 FILLER_75_538 ();
 sg13g2_decap_8 FILLER_75_548 ();
 sg13g2_fill_2 FILLER_75_555 ();
 sg13g2_decap_8 FILLER_75_561 ();
 sg13g2_decap_8 FILLER_75_568 ();
 sg13g2_decap_8 FILLER_75_575 ();
 sg13g2_decap_8 FILLER_75_587 ();
 sg13g2_fill_2 FILLER_75_594 ();
 sg13g2_fill_1 FILLER_75_596 ();
 sg13g2_fill_1 FILLER_75_623 ();
 sg13g2_fill_2 FILLER_75_642 ();
 sg13g2_decap_4 FILLER_75_661 ();
 sg13g2_fill_2 FILLER_75_665 ();
 sg13g2_decap_4 FILLER_75_672 ();
 sg13g2_decap_8 FILLER_75_680 ();
 sg13g2_decap_8 FILLER_75_687 ();
 sg13g2_fill_2 FILLER_75_694 ();
 sg13g2_fill_1 FILLER_75_711 ();
 sg13g2_decap_4 FILLER_75_716 ();
 sg13g2_decap_8 FILLER_75_725 ();
 sg13g2_decap_8 FILLER_75_732 ();
 sg13g2_decap_8 FILLER_75_739 ();
 sg13g2_decap_8 FILLER_75_750 ();
 sg13g2_decap_4 FILLER_75_757 ();
 sg13g2_fill_2 FILLER_75_761 ();
 sg13g2_fill_2 FILLER_75_768 ();
 sg13g2_fill_1 FILLER_75_770 ();
 sg13g2_decap_4 FILLER_75_775 ();
 sg13g2_fill_1 FILLER_75_779 ();
 sg13g2_fill_2 FILLER_75_784 ();
 sg13g2_decap_8 FILLER_75_851 ();
 sg13g2_fill_2 FILLER_75_858 ();
 sg13g2_fill_1 FILLER_75_860 ();
 sg13g2_fill_2 FILLER_75_866 ();
 sg13g2_fill_1 FILLER_75_868 ();
 sg13g2_fill_2 FILLER_75_960 ();
 sg13g2_fill_1 FILLER_75_976 ();
 sg13g2_fill_2 FILLER_75_982 ();
 sg13g2_decap_4 FILLER_75_1010 ();
 sg13g2_fill_1 FILLER_75_1014 ();
 sg13g2_decap_8 FILLER_75_1022 ();
 sg13g2_fill_1 FILLER_75_1029 ();
 sg13g2_fill_1 FILLER_75_1038 ();
 sg13g2_fill_2 FILLER_75_1054 ();
 sg13g2_fill_1 FILLER_75_1062 ();
 sg13g2_fill_1 FILLER_75_1068 ();
 sg13g2_fill_1 FILLER_75_1077 ();
 sg13g2_fill_2 FILLER_75_1083 ();
 sg13g2_fill_1 FILLER_75_1085 ();
 sg13g2_fill_2 FILLER_75_1091 ();
 sg13g2_fill_2 FILLER_75_1096 ();
 sg13g2_fill_2 FILLER_75_1102 ();
 sg13g2_fill_1 FILLER_75_1104 ();
 sg13g2_fill_1 FILLER_75_1115 ();
 sg13g2_decap_4 FILLER_75_1125 ();
 sg13g2_fill_1 FILLER_75_1129 ();
 sg13g2_decap_4 FILLER_75_1134 ();
 sg13g2_decap_4 FILLER_75_1147 ();
 sg13g2_fill_2 FILLER_75_1158 ();
 sg13g2_fill_1 FILLER_75_1160 ();
 sg13g2_fill_1 FILLER_75_1196 ();
 sg13g2_fill_2 FILLER_75_1220 ();
 sg13g2_decap_4 FILLER_75_1232 ();
 sg13g2_fill_2 FILLER_75_1236 ();
 sg13g2_fill_1 FILLER_75_1243 ();
 sg13g2_decap_8 FILLER_75_1247 ();
 sg13g2_decap_8 FILLER_75_1254 ();
 sg13g2_decap_8 FILLER_75_1282 ();
 sg13g2_fill_1 FILLER_75_1289 ();
 sg13g2_fill_1 FILLER_75_1294 ();
 sg13g2_decap_4 FILLER_75_1299 ();
 sg13g2_decap_8 FILLER_75_1337 ();
 sg13g2_decap_8 FILLER_75_1344 ();
 sg13g2_decap_8 FILLER_75_1351 ();
 sg13g2_decap_8 FILLER_75_1358 ();
 sg13g2_fill_2 FILLER_75_1365 ();
 sg13g2_fill_1 FILLER_75_1367 ();
 sg13g2_decap_8 FILLER_75_1407 ();
 sg13g2_decap_4 FILLER_75_1414 ();
 sg13g2_fill_1 FILLER_75_1418 ();
 sg13g2_fill_1 FILLER_75_1422 ();
 sg13g2_decap_8 FILLER_75_1427 ();
 sg13g2_decap_8 FILLER_75_1434 ();
 sg13g2_decap_8 FILLER_75_1441 ();
 sg13g2_decap_8 FILLER_75_1448 ();
 sg13g2_decap_4 FILLER_75_1459 ();
 sg13g2_decap_8 FILLER_75_1467 ();
 sg13g2_fill_2 FILLER_75_1503 ();
 sg13g2_fill_1 FILLER_75_1526 ();
 sg13g2_decap_8 FILLER_75_1553 ();
 sg13g2_decap_8 FILLER_75_1560 ();
 sg13g2_decap_8 FILLER_75_1567 ();
 sg13g2_decap_8 FILLER_75_1574 ();
 sg13g2_decap_8 FILLER_75_1581 ();
 sg13g2_decap_8 FILLER_75_1588 ();
 sg13g2_decap_8 FILLER_75_1595 ();
 sg13g2_decap_8 FILLER_75_1602 ();
 sg13g2_decap_8 FILLER_75_1609 ();
 sg13g2_decap_8 FILLER_75_1616 ();
 sg13g2_decap_8 FILLER_75_1623 ();
 sg13g2_decap_8 FILLER_75_1630 ();
 sg13g2_decap_8 FILLER_75_1637 ();
 sg13g2_decap_8 FILLER_75_1644 ();
 sg13g2_decap_8 FILLER_75_1651 ();
 sg13g2_decap_8 FILLER_75_1658 ();
 sg13g2_decap_8 FILLER_75_1665 ();
 sg13g2_decap_8 FILLER_75_1672 ();
 sg13g2_decap_8 FILLER_75_1679 ();
 sg13g2_decap_8 FILLER_75_1686 ();
 sg13g2_decap_8 FILLER_75_1693 ();
 sg13g2_decap_8 FILLER_75_1700 ();
 sg13g2_decap_8 FILLER_75_1707 ();
 sg13g2_decap_8 FILLER_75_1714 ();
 sg13g2_decap_8 FILLER_75_1721 ();
 sg13g2_decap_8 FILLER_75_1728 ();
 sg13g2_decap_8 FILLER_75_1735 ();
 sg13g2_decap_8 FILLER_75_1742 ();
 sg13g2_decap_8 FILLER_75_1749 ();
 sg13g2_decap_8 FILLER_75_1756 ();
 sg13g2_decap_8 FILLER_75_1763 ();
 sg13g2_decap_4 FILLER_75_1770 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_33 ();
 sg13g2_fill_2 FILLER_76_39 ();
 sg13g2_fill_2 FILLER_76_46 ();
 sg13g2_fill_1 FILLER_76_48 ();
 sg13g2_fill_2 FILLER_76_54 ();
 sg13g2_fill_1 FILLER_76_56 ();
 sg13g2_fill_2 FILLER_76_62 ();
 sg13g2_fill_1 FILLER_76_64 ();
 sg13g2_fill_1 FILLER_76_94 ();
 sg13g2_decap_4 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_109 ();
 sg13g2_fill_2 FILLER_76_114 ();
 sg13g2_fill_1 FILLER_76_116 ();
 sg13g2_fill_2 FILLER_76_131 ();
 sg13g2_fill_1 FILLER_76_158 ();
 sg13g2_fill_1 FILLER_76_164 ();
 sg13g2_fill_1 FILLER_76_169 ();
 sg13g2_fill_2 FILLER_76_208 ();
 sg13g2_fill_1 FILLER_76_219 ();
 sg13g2_fill_1 FILLER_76_233 ();
 sg13g2_fill_2 FILLER_76_278 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_fill_2 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_307 ();
 sg13g2_decap_4 FILLER_76_314 ();
 sg13g2_fill_2 FILLER_76_318 ();
 sg13g2_decap_8 FILLER_76_334 ();
 sg13g2_decap_4 FILLER_76_341 ();
 sg13g2_decap_8 FILLER_76_360 ();
 sg13g2_decap_8 FILLER_76_375 ();
 sg13g2_fill_1 FILLER_76_382 ();
 sg13g2_decap_4 FILLER_76_391 ();
 sg13g2_fill_2 FILLER_76_395 ();
 sg13g2_fill_1 FILLER_76_407 ();
 sg13g2_fill_2 FILLER_76_412 ();
 sg13g2_fill_2 FILLER_76_420 ();
 sg13g2_fill_2 FILLER_76_426 ();
 sg13g2_fill_1 FILLER_76_428 ();
 sg13g2_decap_8 FILLER_76_448 ();
 sg13g2_fill_2 FILLER_76_455 ();
 sg13g2_fill_1 FILLER_76_467 ();
 sg13g2_decap_4 FILLER_76_472 ();
 sg13g2_fill_2 FILLER_76_476 ();
 sg13g2_fill_1 FILLER_76_491 ();
 sg13g2_fill_1 FILLER_76_496 ();
 sg13g2_fill_1 FILLER_76_511 ();
 sg13g2_fill_2 FILLER_76_516 ();
 sg13g2_fill_1 FILLER_76_518 ();
 sg13g2_decap_4 FILLER_76_524 ();
 sg13g2_fill_2 FILLER_76_528 ();
 sg13g2_decap_8 FILLER_76_535 ();
 sg13g2_fill_1 FILLER_76_542 ();
 sg13g2_fill_1 FILLER_76_548 ();
 sg13g2_fill_2 FILLER_76_575 ();
 sg13g2_fill_1 FILLER_76_577 ();
 sg13g2_fill_2 FILLER_76_582 ();
 sg13g2_fill_2 FILLER_76_591 ();
 sg13g2_fill_1 FILLER_76_593 ();
 sg13g2_fill_2 FILLER_76_599 ();
 sg13g2_fill_2 FILLER_76_605 ();
 sg13g2_decap_4 FILLER_76_612 ();
 sg13g2_fill_2 FILLER_76_619 ();
 sg13g2_fill_1 FILLER_76_668 ();
 sg13g2_decap_8 FILLER_76_747 ();
 sg13g2_decap_4 FILLER_76_754 ();
 sg13g2_fill_1 FILLER_76_758 ();
 sg13g2_decap_8 FILLER_76_785 ();
 sg13g2_decap_8 FILLER_76_822 ();
 sg13g2_decap_4 FILLER_76_829 ();
 sg13g2_fill_1 FILLER_76_833 ();
 sg13g2_fill_1 FILLER_76_859 ();
 sg13g2_fill_1 FILLER_76_864 ();
 sg13g2_decap_4 FILLER_76_874 ();
 sg13g2_fill_2 FILLER_76_878 ();
 sg13g2_fill_1 FILLER_76_899 ();
 sg13g2_decap_4 FILLER_76_916 ();
 sg13g2_fill_2 FILLER_76_920 ();
 sg13g2_fill_2 FILLER_76_927 ();
 sg13g2_fill_1 FILLER_76_929 ();
 sg13g2_fill_1 FILLER_76_935 ();
 sg13g2_fill_2 FILLER_76_972 ();
 sg13g2_decap_8 FILLER_76_983 ();
 sg13g2_decap_8 FILLER_76_990 ();
 sg13g2_decap_4 FILLER_76_997 ();
 sg13g2_fill_2 FILLER_76_1008 ();
 sg13g2_fill_1 FILLER_76_1010 ();
 sg13g2_fill_2 FILLER_76_1016 ();
 sg13g2_fill_1 FILLER_76_1025 ();
 sg13g2_fill_1 FILLER_76_1040 ();
 sg13g2_fill_1 FILLER_76_1045 ();
 sg13g2_fill_1 FILLER_76_1051 ();
 sg13g2_fill_1 FILLER_76_1055 ();
 sg13g2_fill_2 FILLER_76_1069 ();
 sg13g2_fill_2 FILLER_76_1086 ();
 sg13g2_fill_2 FILLER_76_1097 ();
 sg13g2_fill_2 FILLER_76_1120 ();
 sg13g2_fill_1 FILLER_76_1122 ();
 sg13g2_decap_8 FILLER_76_1153 ();
 sg13g2_decap_8 FILLER_76_1160 ();
 sg13g2_decap_8 FILLER_76_1167 ();
 sg13g2_fill_2 FILLER_76_1174 ();
 sg13g2_fill_2 FILLER_76_1180 ();
 sg13g2_fill_1 FILLER_76_1182 ();
 sg13g2_decap_8 FILLER_76_1187 ();
 sg13g2_decap_4 FILLER_76_1194 ();
 sg13g2_fill_2 FILLER_76_1198 ();
 sg13g2_fill_1 FILLER_76_1204 ();
 sg13g2_fill_1 FILLER_76_1214 ();
 sg13g2_fill_2 FILLER_76_1220 ();
 sg13g2_decap_8 FILLER_76_1226 ();
 sg13g2_fill_2 FILLER_76_1233 ();
 sg13g2_fill_1 FILLER_76_1235 ();
 sg13g2_decap_8 FILLER_76_1250 ();
 sg13g2_decap_8 FILLER_76_1257 ();
 sg13g2_fill_2 FILLER_76_1269 ();
 sg13g2_decap_4 FILLER_76_1297 ();
 sg13g2_decap_8 FILLER_76_1306 ();
 sg13g2_fill_1 FILLER_76_1313 ();
 sg13g2_decap_8 FILLER_76_1318 ();
 sg13g2_decap_4 FILLER_76_1325 ();
 sg13g2_decap_8 FILLER_76_1333 ();
 sg13g2_fill_2 FILLER_76_1340 ();
 sg13g2_fill_2 FILLER_76_1356 ();
 sg13g2_fill_1 FILLER_76_1358 ();
 sg13g2_decap_8 FILLER_76_1363 ();
 sg13g2_decap_8 FILLER_76_1370 ();
 sg13g2_decap_8 FILLER_76_1377 ();
 sg13g2_decap_8 FILLER_76_1384 ();
 sg13g2_fill_1 FILLER_76_1391 ();
 sg13g2_decap_4 FILLER_76_1397 ();
 sg13g2_decap_8 FILLER_76_1415 ();
 sg13g2_fill_2 FILLER_76_1422 ();
 sg13g2_decap_8 FILLER_76_1443 ();
 sg13g2_decap_8 FILLER_76_1450 ();
 sg13g2_decap_4 FILLER_76_1457 ();
 sg13g2_fill_2 FILLER_76_1476 ();
 sg13g2_fill_1 FILLER_76_1478 ();
 sg13g2_decap_8 FILLER_76_1522 ();
 sg13g2_decap_8 FILLER_76_1529 ();
 sg13g2_decap_8 FILLER_76_1536 ();
 sg13g2_decap_8 FILLER_76_1543 ();
 sg13g2_decap_8 FILLER_76_1550 ();
 sg13g2_decap_8 FILLER_76_1557 ();
 sg13g2_decap_8 FILLER_76_1564 ();
 sg13g2_decap_8 FILLER_76_1571 ();
 sg13g2_decap_8 FILLER_76_1578 ();
 sg13g2_decap_8 FILLER_76_1585 ();
 sg13g2_decap_8 FILLER_76_1592 ();
 sg13g2_decap_8 FILLER_76_1599 ();
 sg13g2_decap_8 FILLER_76_1606 ();
 sg13g2_decap_8 FILLER_76_1613 ();
 sg13g2_decap_8 FILLER_76_1620 ();
 sg13g2_decap_8 FILLER_76_1627 ();
 sg13g2_decap_8 FILLER_76_1634 ();
 sg13g2_decap_8 FILLER_76_1641 ();
 sg13g2_decap_8 FILLER_76_1648 ();
 sg13g2_decap_8 FILLER_76_1655 ();
 sg13g2_decap_8 FILLER_76_1662 ();
 sg13g2_decap_8 FILLER_76_1669 ();
 sg13g2_decap_8 FILLER_76_1676 ();
 sg13g2_decap_8 FILLER_76_1683 ();
 sg13g2_decap_8 FILLER_76_1690 ();
 sg13g2_decap_8 FILLER_76_1697 ();
 sg13g2_decap_8 FILLER_76_1704 ();
 sg13g2_decap_8 FILLER_76_1711 ();
 sg13g2_decap_8 FILLER_76_1718 ();
 sg13g2_decap_8 FILLER_76_1725 ();
 sg13g2_decap_8 FILLER_76_1732 ();
 sg13g2_decap_8 FILLER_76_1739 ();
 sg13g2_decap_8 FILLER_76_1746 ();
 sg13g2_decap_8 FILLER_76_1753 ();
 sg13g2_decap_8 FILLER_76_1760 ();
 sg13g2_decap_8 FILLER_76_1767 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_4 FILLER_77_28 ();
 sg13g2_fill_1 FILLER_77_32 ();
 sg13g2_fill_1 FILLER_77_63 ();
 sg13g2_fill_2 FILLER_77_68 ();
 sg13g2_decap_8 FILLER_77_74 ();
 sg13g2_decap_4 FILLER_77_81 ();
 sg13g2_fill_1 FILLER_77_85 ();
 sg13g2_fill_1 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_101 ();
 sg13g2_decap_8 FILLER_77_108 ();
 sg13g2_decap_4 FILLER_77_115 ();
 sg13g2_decap_8 FILLER_77_124 ();
 sg13g2_fill_2 FILLER_77_131 ();
 sg13g2_fill_1 FILLER_77_133 ();
 sg13g2_fill_2 FILLER_77_138 ();
 sg13g2_fill_1 FILLER_77_140 ();
 sg13g2_fill_1 FILLER_77_175 ();
 sg13g2_fill_2 FILLER_77_203 ();
 sg13g2_fill_1 FILLER_77_228 ();
 sg13g2_fill_2 FILLER_77_264 ();
 sg13g2_fill_2 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_318 ();
 sg13g2_decap_4 FILLER_77_330 ();
 sg13g2_fill_1 FILLER_77_334 ();
 sg13g2_decap_4 FILLER_77_340 ();
 sg13g2_fill_1 FILLER_77_344 ();
 sg13g2_fill_2 FILLER_77_364 ();
 sg13g2_decap_4 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_390 ();
 sg13g2_decap_4 FILLER_77_397 ();
 sg13g2_decap_8 FILLER_77_416 ();
 sg13g2_decap_4 FILLER_77_423 ();
 sg13g2_fill_1 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_437 ();
 sg13g2_fill_1 FILLER_77_444 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_fill_1 FILLER_77_471 ();
 sg13g2_decap_8 FILLER_77_487 ();
 sg13g2_decap_4 FILLER_77_494 ();
 sg13g2_fill_1 FILLER_77_508 ();
 sg13g2_fill_1 FILLER_77_514 ();
 sg13g2_fill_1 FILLER_77_520 ();
 sg13g2_fill_1 FILLER_77_525 ();
 sg13g2_decap_4 FILLER_77_561 ();
 sg13g2_fill_1 FILLER_77_565 ();
 sg13g2_fill_2 FILLER_77_571 ();
 sg13g2_fill_1 FILLER_77_573 ();
 sg13g2_fill_2 FILLER_77_578 ();
 sg13g2_fill_1 FILLER_77_580 ();
 sg13g2_fill_2 FILLER_77_591 ();
 sg13g2_fill_1 FILLER_77_593 ();
 sg13g2_fill_1 FILLER_77_610 ();
 sg13g2_fill_1 FILLER_77_616 ();
 sg13g2_fill_2 FILLER_77_622 ();
 sg13g2_fill_1 FILLER_77_645 ();
 sg13g2_fill_2 FILLER_77_654 ();
 sg13g2_fill_1 FILLER_77_656 ();
 sg13g2_fill_2 FILLER_77_662 ();
 sg13g2_decap_4 FILLER_77_670 ();
 sg13g2_fill_2 FILLER_77_674 ();
 sg13g2_decap_8 FILLER_77_680 ();
 sg13g2_decap_8 FILLER_77_687 ();
 sg13g2_decap_8 FILLER_77_694 ();
 sg13g2_fill_2 FILLER_77_701 ();
 sg13g2_fill_1 FILLER_77_703 ();
 sg13g2_fill_1 FILLER_77_708 ();
 sg13g2_fill_2 FILLER_77_713 ();
 sg13g2_fill_1 FILLER_77_715 ();
 sg13g2_fill_1 FILLER_77_765 ();
 sg13g2_decap_8 FILLER_77_781 ();
 sg13g2_decap_8 FILLER_77_788 ();
 sg13g2_decap_8 FILLER_77_795 ();
 sg13g2_decap_4 FILLER_77_802 ();
 sg13g2_fill_1 FILLER_77_806 ();
 sg13g2_decap_8 FILLER_77_811 ();
 sg13g2_decap_8 FILLER_77_818 ();
 sg13g2_fill_2 FILLER_77_825 ();
 sg13g2_fill_1 FILLER_77_827 ();
 sg13g2_fill_1 FILLER_77_858 ();
 sg13g2_fill_2 FILLER_77_863 ();
 sg13g2_fill_1 FILLER_77_870 ();
 sg13g2_fill_2 FILLER_77_881 ();
 sg13g2_fill_2 FILLER_77_898 ();
 sg13g2_decap_4 FILLER_77_925 ();
 sg13g2_fill_2 FILLER_77_929 ();
 sg13g2_decap_4 FILLER_77_935 ();
 sg13g2_fill_1 FILLER_77_947 ();
 sg13g2_decap_4 FILLER_77_997 ();
 sg13g2_fill_1 FILLER_77_1001 ();
 sg13g2_decap_8 FILLER_77_1006 ();
 sg13g2_fill_1 FILLER_77_1013 ();
 sg13g2_fill_2 FILLER_77_1029 ();
 sg13g2_fill_2 FILLER_77_1036 ();
 sg13g2_fill_1 FILLER_77_1038 ();
 sg13g2_fill_2 FILLER_77_1044 ();
 sg13g2_fill_1 FILLER_77_1046 ();
 sg13g2_fill_2 FILLER_77_1052 ();
 sg13g2_fill_2 FILLER_77_1062 ();
 sg13g2_fill_2 FILLER_77_1101 ();
 sg13g2_fill_1 FILLER_77_1103 ();
 sg13g2_fill_2 FILLER_77_1109 ();
 sg13g2_decap_8 FILLER_77_1114 ();
 sg13g2_fill_2 FILLER_77_1121 ();
 sg13g2_decap_4 FILLER_77_1127 ();
 sg13g2_fill_2 FILLER_77_1140 ();
 sg13g2_fill_1 FILLER_77_1147 ();
 sg13g2_fill_2 FILLER_77_1151 ();
 sg13g2_fill_1 FILLER_77_1153 ();
 sg13g2_decap_8 FILLER_77_1199 ();
 sg13g2_fill_1 FILLER_77_1206 ();
 sg13g2_fill_1 FILLER_77_1231 ();
 sg13g2_decap_8 FILLER_77_1236 ();
 sg13g2_decap_4 FILLER_77_1243 ();
 sg13g2_decap_8 FILLER_77_1251 ();
 sg13g2_decap_8 FILLER_77_1258 ();
 sg13g2_decap_8 FILLER_77_1273 ();
 sg13g2_fill_1 FILLER_77_1280 ();
 sg13g2_fill_1 FILLER_77_1307 ();
 sg13g2_fill_2 FILLER_77_1312 ();
 sg13g2_fill_2 FILLER_77_1318 ();
 sg13g2_fill_1 FILLER_77_1346 ();
 sg13g2_decap_8 FILLER_77_1378 ();
 sg13g2_decap_8 FILLER_77_1385 ();
 sg13g2_fill_2 FILLER_77_1392 ();
 sg13g2_decap_8 FILLER_77_1420 ();
 sg13g2_fill_1 FILLER_77_1427 ();
 sg13g2_fill_2 FILLER_77_1454 ();
 sg13g2_decap_8 FILLER_77_1486 ();
 sg13g2_fill_1 FILLER_77_1493 ();
 sg13g2_decap_8 FILLER_77_1498 ();
 sg13g2_fill_2 FILLER_77_1505 ();
 sg13g2_decap_8 FILLER_77_1550 ();
 sg13g2_decap_8 FILLER_77_1557 ();
 sg13g2_decap_8 FILLER_77_1564 ();
 sg13g2_decap_8 FILLER_77_1571 ();
 sg13g2_decap_8 FILLER_77_1578 ();
 sg13g2_decap_8 FILLER_77_1585 ();
 sg13g2_decap_8 FILLER_77_1592 ();
 sg13g2_decap_8 FILLER_77_1599 ();
 sg13g2_decap_8 FILLER_77_1606 ();
 sg13g2_decap_8 FILLER_77_1613 ();
 sg13g2_decap_8 FILLER_77_1620 ();
 sg13g2_decap_8 FILLER_77_1627 ();
 sg13g2_decap_8 FILLER_77_1634 ();
 sg13g2_decap_8 FILLER_77_1641 ();
 sg13g2_decap_8 FILLER_77_1648 ();
 sg13g2_decap_8 FILLER_77_1655 ();
 sg13g2_decap_8 FILLER_77_1662 ();
 sg13g2_decap_8 FILLER_77_1669 ();
 sg13g2_decap_8 FILLER_77_1676 ();
 sg13g2_decap_8 FILLER_77_1683 ();
 sg13g2_decap_8 FILLER_77_1690 ();
 sg13g2_decap_8 FILLER_77_1697 ();
 sg13g2_decap_8 FILLER_77_1704 ();
 sg13g2_decap_8 FILLER_77_1711 ();
 sg13g2_decap_8 FILLER_77_1718 ();
 sg13g2_decap_8 FILLER_77_1725 ();
 sg13g2_decap_8 FILLER_77_1732 ();
 sg13g2_decap_8 FILLER_77_1739 ();
 sg13g2_decap_8 FILLER_77_1746 ();
 sg13g2_decap_8 FILLER_77_1753 ();
 sg13g2_decap_8 FILLER_77_1760 ();
 sg13g2_decap_8 FILLER_77_1767 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_4 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_43 ();
 sg13g2_decap_8 FILLER_78_50 ();
 sg13g2_decap_4 FILLER_78_57 ();
 sg13g2_fill_2 FILLER_78_61 ();
 sg13g2_fill_1 FILLER_78_93 ();
 sg13g2_decap_4 FILLER_78_103 ();
 sg13g2_fill_2 FILLER_78_146 ();
 sg13g2_fill_2 FILLER_78_185 ();
 sg13g2_fill_2 FILLER_78_255 ();
 sg13g2_decap_8 FILLER_78_302 ();
 sg13g2_fill_1 FILLER_78_309 ();
 sg13g2_fill_2 FILLER_78_314 ();
 sg13g2_fill_1 FILLER_78_354 ();
 sg13g2_decap_8 FILLER_78_365 ();
 sg13g2_fill_1 FILLER_78_372 ();
 sg13g2_fill_1 FILLER_78_377 ();
 sg13g2_decap_8 FILLER_78_388 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_4 FILLER_78_409 ();
 sg13g2_decap_8 FILLER_78_452 ();
 sg13g2_decap_8 FILLER_78_459 ();
 sg13g2_decap_8 FILLER_78_466 ();
 sg13g2_decap_8 FILLER_78_482 ();
 sg13g2_fill_2 FILLER_78_489 ();
 sg13g2_fill_1 FILLER_78_499 ();
 sg13g2_fill_1 FILLER_78_509 ();
 sg13g2_decap_8 FILLER_78_518 ();
 sg13g2_decap_8 FILLER_78_525 ();
 sg13g2_decap_8 FILLER_78_532 ();
 sg13g2_fill_1 FILLER_78_539 ();
 sg13g2_decap_8 FILLER_78_544 ();
 sg13g2_decap_4 FILLER_78_551 ();
 sg13g2_decap_8 FILLER_78_559 ();
 sg13g2_decap_4 FILLER_78_566 ();
 sg13g2_decap_4 FILLER_78_574 ();
 sg13g2_fill_1 FILLER_78_578 ();
 sg13g2_decap_8 FILLER_78_583 ();
 sg13g2_decap_4 FILLER_78_590 ();
 sg13g2_decap_4 FILLER_78_598 ();
 sg13g2_fill_1 FILLER_78_602 ();
 sg13g2_fill_1 FILLER_78_607 ();
 sg13g2_fill_1 FILLER_78_612 ();
 sg13g2_fill_1 FILLER_78_618 ();
 sg13g2_decap_4 FILLER_78_635 ();
 sg13g2_fill_1 FILLER_78_639 ();
 sg13g2_fill_1 FILLER_78_658 ();
 sg13g2_fill_1 FILLER_78_664 ();
 sg13g2_fill_1 FILLER_78_704 ();
 sg13g2_decap_8 FILLER_78_735 ();
 sg13g2_fill_2 FILLER_78_742 ();
 sg13g2_fill_2 FILLER_78_763 ();
 sg13g2_fill_2 FILLER_78_791 ();
 sg13g2_fill_2 FILLER_78_797 ();
 sg13g2_fill_1 FILLER_78_799 ();
 sg13g2_fill_2 FILLER_78_826 ();
 sg13g2_fill_1 FILLER_78_828 ();
 sg13g2_fill_2 FILLER_78_834 ();
 sg13g2_fill_1 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_842 ();
 sg13g2_decap_8 FILLER_78_849 ();
 sg13g2_decap_4 FILLER_78_869 ();
 sg13g2_decap_8 FILLER_78_887 ();
 sg13g2_decap_4 FILLER_78_894 ();
 sg13g2_fill_2 FILLER_78_898 ();
 sg13g2_fill_1 FILLER_78_947 ();
 sg13g2_decap_4 FILLER_78_967 ();
 sg13g2_decap_8 FILLER_78_975 ();
 sg13g2_decap_4 FILLER_78_982 ();
 sg13g2_fill_1 FILLER_78_986 ();
 sg13g2_decap_8 FILLER_78_992 ();
 sg13g2_decap_8 FILLER_78_999 ();
 sg13g2_decap_8 FILLER_78_1006 ();
 sg13g2_fill_2 FILLER_78_1049 ();
 sg13g2_fill_1 FILLER_78_1075 ();
 sg13g2_fill_1 FILLER_78_1116 ();
 sg13g2_fill_2 FILLER_78_1127 ();
 sg13g2_fill_1 FILLER_78_1129 ();
 sg13g2_fill_2 FILLER_78_1140 ();
 sg13g2_fill_2 FILLER_78_1158 ();
 sg13g2_fill_2 FILLER_78_1181 ();
 sg13g2_decap_8 FILLER_78_1198 ();
 sg13g2_fill_2 FILLER_78_1205 ();
 sg13g2_fill_2 FILLER_78_1217 ();
 sg13g2_decap_4 FILLER_78_1224 ();
 sg13g2_fill_2 FILLER_78_1233 ();
 sg13g2_decap_4 FILLER_78_1261 ();
 sg13g2_fill_1 FILLER_78_1291 ();
 sg13g2_fill_2 FILLER_78_1322 ();
 sg13g2_decap_8 FILLER_78_1328 ();
 sg13g2_decap_8 FILLER_78_1335 ();
 sg13g2_fill_2 FILLER_78_1342 ();
 sg13g2_fill_1 FILLER_78_1344 ();
 sg13g2_decap_8 FILLER_78_1357 ();
 sg13g2_decap_8 FILLER_78_1368 ();
 sg13g2_decap_8 FILLER_78_1375 ();
 sg13g2_fill_2 FILLER_78_1382 ();
 sg13g2_decap_8 FILLER_78_1392 ();
 sg13g2_fill_2 FILLER_78_1410 ();
 sg13g2_fill_1 FILLER_78_1417 ();
 sg13g2_decap_8 FILLER_78_1421 ();
 sg13g2_decap_8 FILLER_78_1428 ();
 sg13g2_decap_4 FILLER_78_1435 ();
 sg13g2_fill_2 FILLER_78_1439 ();
 sg13g2_decap_8 FILLER_78_1453 ();
 sg13g2_decap_8 FILLER_78_1460 ();
 sg13g2_decap_8 FILLER_78_1467 ();
 sg13g2_decap_4 FILLER_78_1474 ();
 sg13g2_decap_4 FILLER_78_1503 ();
 sg13g2_fill_2 FILLER_78_1507 ();
 sg13g2_decap_8 FILLER_78_1513 ();
 sg13g2_decap_4 FILLER_78_1524 ();
 sg13g2_fill_2 FILLER_78_1528 ();
 sg13g2_decap_8 FILLER_78_1534 ();
 sg13g2_decap_8 FILLER_78_1541 ();
 sg13g2_decap_8 FILLER_78_1548 ();
 sg13g2_decap_8 FILLER_78_1555 ();
 sg13g2_decap_8 FILLER_78_1562 ();
 sg13g2_decap_8 FILLER_78_1569 ();
 sg13g2_decap_8 FILLER_78_1576 ();
 sg13g2_decap_8 FILLER_78_1583 ();
 sg13g2_decap_8 FILLER_78_1590 ();
 sg13g2_decap_8 FILLER_78_1597 ();
 sg13g2_decap_8 FILLER_78_1604 ();
 sg13g2_decap_8 FILLER_78_1611 ();
 sg13g2_decap_8 FILLER_78_1618 ();
 sg13g2_decap_8 FILLER_78_1625 ();
 sg13g2_decap_8 FILLER_78_1632 ();
 sg13g2_decap_8 FILLER_78_1639 ();
 sg13g2_decap_8 FILLER_78_1646 ();
 sg13g2_decap_8 FILLER_78_1653 ();
 sg13g2_decap_8 FILLER_78_1660 ();
 sg13g2_decap_8 FILLER_78_1667 ();
 sg13g2_decap_8 FILLER_78_1674 ();
 sg13g2_decap_8 FILLER_78_1681 ();
 sg13g2_decap_8 FILLER_78_1688 ();
 sg13g2_decap_8 FILLER_78_1695 ();
 sg13g2_decap_8 FILLER_78_1702 ();
 sg13g2_decap_8 FILLER_78_1709 ();
 sg13g2_decap_8 FILLER_78_1716 ();
 sg13g2_decap_8 FILLER_78_1723 ();
 sg13g2_decap_8 FILLER_78_1730 ();
 sg13g2_decap_8 FILLER_78_1737 ();
 sg13g2_decap_8 FILLER_78_1744 ();
 sg13g2_decap_8 FILLER_78_1751 ();
 sg13g2_decap_8 FILLER_78_1758 ();
 sg13g2_decap_8 FILLER_78_1765 ();
 sg13g2_fill_2 FILLER_78_1772 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_fill_1 FILLER_79_84 ();
 sg13g2_fill_1 FILLER_79_128 ();
 sg13g2_fill_1 FILLER_79_133 ();
 sg13g2_fill_1 FILLER_79_146 ();
 sg13g2_fill_1 FILLER_79_184 ();
 sg13g2_fill_1 FILLER_79_192 ();
 sg13g2_fill_1 FILLER_79_219 ();
 sg13g2_fill_1 FILLER_79_228 ();
 sg13g2_fill_2 FILLER_79_236 ();
 sg13g2_fill_1 FILLER_79_262 ();
 sg13g2_fill_2 FILLER_79_339 ();
 sg13g2_fill_1 FILLER_79_345 ();
 sg13g2_fill_1 FILLER_79_350 ();
 sg13g2_fill_2 FILLER_79_355 ();
 sg13g2_fill_2 FILLER_79_362 ();
 sg13g2_fill_1 FILLER_79_364 ();
 sg13g2_fill_2 FILLER_79_369 ();
 sg13g2_fill_1 FILLER_79_371 ();
 sg13g2_fill_2 FILLER_79_376 ();
 sg13g2_fill_1 FILLER_79_378 ();
 sg13g2_fill_2 FILLER_79_418 ();
 sg13g2_fill_1 FILLER_79_420 ();
 sg13g2_fill_2 FILLER_79_425 ();
 sg13g2_fill_1 FILLER_79_427 ();
 sg13g2_decap_4 FILLER_79_432 ();
 sg13g2_decap_8 FILLER_79_440 ();
 sg13g2_fill_2 FILLER_79_456 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_fill_2 FILLER_79_469 ();
 sg13g2_fill_1 FILLER_79_471 ();
 sg13g2_fill_2 FILLER_79_498 ();
 sg13g2_fill_1 FILLER_79_518 ();
 sg13g2_fill_2 FILLER_79_523 ();
 sg13g2_fill_1 FILLER_79_525 ();
 sg13g2_decap_4 FILLER_79_531 ();
 sg13g2_fill_1 FILLER_79_535 ();
 sg13g2_decap_4 FILLER_79_540 ();
 sg13g2_decap_8 FILLER_79_574 ();
 sg13g2_decap_4 FILLER_79_611 ();
 sg13g2_decap_4 FILLER_79_619 ();
 sg13g2_decap_4 FILLER_79_638 ();
 sg13g2_fill_2 FILLER_79_648 ();
 sg13g2_decap_8 FILLER_79_654 ();
 sg13g2_decap_4 FILLER_79_665 ();
 sg13g2_fill_2 FILLER_79_669 ();
 sg13g2_decap_4 FILLER_79_676 ();
 sg13g2_fill_1 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_690 ();
 sg13g2_fill_2 FILLER_79_697 ();
 sg13g2_fill_1 FILLER_79_699 ();
 sg13g2_fill_1 FILLER_79_715 ();
 sg13g2_fill_2 FILLER_79_720 ();
 sg13g2_decap_8 FILLER_79_726 ();
 sg13g2_decap_4 FILLER_79_733 ();
 sg13g2_fill_2 FILLER_79_737 ();
 sg13g2_decap_4 FILLER_79_765 ();
 sg13g2_fill_1 FILLER_79_769 ();
 sg13g2_fill_2 FILLER_79_774 ();
 sg13g2_fill_2 FILLER_79_780 ();
 sg13g2_fill_2 FILLER_79_786 ();
 sg13g2_fill_1 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_794 ();
 sg13g2_fill_2 FILLER_79_801 ();
 sg13g2_fill_1 FILLER_79_803 ();
 sg13g2_fill_1 FILLER_79_829 ();
 sg13g2_fill_1 FILLER_79_872 ();
 sg13g2_decap_8 FILLER_79_878 ();
 sg13g2_fill_1 FILLER_79_885 ();
 sg13g2_decap_4 FILLER_79_890 ();
 sg13g2_decap_8 FILLER_79_899 ();
 sg13g2_fill_1 FILLER_79_906 ();
 sg13g2_fill_1 FILLER_79_913 ();
 sg13g2_decap_4 FILLER_79_920 ();
 sg13g2_fill_1 FILLER_79_924 ();
 sg13g2_fill_2 FILLER_79_929 ();
 sg13g2_decap_4 FILLER_79_935 ();
 sg13g2_fill_2 FILLER_79_939 ();
 sg13g2_fill_1 FILLER_79_954 ();
 sg13g2_decap_8 FILLER_79_969 ();
 sg13g2_fill_1 FILLER_79_976 ();
 sg13g2_decap_4 FILLER_79_1033 ();
 sg13g2_fill_2 FILLER_79_1037 ();
 sg13g2_decap_4 FILLER_79_1044 ();
 sg13g2_decap_4 FILLER_79_1053 ();
 sg13g2_fill_1 FILLER_79_1057 ();
 sg13g2_fill_2 FILLER_79_1062 ();
 sg13g2_fill_1 FILLER_79_1079 ();
 sg13g2_fill_2 FILLER_79_1089 ();
 sg13g2_decap_8 FILLER_79_1095 ();
 sg13g2_decap_4 FILLER_79_1102 ();
 sg13g2_fill_2 FILLER_79_1106 ();
 sg13g2_decap_8 FILLER_79_1111 ();
 sg13g2_fill_2 FILLER_79_1118 ();
 sg13g2_fill_2 FILLER_79_1135 ();
 sg13g2_decap_8 FILLER_79_1141 ();
 sg13g2_fill_1 FILLER_79_1148 ();
 sg13g2_fill_2 FILLER_79_1173 ();
 sg13g2_fill_1 FILLER_79_1175 ();
 sg13g2_decap_8 FILLER_79_1180 ();
 sg13g2_fill_2 FILLER_79_1187 ();
 sg13g2_fill_1 FILLER_79_1189 ();
 sg13g2_fill_2 FILLER_79_1205 ();
 sg13g2_fill_1 FILLER_79_1207 ();
 sg13g2_decap_4 FILLER_79_1212 ();
 sg13g2_fill_2 FILLER_79_1230 ();
 sg13g2_fill_1 FILLER_79_1232 ();
 sg13g2_decap_4 FILLER_79_1238 ();
 sg13g2_fill_2 FILLER_79_1242 ();
 sg13g2_decap_4 FILLER_79_1248 ();
 sg13g2_decap_8 FILLER_79_1256 ();
 sg13g2_decap_8 FILLER_79_1263 ();
 sg13g2_fill_2 FILLER_79_1274 ();
 sg13g2_decap_8 FILLER_79_1280 ();
 sg13g2_decap_4 FILLER_79_1287 ();
 sg13g2_decap_8 FILLER_79_1295 ();
 sg13g2_decap_8 FILLER_79_1302 ();
 sg13g2_decap_4 FILLER_79_1309 ();
 sg13g2_fill_1 FILLER_79_1313 ();
 sg13g2_fill_1 FILLER_79_1318 ();
 sg13g2_decap_4 FILLER_79_1354 ();
 sg13g2_fill_1 FILLER_79_1358 ();
 sg13g2_decap_4 FILLER_79_1393 ();
 sg13g2_fill_2 FILLER_79_1397 ();
 sg13g2_decap_4 FILLER_79_1403 ();
 sg13g2_decap_4 FILLER_79_1423 ();
 sg13g2_fill_2 FILLER_79_1427 ();
 sg13g2_fill_2 FILLER_79_1476 ();
 sg13g2_fill_1 FILLER_79_1478 ();
 sg13g2_decap_8 FILLER_79_1483 ();
 sg13g2_decap_4 FILLER_79_1490 ();
 sg13g2_fill_2 FILLER_79_1494 ();
 sg13g2_decap_8 FILLER_79_1500 ();
 sg13g2_decap_8 FILLER_79_1507 ();
 sg13g2_decap_8 FILLER_79_1514 ();
 sg13g2_decap_8 FILLER_79_1521 ();
 sg13g2_decap_8 FILLER_79_1528 ();
 sg13g2_decap_8 FILLER_79_1535 ();
 sg13g2_decap_8 FILLER_79_1542 ();
 sg13g2_decap_8 FILLER_79_1549 ();
 sg13g2_decap_8 FILLER_79_1556 ();
 sg13g2_decap_8 FILLER_79_1563 ();
 sg13g2_decap_8 FILLER_79_1570 ();
 sg13g2_decap_8 FILLER_79_1577 ();
 sg13g2_decap_8 FILLER_79_1584 ();
 sg13g2_decap_8 FILLER_79_1591 ();
 sg13g2_decap_8 FILLER_79_1598 ();
 sg13g2_decap_8 FILLER_79_1605 ();
 sg13g2_decap_8 FILLER_79_1612 ();
 sg13g2_decap_8 FILLER_79_1619 ();
 sg13g2_decap_8 FILLER_79_1626 ();
 sg13g2_decap_8 FILLER_79_1633 ();
 sg13g2_decap_8 FILLER_79_1640 ();
 sg13g2_decap_8 FILLER_79_1647 ();
 sg13g2_decap_8 FILLER_79_1654 ();
 sg13g2_decap_8 FILLER_79_1661 ();
 sg13g2_decap_8 FILLER_79_1668 ();
 sg13g2_decap_8 FILLER_79_1675 ();
 sg13g2_decap_8 FILLER_79_1682 ();
 sg13g2_decap_8 FILLER_79_1689 ();
 sg13g2_decap_8 FILLER_79_1696 ();
 sg13g2_decap_8 FILLER_79_1703 ();
 sg13g2_decap_8 FILLER_79_1710 ();
 sg13g2_decap_8 FILLER_79_1717 ();
 sg13g2_decap_8 FILLER_79_1724 ();
 sg13g2_decap_8 FILLER_79_1731 ();
 sg13g2_decap_8 FILLER_79_1738 ();
 sg13g2_decap_8 FILLER_79_1745 ();
 sg13g2_decap_8 FILLER_79_1752 ();
 sg13g2_decap_8 FILLER_79_1759 ();
 sg13g2_decap_8 FILLER_79_1766 ();
 sg13g2_fill_1 FILLER_79_1773 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_1 FILLER_80_70 ();
 sg13g2_decap_4 FILLER_80_87 ();
 sg13g2_fill_1 FILLER_80_161 ();
 sg13g2_fill_2 FILLER_80_286 ();
 sg13g2_fill_2 FILLER_80_295 ();
 sg13g2_fill_2 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_315 ();
 sg13g2_decap_8 FILLER_80_350 ();
 sg13g2_fill_1 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_4 FILLER_80_400 ();
 sg13g2_fill_2 FILLER_80_404 ();
 sg13g2_decap_8 FILLER_80_440 ();
 sg13g2_fill_1 FILLER_80_477 ();
 sg13g2_decap_8 FILLER_80_482 ();
 sg13g2_decap_8 FILLER_80_489 ();
 sg13g2_decap_4 FILLER_80_496 ();
 sg13g2_decap_4 FILLER_80_526 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_decap_8 FILLER_80_563 ();
 sg13g2_decap_8 FILLER_80_570 ();
 sg13g2_decap_8 FILLER_80_577 ();
 sg13g2_fill_1 FILLER_80_584 ();
 sg13g2_decap_8 FILLER_80_589 ();
 sg13g2_decap_4 FILLER_80_596 ();
 sg13g2_decap_8 FILLER_80_604 ();
 sg13g2_fill_1 FILLER_80_611 ();
 sg13g2_decap_8 FILLER_80_642 ();
 sg13g2_fill_2 FILLER_80_649 ();
 sg13g2_fill_1 FILLER_80_651 ();
 sg13g2_decap_8 FILLER_80_678 ();
 sg13g2_decap_8 FILLER_80_685 ();
 sg13g2_decap_4 FILLER_80_692 ();
 sg13g2_fill_1 FILLER_80_696 ();
 sg13g2_decap_8 FILLER_80_738 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_fill_1 FILLER_80_770 ();
 sg13g2_decap_4 FILLER_80_797 ();
 sg13g2_fill_2 FILLER_80_827 ();
 sg13g2_decap_8 FILLER_80_832 ();
 sg13g2_fill_2 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_845 ();
 sg13g2_decap_8 FILLER_80_852 ();
 sg13g2_decap_4 FILLER_80_859 ();
 sg13g2_fill_1 FILLER_80_863 ();
 sg13g2_decap_8 FILLER_80_890 ();
 sg13g2_fill_2 FILLER_80_897 ();
 sg13g2_fill_2 FILLER_80_951 ();
 sg13g2_decap_4 FILLER_80_979 ();
 sg13g2_fill_1 FILLER_80_987 ();
 sg13g2_decap_8 FILLER_80_992 ();
 sg13g2_decap_8 FILLER_80_999 ();
 sg13g2_fill_2 FILLER_80_1006 ();
 sg13g2_fill_1 FILLER_80_1008 ();
 sg13g2_decap_8 FILLER_80_1013 ();
 sg13g2_decap_8 FILLER_80_1020 ();
 sg13g2_decap_8 FILLER_80_1027 ();
 sg13g2_decap_8 FILLER_80_1034 ();
 sg13g2_decap_4 FILLER_80_1041 ();
 sg13g2_fill_2 FILLER_80_1045 ();
 sg13g2_fill_2 FILLER_80_1079 ();
 sg13g2_decap_8 FILLER_80_1111 ();
 sg13g2_decap_8 FILLER_80_1118 ();
 sg13g2_fill_2 FILLER_80_1125 ();
 sg13g2_decap_8 FILLER_80_1153 ();
 sg13g2_decap_4 FILLER_80_1160 ();
 sg13g2_fill_1 FILLER_80_1164 ();
 sg13g2_decap_4 FILLER_80_1195 ();
 sg13g2_fill_2 FILLER_80_1199 ();
 sg13g2_decap_4 FILLER_80_1227 ();
 sg13g2_fill_2 FILLER_80_1231 ();
 sg13g2_decap_4 FILLER_80_1237 ();
 sg13g2_fill_2 FILLER_80_1267 ();
 sg13g2_fill_1 FILLER_80_1269 ();
 sg13g2_decap_8 FILLER_80_1296 ();
 sg13g2_decap_8 FILLER_80_1303 ();
 sg13g2_decap_8 FILLER_80_1310 ();
 sg13g2_decap_8 FILLER_80_1317 ();
 sg13g2_decap_4 FILLER_80_1324 ();
 sg13g2_decap_8 FILLER_80_1332 ();
 sg13g2_decap_4 FILLER_80_1339 ();
 sg13g2_decap_8 FILLER_80_1355 ();
 sg13g2_decap_4 FILLER_80_1362 ();
 sg13g2_fill_2 FILLER_80_1366 ();
 sg13g2_decap_8 FILLER_80_1372 ();
 sg13g2_decap_4 FILLER_80_1379 ();
 sg13g2_decap_8 FILLER_80_1425 ();
 sg13g2_fill_2 FILLER_80_1432 ();
 sg13g2_fill_1 FILLER_80_1434 ();
 sg13g2_fill_1 FILLER_80_1439 ();
 sg13g2_fill_2 FILLER_80_1445 ();
 sg13g2_fill_2 FILLER_80_1454 ();
 sg13g2_decap_8 FILLER_80_1460 ();
 sg13g2_decap_8 FILLER_80_1467 ();
 sg13g2_decap_4 FILLER_80_1474 ();
 sg13g2_fill_2 FILLER_80_1478 ();
 sg13g2_decap_8 FILLER_80_1510 ();
 sg13g2_decap_8 FILLER_80_1517 ();
 sg13g2_decap_8 FILLER_80_1524 ();
 sg13g2_decap_8 FILLER_80_1531 ();
 sg13g2_decap_8 FILLER_80_1538 ();
 sg13g2_decap_8 FILLER_80_1545 ();
 sg13g2_decap_8 FILLER_80_1552 ();
 sg13g2_decap_8 FILLER_80_1559 ();
 sg13g2_decap_8 FILLER_80_1566 ();
 sg13g2_decap_8 FILLER_80_1573 ();
 sg13g2_decap_8 FILLER_80_1580 ();
 sg13g2_decap_8 FILLER_80_1587 ();
 sg13g2_decap_8 FILLER_80_1594 ();
 sg13g2_decap_8 FILLER_80_1601 ();
 sg13g2_decap_8 FILLER_80_1608 ();
 sg13g2_decap_8 FILLER_80_1615 ();
 sg13g2_decap_8 FILLER_80_1622 ();
 sg13g2_decap_8 FILLER_80_1629 ();
 sg13g2_decap_8 FILLER_80_1636 ();
 sg13g2_decap_8 FILLER_80_1643 ();
 sg13g2_decap_8 FILLER_80_1650 ();
 sg13g2_decap_8 FILLER_80_1657 ();
 sg13g2_decap_8 FILLER_80_1664 ();
 sg13g2_decap_8 FILLER_80_1671 ();
 sg13g2_decap_8 FILLER_80_1678 ();
 sg13g2_decap_8 FILLER_80_1685 ();
 sg13g2_decap_8 FILLER_80_1692 ();
 sg13g2_decap_8 FILLER_80_1699 ();
 sg13g2_decap_8 FILLER_80_1706 ();
 sg13g2_decap_8 FILLER_80_1713 ();
 sg13g2_decap_8 FILLER_80_1720 ();
 sg13g2_decap_8 FILLER_80_1727 ();
 sg13g2_decap_8 FILLER_80_1734 ();
 sg13g2_decap_8 FILLER_80_1741 ();
 sg13g2_decap_8 FILLER_80_1748 ();
 sg13g2_decap_8 FILLER_80_1755 ();
 sg13g2_decap_8 FILLER_80_1762 ();
 sg13g2_decap_4 FILLER_80_1769 ();
 sg13g2_fill_1 FILLER_80_1773 ();
endmodule
